magic
tech sky130A
magscale 1 2
timestamp 1605730173
<< checkpaint >>
rect -1260 -1260 586176 705260
<< locali >>
rect 288761 700859 288795 701029
rect 229605 699771 229639 699873
rect 239265 699703 239299 699873
rect 259229 699703 259263 699873
rect 264105 699703 264139 699873
rect 278549 699703 278583 699941
rect 278641 699703 278675 699873
rect 287381 699771 287415 699941
rect 290049 699907 290083 701097
rect 292383 700961 292533 700995
rect 296305 700927 296339 701097
rect 292291 700825 292475 700859
rect 292257 699839 292291 700213
rect 292349 700043 292383 700213
rect 292441 700043 292475 700825
rect 294591 699941 294741 699975
rect 296121 699839 296155 700009
rect 296213 699907 296247 700893
rect 292257 699805 292625 699839
rect 287381 699737 287473 699771
rect 288853 699737 289037 699771
rect 291613 699737 291889 699771
rect 288853 699703 288887 699737
rect 291613 699703 291647 699737
rect 378737 685899 378771 695453
rect 508457 685899 508491 695453
rect 314153 666587 314187 676073
rect 378645 666587 378679 676073
rect 443873 666587 443907 676073
rect 508365 666587 508399 676073
rect 573593 666587 573627 676073
rect 314153 627963 314187 637449
rect 443873 627963 443907 637449
rect 573593 627963 573627 637449
rect 443689 601579 443723 608549
rect 573409 601579 573443 608549
rect 313877 589339 313911 598825
rect 443873 589339 443907 598825
rect 573593 589339 573627 598825
rect 378645 579683 378679 589237
rect 508365 579683 508399 589237
rect 313969 570027 314003 579581
rect 378737 562955 378771 569857
rect 508457 562955 508491 569857
rect 443505 550647 443539 553401
rect 573225 550647 573259 553401
rect 443505 531335 443539 534089
rect 573225 531335 573259 534089
rect 443597 524331 443631 531233
rect 573317 524331 573351 531233
rect 443505 485707 443539 485877
rect 573225 485707 573259 485877
rect 268889 463131 268923 463641
rect 283701 463063 283735 463233
rect 284713 463233 284897 463267
rect 284713 463199 284747 463233
rect 291613 462179 291647 463097
rect 292625 462315 292659 463097
rect 301273 462179 301307 463097
rect 302285 462247 302319 463165
rect 302929 462179 302963 463709
rect 443597 463199 443631 471937
rect 573317 463063 573351 471937
rect 225373 459867 225407 460037
rect 7333 459527 7367 459765
rect 7425 459595 7459 459765
rect 16993 459595 17027 459765
rect 17085 459595 17119 459765
rect 26653 459527 26687 459765
rect 26745 459595 26779 459765
rect 36313 459595 36347 459765
rect 36405 459595 36439 459765
rect 45973 459527 46007 459765
rect 46065 459595 46099 459765
rect 55633 459595 55667 459765
rect 55725 459595 55759 459765
rect 65293 459527 65327 459765
rect 65385 459595 65419 459765
rect 74953 459595 74987 459765
rect 75045 459595 75079 459765
rect 84613 459527 84647 459765
rect 84705 459595 84739 459765
rect 94273 459595 94307 459765
rect 94365 459595 94399 459765
rect 103933 459527 103967 459765
rect 104025 459595 104059 459765
rect 113593 459595 113627 459765
rect 113685 459595 113719 459765
rect 123253 459527 123287 459765
rect 123345 459595 123379 459765
rect 132913 459595 132947 459765
rect 133005 459595 133039 459765
rect 142573 459527 142607 459765
rect 142665 459595 142699 459765
rect 152233 459595 152267 459765
rect 152325 459595 152359 459765
rect 161893 459527 161927 459765
rect 161985 459595 162019 459765
rect 171553 459595 171587 459765
rect 171645 459595 171679 459765
rect 181213 459527 181247 459765
rect 181305 459595 181339 459765
rect 190873 459595 190907 459765
rect 190965 459595 190999 459765
rect 200533 459527 200567 459765
rect 200625 459595 200659 459765
rect 210193 459595 210227 459765
rect 210285 459595 210319 459765
rect 229513 459595 229547 459833
rect 234297 458235 234331 459629
rect 235067 459561 235125 459595
rect 242025 459459 242059 459629
rect 250121 458915 250155 459629
rect 251593 459459 251627 459561
rect 251685 459391 251719 459493
rect 256377 458439 256411 459629
rect 261253 459391 261287 459629
rect 261345 459459 261379 459697
rect 270913 459459 270947 459561
rect 280665 459527 280699 459697
rect 293027 459629 293211 459663
rect 290233 459527 290267 459629
rect 293177 459595 293211 459629
rect 312347 459629 312405 459663
rect 299985 459459 300019 459561
rect 309553 459459 309587 459629
rect 323537 458847 323571 459629
rect 327493 458711 327527 459629
rect 329517 458779 329551 459629
rect 331725 458371 331759 459629
rect 337797 458303 337831 459629
rect 345617 458507 345651 459629
rect 26745 337739 26779 337909
rect 36313 337603 36347 337909
rect 36405 337603 36439 337977
rect 113685 337603 113719 338113
rect 17085 337195 17119 337365
rect 55725 337195 55759 337569
rect 75045 336991 75079 337569
rect 94365 336855 94399 337569
rect 101081 336651 101115 336821
rect 103841 336651 103875 337569
rect 113777 337399 113811 337569
rect 113719 337365 113811 337399
rect 113869 336651 113903 337365
rect 116261 336447 116295 337501
rect 119205 337399 119239 338249
rect 119297 337399 119331 338113
rect 128957 337603 128991 338181
rect 129417 337943 129451 338113
rect 129509 337739 129543 337909
rect 123989 337399 124023 337569
rect 133189 337467 133223 337569
rect 138341 337399 138375 338181
rect 142665 337943 142699 338113
rect 152325 337943 152359 338113
rect 161985 337943 162019 338113
rect 171645 337943 171679 338113
rect 181305 337943 181339 338113
rect 190965 337943 190999 338113
rect 200625 337943 200659 338113
rect 210285 337943 210319 338113
rect 219945 337943 219979 338113
rect 142515 337909 142607 337943
rect 152175 337909 152267 337943
rect 161835 337909 161927 337943
rect 171495 337909 171587 337943
rect 181155 337909 181247 337943
rect 190815 337909 190907 337943
rect 200475 337909 200567 337943
rect 210135 337909 210227 337943
rect 219795 337909 219887 337943
rect 142573 337739 142607 337909
rect 142757 337739 142791 337909
rect 142699 337705 142791 337739
rect 152233 337739 152267 337909
rect 152417 337739 152451 337909
rect 152359 337705 152451 337739
rect 161893 337739 161927 337909
rect 162077 337739 162111 337909
rect 162019 337705 162111 337739
rect 171553 337739 171587 337909
rect 171737 337739 171771 337909
rect 171679 337705 171771 337739
rect 181213 337739 181247 337909
rect 181397 337739 181431 337909
rect 181339 337705 181431 337739
rect 190873 337739 190907 337909
rect 191057 337739 191091 337909
rect 190999 337705 191091 337739
rect 200533 337739 200567 337909
rect 200717 337739 200751 337909
rect 200659 337705 200751 337739
rect 210193 337739 210227 337909
rect 210377 337739 210411 337909
rect 210319 337705 210411 337739
rect 219853 337739 219887 337909
rect 220037 337739 220071 337909
rect 219979 337705 220071 337739
rect 138341 337365 138433 337399
rect 142389 336651 142423 337637
rect 142481 337569 142573 337603
rect 142481 337399 142515 337569
rect 142849 336651 142883 337637
rect 152049 336651 152083 337637
rect 152359 337569 152451 337603
rect 152417 337399 152451 337569
rect 152509 336651 152543 337637
rect 161709 336651 161743 337637
rect 161801 337569 161893 337603
rect 161801 337399 161835 337569
rect 162169 336651 162203 337637
rect 171369 336651 171403 337637
rect 171679 337569 171771 337603
rect 171737 337399 171771 337569
rect 171829 336651 171863 337637
rect 181029 336651 181063 337637
rect 181121 337569 181213 337603
rect 181121 337399 181155 337569
rect 181489 336651 181523 337637
rect 190689 336651 190723 337637
rect 190999 337569 191091 337603
rect 191057 337399 191091 337569
rect 191149 336651 191183 337637
rect 200349 336651 200383 337637
rect 200441 337569 200533 337603
rect 200441 337399 200475 337569
rect 200809 336651 200843 337637
rect 210009 336651 210043 337637
rect 210319 337569 210411 337603
rect 210377 337399 210411 337569
rect 210469 336651 210503 337637
rect 219669 336651 219703 337637
rect 219761 337569 219853 337603
rect 219761 337399 219795 337569
rect 220129 336651 220163 337637
rect 225465 337603 225499 338181
rect 225557 337603 225591 338113
rect 226753 337399 226787 338113
rect 230157 338011 230191 338249
rect 230249 337739 230283 337977
rect 234757 337739 234791 338249
rect 230341 337467 230375 337705
rect 230007 337433 230375 337467
rect 245337 336855 245371 337161
rect 152233 327131 152267 334645
rect 170173 327131 170207 327777
rect 214333 327131 214367 331993
rect 259045 331211 259079 331381
rect 259137 331143 259171 338045
rect 266773 337059 266807 337637
rect 270913 333251 270947 337909
rect 278549 337671 278583 338045
rect 280699 337977 280791 338011
rect 280757 337739 280791 337977
rect 314187 337501 314279 337535
rect 308449 337127 308483 337365
rect 314245 337127 314279 337501
rect 315073 336991 315107 337705
rect 317097 337059 317131 337637
rect 317189 337467 317223 337909
rect 318201 337195 318235 337501
rect 321973 337127 322007 337569
rect 229881 321419 229915 328389
rect 235493 318903 235527 328389
rect 235677 318903 235711 321929
rect 268613 321419 268647 328389
rect 276525 324411 276559 333897
rect 278733 326859 278767 331925
rect 279837 327131 279871 334305
rect 284989 331143 285023 336413
rect 285357 328491 285391 331449
rect 318661 321419 318695 328389
rect 261253 320263 261287 320637
rect 276985 318699 277019 318869
rect 135673 307819 135707 317373
rect 152233 307819 152267 317373
rect 170173 307819 170207 317373
rect 190873 307819 190907 309757
rect 214333 307819 214367 317373
rect 235493 311831 235527 318665
rect 268705 311627 268739 311933
rect 285265 309179 285299 318665
rect 285633 309179 285667 318665
rect 318937 314075 318971 318665
rect 309185 309179 309219 311797
rect 319121 309859 319155 318665
rect 319949 317475 319983 335257
rect 371929 331143 371963 337909
rect 328137 317475 328171 327029
rect 371929 321419 371963 328389
rect 373033 318699 373067 327029
rect 331173 309247 331207 311933
rect 225373 299523 225407 309077
rect 259321 299523 259355 309077
rect 357945 299523 357979 309077
rect 371837 302175 371871 309077
rect 385545 307819 385579 317373
rect 392445 307819 392479 317373
rect 235677 297415 235711 299421
rect 275513 296939 275547 299489
rect 272661 295239 272695 295545
rect 272753 295307 272787 295477
rect 91513 280279 91547 286297
rect 235493 282795 235527 285277
rect 259413 280279 259447 289765
rect 276617 285719 276651 295205
rect 276709 285719 276743 295273
rect 309185 289867 309219 299421
rect 319949 292451 319983 297993
rect 268705 282795 268739 284937
rect 271465 282795 271499 283033
rect 276709 280007 276743 285141
rect 276801 280075 276835 280449
rect 340925 280279 340959 289765
rect 341109 282795 341143 282965
rect 358037 280347 358071 289697
rect 371929 282795 371963 289697
rect 553905 280279 553939 289697
rect 242117 277355 242151 278817
rect 246625 277355 246659 278817
rect 259321 270555 259355 273309
rect 91513 260899 91547 270453
rect 225373 260899 225407 270453
rect 242761 267563 242795 269705
rect 285173 269127 285207 279837
rect 285265 270555 285299 279837
rect 309185 270555 309219 280041
rect 331265 270555 331299 280041
rect 372941 278783 372975 280245
rect 235585 253827 235619 260797
rect 242853 255323 242887 264809
rect 273029 255323 273063 256853
rect 91513 241655 91547 251141
rect 225373 241655 225407 251141
rect 229973 244171 230007 251141
rect 242577 245667 242611 255221
rect 246533 249815 246567 254133
rect 242761 241995 242795 246789
rect 235493 230503 235527 240057
rect 242485 227783 242519 237337
rect 273029 236011 273063 253861
rect 275605 245667 275639 255221
rect 285265 251243 285299 260729
rect 285633 251243 285667 260797
rect 305045 249815 305079 259369
rect 320041 258111 320075 263585
rect 357945 260899 357979 270453
rect 535965 269127 535999 271133
rect 553905 260967 553939 270453
rect 328321 253895 328355 256649
rect 331265 251243 331299 260797
rect 341109 251243 341143 260797
rect 285357 244171 285391 244341
rect 357945 241655 357979 251141
rect 553905 241655 553939 251141
rect 272845 231591 272879 235909
rect 268705 222207 268739 227001
rect 275697 224995 275731 234549
rect 276525 227783 276559 232577
rect 285357 231931 285391 236725
rect 309185 234379 309219 241417
rect 272937 217991 272971 224893
rect 242485 207043 242519 216597
rect 275605 215339 275639 224825
rect 272845 210443 272879 215237
rect 275605 210443 275639 211225
rect 276709 211191 276743 220745
rect 285265 219487 285299 224961
rect 320041 220983 320075 224961
rect 328321 211191 328355 235909
rect 341017 215271 341051 220745
rect 373217 212483 373251 220745
rect 229973 205547 230007 205785
rect 235493 203031 235527 205717
rect 268705 205547 268739 207689
rect 271465 205547 271499 205717
rect 235585 195755 235619 202793
rect 242485 189091 242519 198645
rect 275697 197387 275731 197557
rect 276985 189091 277019 198101
rect 279837 190519 279871 200073
rect 285081 198747 285115 208233
rect 309093 205547 309127 205717
rect 328413 204935 328447 209729
rect 341109 205547 341143 205785
rect 357945 203031 357979 212449
rect 320041 195959 320075 200073
rect 328413 195755 328447 200005
rect 341109 193375 341143 202793
rect 372021 191267 372055 200073
rect 373033 190587 373067 200073
rect 552433 196299 552467 201433
rect 229881 176579 229915 182121
rect 242853 182019 242887 188989
rect 309001 183583 309035 186337
rect 341109 183651 341143 186337
rect 552433 183515 552467 191777
rect 235493 166923 235527 167161
rect 135673 153255 135707 162809
rect 152233 153255 152267 162809
rect 170173 153255 170207 162809
rect 190873 153255 190907 162809
rect 214333 153255 214367 162809
rect 230065 157131 230099 162809
rect 235493 157131 235527 159273
rect 242485 157947 242519 162809
rect 242669 157131 242703 164169
rect 246625 153255 246659 162809
rect 246901 161483 246935 169269
rect 246809 157131 246843 159477
rect 259321 157335 259355 164169
rect 273029 163523 273063 168317
rect 275605 163523 275639 173213
rect 278825 171139 278859 180761
rect 285173 172567 285207 182121
rect 328321 176579 328355 182121
rect 268521 157131 268555 161245
rect 268705 147611 268739 154377
rect 273029 147679 273063 157301
rect 275605 147679 275639 157301
rect 135673 133943 135707 143429
rect 152233 133943 152267 143429
rect 170173 133943 170207 143429
rect 190873 133943 190907 143429
rect 214333 133943 214367 143429
rect 225373 135371 225407 144857
rect 273029 139451 273063 143701
rect 278733 142171 278767 149821
rect 259413 128299 259447 135201
rect 268705 128299 268739 135201
rect 271465 128503 271499 137921
rect 279745 129795 279779 139349
rect 285081 137887 285115 156757
rect 285265 138091 285299 157369
rect 305137 157335 305171 164169
rect 371929 161483 371963 179333
rect 385545 153255 385579 162809
rect 392445 153255 392479 162809
rect 529065 153255 529099 162809
rect 535965 153255 535999 162809
rect 552525 153255 552559 162809
rect 553905 154683 553939 164169
rect 571845 153255 571879 162809
rect 373125 145163 373159 153153
rect 285633 137955 285667 144857
rect 285449 135303 285483 135541
rect 309093 134691 309127 140709
rect 319949 133943 319983 143497
rect 328413 133943 328447 143497
rect 371929 128299 371963 135201
rect 385545 133943 385579 143497
rect 392445 133943 392479 143497
rect 529065 133943 529099 143497
rect 535965 133943 535999 143497
rect 552249 133943 552283 143497
rect 553905 135371 553939 144857
rect 571845 133943 571879 143497
rect 91513 106335 91547 115753
rect 135673 114563 135707 124117
rect 152233 114563 152267 124117
rect 170173 114563 170207 124117
rect 190873 114563 190907 124117
rect 214333 114563 214367 124117
rect 229789 114699 229823 118745
rect 242853 116739 242887 125545
rect 235585 108987 235619 115753
rect 135673 95319 135707 104805
rect 152233 95319 152267 104805
rect 170173 95319 170207 104805
rect 190873 95319 190907 104805
rect 214333 95319 214367 104805
rect 229823 103445 229915 103479
rect 229881 85595 229915 103445
rect 235493 96679 235527 106233
rect 242669 104907 242703 111129
rect 242853 110551 242887 114461
rect 272845 111843 272879 121397
rect 285633 111299 285667 120037
rect 305137 118507 305171 125545
rect 309001 119391 309035 125545
rect 341109 116059 341143 125545
rect 552249 125443 552283 133705
rect 235585 89675 235619 96577
rect 242025 93891 242059 101405
rect 275513 100759 275547 106301
rect 320133 104907 320167 109021
rect 328413 104907 328447 109021
rect 357945 106335 357979 115753
rect 373125 114563 373159 124117
rect 385545 114563 385579 124117
rect 392445 114563 392479 124117
rect 529065 114563 529099 124117
rect 535965 114563 535999 124117
rect 571845 114563 571879 124117
rect 285265 102187 285299 102357
rect 305045 99331 305079 104805
rect 246533 88451 246567 90049
rect 268705 89675 268739 96577
rect 308909 93891 308943 103445
rect 319949 93891 319983 103445
rect 373125 95319 373159 104805
rect 385545 95319 385579 104805
rect 392445 95319 392479 104805
rect 529065 95319 529099 104805
rect 535965 95319 535999 104805
rect 242485 86887 242519 87193
rect 91513 67643 91547 77129
rect 135673 75939 135707 85493
rect 152233 75939 152267 85493
rect 170173 75939 170207 85493
rect 190873 75939 190907 85493
rect 214333 75939 214367 85493
rect 242485 85323 242519 85493
rect 229973 79883 230007 80121
rect 271373 80087 271407 81481
rect 235493 67643 235527 77129
rect 246717 66283 246751 70465
rect 91513 48331 91547 57885
rect 135673 56695 135707 66181
rect 152233 56695 152267 66181
rect 170173 56695 170207 66181
rect 190873 56695 190907 66181
rect 214333 56695 214367 66181
rect 271465 63563 271499 76585
rect 276617 73219 276651 82773
rect 285265 77979 285299 82773
rect 305137 79883 305171 86921
rect 319949 75939 319983 85493
rect 341109 77435 341143 86921
rect 371929 85595 371963 95081
rect 552525 93891 552559 103445
rect 553905 96747 553939 109701
rect 571845 95319 571879 104805
rect 552433 86887 552467 87125
rect 279929 74443 279963 74613
rect 275605 63563 275639 73117
rect 341109 67643 341143 77129
rect 357945 67643 357979 77129
rect 373125 75939 373159 85493
rect 385545 75939 385579 85493
rect 392445 75939 392479 85493
rect 529065 75939 529099 85493
rect 535965 75939 535999 85493
rect 552341 77163 552375 85493
rect 571845 75939 571879 85493
rect 235401 48331 235435 57885
rect 91513 29019 91547 38505
rect 135673 37315 135707 46869
rect 152233 37315 152267 46869
rect 170173 37315 170207 46869
rect 190873 37315 190907 46869
rect 214333 37315 214367 46869
rect 225373 37315 225407 46869
rect 242485 45611 242519 63461
rect 277077 62747 277111 67609
rect 246901 45611 246935 55165
rect 272845 48331 272879 57885
rect 275605 52479 275639 57953
rect 259321 38743 259355 48229
rect 272845 37315 272879 46869
rect 275605 42823 275639 46937
rect 276525 44183 276559 57273
rect 278641 55267 278675 64821
rect 279745 55267 279779 64821
rect 285265 56491 285299 64821
rect 308909 56695 308943 66181
rect 320133 56695 320167 66181
rect 331265 62815 331299 67541
rect 357945 48331 357979 57885
rect 371929 55267 371963 64821
rect 385545 56695 385579 66181
rect 392445 56695 392479 66181
rect 529065 56695 529099 66181
rect 535965 56695 535999 66181
rect 552525 56695 552559 66181
rect 571845 56695 571879 66181
rect 278733 45611 278767 48297
rect 235493 29019 235527 31773
rect 91513 9707 91547 19261
rect 135305 18071 135339 27557
rect 151865 18071 151899 27557
rect 169713 18071 169747 27557
rect 225097 18071 225131 27557
rect 242577 22695 242611 27557
rect 254813 21403 254847 28917
rect 268429 26027 268463 26197
rect 272845 18071 272879 27557
rect 273029 26027 273063 26197
rect 275605 24871 275639 37961
rect 285725 29019 285759 42041
rect 319949 37315 319983 46869
rect 320317 31875 320351 38505
rect 328229 37315 328263 46869
rect 341017 29019 341051 31841
rect 357945 29019 357979 38505
rect 385545 37315 385579 46869
rect 392445 46699 392479 46869
rect 529065 37315 529099 46869
rect 535965 37315 535999 46869
rect 552525 37315 552559 46869
rect 553813 38403 553847 46869
rect 571845 37315 571879 46869
rect 278825 26299 278859 27625
rect 285173 19363 285207 28917
rect 285725 19363 285759 24157
rect 305137 18071 305171 27557
rect 123345 10523 123379 11033
rect 128957 10795 128991 11101
rect 129049 10999 129083 11169
rect 128865 10183 128899 10761
rect 133557 10251 133591 10693
rect 133649 10455 133683 10965
rect 133741 10523 133775 10625
rect 133833 10455 133867 11033
rect 133925 10387 133959 10489
rect 133649 10353 133959 10387
rect 133649 10183 133683 10353
rect 128865 10149 128957 10183
rect 133407 10149 133683 10183
rect 138157 9639 138191 10149
rect 138249 10115 138283 11101
rect 138375 10489 138467 10523
rect 138433 10183 138467 10489
rect 138525 10183 138559 11033
rect 147909 10727 147943 11101
rect 148093 10795 148127 11033
rect 148185 10727 148219 11033
rect 148277 10795 148311 11169
rect 143343 10693 143527 10727
rect 148369 10727 148403 11101
rect 152877 10761 153153 10795
rect 152877 10727 152911 10761
rect 143493 10659 143527 10693
rect 148001 10251 148035 10693
rect 143217 10115 143251 10217
rect 147817 10217 148035 10251
rect 157661 10251 157695 11033
rect 147817 10115 147851 10217
rect 157753 10183 157787 11169
rect 138249 10081 138341 10115
rect 143217 10081 143401 10115
rect 147909 9639 147943 10081
rect 138157 9605 138341 9639
rect 138525 9605 138709 9639
rect 148001 9639 148035 10149
rect 138525 9571 138559 9605
rect 148093 9571 148127 10149
rect 18465 8959 18499 9129
rect 28033 8959 28067 9129
rect 36405 9027 36439 9129
rect 31529 8891 31563 8993
rect 37785 8619 37819 8925
rect 42661 8891 42695 9129
rect 47353 8619 47387 8925
rect 54253 8891 54287 9129
rect 65385 9027 65419 9129
rect 75045 9027 75079 9129
rect 57105 8823 57139 8925
rect 66673 8823 66707 8925
rect 68145 8823 68179 8925
rect 81209 8891 81243 9129
rect 85717 8993 85993 9027
rect 85717 8823 85751 8993
rect 92893 8891 92927 9129
rect 104025 9027 104059 9129
rect 113685 9027 113719 9129
rect 116261 9027 116295 9129
rect 148093 9027 148127 9333
rect 85935 8857 85993 8891
rect 115065 8619 115099 8925
rect 124633 8619 124667 8925
rect 134385 8823 134419 8925
rect 138525 8823 138559 8925
rect 140089 8891 140123 8993
rect 148277 8891 148311 9605
rect 140089 8857 140273 8891
rect 157845 8891 157879 11033
rect 167597 10251 167631 11033
rect 176705 10795 176739 11305
rect 172381 10659 172415 10693
rect 172231 10625 172415 10659
rect 176797 10659 176831 11033
rect 176889 10727 176923 11101
rect 177073 10795 177107 11169
rect 179189 11135 179223 11305
rect 186917 10795 186951 11033
rect 187009 10727 187043 11101
rect 191517 10761 191793 10795
rect 191517 10727 191551 10761
rect 176981 10659 177015 10693
rect 176797 10625 177015 10659
rect 167539 10217 167631 10251
rect 196209 10183 196243 11033
rect 138467 8789 138559 8823
rect 162537 8551 162571 9605
rect 196577 9027 196611 11033
rect 225557 10115 225591 11101
rect 230065 10829 230375 10863
rect 230065 10795 230099 10829
rect 230157 10659 230191 10761
rect 230341 10727 230375 10829
rect 232399 10217 232457 10251
rect 234757 9095 234791 11237
rect 235493 10795 235527 11033
rect 235159 10693 235343 10727
rect 234941 10183 234975 10693
rect 235309 10251 235343 10693
rect 235401 10183 235435 10761
rect 238345 10659 238379 11169
rect 244877 9707 244911 10149
rect 244969 9571 245003 9673
rect 244785 9537 245003 9571
rect 244785 9503 244819 9537
rect 244877 9367 244911 9469
rect 244819 9333 244911 9367
rect 254353 9163 254387 9673
rect 254537 9639 254571 10081
rect 162629 8823 162663 8993
rect 162905 8619 162939 8857
rect 172289 8619 172323 8993
rect 181949 8619 181983 8993
rect 191609 8619 191643 8993
rect 201269 8619 201303 8993
rect 177165 5899 177199 8313
rect 186641 7803 186675 8381
rect 186733 5831 186767 7769
rect 195013 7735 195047 8313
rect 196393 7871 196427 8381
rect 210929 8347 210963 8993
rect 215897 8347 215931 8993
rect 254629 8823 254663 9877
rect 254721 8891 254755 9673
rect 254479 8789 254663 8823
rect 254813 8823 254847 9673
rect 259137 9503 259171 9877
rect 308265 9707 308299 19261
rect 331265 10251 331299 11169
rect 331449 10183 331483 11305
rect 331541 10795 331575 11237
rect 331541 10115 331575 10149
rect 331449 10081 331575 10115
rect 331449 10047 331483 10081
rect 331633 10047 331667 10761
rect 331725 10659 331759 11033
rect 331909 10727 331943 11101
rect 333749 10999 333783 11305
rect 340925 10727 340959 11305
rect 341017 11135 341051 11169
rect 341017 11101 341235 11135
rect 341109 10659 341143 11033
rect 341201 10659 341235 11101
rect 341293 10727 341327 11237
rect 331207 10013 331483 10047
rect 331575 10013 331667 10047
rect 350677 9469 350895 9503
rect 350677 9367 350711 9469
rect 225189 8381 225373 8415
rect 225189 8347 225223 8381
rect 341201 8279 341235 9061
rect 215897 6171 215931 6273
rect 215839 6137 215931 6171
rect 36405 3179 36439 3485
rect 44777 3383 44811 3621
rect 40177 3111 40211 3349
rect 45881 3111 45915 3417
rect 45973 3179 46007 3485
rect 56277 3179 56311 3485
rect 56369 3111 56403 3417
rect 65201 3111 65235 3485
rect 65293 3179 65327 3485
rect 75045 2975 75079 3485
rect 75137 2907 75171 3417
rect 84521 2907 84555 3417
rect 84613 2975 84647 3485
rect 93721 2907 93755 3485
rect 103933 2975 103967 3485
rect 103875 2941 103967 2975
rect 108625 2839 108659 2873
rect 108625 2805 108809 2839
rect 112799 2805 113409 2839
rect 113501 2635 113535 2873
rect 113685 2635 113719 2805
rect 123345 2635 123379 4165
rect 128957 3519 128991 4165
rect 133005 3995 133039 4165
rect 134293 3995 134327 4165
rect 138433 3519 138467 3961
rect 128255 3485 128899 3519
rect 138375 3485 138467 3519
rect 138801 3519 138835 4233
rect 147909 4233 148127 4267
rect 147909 4199 147943 4233
rect 138893 3519 138927 3621
rect 128865 3451 128899 3485
rect 128865 3417 129049 3451
rect 132821 2635 132855 3417
rect 132913 2805 133315 2839
rect 132913 2567 132947 2805
rect 133281 2567 133315 2805
rect 133373 2635 133407 3417
rect 142389 2635 142423 3417
rect 142573 2567 142607 3417
rect 142757 2635 142791 3621
rect 148001 3519 148035 4165
rect 148093 3519 148127 4233
rect 152233 3655 152267 4165
rect 148495 3621 149565 3655
rect 152141 2635 152175 3621
rect 157753 3519 157787 4233
rect 157845 3519 157879 4233
rect 167505 4233 167723 4267
rect 159133 3655 159167 4165
rect 167505 3655 167539 4233
rect 167689 4199 167723 4233
rect 177165 4233 177441 4267
rect 162755 3621 163365 3655
rect 166343 3621 167413 3655
rect 167597 3655 167631 4165
rect 152325 2567 152359 3417
rect 152509 2635 152543 3417
rect 161617 2635 161651 3485
rect 161893 2567 161927 3485
rect 162077 2635 162111 3621
rect 171461 2635 171495 4165
rect 171737 2635 171771 4165
rect 176889 3587 176923 4165
rect 176981 3655 177015 4165
rect 177073 3587 177107 3621
rect 176889 3553 177107 3587
rect 177165 3519 177199 4233
rect 177257 3519 177291 4165
rect 181121 2635 181155 3621
rect 181247 3553 181489 3587
rect 186733 3519 186767 4165
rect 181397 2635 181431 3485
rect 186951 3077 187043 3111
rect 187009 3043 187043 3077
rect 187101 2907 187135 3417
rect 186951 2873 187135 2907
rect 186825 2839 186859 2873
rect 186825 2805 187009 2839
rect 190781 2635 190815 4165
rect 190965 2567 190999 4233
rect 191057 2635 191091 4165
rect 196117 2635 196151 5661
rect 229329 5117 229547 5151
rect 229329 5083 229363 5117
rect 220497 4743 220531 4981
rect 220681 4811 220715 5049
rect 227581 5015 227615 5049
rect 227581 4981 227765 5015
rect 220773 4743 220807 4777
rect 220497 4709 220807 4743
rect 196243 3009 196577 3043
rect 196209 2635 196243 2873
rect 196301 2873 196485 2907
rect 196301 2839 196335 2873
rect 198509 2635 198543 2941
rect 200257 2635 200291 4165
rect 200533 2805 200659 2839
rect 200533 2567 200567 2805
rect 200625 2567 200659 2805
rect 200717 2635 200751 4165
rect 206145 3519 206179 4233
rect 215897 3655 215931 4233
rect 217461 3995 217495 4233
rect 218565 3995 218599 4233
rect 220497 4233 220681 4267
rect 220497 4199 220531 4233
rect 219703 3961 219795 3995
rect 205961 3077 206053 3111
rect 205961 3043 205995 3077
rect 205903 2941 206145 2975
rect 209917 2635 209951 3417
rect 210193 2567 210227 3417
rect 210377 2635 210411 3621
rect 219761 2635 219795 3961
rect 219853 3587 219887 3961
rect 219945 3655 219979 3961
rect 219853 3553 219979 3587
rect 219945 2567 219979 3553
rect 225407 3417 225465 3451
rect 229421 2635 229455 5049
rect 229513 5015 229547 5117
rect 229513 4981 229789 5015
rect 229697 2567 229731 4029
rect 232917 3995 232951 7837
rect 230341 3723 230375 3961
rect 234975 3893 235067 3927
rect 235033 3587 235067 3893
rect 235217 595 235251 6273
rect 245061 5287 245095 6273
rect 254169 5287 254203 6273
rect 254353 4063 254387 5185
rect 259045 4743 259079 6341
rect 272845 6171 272879 8245
rect 341293 8075 341327 9129
rect 322157 6987 322191 7157
rect 264197 5389 264415 5423
rect 264197 5355 264231 5389
rect 264381 5355 264415 5389
rect 264381 5321 264507 5355
rect 259263 5253 259447 5287
rect 263955 5253 264047 5287
rect 259413 5219 259447 5253
rect 264013 4743 264047 5253
rect 263921 4131 263955 4709
rect 264289 4131 264323 5321
rect 264473 4539 264507 5321
rect 302561 5287 302595 5593
rect 235309 3587 235343 3689
rect 249569 3519 249603 3689
rect 264565 3383 264599 4641
rect 267509 4471 267543 4573
rect 267417 4131 267451 4437
rect 268889 4199 268923 4573
rect 301089 4131 301123 4777
rect 301181 4063 301215 5117
rect 302653 5083 302687 5253
rect 302595 5049 302687 5083
rect 302745 5117 302837 5151
rect 307471 5117 307747 5151
rect 302745 4811 302779 5117
rect 302837 4607 302871 4777
rect 307621 4675 307655 4981
rect 307713 4675 307747 5117
rect 312129 5083 312163 5661
rect 312221 5355 312255 5729
rect 312313 5559 312347 6069
rect 312313 4675 312347 5321
rect 312497 5219 312531 5661
rect 312681 5287 312715 5729
rect 314613 5695 314647 6273
rect 317189 5763 317223 6341
rect 321789 6239 321823 6885
rect 323813 6443 323847 7225
rect 336509 6987 336543 7837
rect 339637 7531 339671 7905
rect 339637 7497 340925 7531
rect 341293 7395 341327 7497
rect 341235 7361 341327 7395
rect 321881 6375 321915 6409
rect 321881 6341 322065 6375
rect 328723 6273 328873 6307
rect 345341 5389 346479 5423
rect 312405 4947 312439 5185
rect 317097 5083 317131 5253
rect 317281 5151 317315 5321
rect 341385 5287 341419 5321
rect 341327 5253 341419 5287
rect 345341 5287 345375 5389
rect 346445 5355 346479 5389
rect 332461 5151 332495 5253
rect 317373 5083 317407 5117
rect 317097 5049 317407 5083
rect 346077 5151 346111 5253
rect 346077 5117 346261 5151
rect 312405 4913 312623 4947
rect 312255 4641 312347 4675
rect 302779 4573 302871 4607
rect 302653 4267 302687 4505
rect 302595 4233 302687 4267
rect 312405 4131 312439 4709
rect 283977 3927 284011 4029
rect 302469 4097 302653 4131
rect 283977 3893 284161 3927
rect 278733 3587 278767 3621
rect 268889 2839 268923 3553
rect 278549 3553 278767 3587
rect 278549 3519 278583 3553
rect 278641 3451 278675 3485
rect 275697 3043 275731 3417
rect 278457 3417 278675 3451
rect 278457 3043 278491 3417
rect 298513 3383 298547 3893
rect 299709 3723 299743 4029
rect 302469 3995 302503 4097
rect 312497 4063 312531 4709
rect 312589 4063 312623 4913
rect 332369 4607 332403 5117
rect 345433 4675 345467 5049
rect 346353 4811 346387 5321
rect 322893 3927 322927 4097
rect 324181 3927 324215 4165
rect 325929 3961 326331 3995
rect 325929 3927 325963 3961
rect 300997 3451 301031 3553
rect 326021 3519 326055 3893
rect 326297 3519 326331 3961
rect 331541 3723 331575 4233
rect 331633 3723 331667 4165
rect 341385 3519 341419 4505
rect 278549 3043 278583 3349
rect 298605 2839 298639 3349
rect 301089 3179 301123 3417
rect 309093 595 309127 2805
rect 326205 2635 326239 3485
rect 345617 2567 345651 4505
rect 346169 4267 346203 4437
rect 346261 4267 346295 4777
rect 346537 4539 346571 9333
rect 350769 9163 350803 9401
rect 350861 9299 350895 9469
rect 350953 9367 350987 11237
rect 351079 9401 351171 9435
rect 350861 9265 350987 9299
rect 350769 9129 350861 9163
rect 350677 7871 350711 9129
rect 350953 9095 350987 9265
rect 351137 9163 351171 9401
rect 350769 7939 350803 9061
rect 351045 8959 351079 9129
rect 351321 9027 351355 11169
rect 355921 9095 355955 9333
rect 356013 9027 356047 9333
rect 355771 8993 356047 9027
rect 351045 8925 351137 8959
rect 355553 8449 355737 8483
rect 355553 8415 355587 8449
rect 373125 8415 373159 17833
rect 409097 10523 409131 11101
rect 418481 10523 418515 11101
rect 418573 10523 418607 11033
rect 418757 10591 418791 11101
rect 418665 10523 418699 10557
rect 423357 10523 423391 10557
rect 418665 10489 418791 10523
rect 423357 10489 423541 10523
rect 418665 9639 418699 10421
rect 418757 9571 418791 10489
rect 529065 9707 529099 27557
rect 535965 9707 535999 27557
rect 541485 9707 541519 19261
rect 552525 9707 552559 27557
rect 560805 9707 560839 19261
rect 571845 9707 571879 27557
rect 428325 9503 428359 9673
rect 350861 7973 350953 8007
rect 350861 7871 350895 7973
rect 350677 7837 350895 7871
rect 357979 7429 358129 7463
rect 346939 7361 346997 7395
rect 424185 6851 424219 7361
rect 433753 6851 433787 7361
rect 457305 6783 457339 7701
rect 457397 6851 457431 7769
rect 457489 7735 457523 8381
rect 457581 7803 457615 8313
rect 473899 7497 474049 7531
rect 462825 6715 462859 7361
rect 473991 7361 474141 7395
rect 472393 6715 472427 7361
rect 473991 7225 474141 7259
rect 357979 6341 358129 6375
rect 346939 6273 346997 6307
rect 424185 6103 424219 6273
rect 370767 5593 370951 5627
rect 350769 2567 350803 3485
rect 355093 3009 355403 3043
rect 355093 2975 355127 3009
rect 355369 2975 355403 3009
rect 355277 2635 355311 2941
rect 360705 2839 360739 3485
rect 370365 2839 370399 3485
rect 370457 3111 370491 3553
rect 370825 3179 370859 5525
rect 370917 3247 370951 5593
rect 505881 5083 505915 5525
rect 370917 3213 374815 3247
rect 370825 3145 374723 3179
rect 370457 3077 374631 3111
rect 360705 2805 364695 2839
rect 364661 2635 364695 2805
rect 364753 2567 364787 2805
rect 370365 2805 374355 2839
rect 364937 2635 364971 2805
rect 374321 2635 374355 2805
rect 374597 2635 374631 3077
rect 374689 2499 374723 3145
rect 374781 2431 374815 3213
rect 383981 2635 384015 3553
rect 384073 2567 384107 3553
rect 390053 2635 390087 3417
rect 418757 3043 418791 4097
rect 505605 4063 505639 4981
rect 505697 4131 505731 4981
rect 505789 3995 505823 5049
rect 515173 5015 515207 5593
rect 515081 4131 515115 4981
rect 529525 4267 529559 4777
rect 534585 4675 534619 4777
rect 559459 4709 559517 4743
rect 529617 4267 529651 4573
rect 538725 4471 538759 4641
rect 549857 4607 549891 4641
rect 549799 4573 549891 4607
rect 548293 4471 548327 4573
rect 515265 4131 515299 4165
rect 515265 4097 515449 4131
rect 420873 595 420907 2805
<< viali >>
rect 290049 701097 290083 701131
rect 288761 701029 288795 701063
rect 288761 700825 288795 700859
rect 278549 699941 278583 699975
rect 229605 699873 229639 699907
rect 229605 699737 229639 699771
rect 239265 699873 239299 699907
rect 239265 699669 239299 699703
rect 259229 699873 259263 699907
rect 259229 699669 259263 699703
rect 264105 699873 264139 699907
rect 264105 699669 264139 699703
rect 287381 699941 287415 699975
rect 278549 699669 278583 699703
rect 278641 699873 278675 699907
rect 296305 701097 296339 701131
rect 292349 700961 292383 700995
rect 292533 700961 292567 700995
rect 296213 700893 296247 700927
rect 296305 700893 296339 700927
rect 292257 700825 292291 700859
rect 290049 699873 290083 699907
rect 292257 700213 292291 700247
rect 292349 700213 292383 700247
rect 292349 700009 292383 700043
rect 292441 700009 292475 700043
rect 296121 700009 296155 700043
rect 294557 699941 294591 699975
rect 294741 699941 294775 699975
rect 296213 699873 296247 699907
rect 292625 699805 292659 699839
rect 296121 699805 296155 699839
rect 287473 699737 287507 699771
rect 289037 699737 289071 699771
rect 291889 699737 291923 699771
rect 278641 699669 278675 699703
rect 288853 699669 288887 699703
rect 291613 699669 291647 699703
rect 378737 695453 378771 695487
rect 378737 685865 378771 685899
rect 508457 695453 508491 695487
rect 508457 685865 508491 685899
rect 314153 676073 314187 676107
rect 314153 666553 314187 666587
rect 378645 676073 378679 676107
rect 378645 666553 378679 666587
rect 443873 676073 443907 676107
rect 443873 666553 443907 666587
rect 508365 676073 508399 676107
rect 508365 666553 508399 666587
rect 573593 676073 573627 676107
rect 573593 666553 573627 666587
rect 314153 637449 314187 637483
rect 314153 627929 314187 627963
rect 443873 637449 443907 637483
rect 443873 627929 443907 627963
rect 573593 637449 573627 637483
rect 573593 627929 573627 627963
rect 443689 608549 443723 608583
rect 443689 601545 443723 601579
rect 573409 608549 573443 608583
rect 573409 601545 573443 601579
rect 313877 598825 313911 598859
rect 313877 589305 313911 589339
rect 443873 598825 443907 598859
rect 443873 589305 443907 589339
rect 573593 598825 573627 598859
rect 573593 589305 573627 589339
rect 378645 589237 378679 589271
rect 378645 579649 378679 579683
rect 508365 589237 508399 589271
rect 508365 579649 508399 579683
rect 313969 579581 314003 579615
rect 313969 569993 314003 570027
rect 378737 569857 378771 569891
rect 378737 562921 378771 562955
rect 508457 569857 508491 569891
rect 508457 562921 508491 562955
rect 443505 553401 443539 553435
rect 443505 550613 443539 550647
rect 573225 553401 573259 553435
rect 573225 550613 573259 550647
rect 443505 534089 443539 534123
rect 443505 531301 443539 531335
rect 573225 534089 573259 534123
rect 573225 531301 573259 531335
rect 443597 531233 443631 531267
rect 443597 524297 443631 524331
rect 573317 531233 573351 531267
rect 573317 524297 573351 524331
rect 443505 485877 443539 485911
rect 443505 485673 443539 485707
rect 573225 485877 573259 485911
rect 573225 485673 573259 485707
rect 443597 471937 443631 471971
rect 302929 463709 302963 463743
rect 268889 463641 268923 463675
rect 268889 463097 268923 463131
rect 283701 463233 283735 463267
rect 284897 463233 284931 463267
rect 284713 463165 284747 463199
rect 302285 463165 302319 463199
rect 283701 463029 283735 463063
rect 291613 463097 291647 463131
rect 292625 463097 292659 463131
rect 292625 462281 292659 462315
rect 301273 463097 301307 463131
rect 291613 462145 291647 462179
rect 302285 462213 302319 462247
rect 301273 462145 301307 462179
rect 443597 463165 443631 463199
rect 573317 471937 573351 471971
rect 573317 463029 573351 463063
rect 302929 462145 302963 462179
rect 225373 460037 225407 460071
rect 225373 459833 225407 459867
rect 229513 459833 229547 459867
rect 7333 459765 7367 459799
rect 7425 459765 7459 459799
rect 7425 459561 7459 459595
rect 16993 459765 17027 459799
rect 16993 459561 17027 459595
rect 17085 459765 17119 459799
rect 17085 459561 17119 459595
rect 26653 459765 26687 459799
rect 7333 459493 7367 459527
rect 26745 459765 26779 459799
rect 26745 459561 26779 459595
rect 36313 459765 36347 459799
rect 36313 459561 36347 459595
rect 36405 459765 36439 459799
rect 36405 459561 36439 459595
rect 45973 459765 46007 459799
rect 26653 459493 26687 459527
rect 46065 459765 46099 459799
rect 46065 459561 46099 459595
rect 55633 459765 55667 459799
rect 55633 459561 55667 459595
rect 55725 459765 55759 459799
rect 55725 459561 55759 459595
rect 65293 459765 65327 459799
rect 45973 459493 46007 459527
rect 65385 459765 65419 459799
rect 65385 459561 65419 459595
rect 74953 459765 74987 459799
rect 74953 459561 74987 459595
rect 75045 459765 75079 459799
rect 75045 459561 75079 459595
rect 84613 459765 84647 459799
rect 65293 459493 65327 459527
rect 84705 459765 84739 459799
rect 84705 459561 84739 459595
rect 94273 459765 94307 459799
rect 94273 459561 94307 459595
rect 94365 459765 94399 459799
rect 94365 459561 94399 459595
rect 103933 459765 103967 459799
rect 84613 459493 84647 459527
rect 104025 459765 104059 459799
rect 104025 459561 104059 459595
rect 113593 459765 113627 459799
rect 113593 459561 113627 459595
rect 113685 459765 113719 459799
rect 113685 459561 113719 459595
rect 123253 459765 123287 459799
rect 103933 459493 103967 459527
rect 123345 459765 123379 459799
rect 123345 459561 123379 459595
rect 132913 459765 132947 459799
rect 132913 459561 132947 459595
rect 133005 459765 133039 459799
rect 133005 459561 133039 459595
rect 142573 459765 142607 459799
rect 123253 459493 123287 459527
rect 142665 459765 142699 459799
rect 142665 459561 142699 459595
rect 152233 459765 152267 459799
rect 152233 459561 152267 459595
rect 152325 459765 152359 459799
rect 152325 459561 152359 459595
rect 161893 459765 161927 459799
rect 142573 459493 142607 459527
rect 161985 459765 162019 459799
rect 161985 459561 162019 459595
rect 171553 459765 171587 459799
rect 171553 459561 171587 459595
rect 171645 459765 171679 459799
rect 171645 459561 171679 459595
rect 181213 459765 181247 459799
rect 161893 459493 161927 459527
rect 181305 459765 181339 459799
rect 181305 459561 181339 459595
rect 190873 459765 190907 459799
rect 190873 459561 190907 459595
rect 190965 459765 190999 459799
rect 190965 459561 190999 459595
rect 200533 459765 200567 459799
rect 181213 459493 181247 459527
rect 200625 459765 200659 459799
rect 200625 459561 200659 459595
rect 210193 459765 210227 459799
rect 210193 459561 210227 459595
rect 210285 459765 210319 459799
rect 210285 459561 210319 459595
rect 261345 459697 261379 459731
rect 229513 459561 229547 459595
rect 234297 459629 234331 459663
rect 200533 459493 200567 459527
rect 242025 459629 242059 459663
rect 235033 459561 235067 459595
rect 235125 459561 235159 459595
rect 242025 459425 242059 459459
rect 250121 459629 250155 459663
rect 256377 459629 256411 459663
rect 251593 459561 251627 459595
rect 251593 459425 251627 459459
rect 251685 459493 251719 459527
rect 251685 459357 251719 459391
rect 250121 458881 250155 458915
rect 261253 459629 261287 459663
rect 280665 459697 280699 459731
rect 261345 459425 261379 459459
rect 270913 459561 270947 459595
rect 280665 459493 280699 459527
rect 290233 459629 290267 459663
rect 292993 459629 293027 459663
rect 309553 459629 309587 459663
rect 312313 459629 312347 459663
rect 312405 459629 312439 459663
rect 323537 459629 323571 459663
rect 293177 459561 293211 459595
rect 299985 459561 300019 459595
rect 290233 459493 290267 459527
rect 270913 459425 270947 459459
rect 299985 459425 300019 459459
rect 309553 459425 309587 459459
rect 261253 459357 261287 459391
rect 323537 458813 323571 458847
rect 327493 459629 327527 459663
rect 329517 459629 329551 459663
rect 329517 458745 329551 458779
rect 331725 459629 331759 459663
rect 327493 458677 327527 458711
rect 256377 458405 256411 458439
rect 331725 458337 331759 458371
rect 337797 459629 337831 459663
rect 345617 459629 345651 459663
rect 345617 458473 345651 458507
rect 337797 458269 337831 458303
rect 234297 458201 234331 458235
rect 119205 338249 119239 338283
rect 113685 338113 113719 338147
rect 36405 337977 36439 338011
rect 26745 337909 26779 337943
rect 26745 337705 26779 337739
rect 36313 337909 36347 337943
rect 36313 337569 36347 337603
rect 36405 337569 36439 337603
rect 55725 337569 55759 337603
rect 17085 337365 17119 337399
rect 17085 337161 17119 337195
rect 55725 337161 55759 337195
rect 75045 337569 75079 337603
rect 75045 336957 75079 336991
rect 94365 337569 94399 337603
rect 103841 337569 103875 337603
rect 113685 337569 113719 337603
rect 113777 337569 113811 337603
rect 94365 336821 94399 336855
rect 101081 336821 101115 336855
rect 101081 336617 101115 336651
rect 116261 337501 116295 337535
rect 113685 337365 113719 337399
rect 113869 337365 113903 337399
rect 103841 336617 103875 336651
rect 113869 336617 113903 336651
rect 230157 338249 230191 338283
rect 128957 338181 128991 338215
rect 119205 337365 119239 337399
rect 119297 338113 119331 338147
rect 138341 338181 138375 338215
rect 129417 338113 129451 338147
rect 129417 337909 129451 337943
rect 129509 337909 129543 337943
rect 129509 337705 129543 337739
rect 119297 337365 119331 337399
rect 123989 337569 124023 337603
rect 128957 337569 128991 337603
rect 133189 337569 133223 337603
rect 133189 337433 133223 337467
rect 123989 337365 124023 337399
rect 225465 338181 225499 338215
rect 142665 338113 142699 338147
rect 152325 338113 152359 338147
rect 161985 338113 162019 338147
rect 171645 338113 171679 338147
rect 181305 338113 181339 338147
rect 190965 338113 190999 338147
rect 200625 338113 200659 338147
rect 210285 338113 210319 338147
rect 219945 338113 219979 338147
rect 142481 337909 142515 337943
rect 142665 337909 142699 337943
rect 142757 337909 142791 337943
rect 152141 337909 152175 337943
rect 152325 337909 152359 337943
rect 152417 337909 152451 337943
rect 161801 337909 161835 337943
rect 161985 337909 162019 337943
rect 162077 337909 162111 337943
rect 171461 337909 171495 337943
rect 171645 337909 171679 337943
rect 171737 337909 171771 337943
rect 181121 337909 181155 337943
rect 181305 337909 181339 337943
rect 181397 337909 181431 337943
rect 190781 337909 190815 337943
rect 190965 337909 190999 337943
rect 191057 337909 191091 337943
rect 200441 337909 200475 337943
rect 200625 337909 200659 337943
rect 200717 337909 200751 337943
rect 210101 337909 210135 337943
rect 210285 337909 210319 337943
rect 210377 337909 210411 337943
rect 219761 337909 219795 337943
rect 219945 337909 219979 337943
rect 220037 337909 220071 337943
rect 142573 337705 142607 337739
rect 142665 337705 142699 337739
rect 152233 337705 152267 337739
rect 152325 337705 152359 337739
rect 161893 337705 161927 337739
rect 161985 337705 162019 337739
rect 171553 337705 171587 337739
rect 171645 337705 171679 337739
rect 181213 337705 181247 337739
rect 181305 337705 181339 337739
rect 190873 337705 190907 337739
rect 190965 337705 190999 337739
rect 200533 337705 200567 337739
rect 200625 337705 200659 337739
rect 210193 337705 210227 337739
rect 210285 337705 210319 337739
rect 219853 337705 219887 337739
rect 219945 337705 219979 337739
rect 142389 337637 142423 337671
rect 138433 337365 138467 337399
rect 142849 337637 142883 337671
rect 142573 337569 142607 337603
rect 142481 337365 142515 337399
rect 142389 336617 142423 336651
rect 142849 336617 142883 336651
rect 152049 337637 152083 337671
rect 152509 337637 152543 337671
rect 152325 337569 152359 337603
rect 152417 337365 152451 337399
rect 152049 336617 152083 336651
rect 152509 336617 152543 336651
rect 161709 337637 161743 337671
rect 162169 337637 162203 337671
rect 161893 337569 161927 337603
rect 161801 337365 161835 337399
rect 161709 336617 161743 336651
rect 162169 336617 162203 336651
rect 171369 337637 171403 337671
rect 171829 337637 171863 337671
rect 171645 337569 171679 337603
rect 171737 337365 171771 337399
rect 171369 336617 171403 336651
rect 171829 336617 171863 336651
rect 181029 337637 181063 337671
rect 181489 337637 181523 337671
rect 181213 337569 181247 337603
rect 181121 337365 181155 337399
rect 181029 336617 181063 336651
rect 181489 336617 181523 336651
rect 190689 337637 190723 337671
rect 191149 337637 191183 337671
rect 190965 337569 190999 337603
rect 191057 337365 191091 337399
rect 190689 336617 190723 336651
rect 191149 336617 191183 336651
rect 200349 337637 200383 337671
rect 200809 337637 200843 337671
rect 200533 337569 200567 337603
rect 200441 337365 200475 337399
rect 200349 336617 200383 336651
rect 200809 336617 200843 336651
rect 210009 337637 210043 337671
rect 210469 337637 210503 337671
rect 210285 337569 210319 337603
rect 210377 337365 210411 337399
rect 210009 336617 210043 336651
rect 210469 336617 210503 336651
rect 219669 337637 219703 337671
rect 220129 337637 220163 337671
rect 219853 337569 219887 337603
rect 219761 337365 219795 337399
rect 219669 336617 219703 336651
rect 225465 337569 225499 337603
rect 225557 338113 225591 338147
rect 225557 337569 225591 337603
rect 226753 338113 226787 338147
rect 234757 338249 234791 338283
rect 230157 337977 230191 338011
rect 230249 337977 230283 338011
rect 230249 337705 230283 337739
rect 230341 337705 230375 337739
rect 234757 337705 234791 337739
rect 259137 338045 259171 338079
rect 229973 337433 230007 337467
rect 226753 337365 226787 337399
rect 245337 337161 245371 337195
rect 245337 336821 245371 336855
rect 220129 336617 220163 336651
rect 116261 336413 116295 336447
rect 152233 334645 152267 334679
rect 214333 331993 214367 332027
rect 152233 327097 152267 327131
rect 170173 327777 170207 327811
rect 170173 327097 170207 327131
rect 259045 331381 259079 331415
rect 259045 331177 259079 331211
rect 278549 338045 278583 338079
rect 270913 337909 270947 337943
rect 266773 337637 266807 337671
rect 266773 337025 266807 337059
rect 280665 337977 280699 338011
rect 317189 337909 317223 337943
rect 280757 337705 280791 337739
rect 315073 337705 315107 337739
rect 278549 337637 278583 337671
rect 314153 337501 314187 337535
rect 308449 337365 308483 337399
rect 308449 337093 308483 337127
rect 314245 337093 314279 337127
rect 317097 337637 317131 337671
rect 371929 337909 371963 337943
rect 321973 337569 322007 337603
rect 317189 337433 317223 337467
rect 318201 337501 318235 337535
rect 318201 337161 318235 337195
rect 321973 337093 322007 337127
rect 317097 337025 317131 337059
rect 315073 336957 315107 336991
rect 284989 336413 285023 336447
rect 279837 334305 279871 334339
rect 270913 333217 270947 333251
rect 276525 333897 276559 333931
rect 259137 331109 259171 331143
rect 214333 327097 214367 327131
rect 229881 328389 229915 328423
rect 229881 321385 229915 321419
rect 235493 328389 235527 328423
rect 268613 328389 268647 328423
rect 235493 318869 235527 318903
rect 235677 321929 235711 321963
rect 278733 331925 278767 331959
rect 319949 335257 319983 335291
rect 284989 331109 285023 331143
rect 285357 331449 285391 331483
rect 285357 328457 285391 328491
rect 279837 327097 279871 327131
rect 318661 328389 318695 328423
rect 278733 326825 278767 326859
rect 276525 324377 276559 324411
rect 268613 321385 268647 321419
rect 318661 321385 318695 321419
rect 261253 320637 261287 320671
rect 261253 320229 261287 320263
rect 235677 318869 235711 318903
rect 276985 318869 277019 318903
rect 235493 318665 235527 318699
rect 276985 318665 277019 318699
rect 285265 318665 285299 318699
rect 135673 317373 135707 317407
rect 135673 307785 135707 307819
rect 152233 317373 152267 317407
rect 152233 307785 152267 307819
rect 170173 317373 170207 317407
rect 214333 317373 214367 317407
rect 170173 307785 170207 307819
rect 190873 309757 190907 309791
rect 190873 307785 190907 307819
rect 235493 311797 235527 311831
rect 268705 311933 268739 311967
rect 268705 311593 268739 311627
rect 285265 309145 285299 309179
rect 285633 318665 285667 318699
rect 318937 318665 318971 318699
rect 318937 314041 318971 314075
rect 319121 318665 319155 318699
rect 285633 309145 285667 309179
rect 309185 311797 309219 311831
rect 371929 331109 371963 331143
rect 371929 328389 371963 328423
rect 319949 317441 319983 317475
rect 328137 327029 328171 327063
rect 371929 321385 371963 321419
rect 373033 327029 373067 327063
rect 373033 318665 373067 318699
rect 328137 317441 328171 317475
rect 385545 317373 385579 317407
rect 319121 309825 319155 309859
rect 331173 311933 331207 311967
rect 331173 309213 331207 309247
rect 309185 309145 309219 309179
rect 214333 307785 214367 307819
rect 225373 309077 225407 309111
rect 225373 299489 225407 299523
rect 259321 309077 259355 309111
rect 357945 309077 357979 309111
rect 371837 309077 371871 309111
rect 385545 307785 385579 307819
rect 392445 317373 392479 317407
rect 392445 307785 392479 307819
rect 371837 302141 371871 302175
rect 259321 299489 259355 299523
rect 275513 299489 275547 299523
rect 357945 299489 357979 299523
rect 235677 299421 235711 299455
rect 235677 297381 235711 297415
rect 275513 296905 275547 296939
rect 309185 299421 309219 299455
rect 272661 295545 272695 295579
rect 272753 295477 272787 295511
rect 272753 295273 272787 295307
rect 276709 295273 276743 295307
rect 272661 295205 272695 295239
rect 276617 295205 276651 295239
rect 259413 289765 259447 289799
rect 91513 286297 91547 286331
rect 235493 285277 235527 285311
rect 235493 282761 235527 282795
rect 91513 280245 91547 280279
rect 276617 285685 276651 285719
rect 319949 297993 319983 298027
rect 319949 292417 319983 292451
rect 309185 289833 309219 289867
rect 276709 285685 276743 285719
rect 340925 289765 340959 289799
rect 276709 285141 276743 285175
rect 268705 284937 268739 284971
rect 268705 282761 268739 282795
rect 271465 283033 271499 283067
rect 271465 282761 271499 282795
rect 259413 280245 259447 280279
rect 276801 280449 276835 280483
rect 358037 289697 358071 289731
rect 341109 282965 341143 282999
rect 341109 282761 341143 282795
rect 371929 289697 371963 289731
rect 371929 282761 371963 282795
rect 553905 289697 553939 289731
rect 358037 280313 358071 280347
rect 340925 280245 340959 280279
rect 372941 280245 372975 280279
rect 553905 280245 553939 280279
rect 276801 280041 276835 280075
rect 309185 280041 309219 280075
rect 276709 279973 276743 280007
rect 285173 279837 285207 279871
rect 242117 278817 242151 278851
rect 242117 277321 242151 277355
rect 246625 278817 246659 278851
rect 246625 277321 246659 277355
rect 259321 273309 259355 273343
rect 259321 270521 259355 270555
rect 91513 270453 91547 270487
rect 91513 260865 91547 260899
rect 225373 270453 225407 270487
rect 242761 269705 242795 269739
rect 285265 279837 285299 279871
rect 285265 270521 285299 270555
rect 309185 270521 309219 270555
rect 331265 280041 331299 280075
rect 372941 278749 372975 278783
rect 331265 270521 331299 270555
rect 535965 271133 535999 271167
rect 285173 269093 285207 269127
rect 357945 270453 357979 270487
rect 242761 267529 242795 267563
rect 225373 260865 225407 260899
rect 242853 264809 242887 264843
rect 235585 260797 235619 260831
rect 320041 263585 320075 263619
rect 285633 260797 285667 260831
rect 285265 260729 285299 260763
rect 242853 255289 242887 255323
rect 273029 256853 273063 256887
rect 273029 255289 273063 255323
rect 235585 253793 235619 253827
rect 242577 255221 242611 255255
rect 91513 251141 91547 251175
rect 91513 241621 91547 241655
rect 225373 251141 225407 251175
rect 229973 251141 230007 251175
rect 275605 255221 275639 255255
rect 246533 254133 246567 254167
rect 246533 249781 246567 249815
rect 273029 253861 273063 253895
rect 242577 245633 242611 245667
rect 242761 246789 242795 246823
rect 229973 244137 230007 244171
rect 242761 241961 242795 241995
rect 225373 241621 225407 241655
rect 235493 240057 235527 240091
rect 235493 230469 235527 230503
rect 242485 237337 242519 237371
rect 285265 251209 285299 251243
rect 285633 251209 285667 251243
rect 305045 259369 305079 259403
rect 535965 269093 535999 269127
rect 553905 270453 553939 270487
rect 553905 260933 553939 260967
rect 357945 260865 357979 260899
rect 320041 258077 320075 258111
rect 331265 260797 331299 260831
rect 328321 256649 328355 256683
rect 328321 253861 328355 253895
rect 331265 251209 331299 251243
rect 341109 260797 341143 260831
rect 341109 251209 341143 251243
rect 305045 249781 305079 249815
rect 357945 251141 357979 251175
rect 275605 245633 275639 245667
rect 285357 244341 285391 244375
rect 285357 244137 285391 244171
rect 357945 241621 357979 241655
rect 553905 251141 553939 251175
rect 553905 241621 553939 241655
rect 309185 241417 309219 241451
rect 273029 235977 273063 236011
rect 285357 236725 285391 236759
rect 272845 235909 272879 235943
rect 272845 231557 272879 231591
rect 275697 234549 275731 234583
rect 242485 227749 242519 227783
rect 268705 227001 268739 227035
rect 276525 232577 276559 232611
rect 309185 234345 309219 234379
rect 328321 235909 328355 235943
rect 285357 231897 285391 231931
rect 276525 227749 276559 227783
rect 275697 224961 275731 224995
rect 285265 224961 285299 224995
rect 268705 222173 268739 222207
rect 272937 224893 272971 224927
rect 272937 217957 272971 217991
rect 275605 224825 275639 224859
rect 242485 216597 242519 216631
rect 275605 215305 275639 215339
rect 276709 220745 276743 220779
rect 272845 215237 272879 215271
rect 272845 210409 272879 210443
rect 275605 211225 275639 211259
rect 320041 224961 320075 224995
rect 320041 220949 320075 220983
rect 285265 219453 285299 219487
rect 276709 211157 276743 211191
rect 341017 220745 341051 220779
rect 341017 215237 341051 215271
rect 373217 220745 373251 220779
rect 328321 211157 328355 211191
rect 357945 212449 357979 212483
rect 373217 212449 373251 212483
rect 275605 210409 275639 210443
rect 328413 209729 328447 209763
rect 285081 208233 285115 208267
rect 242485 207009 242519 207043
rect 268705 207689 268739 207723
rect 229973 205785 230007 205819
rect 229973 205513 230007 205547
rect 235493 205717 235527 205751
rect 268705 205513 268739 205547
rect 271465 205717 271499 205751
rect 271465 205513 271499 205547
rect 235493 202997 235527 203031
rect 235585 202793 235619 202827
rect 279837 200073 279871 200107
rect 235585 195721 235619 195755
rect 242485 198645 242519 198679
rect 276985 198101 277019 198135
rect 275697 197557 275731 197591
rect 275697 197353 275731 197387
rect 242485 189057 242519 189091
rect 309093 205717 309127 205751
rect 309093 205513 309127 205547
rect 341109 205785 341143 205819
rect 341109 205513 341143 205547
rect 328413 204901 328447 204935
rect 357945 202997 357979 203031
rect 341109 202793 341143 202827
rect 285081 198713 285115 198747
rect 320041 200073 320075 200107
rect 320041 195925 320075 195959
rect 328413 200005 328447 200039
rect 328413 195721 328447 195755
rect 552433 201433 552467 201467
rect 341109 193341 341143 193375
rect 372021 200073 372055 200107
rect 372021 191233 372055 191267
rect 373033 200073 373067 200107
rect 552433 196265 552467 196299
rect 373033 190553 373067 190587
rect 552433 191777 552467 191811
rect 279837 190485 279871 190519
rect 276985 189057 277019 189091
rect 242853 188989 242887 189023
rect 229881 182121 229915 182155
rect 309001 186337 309035 186371
rect 341109 186337 341143 186371
rect 341109 183617 341143 183651
rect 309001 183549 309035 183583
rect 552433 183481 552467 183515
rect 242853 181985 242887 182019
rect 285173 182121 285207 182155
rect 229881 176545 229915 176579
rect 278825 180761 278859 180795
rect 275605 173213 275639 173247
rect 246901 169269 246935 169303
rect 235493 167161 235527 167195
rect 235493 166889 235527 166923
rect 242669 164169 242703 164203
rect 135673 162809 135707 162843
rect 135673 153221 135707 153255
rect 152233 162809 152267 162843
rect 152233 153221 152267 153255
rect 170173 162809 170207 162843
rect 170173 153221 170207 153255
rect 190873 162809 190907 162843
rect 190873 153221 190907 153255
rect 214333 162809 214367 162843
rect 230065 162809 230099 162843
rect 242485 162809 242519 162843
rect 230065 157097 230099 157131
rect 235493 159273 235527 159307
rect 242485 157913 242519 157947
rect 235493 157097 235527 157131
rect 242669 157097 242703 157131
rect 246625 162809 246659 162843
rect 214333 153221 214367 153255
rect 273029 168317 273063 168351
rect 246901 161449 246935 161483
rect 259321 164169 259355 164203
rect 246809 159477 246843 159511
rect 273029 163489 273063 163523
rect 328321 182121 328355 182155
rect 328321 176545 328355 176579
rect 371929 179333 371963 179367
rect 285173 172533 285207 172567
rect 278825 171105 278859 171139
rect 275605 163489 275639 163523
rect 305137 164169 305171 164203
rect 259321 157301 259355 157335
rect 268521 161245 268555 161279
rect 246809 157097 246843 157131
rect 285265 157369 285299 157403
rect 268521 157097 268555 157131
rect 273029 157301 273063 157335
rect 246625 153221 246659 153255
rect 268705 154377 268739 154411
rect 273029 147645 273063 147679
rect 275605 157301 275639 157335
rect 285081 156757 285115 156791
rect 275605 147645 275639 147679
rect 278733 149821 278767 149855
rect 268705 147577 268739 147611
rect 225373 144857 225407 144891
rect 135673 143429 135707 143463
rect 135673 133909 135707 133943
rect 152233 143429 152267 143463
rect 152233 133909 152267 133943
rect 170173 143429 170207 143463
rect 170173 133909 170207 133943
rect 190873 143429 190907 143463
rect 190873 133909 190907 133943
rect 214333 143429 214367 143463
rect 273029 143701 273063 143735
rect 278733 142137 278767 142171
rect 273029 139417 273063 139451
rect 279745 139349 279779 139383
rect 225373 135337 225407 135371
rect 271465 137921 271499 137955
rect 214333 133909 214367 133943
rect 259413 135201 259447 135235
rect 259413 128265 259447 128299
rect 268705 135201 268739 135235
rect 553905 164169 553939 164203
rect 371929 161449 371963 161483
rect 385545 162809 385579 162843
rect 305137 157301 305171 157335
rect 385545 153221 385579 153255
rect 392445 162809 392479 162843
rect 392445 153221 392479 153255
rect 529065 162809 529099 162843
rect 529065 153221 529099 153255
rect 535965 162809 535999 162843
rect 535965 153221 535999 153255
rect 552525 162809 552559 162843
rect 553905 154649 553939 154683
rect 571845 162809 571879 162843
rect 552525 153221 552559 153255
rect 571845 153221 571879 153255
rect 373125 153153 373159 153187
rect 373125 145129 373159 145163
rect 285265 138057 285299 138091
rect 285633 144857 285667 144891
rect 553905 144857 553939 144891
rect 319949 143497 319983 143531
rect 285633 137921 285667 137955
rect 309093 140709 309127 140743
rect 285081 137853 285115 137887
rect 285449 135541 285483 135575
rect 285449 135269 285483 135303
rect 309093 134657 309127 134691
rect 319949 133909 319983 133943
rect 328413 143497 328447 143531
rect 385545 143497 385579 143531
rect 328413 133909 328447 133943
rect 371929 135201 371963 135235
rect 279745 129761 279779 129795
rect 271465 128469 271499 128503
rect 268705 128265 268739 128299
rect 385545 133909 385579 133943
rect 392445 143497 392479 143531
rect 392445 133909 392479 133943
rect 529065 143497 529099 143531
rect 529065 133909 529099 133943
rect 535965 143497 535999 143531
rect 535965 133909 535999 133943
rect 552249 143497 552283 143531
rect 553905 135337 553939 135371
rect 571845 143497 571879 143531
rect 552249 133909 552283 133943
rect 571845 133909 571879 133943
rect 371929 128265 371963 128299
rect 552249 133705 552283 133739
rect 242853 125545 242887 125579
rect 135673 124117 135707 124151
rect 91513 115753 91547 115787
rect 135673 114529 135707 114563
rect 152233 124117 152267 124151
rect 152233 114529 152267 114563
rect 170173 124117 170207 124151
rect 170173 114529 170207 114563
rect 190873 124117 190907 124151
rect 190873 114529 190907 114563
rect 214333 124117 214367 124151
rect 229789 118745 229823 118779
rect 305137 125545 305171 125579
rect 242853 116705 242887 116739
rect 272845 121397 272879 121431
rect 229789 114665 229823 114699
rect 235585 115753 235619 115787
rect 214333 114529 214367 114563
rect 242853 114461 242887 114495
rect 235585 108953 235619 108987
rect 242669 111129 242703 111163
rect 91513 106301 91547 106335
rect 235493 106233 235527 106267
rect 135673 104805 135707 104839
rect 135673 95285 135707 95319
rect 152233 104805 152267 104839
rect 152233 95285 152267 95319
rect 170173 104805 170207 104839
rect 170173 95285 170207 95319
rect 190873 104805 190907 104839
rect 190873 95285 190907 95319
rect 214333 104805 214367 104839
rect 229789 103445 229823 103479
rect 214333 95285 214367 95319
rect 272845 111809 272879 111843
rect 285633 120037 285667 120071
rect 309001 125545 309035 125579
rect 309001 119357 309035 119391
rect 341109 125545 341143 125579
rect 305137 118473 305171 118507
rect 552249 125409 552283 125443
rect 341109 116025 341143 116059
rect 373125 124117 373159 124151
rect 285633 111265 285667 111299
rect 357945 115753 357979 115787
rect 242853 110517 242887 110551
rect 320133 109021 320167 109055
rect 242669 104873 242703 104907
rect 275513 106301 275547 106335
rect 235493 96645 235527 96679
rect 242025 101405 242059 101439
rect 235585 96577 235619 96611
rect 320133 104873 320167 104907
rect 328413 109021 328447 109055
rect 373125 114529 373159 114563
rect 385545 124117 385579 124151
rect 385545 114529 385579 114563
rect 392445 124117 392479 124151
rect 392445 114529 392479 114563
rect 529065 124117 529099 124151
rect 529065 114529 529099 114563
rect 535965 124117 535999 124151
rect 535965 114529 535999 114563
rect 571845 124117 571879 124151
rect 571845 114529 571879 114563
rect 357945 106301 357979 106335
rect 553905 109701 553939 109735
rect 328413 104873 328447 104907
rect 305045 104805 305079 104839
rect 285265 102357 285299 102391
rect 285265 102153 285299 102187
rect 275513 100725 275547 100759
rect 373125 104805 373159 104839
rect 305045 99297 305079 99331
rect 308909 103445 308943 103479
rect 242025 93857 242059 93891
rect 268705 96577 268739 96611
rect 235585 89641 235619 89675
rect 246533 90049 246567 90083
rect 308909 93857 308943 93891
rect 319949 103445 319983 103479
rect 373125 95285 373159 95319
rect 385545 104805 385579 104839
rect 385545 95285 385579 95319
rect 392445 104805 392479 104839
rect 392445 95285 392479 95319
rect 529065 104805 529099 104839
rect 529065 95285 529099 95319
rect 535965 104805 535999 104839
rect 535965 95285 535999 95319
rect 552525 103445 552559 103479
rect 319949 93857 319983 93891
rect 371929 95081 371963 95115
rect 268705 89641 268739 89675
rect 246533 88417 246567 88451
rect 242485 87193 242519 87227
rect 242485 86853 242519 86887
rect 305137 86921 305171 86955
rect 229881 85561 229915 85595
rect 135673 85493 135707 85527
rect 91513 77129 91547 77163
rect 135673 75905 135707 75939
rect 152233 85493 152267 85527
rect 152233 75905 152267 75939
rect 170173 85493 170207 85527
rect 170173 75905 170207 75939
rect 190873 85493 190907 85527
rect 190873 75905 190907 75939
rect 214333 85493 214367 85527
rect 242485 85493 242519 85527
rect 242485 85289 242519 85323
rect 276617 82773 276651 82807
rect 271373 81481 271407 81515
rect 229973 80121 230007 80155
rect 271373 80053 271407 80087
rect 229973 79849 230007 79883
rect 214333 75905 214367 75939
rect 235493 77129 235527 77163
rect 91513 67609 91547 67643
rect 271465 76585 271499 76619
rect 235493 67609 235527 67643
rect 246717 70465 246751 70499
rect 246717 66249 246751 66283
rect 135673 66181 135707 66215
rect 91513 57885 91547 57919
rect 135673 56661 135707 56695
rect 152233 66181 152267 66215
rect 152233 56661 152267 56695
rect 170173 66181 170207 66215
rect 170173 56661 170207 56695
rect 190873 66181 190907 66215
rect 190873 56661 190907 56695
rect 214333 66181 214367 66215
rect 285265 82773 285299 82807
rect 341109 86921 341143 86955
rect 305137 79849 305171 79883
rect 319949 85493 319983 85527
rect 285265 77945 285299 77979
rect 553905 96713 553939 96747
rect 571845 104805 571879 104839
rect 571845 95285 571879 95319
rect 552525 93857 552559 93891
rect 552433 87125 552467 87159
rect 552433 86853 552467 86887
rect 371929 85561 371963 85595
rect 341109 77401 341143 77435
rect 373125 85493 373159 85527
rect 319949 75905 319983 75939
rect 341109 77129 341143 77163
rect 279929 74613 279963 74647
rect 279929 74409 279963 74443
rect 276617 73185 276651 73219
rect 271465 63529 271499 63563
rect 275605 73117 275639 73151
rect 275605 63529 275639 63563
rect 277077 67609 277111 67643
rect 341109 67609 341143 67643
rect 357945 77129 357979 77163
rect 373125 75905 373159 75939
rect 385545 85493 385579 85527
rect 385545 75905 385579 75939
rect 392445 85493 392479 85527
rect 392445 75905 392479 75939
rect 529065 85493 529099 85527
rect 529065 75905 529099 75939
rect 535965 85493 535999 85527
rect 552341 85493 552375 85527
rect 552341 77129 552375 77163
rect 571845 85493 571879 85527
rect 535965 75905 535999 75939
rect 571845 75905 571879 75939
rect 357945 67609 357979 67643
rect 242485 63461 242519 63495
rect 214333 56661 214367 56695
rect 235401 57885 235435 57919
rect 91513 48297 91547 48331
rect 235401 48297 235435 48331
rect 135673 46869 135707 46903
rect 91513 38505 91547 38539
rect 135673 37281 135707 37315
rect 152233 46869 152267 46903
rect 152233 37281 152267 37315
rect 170173 46869 170207 46903
rect 170173 37281 170207 37315
rect 190873 46869 190907 46903
rect 190873 37281 190907 37315
rect 214333 46869 214367 46903
rect 214333 37281 214367 37315
rect 225373 46869 225407 46903
rect 331265 67541 331299 67575
rect 308909 66181 308943 66215
rect 277077 62713 277111 62747
rect 278641 64821 278675 64855
rect 275605 57953 275639 57987
rect 272845 57885 272879 57919
rect 242485 45577 242519 45611
rect 246901 55165 246935 55199
rect 275605 52445 275639 52479
rect 276525 57273 276559 57307
rect 272845 48297 272879 48331
rect 246901 45577 246935 45611
rect 259321 48229 259355 48263
rect 275605 46937 275639 46971
rect 259321 38709 259355 38743
rect 272845 46869 272879 46903
rect 225373 37281 225407 37315
rect 278641 55233 278675 55267
rect 279745 64821 279779 64855
rect 285265 64821 285299 64855
rect 308909 56661 308943 56695
rect 320133 66181 320167 66215
rect 385545 66181 385579 66215
rect 331265 62781 331299 62815
rect 371929 64821 371963 64855
rect 320133 56661 320167 56695
rect 357945 57885 357979 57919
rect 285265 56457 285299 56491
rect 279745 55233 279779 55267
rect 385545 56661 385579 56695
rect 392445 66181 392479 66215
rect 392445 56661 392479 56695
rect 529065 66181 529099 66215
rect 529065 56661 529099 56695
rect 535965 66181 535999 66215
rect 535965 56661 535999 56695
rect 552525 66181 552559 66215
rect 552525 56661 552559 56695
rect 571845 66181 571879 66215
rect 571845 56661 571879 56695
rect 371929 55233 371963 55267
rect 278733 48297 278767 48331
rect 357945 48297 357979 48331
rect 278733 45577 278767 45611
rect 319949 46869 319983 46903
rect 276525 44149 276559 44183
rect 275605 42789 275639 42823
rect 285725 42041 285759 42075
rect 272845 37281 272879 37315
rect 275605 37961 275639 37995
rect 91513 28985 91547 29019
rect 235493 31773 235527 31807
rect 235493 28985 235527 29019
rect 254813 28917 254847 28951
rect 135305 27557 135339 27591
rect 91513 19261 91547 19295
rect 135305 18037 135339 18071
rect 151865 27557 151899 27591
rect 151865 18037 151899 18071
rect 169713 27557 169747 27591
rect 169713 18037 169747 18071
rect 225097 27557 225131 27591
rect 242577 27557 242611 27591
rect 242577 22661 242611 22695
rect 272845 27557 272879 27591
rect 268429 26197 268463 26231
rect 268429 25993 268463 26027
rect 254813 21369 254847 21403
rect 225097 18037 225131 18071
rect 273029 26197 273063 26231
rect 273029 25993 273063 26027
rect 328229 46869 328263 46903
rect 319949 37281 319983 37315
rect 320317 38505 320351 38539
rect 385545 46869 385579 46903
rect 328229 37281 328263 37315
rect 357945 38505 357979 38539
rect 320317 31841 320351 31875
rect 341017 31841 341051 31875
rect 285725 28985 285759 29019
rect 341017 28985 341051 29019
rect 392445 46869 392479 46903
rect 392445 46665 392479 46699
rect 529065 46869 529099 46903
rect 385545 37281 385579 37315
rect 529065 37281 529099 37315
rect 535965 46869 535999 46903
rect 535965 37281 535999 37315
rect 552525 46869 552559 46903
rect 553813 46869 553847 46903
rect 553813 38369 553847 38403
rect 571845 46869 571879 46903
rect 552525 37281 552559 37315
rect 571845 37281 571879 37315
rect 357945 28985 357979 29019
rect 285173 28917 285207 28951
rect 278825 27625 278859 27659
rect 278825 26265 278859 26299
rect 275605 24837 275639 24871
rect 305137 27557 305171 27591
rect 285173 19329 285207 19363
rect 285725 24157 285759 24191
rect 285725 19329 285759 19363
rect 272845 18037 272879 18071
rect 529065 27557 529099 27591
rect 305137 18037 305171 18071
rect 308265 19261 308299 19295
rect 176705 11305 176739 11339
rect 129049 11169 129083 11203
rect 128957 11101 128991 11135
rect 123345 11033 123379 11067
rect 148277 11169 148311 11203
rect 138249 11101 138283 11135
rect 133833 11033 133867 11067
rect 129049 10965 129083 10999
rect 133649 10965 133683 10999
rect 123345 10489 123379 10523
rect 128865 10761 128899 10795
rect 128957 10761 128991 10795
rect 133557 10693 133591 10727
rect 133741 10625 133775 10659
rect 133741 10489 133775 10523
rect 133649 10421 133683 10455
rect 133833 10421 133867 10455
rect 133925 10489 133959 10523
rect 133557 10217 133591 10251
rect 128957 10149 128991 10183
rect 133373 10149 133407 10183
rect 138157 10149 138191 10183
rect 91513 9673 91547 9707
rect 147909 11101 147943 11135
rect 138525 11033 138559 11067
rect 138341 10489 138375 10523
rect 138433 10149 138467 10183
rect 148093 11033 148127 11067
rect 148093 10761 148127 10795
rect 148185 11033 148219 11067
rect 157753 11169 157787 11203
rect 148277 10761 148311 10795
rect 148369 11101 148403 11135
rect 143309 10693 143343 10727
rect 147909 10693 147943 10727
rect 148001 10693 148035 10727
rect 148185 10693 148219 10727
rect 157661 11033 157695 11067
rect 148369 10693 148403 10727
rect 153153 10761 153187 10795
rect 152877 10693 152911 10727
rect 143493 10625 143527 10659
rect 138525 10149 138559 10183
rect 143217 10217 143251 10251
rect 157661 10217 157695 10251
rect 148001 10149 148035 10183
rect 138341 10081 138375 10115
rect 143401 10081 143435 10115
rect 147817 10081 147851 10115
rect 147909 10081 147943 10115
rect 138341 9605 138375 9639
rect 138709 9605 138743 9639
rect 147909 9605 147943 9639
rect 148001 9605 148035 9639
rect 148093 10149 148127 10183
rect 157753 10149 157787 10183
rect 157845 11033 157879 11067
rect 138525 9537 138559 9571
rect 148093 9537 148127 9571
rect 148277 9605 148311 9639
rect 148093 9333 148127 9367
rect 18465 9129 18499 9163
rect 18465 8925 18499 8959
rect 28033 9129 28067 9163
rect 36405 9129 36439 9163
rect 28033 8925 28067 8959
rect 31529 8993 31563 9027
rect 36405 8993 36439 9027
rect 42661 9129 42695 9163
rect 31529 8857 31563 8891
rect 37785 8925 37819 8959
rect 54253 9129 54287 9163
rect 42661 8857 42695 8891
rect 47353 8925 47387 8959
rect 37785 8585 37819 8619
rect 65385 9129 65419 9163
rect 65385 8993 65419 9027
rect 75045 9129 75079 9163
rect 75045 8993 75079 9027
rect 81209 9129 81243 9163
rect 54253 8857 54287 8891
rect 57105 8925 57139 8959
rect 57105 8789 57139 8823
rect 66673 8925 66707 8959
rect 66673 8789 66707 8823
rect 68145 8925 68179 8959
rect 92893 9129 92927 9163
rect 81209 8857 81243 8891
rect 85993 8993 86027 9027
rect 68145 8789 68179 8823
rect 104025 9129 104059 9163
rect 104025 8993 104059 9027
rect 113685 9129 113719 9163
rect 113685 8993 113719 9027
rect 116261 9129 116295 9163
rect 116261 8993 116295 9027
rect 140089 8993 140123 9027
rect 148093 8993 148127 9027
rect 85901 8857 85935 8891
rect 85993 8857 86027 8891
rect 92893 8857 92927 8891
rect 115065 8925 115099 8959
rect 85717 8789 85751 8823
rect 47353 8585 47387 8619
rect 115065 8585 115099 8619
rect 124633 8925 124667 8959
rect 134385 8925 134419 8959
rect 138525 8925 138559 8959
rect 140273 8857 140307 8891
rect 148277 8857 148311 8891
rect 167597 11033 167631 11067
rect 179189 11305 179223 11339
rect 177073 11169 177107 11203
rect 176889 11101 176923 11135
rect 176705 10761 176739 10795
rect 176797 11033 176831 11067
rect 172381 10693 172415 10727
rect 172197 10625 172231 10659
rect 234757 11237 234791 11271
rect 179189 11101 179223 11135
rect 187009 11101 187043 11135
rect 177073 10761 177107 10795
rect 186917 11033 186951 11067
rect 186917 10761 186951 10795
rect 225557 11101 225591 11135
rect 196209 11033 196243 11067
rect 176889 10693 176923 10727
rect 176981 10693 177015 10727
rect 187009 10693 187043 10727
rect 191793 10761 191827 10795
rect 191517 10693 191551 10727
rect 167505 10217 167539 10251
rect 196209 10149 196243 10183
rect 196577 11033 196611 11067
rect 157845 8857 157879 8891
rect 162537 9605 162571 9639
rect 134385 8789 134419 8823
rect 138433 8789 138467 8823
rect 124633 8585 124667 8619
rect 230065 10761 230099 10795
rect 230157 10761 230191 10795
rect 230341 10693 230375 10727
rect 230157 10625 230191 10659
rect 232365 10217 232399 10251
rect 232457 10217 232491 10251
rect 225557 10081 225591 10115
rect 238345 11169 238379 11203
rect 235493 11033 235527 11067
rect 235401 10761 235435 10795
rect 235493 10761 235527 10795
rect 234941 10693 234975 10727
rect 235125 10693 235159 10727
rect 235309 10217 235343 10251
rect 234941 10149 234975 10183
rect 238345 10625 238379 10659
rect 235401 10149 235435 10183
rect 244877 10149 244911 10183
rect 254537 10081 254571 10115
rect 244877 9673 244911 9707
rect 244969 9673 245003 9707
rect 254353 9673 254387 9707
rect 244785 9469 244819 9503
rect 244877 9469 244911 9503
rect 244785 9333 244819 9367
rect 254537 9605 254571 9639
rect 254629 9877 254663 9911
rect 254353 9129 254387 9163
rect 234757 9061 234791 9095
rect 162629 8993 162663 9027
rect 172289 8993 172323 9027
rect 162629 8789 162663 8823
rect 162905 8857 162939 8891
rect 162905 8585 162939 8619
rect 172289 8585 172323 8619
rect 181949 8993 181983 9027
rect 181949 8585 181983 8619
rect 191609 8993 191643 9027
rect 196577 8993 196611 9027
rect 201269 8993 201303 9027
rect 191609 8585 191643 8619
rect 201269 8585 201303 8619
rect 210929 8993 210963 9027
rect 162537 8517 162571 8551
rect 186641 8381 186675 8415
rect 177165 8313 177199 8347
rect 196393 8381 196427 8415
rect 195013 8313 195047 8347
rect 186641 7769 186675 7803
rect 186733 7769 186767 7803
rect 177165 5865 177199 5899
rect 210929 8313 210963 8347
rect 215897 8993 215931 9027
rect 259137 9877 259171 9911
rect 254721 9673 254755 9707
rect 254721 8857 254755 8891
rect 254813 9673 254847 9707
rect 254445 8789 254479 8823
rect 373125 17833 373159 17867
rect 331449 11305 331483 11339
rect 331265 11169 331299 11203
rect 331265 10217 331299 10251
rect 333749 11305 333783 11339
rect 331541 11237 331575 11271
rect 331909 11101 331943 11135
rect 331725 11033 331759 11067
rect 331541 10761 331575 10795
rect 331633 10761 331667 10795
rect 331449 10149 331483 10183
rect 331541 10149 331575 10183
rect 333749 10965 333783 10999
rect 340925 11305 340959 11339
rect 331909 10693 331943 10727
rect 341293 11237 341327 11271
rect 341017 11169 341051 11203
rect 340925 10693 340959 10727
rect 341109 11033 341143 11067
rect 331725 10625 331759 10659
rect 341109 10625 341143 10659
rect 341293 10693 341327 10727
rect 350953 11237 350987 11271
rect 341201 10625 341235 10659
rect 331173 10013 331207 10047
rect 331541 10013 331575 10047
rect 308265 9673 308299 9707
rect 259137 9469 259171 9503
rect 346537 9333 346571 9367
rect 350677 9333 350711 9367
rect 350769 9401 350803 9435
rect 341293 9129 341327 9163
rect 254813 8789 254847 8823
rect 341201 9061 341235 9095
rect 215897 8313 215931 8347
rect 225373 8381 225407 8415
rect 225189 8313 225223 8347
rect 272845 8245 272879 8279
rect 341201 8245 341235 8279
rect 196393 7837 196427 7871
rect 232917 7837 232951 7871
rect 195013 7701 195047 7735
rect 215897 6273 215931 6307
rect 215805 6137 215839 6171
rect 186733 5797 186767 5831
rect 196117 5661 196151 5695
rect 138801 4233 138835 4267
rect 123345 4165 123379 4199
rect 44777 3621 44811 3655
rect 36405 3485 36439 3519
rect 45973 3485 46007 3519
rect 36405 3145 36439 3179
rect 40177 3349 40211 3383
rect 44777 3349 44811 3383
rect 45881 3417 45915 3451
rect 40177 3077 40211 3111
rect 45973 3145 46007 3179
rect 56277 3485 56311 3519
rect 65201 3485 65235 3519
rect 56277 3145 56311 3179
rect 56369 3417 56403 3451
rect 45881 3077 45915 3111
rect 56369 3077 56403 3111
rect 65293 3485 65327 3519
rect 65293 3145 65327 3179
rect 75045 3485 75079 3519
rect 65201 3077 65235 3111
rect 84613 3485 84647 3519
rect 75045 2941 75079 2975
rect 75137 3417 75171 3451
rect 75137 2873 75171 2907
rect 84521 3417 84555 3451
rect 84613 2941 84647 2975
rect 93721 3485 93755 3519
rect 84521 2873 84555 2907
rect 103933 3485 103967 3519
rect 103841 2941 103875 2975
rect 93721 2873 93755 2907
rect 108625 2873 108659 2907
rect 113501 2873 113535 2907
rect 108809 2805 108843 2839
rect 112765 2805 112799 2839
rect 113409 2805 113443 2839
rect 113501 2601 113535 2635
rect 113685 2805 113719 2839
rect 113685 2601 113719 2635
rect 128957 4165 128991 4199
rect 133005 4165 133039 4199
rect 133005 3961 133039 3995
rect 134293 4165 134327 4199
rect 134293 3961 134327 3995
rect 138433 3961 138467 3995
rect 128221 3485 128255 3519
rect 128957 3485 128991 3519
rect 138341 3485 138375 3519
rect 147909 4165 147943 4199
rect 148001 4165 148035 4199
rect 138801 3485 138835 3519
rect 138893 3621 138927 3655
rect 138893 3485 138927 3519
rect 142757 3621 142791 3655
rect 129049 3417 129083 3451
rect 132821 3417 132855 3451
rect 123345 2601 123379 2635
rect 133373 3417 133407 3451
rect 132821 2601 132855 2635
rect 132913 2533 132947 2567
rect 133373 2601 133407 2635
rect 142389 3417 142423 3451
rect 142389 2601 142423 2635
rect 142573 3417 142607 3451
rect 133281 2533 133315 2567
rect 148001 3485 148035 3519
rect 157753 4233 157787 4267
rect 152233 4165 152267 4199
rect 148461 3621 148495 3655
rect 149565 3621 149599 3655
rect 152141 3621 152175 3655
rect 152233 3621 152267 3655
rect 148093 3485 148127 3519
rect 142757 2601 142791 2635
rect 157753 3485 157787 3519
rect 157845 4233 157879 4267
rect 159133 4165 159167 4199
rect 177441 4233 177475 4267
rect 190965 4233 190999 4267
rect 159133 3621 159167 3655
rect 162077 3621 162111 3655
rect 162721 3621 162755 3655
rect 163365 3621 163399 3655
rect 166309 3621 166343 3655
rect 167413 3621 167447 3655
rect 167505 3621 167539 3655
rect 167597 4165 167631 4199
rect 167689 4165 167723 4199
rect 171461 4165 171495 4199
rect 167597 3621 167631 3655
rect 157845 3485 157879 3519
rect 161617 3485 161651 3519
rect 152141 2601 152175 2635
rect 152325 3417 152359 3451
rect 142573 2533 142607 2567
rect 152509 3417 152543 3451
rect 152509 2601 152543 2635
rect 161617 2601 161651 2635
rect 161893 3485 161927 3519
rect 152325 2533 152359 2567
rect 162077 2601 162111 2635
rect 171461 2601 171495 2635
rect 171737 4165 171771 4199
rect 176889 4165 176923 4199
rect 176981 4165 177015 4199
rect 176981 3621 177015 3655
rect 177073 3621 177107 3655
rect 177165 3485 177199 3519
rect 177257 4165 177291 4199
rect 186733 4165 186767 4199
rect 177257 3485 177291 3519
rect 181121 3621 181155 3655
rect 171737 2601 171771 2635
rect 181213 3553 181247 3587
rect 181489 3553 181523 3587
rect 181121 2601 181155 2635
rect 181397 3485 181431 3519
rect 186733 3485 186767 3519
rect 190781 4165 190815 4199
rect 187101 3417 187135 3451
rect 186917 3077 186951 3111
rect 187009 3009 187043 3043
rect 186825 2873 186859 2907
rect 186917 2873 186951 2907
rect 187009 2805 187043 2839
rect 181397 2601 181431 2635
rect 190781 2601 190815 2635
rect 161893 2533 161927 2567
rect 191057 4165 191091 4199
rect 191057 2601 191091 2635
rect 220681 5049 220715 5083
rect 220497 4981 220531 5015
rect 227581 5049 227615 5083
rect 229329 5049 229363 5083
rect 229421 5049 229455 5083
rect 227765 4981 227799 5015
rect 220681 4777 220715 4811
rect 220773 4777 220807 4811
rect 206145 4233 206179 4267
rect 200257 4165 200291 4199
rect 196209 3009 196243 3043
rect 196577 3009 196611 3043
rect 198509 2941 198543 2975
rect 196117 2601 196151 2635
rect 196209 2873 196243 2907
rect 196485 2873 196519 2907
rect 196301 2805 196335 2839
rect 196209 2601 196243 2635
rect 198509 2601 198543 2635
rect 200717 4165 200751 4199
rect 200257 2601 200291 2635
rect 190965 2533 190999 2567
rect 200533 2533 200567 2567
rect 215897 4233 215931 4267
rect 217461 4233 217495 4267
rect 217461 3961 217495 3995
rect 218565 4233 218599 4267
rect 220681 4233 220715 4267
rect 220497 4165 220531 4199
rect 218565 3961 218599 3995
rect 219669 3961 219703 3995
rect 206145 3485 206179 3519
rect 210377 3621 210411 3655
rect 215897 3621 215931 3655
rect 209917 3417 209951 3451
rect 206053 3077 206087 3111
rect 205961 3009 205995 3043
rect 205869 2941 205903 2975
rect 206145 2941 206179 2975
rect 200717 2601 200751 2635
rect 209917 2601 209951 2635
rect 210193 3417 210227 3451
rect 200625 2533 200659 2567
rect 210377 2601 210411 2635
rect 219853 3961 219887 3995
rect 219945 3961 219979 3995
rect 219945 3621 219979 3655
rect 219761 2601 219795 2635
rect 210193 2533 210227 2567
rect 225373 3417 225407 3451
rect 225465 3417 225499 3451
rect 229789 4981 229823 5015
rect 229421 2601 229455 2635
rect 229697 4029 229731 4063
rect 219945 2533 219979 2567
rect 259045 6341 259079 6375
rect 230341 3961 230375 3995
rect 232917 3961 232951 3995
rect 235217 6273 235251 6307
rect 234941 3893 234975 3927
rect 230341 3689 230375 3723
rect 235033 3553 235067 3587
rect 229697 2533 229731 2567
rect 245061 6273 245095 6307
rect 245061 5253 245095 5287
rect 254169 6273 254203 6307
rect 254169 5253 254203 5287
rect 254353 5185 254387 5219
rect 341293 8041 341327 8075
rect 339637 7905 339671 7939
rect 336509 7837 336543 7871
rect 323813 7225 323847 7259
rect 322157 7157 322191 7191
rect 322157 6953 322191 6987
rect 321789 6885 321823 6919
rect 317189 6341 317223 6375
rect 272845 6137 272879 6171
rect 314613 6273 314647 6307
rect 312313 6069 312347 6103
rect 312221 5729 312255 5763
rect 312129 5661 312163 5695
rect 302561 5593 302595 5627
rect 264197 5321 264231 5355
rect 264289 5321 264323 5355
rect 259229 5253 259263 5287
rect 263921 5253 263955 5287
rect 259413 5185 259447 5219
rect 259045 4709 259079 4743
rect 263921 4709 263955 4743
rect 264013 4709 264047 4743
rect 263921 4097 263955 4131
rect 302561 5253 302595 5287
rect 302653 5253 302687 5287
rect 301181 5117 301215 5151
rect 301089 4777 301123 4811
rect 264473 4505 264507 4539
rect 264565 4641 264599 4675
rect 264289 4097 264323 4131
rect 254353 4029 254387 4063
rect 235309 3689 235343 3723
rect 235309 3553 235343 3587
rect 249569 3689 249603 3723
rect 249569 3485 249603 3519
rect 267509 4573 267543 4607
rect 267417 4437 267451 4471
rect 267509 4437 267543 4471
rect 268889 4573 268923 4607
rect 268889 4165 268923 4199
rect 267417 4097 267451 4131
rect 301089 4097 301123 4131
rect 302561 5049 302595 5083
rect 302837 5117 302871 5151
rect 307437 5117 307471 5151
rect 307621 4981 307655 5015
rect 302745 4777 302779 4811
rect 302837 4777 302871 4811
rect 307621 4641 307655 4675
rect 312681 5729 312715 5763
rect 312313 5525 312347 5559
rect 312497 5661 312531 5695
rect 312221 5321 312255 5355
rect 312313 5321 312347 5355
rect 312129 5049 312163 5083
rect 340925 7497 340959 7531
rect 341293 7497 341327 7531
rect 341201 7361 341235 7395
rect 336509 6953 336543 6987
rect 321881 6409 321915 6443
rect 323813 6409 323847 6443
rect 322065 6341 322099 6375
rect 328689 6273 328723 6307
rect 328873 6273 328907 6307
rect 321789 6205 321823 6239
rect 317189 5729 317223 5763
rect 314613 5661 314647 5695
rect 317281 5321 317315 5355
rect 312681 5253 312715 5287
rect 317097 5253 317131 5287
rect 312405 5185 312439 5219
rect 312497 5185 312531 5219
rect 341385 5321 341419 5355
rect 332461 5253 332495 5287
rect 341293 5253 341327 5287
rect 346353 5321 346387 5355
rect 346445 5321 346479 5355
rect 345341 5253 345375 5287
rect 346077 5253 346111 5287
rect 317281 5117 317315 5151
rect 317373 5117 317407 5151
rect 332369 5117 332403 5151
rect 332461 5117 332495 5151
rect 346261 5117 346295 5151
rect 307713 4641 307747 4675
rect 312221 4641 312255 4675
rect 312405 4709 312439 4743
rect 302745 4573 302779 4607
rect 302653 4505 302687 4539
rect 302561 4233 302595 4267
rect 283977 4029 284011 4063
rect 299709 4029 299743 4063
rect 301181 4029 301215 4063
rect 302653 4097 302687 4131
rect 312405 4097 312439 4131
rect 312497 4709 312531 4743
rect 284161 3893 284195 3927
rect 298513 3893 298547 3927
rect 278733 3621 278767 3655
rect 264565 3349 264599 3383
rect 268889 3553 268923 3587
rect 278549 3485 278583 3519
rect 278641 3485 278675 3519
rect 275697 3417 275731 3451
rect 275697 3009 275731 3043
rect 312497 4029 312531 4063
rect 345433 5049 345467 5083
rect 345433 4641 345467 4675
rect 346261 4777 346295 4811
rect 346353 4777 346387 4811
rect 332369 4573 332403 4607
rect 341385 4505 341419 4539
rect 331541 4233 331575 4267
rect 324181 4165 324215 4199
rect 312589 4029 312623 4063
rect 322893 4097 322927 4131
rect 302469 3961 302503 3995
rect 322893 3893 322927 3927
rect 324181 3893 324215 3927
rect 325929 3893 325963 3927
rect 326021 3893 326055 3927
rect 299709 3689 299743 3723
rect 300997 3553 301031 3587
rect 331541 3689 331575 3723
rect 331633 4165 331667 4199
rect 331633 3689 331667 3723
rect 326021 3485 326055 3519
rect 326205 3485 326239 3519
rect 326297 3485 326331 3519
rect 341385 3485 341419 3519
rect 345617 4505 345651 4539
rect 300997 3417 301031 3451
rect 301089 3417 301123 3451
rect 278457 3009 278491 3043
rect 278549 3349 278583 3383
rect 298513 3349 298547 3383
rect 298605 3349 298639 3383
rect 278549 3009 278583 3043
rect 268889 2805 268923 2839
rect 301089 3145 301123 3179
rect 298605 2805 298639 2839
rect 309093 2805 309127 2839
rect 235217 561 235251 595
rect 326205 2601 326239 2635
rect 346169 4437 346203 4471
rect 346169 4233 346203 4267
rect 351321 11169 351355 11203
rect 351045 9401 351079 9435
rect 350953 9333 350987 9367
rect 350677 9129 350711 9163
rect 350861 9129 350895 9163
rect 350769 9061 350803 9095
rect 350953 9061 350987 9095
rect 351045 9129 351079 9163
rect 351137 9129 351171 9163
rect 355921 9333 355955 9367
rect 355921 9061 355955 9095
rect 356013 9333 356047 9367
rect 351321 8993 351355 9027
rect 355737 8993 355771 9027
rect 351137 8925 351171 8959
rect 355737 8449 355771 8483
rect 355553 8381 355587 8415
rect 409097 11101 409131 11135
rect 409097 10489 409131 10523
rect 418481 11101 418515 11135
rect 418757 11101 418791 11135
rect 418481 10489 418515 10523
rect 418573 11033 418607 11067
rect 418573 10489 418607 10523
rect 418665 10557 418699 10591
rect 418757 10557 418791 10591
rect 423357 10557 423391 10591
rect 423541 10489 423575 10523
rect 418665 10421 418699 10455
rect 418665 9605 418699 9639
rect 418757 9537 418791 9571
rect 428325 9673 428359 9707
rect 529065 9673 529099 9707
rect 535965 27557 535999 27591
rect 552525 27557 552559 27591
rect 535965 9673 535999 9707
rect 541485 19261 541519 19295
rect 541485 9673 541519 9707
rect 571845 27557 571879 27591
rect 552525 9673 552559 9707
rect 560805 19261 560839 19295
rect 560805 9673 560839 9707
rect 571845 9673 571879 9707
rect 428325 9469 428359 9503
rect 373125 8381 373159 8415
rect 457489 8381 457523 8415
rect 350769 7905 350803 7939
rect 350953 7973 350987 8007
rect 457397 7769 457431 7803
rect 457305 7701 457339 7735
rect 357945 7429 357979 7463
rect 358129 7429 358163 7463
rect 346905 7361 346939 7395
rect 346997 7361 347031 7395
rect 424185 7361 424219 7395
rect 424185 6817 424219 6851
rect 433753 7361 433787 7395
rect 433753 6817 433787 6851
rect 457581 8313 457615 8347
rect 457581 7769 457615 7803
rect 457489 7701 457523 7735
rect 473865 7497 473899 7531
rect 474049 7497 474083 7531
rect 457397 6817 457431 6851
rect 462825 7361 462859 7395
rect 457305 6749 457339 6783
rect 462825 6681 462859 6715
rect 472393 7361 472427 7395
rect 473957 7361 473991 7395
rect 474141 7361 474175 7395
rect 473957 7225 473991 7259
rect 474141 7225 474175 7259
rect 472393 6681 472427 6715
rect 357945 6341 357979 6375
rect 358129 6341 358163 6375
rect 346905 6273 346939 6307
rect 346997 6273 347031 6307
rect 424185 6273 424219 6307
rect 424185 6069 424219 6103
rect 370733 5593 370767 5627
rect 346537 4505 346571 4539
rect 370825 5525 370859 5559
rect 346261 4233 346295 4267
rect 370457 3553 370491 3587
rect 345617 2533 345651 2567
rect 350769 3485 350803 3519
rect 360705 3485 360739 3519
rect 355093 2941 355127 2975
rect 355277 2941 355311 2975
rect 355369 2941 355403 2975
rect 370365 3485 370399 3519
rect 515173 5593 515207 5627
rect 505881 5525 505915 5559
rect 505789 5049 505823 5083
rect 505881 5049 505915 5083
rect 505605 4981 505639 5015
rect 418757 4097 418791 4131
rect 383981 3553 384015 3587
rect 355277 2601 355311 2635
rect 364661 2601 364695 2635
rect 364753 2805 364787 2839
rect 350769 2533 350803 2567
rect 364937 2805 364971 2839
rect 364937 2601 364971 2635
rect 374321 2601 374355 2635
rect 374597 2601 374631 2635
rect 364753 2533 364787 2567
rect 374689 2465 374723 2499
rect 383981 2601 384015 2635
rect 384073 3553 384107 3587
rect 390053 3417 390087 3451
rect 505697 4981 505731 5015
rect 505697 4097 505731 4131
rect 505605 4029 505639 4063
rect 515081 4981 515115 5015
rect 515173 4981 515207 5015
rect 529525 4777 529559 4811
rect 534585 4777 534619 4811
rect 559425 4709 559459 4743
rect 559517 4709 559551 4743
rect 534585 4641 534619 4675
rect 538725 4641 538759 4675
rect 529525 4233 529559 4267
rect 529617 4573 529651 4607
rect 549857 4641 549891 4675
rect 538725 4437 538759 4471
rect 548293 4573 548327 4607
rect 549765 4573 549799 4607
rect 548293 4437 548327 4471
rect 529617 4233 529651 4267
rect 515081 4097 515115 4131
rect 515265 4165 515299 4199
rect 515449 4097 515483 4131
rect 505789 3961 505823 3995
rect 418757 3009 418791 3043
rect 390053 2601 390087 2635
rect 420873 2805 420907 2839
rect 384073 2533 384107 2567
rect 374781 2397 374815 2431
rect 309093 561 309127 595
rect 420873 561 420907 595
<< metal1 >>
rect 1600 701712 583316 701808
rect 1600 701168 583316 701264
rect 290037 701131 290095 701137
rect 290037 701097 290049 701131
rect 290083 701128 290095 701131
rect 296293 701131 296351 701137
rect 296293 701128 296305 701131
rect 290083 701100 296305 701128
rect 290083 701097 290095 701100
rect 290037 701091 290095 701097
rect 296293 701097 296305 701100
rect 296339 701097 296351 701131
rect 296293 701091 296351 701097
rect 288749 701063 288807 701069
rect 288749 701029 288761 701063
rect 288795 701060 288807 701063
rect 288795 701032 292472 701060
rect 288795 701029 288807 701032
rect 288749 701023 288807 701029
rect 119374 700952 119380 701004
rect 119432 700992 119438 701004
rect 292337 700995 292395 701001
rect 292337 700992 292349 700995
rect 119432 700964 292349 700992
rect 119432 700952 119438 700964
rect 292337 700961 292349 700964
rect 292383 700961 292395 700995
rect 292337 700955 292395 700961
rect 249186 700884 249192 700936
rect 249244 700924 249250 700936
rect 250198 700924 250204 700936
rect 249244 700896 250204 700924
rect 249244 700884 249250 700896
rect 250198 700884 250204 700896
rect 250256 700884 250262 700936
rect 284698 700884 284704 700936
rect 284756 700924 284762 700936
rect 292444 700924 292472 701032
rect 292521 700995 292579 701001
rect 292521 700961 292533 700995
rect 292567 700992 292579 700995
rect 299970 700992 299976 701004
rect 292567 700964 299976 700992
rect 292567 700961 292579 700964
rect 292521 700955 292579 700961
rect 299970 700952 299976 700964
rect 300028 700952 300034 701004
rect 296201 700927 296259 700933
rect 296201 700924 296213 700927
rect 284756 700896 292380 700924
rect 292444 700896 296213 700924
rect 284756 700884 284762 700896
rect 184234 700816 184240 700868
rect 184292 700856 184298 700868
rect 185338 700856 185344 700868
rect 184292 700828 185344 700856
rect 184292 700816 184298 700828
rect 185338 700816 185344 700828
rect 185396 700816 185402 700868
rect 286078 700816 286084 700868
rect 286136 700856 286142 700868
rect 288749 700859 288807 700865
rect 288749 700856 288761 700859
rect 286136 700828 288761 700856
rect 286136 700816 286142 700828
rect 288749 700825 288761 700828
rect 288795 700825 288807 700859
rect 288749 700819 288807 700825
rect 288838 700816 288844 700868
rect 288896 700856 288902 700868
rect 292245 700859 292303 700865
rect 292245 700856 292257 700859
rect 288896 700828 292257 700856
rect 288896 700816 288902 700828
rect 292245 700825 292257 700828
rect 292291 700825 292303 700859
rect 292352 700856 292380 700896
rect 296201 700893 296213 700896
rect 296247 700893 296259 700927
rect 296201 700887 296259 700893
rect 296293 700927 296351 700933
rect 296293 700893 296305 700927
rect 296339 700924 296351 700927
rect 465478 700924 465484 700936
rect 296339 700896 465484 700924
rect 296339 700893 296351 700896
rect 296293 700887 296351 700893
rect 465478 700884 465484 700896
rect 465536 700884 465542 700936
rect 487098 700856 487104 700868
rect 292352 700828 487104 700856
rect 292245 700819 292303 700825
rect 487098 700816 487104 700828
rect 487156 700816 487162 700868
rect 97754 700748 97760 700800
rect 97812 700788 97818 700800
rect 301350 700788 301356 700800
rect 97812 700760 301356 700788
rect 97812 700748 97818 700760
rect 301350 700748 301356 700760
rect 301408 700748 301414 700800
rect 1600 700624 583316 700720
rect 76134 700544 76140 700596
rect 76192 700584 76198 700596
rect 301442 700584 301448 700596
rect 76192 700556 301448 700584
rect 76192 700544 76198 700556
rect 301442 700544 301448 700556
rect 301500 700544 301506 700596
rect 54514 700476 54520 700528
rect 54572 700516 54578 700528
rect 302730 700516 302736 700528
rect 54572 700488 302736 700516
rect 54572 700476 54578 700488
rect 302730 700476 302736 700488
rect 302788 700476 302794 700528
rect 280558 700408 280564 700460
rect 280616 700448 280622 700460
rect 530338 700448 530344 700460
rect 280616 700420 530344 700448
rect 280616 700408 280622 700420
rect 530338 700408 530344 700420
rect 530396 700408 530402 700460
rect 280466 700340 280472 700392
rect 280524 700380 280530 700392
rect 551958 700380 551964 700392
rect 280524 700352 551964 700380
rect 280524 700340 280530 700352
rect 551958 700340 551964 700352
rect 552016 700340 552022 700392
rect 32894 700272 32900 700324
rect 32952 700312 32958 700324
rect 305490 700312 305496 700324
rect 32952 700284 305496 700312
rect 32952 700272 32958 700284
rect 305490 700272 305496 700284
rect 305548 700272 305554 700324
rect 140994 700204 141000 700256
rect 141052 700244 141058 700256
rect 292245 700247 292303 700253
rect 292245 700244 292257 700247
rect 141052 700216 292257 700244
rect 141052 700204 141058 700216
rect 292245 700213 292257 700216
rect 292291 700213 292303 700247
rect 292245 700207 292303 700213
rect 292337 700247 292395 700253
rect 292337 700213 292349 700247
rect 292383 700244 292395 700247
rect 298590 700244 298596 700256
rect 292383 700216 298596 700244
rect 292383 700213 292395 700216
rect 292337 700207 292395 700213
rect 298590 700204 298596 700216
rect 298648 700204 298654 700256
rect 1600 700080 583316 700176
rect 162614 700000 162620 700052
rect 162672 700040 162678 700052
rect 292337 700043 292395 700049
rect 292337 700040 292349 700043
rect 162672 700012 292349 700040
rect 162672 700000 162678 700012
rect 292337 700009 292349 700012
rect 292383 700009 292395 700043
rect 292337 700003 292395 700009
rect 292429 700043 292487 700049
rect 292429 700009 292441 700043
rect 292475 700040 292487 700043
rect 296109 700043 296167 700049
rect 296109 700040 296121 700043
rect 292475 700012 296121 700040
rect 292475 700009 292487 700012
rect 292429 700003 292487 700009
rect 296109 700009 296121 700012
rect 296155 700009 296167 700043
rect 296109 700003 296167 700009
rect 270806 699932 270812 699984
rect 270864 699972 270870 699984
rect 278537 699975 278595 699981
rect 270864 699944 278488 699972
rect 270864 699932 270870 699944
rect 229593 699907 229651 699913
rect 229593 699873 229605 699907
rect 229639 699904 229651 699907
rect 239253 699907 239311 699913
rect 239253 699904 239265 699907
rect 229639 699876 239265 699904
rect 229639 699873 229651 699876
rect 229593 699867 229651 699873
rect 239253 699873 239265 699876
rect 239299 699873 239311 699907
rect 239253 699867 239311 699873
rect 259217 699907 259275 699913
rect 259217 699873 259229 699907
rect 259263 699904 259275 699907
rect 264093 699907 264151 699913
rect 264093 699904 264105 699907
rect 259263 699876 264105 699904
rect 259263 699873 259275 699876
rect 259217 699867 259275 699873
rect 264093 699873 264105 699876
rect 264139 699873 264151 699907
rect 278460 699904 278488 699944
rect 278537 699941 278549 699975
rect 278583 699972 278595 699975
rect 287369 699975 287427 699981
rect 287369 699972 287381 699975
rect 278583 699944 287381 699972
rect 278583 699941 278595 699944
rect 278537 699935 278595 699941
rect 287369 699941 287381 699944
rect 287415 699941 287427 699975
rect 287369 699935 287427 699941
rect 287458 699932 287464 699984
rect 287516 699972 287522 699984
rect 294545 699975 294603 699981
rect 294545 699972 294557 699975
rect 287516 699944 294557 699972
rect 287516 699932 287522 699944
rect 294545 699941 294557 699944
rect 294591 699941 294603 699975
rect 294545 699935 294603 699941
rect 294729 699975 294787 699981
rect 294729 699941 294741 699975
rect 294775 699972 294787 699975
rect 422238 699972 422244 699984
rect 294775 699944 422244 699972
rect 294775 699941 294787 699944
rect 294729 699935 294787 699941
rect 422238 699932 422244 699944
rect 422296 699932 422302 699984
rect 278629 699907 278687 699913
rect 278629 699904 278641 699907
rect 278460 699876 278641 699904
rect 264093 699867 264151 699873
rect 278629 699873 278641 699876
rect 278675 699873 278687 699907
rect 278629 699867 278687 699873
rect 283318 699864 283324 699916
rect 283376 699904 283382 699916
rect 290037 699907 290095 699913
rect 290037 699904 290049 699907
rect 283376 699876 290049 699904
rect 283376 699864 283382 699876
rect 290037 699873 290049 699876
rect 290083 699873 290095 699907
rect 294450 699904 294456 699916
rect 290037 699867 290095 699873
rect 290144 699876 294456 699904
rect 205946 699796 205952 699848
rect 206004 699836 206010 699848
rect 290144 699836 290172 699876
rect 294450 699864 294456 699876
rect 294508 699864 294514 699916
rect 296201 699907 296259 699913
rect 296201 699873 296213 699907
rect 296247 699904 296259 699907
rect 400618 699904 400624 699916
rect 296247 699876 400624 699904
rect 296247 699873 296259 699876
rect 296201 699867 296259 699873
rect 400618 699864 400624 699876
rect 400676 699864 400682 699916
rect 206004 699808 290172 699836
rect 206004 699796 206010 699808
rect 290218 699796 290224 699848
rect 290276 699836 290282 699848
rect 292518 699836 292524 699848
rect 290276 699808 292524 699836
rect 290276 699796 290282 699808
rect 292518 699796 292524 699808
rect 292576 699796 292582 699848
rect 292613 699839 292671 699845
rect 292613 699805 292625 699839
rect 292659 699836 292671 699839
rect 296109 699839 296167 699845
rect 292659 699808 296060 699836
rect 292659 699805 292671 699808
rect 292613 699799 292671 699805
rect 227566 699728 227572 699780
rect 227624 699768 227630 699780
rect 229593 699771 229651 699777
rect 229593 699768 229605 699771
rect 227624 699740 229605 699768
rect 227624 699728 227630 699740
rect 229593 699737 229605 699740
rect 229639 699737 229651 699771
rect 229593 699731 229651 699737
rect 287461 699771 287519 699777
rect 287461 699737 287473 699771
rect 287507 699768 287519 699771
rect 289025 699771 289083 699777
rect 287507 699740 288976 699768
rect 287507 699737 287519 699740
rect 287461 699731 287519 699737
rect 239253 699703 239311 699709
rect 239253 699669 239265 699703
rect 239299 699700 239311 699703
rect 259217 699703 259275 699709
rect 259217 699700 259229 699703
rect 239299 699672 259229 699700
rect 239299 699669 239311 699672
rect 239253 699663 239311 699669
rect 259217 699669 259229 699672
rect 259263 699669 259275 699703
rect 259217 699663 259275 699669
rect 264093 699703 264151 699709
rect 264093 699669 264105 699703
rect 264139 699700 264151 699703
rect 278537 699703 278595 699709
rect 278537 699700 278549 699703
rect 264139 699672 278549 699700
rect 264139 699669 264151 699672
rect 264093 699663 264151 699669
rect 278537 699669 278549 699672
rect 278583 699669 278595 699703
rect 278537 699663 278595 699669
rect 278629 699703 278687 699709
rect 278629 699669 278641 699703
rect 278675 699700 278687 699703
rect 288841 699703 288899 699709
rect 288841 699700 288853 699703
rect 278675 699672 288853 699700
rect 278675 699669 278687 699672
rect 278629 699663 278687 699669
rect 288841 699669 288853 699672
rect 288887 699669 288899 699703
rect 288948 699700 288976 699740
rect 289025 699737 289037 699771
rect 289071 699768 289083 699771
rect 291782 699768 291788 699780
rect 289071 699740 291788 699768
rect 289071 699737 289083 699740
rect 289025 699731 289083 699737
rect 291782 699728 291788 699740
rect 291840 699728 291846 699780
rect 291877 699771 291935 699777
rect 291877 699737 291889 699771
rect 291923 699768 291935 699771
rect 295922 699768 295928 699780
rect 291923 699740 295928 699768
rect 291923 699737 291935 699740
rect 291877 699731 291935 699737
rect 295922 699728 295928 699740
rect 295980 699728 295986 699780
rect 296032 699768 296060 699808
rect 296109 699805 296121 699839
rect 296155 699836 296167 699839
rect 335666 699836 335672 699848
rect 296155 699808 335672 699836
rect 296155 699805 296167 699808
rect 296109 699799 296167 699805
rect 335666 699796 335672 699808
rect 335724 699796 335730 699848
rect 297210 699768 297216 699780
rect 296032 699740 297216 699768
rect 297210 699728 297216 699740
rect 297268 699728 297274 699780
rect 291601 699703 291659 699709
rect 291601 699700 291613 699703
rect 288948 699672 291613 699700
rect 288841 699663 288899 699669
rect 291601 699669 291613 699672
rect 291647 699669 291659 699703
rect 291601 699663 291659 699669
rect 291690 699660 291696 699712
rect 291748 699700 291754 699712
rect 292426 699700 292432 699712
rect 291748 699672 292432 699700
rect 291748 699660 291754 699672
rect 292426 699660 292432 699672
rect 292484 699660 292490 699712
rect 292518 699660 292524 699712
rect 292576 699700 292582 699712
rect 357286 699700 357292 699712
rect 292576 699672 357292 699700
rect 292576 699660 292582 699672
rect 357286 699660 357292 699672
rect 357344 699660 357350 699712
rect 1600 699536 583316 699632
rect 1600 698992 583316 699088
rect 1600 698448 583316 698544
rect 1600 697904 583316 698000
rect 1600 697360 583316 697456
rect 1600 696816 583316 696912
rect 1600 696272 583316 696368
rect 1600 695728 583316 695824
rect 276418 695512 276424 695564
rect 276476 695552 276482 695564
rect 580110 695552 580116 695564
rect 276476 695524 580116 695552
rect 276476 695512 276482 695524
rect 580110 695512 580116 695524
rect 580168 695512 580174 695564
rect 378722 695484 378728 695496
rect 378683 695456 378728 695484
rect 378722 695444 378728 695456
rect 378780 695444 378786 695496
rect 508442 695484 508448 695496
rect 508403 695456 508448 695484
rect 508442 695444 508448 695456
rect 508500 695444 508506 695496
rect 1600 695184 583316 695280
rect 1600 694640 583316 694736
rect 3730 694220 3736 694272
rect 3788 694260 3794 694272
rect 305582 694260 305588 694272
rect 3788 694232 305588 694260
rect 3788 694220 3794 694232
rect 305582 694220 305588 694232
rect 305640 694220 305646 694272
rect 1600 694096 583316 694192
rect 1600 693552 583316 693648
rect 1600 693008 583316 693104
rect 1600 692464 583316 692560
rect 1600 691920 583316 692016
rect 1600 691376 583316 691472
rect 1600 690832 583316 690928
rect 1600 690288 583316 690384
rect 1600 689744 583316 689840
rect 1600 689200 583316 689296
rect 1600 688656 583316 688752
rect 314046 688576 314052 688628
rect 314104 688616 314110 688628
rect 314230 688616 314236 688628
rect 314104 688588 314236 688616
rect 314104 688576 314110 688588
rect 314230 688576 314236 688588
rect 314288 688576 314294 688628
rect 443766 688576 443772 688628
rect 443824 688616 443830 688628
rect 443950 688616 443956 688628
rect 443824 688588 443956 688616
rect 443824 688576 443830 688588
rect 443950 688576 443956 688588
rect 444008 688576 444014 688628
rect 573486 688576 573492 688628
rect 573544 688616 573550 688628
rect 573670 688616 573676 688628
rect 573544 688588 573676 688616
rect 573544 688576 573550 688588
rect 573670 688576 573676 688588
rect 573728 688576 573734 688628
rect 1600 688112 583316 688208
rect 1600 687568 583316 687664
rect 1600 687024 583316 687120
rect 1600 686480 583316 686576
rect 1600 685936 583316 686032
rect 378725 685899 378783 685905
rect 378725 685865 378737 685899
rect 378771 685896 378783 685899
rect 378814 685896 378820 685908
rect 378771 685868 378820 685896
rect 378771 685865 378783 685868
rect 378725 685859 378783 685865
rect 378814 685856 378820 685868
rect 378872 685856 378878 685908
rect 508445 685899 508503 685905
rect 508445 685865 508457 685899
rect 508491 685896 508503 685899
rect 508534 685896 508540 685908
rect 508491 685868 508540 685896
rect 508491 685865 508503 685868
rect 508445 685859 508503 685865
rect 508534 685856 508540 685868
rect 508592 685856 508598 685908
rect 1600 685392 583316 685488
rect 1600 684848 583316 684944
rect 1600 684304 583316 684400
rect 1600 683760 583316 683856
rect 1600 683216 583316 683312
rect 1600 682672 583316 682768
rect 1600 682128 583316 682224
rect 1600 681584 583316 681680
rect 1600 681040 583316 681136
rect 1600 680496 583316 680592
rect 277798 680348 277804 680400
rect 277856 680388 277862 680400
rect 580110 680388 580116 680400
rect 277856 680360 580116 680388
rect 277856 680348 277862 680360
rect 580110 680348 580116 680360
rect 580168 680348 580174 680400
rect 1600 679952 583316 680048
rect 1600 679408 583316 679504
rect 1600 678864 583316 678960
rect 1600 678320 583316 678416
rect 1600 677776 583316 677872
rect 3914 677560 3920 677612
rect 3972 677600 3978 677612
rect 308250 677600 308256 677612
rect 3972 677572 308256 677600
rect 3972 677560 3978 677572
rect 308250 677560 308256 677572
rect 308308 677560 308314 677612
rect 1600 677232 583316 677328
rect 1600 676688 583316 676784
rect 1600 676144 583316 676240
rect 314138 676104 314144 676116
rect 314099 676076 314144 676104
rect 314138 676064 314144 676076
rect 314196 676064 314202 676116
rect 378630 676104 378636 676116
rect 378591 676076 378636 676104
rect 378630 676064 378636 676076
rect 378688 676064 378694 676116
rect 443858 676104 443864 676116
rect 443819 676076 443864 676104
rect 443858 676064 443864 676076
rect 443916 676064 443922 676116
rect 508350 676104 508356 676116
rect 508311 676076 508356 676104
rect 508350 676064 508356 676076
rect 508408 676064 508414 676116
rect 573578 676104 573584 676116
rect 573539 676076 573584 676104
rect 573578 676064 573584 676076
rect 573636 676064 573642 676116
rect 1600 675600 583316 675696
rect 1600 675056 583316 675152
rect 1600 674512 583316 674608
rect 1600 673968 583316 674064
rect 1600 673424 583316 673520
rect 1600 672880 583316 672976
rect 1600 672336 583316 672432
rect 1600 671792 583316 671888
rect 1600 671248 583316 671344
rect 1600 670704 583316 670800
rect 1600 670160 583316 670256
rect 1600 669616 583316 669712
rect 1600 669072 583316 669168
rect 1600 668528 583316 668624
rect 1600 667984 583316 668080
rect 1600 667440 583316 667536
rect 1600 666896 583316 666992
rect 314141 666587 314199 666593
rect 314141 666553 314153 666587
rect 314187 666584 314199 666587
rect 314230 666584 314236 666596
rect 314187 666556 314236 666584
rect 314187 666553 314199 666556
rect 314141 666547 314199 666553
rect 314230 666544 314236 666556
rect 314288 666544 314294 666596
rect 378633 666587 378691 666593
rect 378633 666553 378645 666587
rect 378679 666584 378691 666587
rect 378722 666584 378728 666596
rect 378679 666556 378728 666584
rect 378679 666553 378691 666556
rect 378633 666547 378691 666553
rect 378722 666544 378728 666556
rect 378780 666544 378786 666596
rect 443861 666587 443919 666593
rect 443861 666553 443873 666587
rect 443907 666584 443919 666587
rect 443950 666584 443956 666596
rect 443907 666556 443956 666584
rect 443907 666553 443919 666556
rect 443861 666547 443919 666553
rect 443950 666544 443956 666556
rect 444008 666544 444014 666596
rect 508353 666587 508411 666593
rect 508353 666553 508365 666587
rect 508399 666584 508411 666587
rect 508442 666584 508448 666596
rect 508399 666556 508448 666584
rect 508399 666553 508411 666556
rect 508353 666547 508411 666553
rect 508442 666544 508448 666556
rect 508500 666544 508506 666596
rect 573581 666587 573639 666593
rect 573581 666553 573593 666587
rect 573627 666584 573639 666587
rect 573670 666584 573676 666596
rect 573627 666556 573676 666584
rect 573627 666553 573639 666556
rect 573581 666547 573639 666553
rect 573670 666544 573676 666556
rect 573728 666544 573734 666596
rect 1600 666352 583316 666448
rect 1600 665808 583316 665904
rect 1600 665264 583316 665360
rect 1600 664720 583316 664816
rect 1600 664176 583316 664272
rect 275038 663756 275044 663808
rect 275096 663796 275102 663808
rect 580110 663796 580116 663808
rect 275096 663768 580116 663796
rect 275096 663756 275102 663768
rect 580110 663756 580116 663768
rect 580168 663756 580174 663808
rect 1600 663632 583316 663728
rect 1600 663088 583316 663184
rect 1600 662544 583316 662640
rect 1600 662000 583316 662096
rect 1600 661456 583316 661552
rect 3914 661036 3920 661088
rect 3972 661076 3978 661088
rect 306870 661076 306876 661088
rect 3972 661048 306876 661076
rect 3972 661036 3978 661048
rect 306870 661036 306876 661048
rect 306928 661036 306934 661088
rect 1600 660912 583316 661008
rect 1600 660368 583316 660464
rect 1600 659824 583316 659920
rect 378722 659676 378728 659728
rect 378780 659716 378786 659728
rect 378814 659716 378820 659728
rect 378780 659688 378820 659716
rect 378780 659676 378786 659688
rect 378814 659676 378820 659688
rect 378872 659676 378878 659728
rect 508442 659676 508448 659728
rect 508500 659716 508506 659728
rect 508534 659716 508540 659728
rect 508500 659688 508540 659716
rect 508500 659676 508506 659688
rect 508534 659676 508540 659688
rect 508592 659676 508598 659728
rect 1600 659280 583316 659376
rect 1600 658736 583316 658832
rect 1600 658192 583316 658288
rect 1600 657648 583316 657744
rect 1600 657104 583316 657200
rect 1600 656560 583316 656656
rect 1600 656016 583316 656112
rect 1600 655472 583316 655568
rect 1600 654928 583316 655024
rect 1600 654384 583316 654480
rect 378630 654100 378636 654152
rect 378688 654140 378694 654152
rect 378814 654140 378820 654152
rect 378688 654112 378820 654140
rect 378688 654100 378694 654112
rect 378814 654100 378820 654112
rect 378872 654100 378878 654152
rect 508350 654100 508356 654152
rect 508408 654140 508414 654152
rect 508534 654140 508540 654152
rect 508408 654112 508540 654140
rect 508408 654100 508414 654112
rect 508534 654100 508540 654112
rect 508592 654100 508598 654152
rect 1600 653840 583316 653936
rect 1600 653296 583316 653392
rect 1600 652752 583316 652848
rect 1600 652208 583316 652304
rect 1600 651664 583316 651760
rect 1600 651120 583316 651216
rect 1600 650576 583316 650672
rect 1600 650032 583316 650128
rect 1600 649488 583316 649584
rect 1600 648944 583316 649040
rect 273658 648592 273664 648644
rect 273716 648632 273722 648644
rect 580110 648632 580116 648644
rect 273716 648604 580116 648632
rect 273716 648592 273722 648604
rect 580110 648592 580116 648604
rect 580168 648592 580174 648644
rect 1600 648400 583316 648496
rect 1600 647856 583316 647952
rect 1600 647312 583316 647408
rect 313954 647232 313960 647284
rect 314012 647272 314018 647284
rect 314046 647272 314052 647284
rect 314012 647244 314052 647272
rect 314012 647232 314018 647244
rect 314046 647232 314052 647244
rect 314104 647232 314110 647284
rect 443674 647232 443680 647284
rect 443732 647272 443738 647284
rect 443766 647272 443772 647284
rect 443732 647244 443772 647272
rect 443732 647232 443738 647244
rect 443766 647232 443772 647244
rect 443824 647232 443830 647284
rect 573394 647232 573400 647284
rect 573452 647272 573458 647284
rect 573486 647272 573492 647284
rect 573452 647244 573492 647272
rect 573452 647232 573458 647244
rect 573486 647232 573492 647244
rect 573544 647232 573550 647284
rect 1600 646768 583316 646864
rect 1600 646224 583316 646320
rect 1600 645680 583316 645776
rect 1600 645136 583316 645232
rect 1600 644592 583316 644688
rect 3546 644444 3552 644496
rect 3604 644484 3610 644496
rect 309630 644484 309636 644496
rect 3604 644456 309636 644484
rect 3604 644444 3610 644456
rect 309630 644444 309636 644456
rect 309688 644444 309694 644496
rect 1600 644048 583316 644144
rect 1600 643504 583316 643600
rect 1600 642960 583316 643056
rect 1600 642416 583316 642512
rect 1600 641872 583316 641968
rect 1600 641328 583316 641424
rect 1600 640784 583316 640880
rect 1600 640240 583316 640336
rect 1600 639696 583316 639792
rect 1600 639152 583316 639248
rect 1600 638608 583316 638704
rect 1600 638064 583316 638160
rect 1600 637520 583316 637616
rect 314138 637480 314144 637492
rect 314099 637452 314144 637480
rect 314138 637440 314144 637452
rect 314196 637440 314202 637492
rect 443858 637480 443864 637492
rect 443819 637452 443864 637480
rect 443858 637440 443864 637452
rect 443916 637440 443922 637492
rect 573578 637480 573584 637492
rect 573539 637452 573584 637480
rect 573578 637440 573584 637452
rect 573636 637440 573642 637492
rect 1600 636976 583316 637072
rect 1600 636432 583316 636528
rect 1600 635888 583316 635984
rect 1600 635344 583316 635440
rect 1600 634800 583316 634896
rect 1600 634256 583316 634352
rect 1600 633712 583316 633808
rect 274946 633428 274952 633480
rect 275004 633468 275010 633480
rect 580110 633468 580116 633480
rect 275004 633440 580116 633468
rect 275004 633428 275010 633440
rect 580110 633428 580116 633440
rect 580168 633428 580174 633480
rect 1600 633168 583316 633264
rect 1600 632624 583316 632720
rect 1600 632080 583316 632176
rect 1600 631536 583316 631632
rect 1600 630992 583316 631088
rect 1600 630448 583316 630544
rect 1600 629904 583316 630000
rect 1600 629360 583316 629456
rect 1600 628816 583316 628912
rect 1600 628272 583316 628368
rect 3914 627920 3920 627972
rect 3972 627960 3978 627972
rect 311010 627960 311016 627972
rect 3972 627932 311016 627960
rect 3972 627920 3978 627932
rect 311010 627920 311016 627932
rect 311068 627920 311074 627972
rect 314141 627963 314199 627969
rect 314141 627929 314153 627963
rect 314187 627960 314199 627963
rect 314230 627960 314236 627972
rect 314187 627932 314236 627960
rect 314187 627929 314199 627932
rect 314141 627923 314199 627929
rect 314230 627920 314236 627932
rect 314288 627920 314294 627972
rect 443861 627963 443919 627969
rect 443861 627929 443873 627963
rect 443907 627960 443919 627963
rect 443950 627960 443956 627972
rect 443907 627932 443956 627960
rect 443907 627929 443919 627932
rect 443861 627923 443919 627929
rect 443950 627920 443956 627932
rect 444008 627920 444014 627972
rect 573581 627963 573639 627969
rect 573581 627929 573593 627963
rect 573627 627960 573639 627963
rect 573670 627960 573676 627972
rect 573627 627932 573676 627960
rect 573627 627929 573639 627932
rect 573581 627923 573639 627929
rect 573670 627920 573676 627932
rect 573728 627920 573734 627972
rect 1600 627728 583316 627824
rect 1600 627184 583316 627280
rect 1600 626640 583316 626736
rect 1600 626096 583316 626192
rect 1600 625552 583316 625648
rect 1600 625008 583316 625104
rect 1600 624464 583316 624560
rect 1600 623920 583316 624016
rect 1600 623376 583316 623472
rect 1600 622832 583316 622928
rect 1600 622288 583316 622384
rect 1600 621744 583316 621840
rect 1600 621200 583316 621296
rect 1600 620656 583316 620752
rect 1600 620112 583316 620208
rect 1600 619568 583316 619664
rect 1600 619024 583316 619120
rect 1600 618480 583316 618576
rect 314046 618264 314052 618316
rect 314104 618304 314110 618316
rect 314230 618304 314236 618316
rect 314104 618276 314236 618304
rect 314104 618264 314110 618276
rect 314230 618264 314236 618276
rect 314288 618264 314294 618316
rect 443766 618264 443772 618316
rect 443824 618304 443830 618316
rect 443950 618304 443956 618316
rect 443824 618276 443956 618304
rect 443824 618264 443830 618276
rect 443950 618264 443956 618276
rect 444008 618264 444014 618316
rect 573486 618264 573492 618316
rect 573544 618304 573550 618316
rect 573670 618304 573676 618316
rect 573544 618276 573676 618304
rect 573544 618264 573550 618276
rect 573670 618264 573676 618276
rect 573728 618264 573734 618316
rect 573486 618128 573492 618180
rect 573544 618168 573550 618180
rect 573762 618168 573768 618180
rect 573544 618140 573768 618168
rect 573544 618128 573550 618140
rect 573762 618128 573768 618140
rect 573820 618128 573826 618180
rect 1600 617936 583316 618032
rect 1600 617392 583316 617488
rect 272278 616972 272284 617024
rect 272336 617012 272342 617024
rect 580110 617012 580116 617024
rect 272336 616984 580116 617012
rect 272336 616972 272342 616984
rect 580110 616972 580116 616984
rect 580168 616972 580174 617024
rect 1600 616848 583316 616944
rect 1600 616304 583316 616400
rect 1600 615760 583316 615856
rect 378630 615476 378636 615528
rect 378688 615516 378694 615528
rect 378814 615516 378820 615528
rect 378688 615488 378820 615516
rect 378688 615476 378694 615488
rect 378814 615476 378820 615488
rect 378872 615476 378878 615528
rect 508350 615476 508356 615528
rect 508408 615516 508414 615528
rect 508534 615516 508540 615528
rect 508408 615488 508540 615516
rect 508408 615476 508414 615488
rect 508534 615476 508540 615488
rect 508592 615476 508598 615528
rect 1600 615216 583316 615312
rect 1600 614672 583316 614768
rect 1600 614128 583316 614224
rect 1600 613584 583316 613680
rect 1600 613040 583316 613136
rect 1600 612496 583316 612592
rect 1600 611952 583316 612048
rect 1600 611408 583316 611504
rect 3822 611328 3828 611380
rect 3880 611368 3886 611380
rect 309722 611368 309728 611380
rect 3880 611340 309728 611368
rect 3880 611328 3886 611340
rect 309722 611328 309728 611340
rect 309780 611328 309786 611380
rect 1600 610864 583316 610960
rect 1600 610320 583316 610416
rect 1600 609776 583316 609872
rect 1600 609232 583316 609328
rect 1600 608688 583316 608784
rect 313770 608608 313776 608660
rect 313828 608648 313834 608660
rect 313954 608648 313960 608660
rect 313828 608620 313960 608648
rect 313828 608608 313834 608620
rect 313954 608608 313960 608620
rect 314012 608608 314018 608660
rect 443674 608580 443680 608592
rect 443635 608552 443680 608580
rect 443674 608540 443680 608552
rect 443732 608540 443738 608592
rect 573394 608580 573400 608592
rect 573355 608552 573400 608580
rect 573394 608540 573400 608552
rect 573452 608540 573458 608592
rect 1600 608144 583316 608240
rect 1600 607600 583316 607696
rect 1600 607056 583316 607152
rect 1600 606512 583316 606608
rect 1600 605968 583316 606064
rect 1600 605424 583316 605520
rect 1600 604880 583316 604976
rect 1600 604336 583316 604432
rect 1600 603792 583316 603888
rect 1600 603248 583316 603344
rect 1600 602704 583316 602800
rect 1600 602160 583316 602256
rect 270898 601740 270904 601792
rect 270956 601780 270962 601792
rect 580110 601780 580116 601792
rect 270956 601752 580116 601780
rect 270956 601740 270962 601752
rect 580110 601740 580116 601752
rect 580168 601740 580174 601792
rect 1600 601616 583316 601712
rect 443677 601579 443735 601585
rect 443677 601545 443689 601579
rect 443723 601576 443735 601579
rect 443858 601576 443864 601588
rect 443723 601548 443864 601576
rect 443723 601545 443735 601548
rect 443677 601539 443735 601545
rect 443858 601536 443864 601548
rect 443916 601536 443922 601588
rect 573397 601579 573455 601585
rect 573397 601545 573409 601579
rect 573443 601576 573455 601579
rect 573578 601576 573584 601588
rect 573443 601548 573584 601576
rect 573443 601545 573455 601548
rect 573397 601539 573455 601545
rect 573578 601536 573584 601548
rect 573636 601536 573642 601588
rect 1600 601072 583316 601168
rect 1600 600528 583316 600624
rect 1600 599984 583316 600080
rect 1600 599440 583316 599536
rect 1600 598896 583316 598992
rect 313862 598856 313868 598868
rect 313823 598828 313868 598856
rect 313862 598816 313868 598828
rect 313920 598816 313926 598868
rect 443858 598856 443864 598868
rect 443819 598828 443864 598856
rect 443858 598816 443864 598828
rect 443916 598816 443922 598868
rect 573578 598856 573584 598868
rect 573539 598828 573584 598856
rect 573578 598816 573584 598828
rect 573636 598816 573642 598868
rect 1600 598352 583316 598448
rect 1600 597808 583316 597904
rect 1600 597264 583316 597360
rect 1600 596720 583316 596816
rect 1600 596176 583316 596272
rect 1600 595632 583316 595728
rect 1600 595088 583316 595184
rect 3914 594804 3920 594856
rect 3972 594844 3978 594856
rect 312390 594844 312396 594856
rect 3972 594816 312396 594844
rect 3972 594804 3978 594816
rect 312390 594804 312396 594816
rect 312448 594804 312454 594856
rect 1600 594544 583316 594640
rect 1600 594000 583316 594096
rect 1600 593456 583316 593552
rect 1600 592912 583316 593008
rect 1600 592368 583316 592464
rect 1600 591824 583316 591920
rect 1600 591280 583316 591376
rect 1600 590736 583316 590832
rect 1600 590192 583316 590288
rect 1600 589648 583316 589744
rect 313865 589339 313923 589345
rect 313865 589305 313877 589339
rect 313911 589336 313923 589339
rect 314046 589336 314052 589348
rect 313911 589308 314052 589336
rect 313911 589305 313923 589308
rect 313865 589299 313923 589305
rect 314046 589296 314052 589308
rect 314104 589296 314110 589348
rect 443861 589339 443919 589345
rect 443861 589305 443873 589339
rect 443907 589336 443919 589339
rect 443950 589336 443956 589348
rect 443907 589308 443956 589336
rect 443907 589305 443919 589308
rect 443861 589299 443919 589305
rect 443950 589296 443956 589308
rect 444008 589296 444014 589348
rect 573581 589339 573639 589345
rect 573581 589305 573593 589339
rect 573627 589336 573639 589339
rect 573670 589336 573676 589348
rect 573627 589308 573676 589336
rect 573627 589305 573639 589308
rect 573581 589299 573639 589305
rect 573670 589296 573676 589308
rect 573728 589296 573734 589348
rect 378633 589271 378691 589277
rect 378633 589237 378645 589271
rect 378679 589268 378691 589271
rect 378722 589268 378728 589280
rect 378679 589240 378728 589268
rect 378679 589237 378691 589240
rect 378633 589231 378691 589237
rect 378722 589228 378728 589240
rect 378780 589228 378786 589280
rect 508353 589271 508411 589277
rect 508353 589237 508365 589271
rect 508399 589268 508411 589271
rect 508442 589268 508448 589280
rect 508399 589240 508448 589268
rect 508399 589237 508411 589240
rect 508353 589231 508411 589237
rect 508442 589228 508448 589240
rect 508500 589228 508506 589280
rect 1600 589104 583316 589200
rect 1600 588560 583316 588656
rect 1600 588016 583316 588112
rect 1600 587472 583316 587568
rect 1600 586928 583316 587024
rect 270806 586508 270812 586560
rect 270864 586548 270870 586560
rect 580110 586548 580116 586560
rect 270864 586520 580116 586548
rect 270864 586508 270870 586520
rect 580110 586508 580116 586520
rect 580168 586508 580174 586560
rect 1600 586384 583316 586480
rect 1600 585840 583316 585936
rect 1600 585296 583316 585392
rect 1600 584752 583316 584848
rect 1600 584208 583316 584304
rect 1600 583664 583316 583760
rect 1600 583120 583316 583216
rect 1600 582576 583316 582672
rect 443950 582468 443956 582480
rect 443876 582440 443956 582468
rect 314046 582360 314052 582412
rect 314104 582360 314110 582412
rect 314064 582332 314092 582360
rect 443876 582344 443904 582440
rect 443950 582428 443956 582440
rect 444008 582428 444014 582480
rect 573670 582468 573676 582480
rect 573596 582440 573676 582468
rect 573596 582344 573624 582440
rect 573670 582428 573676 582440
rect 573728 582428 573734 582480
rect 314138 582332 314144 582344
rect 314064 582304 314144 582332
rect 314138 582292 314144 582304
rect 314196 582292 314202 582344
rect 443858 582292 443864 582344
rect 443916 582292 443922 582344
rect 573578 582292 573584 582344
rect 573636 582292 573642 582344
rect 1600 582032 583316 582128
rect 1600 581488 583316 581584
rect 1600 580944 583316 581040
rect 1600 580400 583316 580496
rect 1600 579856 583316 579952
rect 378630 579680 378636 579692
rect 378591 579652 378636 579680
rect 378630 579640 378636 579652
rect 378688 579640 378694 579692
rect 508350 579680 508356 579692
rect 508311 579652 508356 579680
rect 508350 579640 508356 579652
rect 508408 579640 508414 579692
rect 313957 579615 314015 579621
rect 313957 579581 313969 579615
rect 314003 579612 314015 579615
rect 314138 579612 314144 579624
rect 314003 579584 314144 579612
rect 314003 579581 314015 579584
rect 313957 579575 314015 579581
rect 314138 579572 314144 579584
rect 314196 579572 314202 579624
rect 1600 579312 583316 579408
rect 1600 578768 583316 578864
rect 1600 578224 583316 578320
rect 1600 577680 583316 577776
rect 1600 577136 583316 577232
rect 3730 576852 3736 576904
rect 3788 576892 3794 576904
rect 313862 576892 313868 576904
rect 3788 576864 313868 576892
rect 3788 576852 3794 576864
rect 313862 576852 313868 576864
rect 313920 576852 313926 576904
rect 1600 576592 583316 576688
rect 1600 576048 583316 576144
rect 1600 575504 583316 575600
rect 1600 574960 583316 575056
rect 1600 574416 583316 574512
rect 1600 573872 583316 573968
rect 1600 573328 583316 573424
rect 1600 572784 583316 572880
rect 1600 572240 583316 572336
rect 1600 571696 583316 571792
rect 1600 571152 583316 571248
rect 1600 570608 583316 570704
rect 1600 570064 583316 570160
rect 313954 570024 313960 570036
rect 313915 569996 313960 570024
rect 313954 569984 313960 569996
rect 314012 569984 314018 570036
rect 269518 569916 269524 569968
rect 269576 569956 269582 569968
rect 580110 569956 580116 569968
rect 269576 569928 580116 569956
rect 269576 569916 269582 569928
rect 580110 569916 580116 569928
rect 580168 569916 580174 569968
rect 378722 569888 378728 569900
rect 378683 569860 378728 569888
rect 378722 569848 378728 569860
rect 378780 569848 378786 569900
rect 508442 569888 508448 569900
rect 508403 569860 508448 569888
rect 508442 569848 508448 569860
rect 508500 569848 508506 569900
rect 1600 569520 583316 569616
rect 1600 568976 583316 569072
rect 1600 568432 583316 568528
rect 1600 567888 583316 567984
rect 1600 567344 583316 567440
rect 1600 566800 583316 566896
rect 1600 566256 583316 566352
rect 1600 565712 583316 565808
rect 1600 565168 583316 565264
rect 1600 564624 583316 564720
rect 1600 564080 583316 564176
rect 1600 563536 583316 563632
rect 1600 562992 583316 563088
rect 378725 562955 378783 562961
rect 378725 562921 378737 562955
rect 378771 562952 378783 562955
rect 378906 562952 378912 562964
rect 378771 562924 378912 562952
rect 378771 562921 378783 562924
rect 378725 562915 378783 562921
rect 378906 562912 378912 562924
rect 378964 562912 378970 562964
rect 508445 562955 508503 562961
rect 508445 562921 508457 562955
rect 508491 562952 508503 562955
rect 508626 562952 508632 562964
rect 508491 562924 508632 562952
rect 508491 562921 508503 562924
rect 508445 562915 508503 562921
rect 508626 562912 508632 562924
rect 508684 562912 508690 562964
rect 1600 562448 583316 562544
rect 1600 561904 583316 562000
rect 1600 561360 583316 561456
rect 1600 560816 583316 560912
rect 3914 560396 3920 560448
rect 3972 560436 3978 560448
rect 313954 560436 313960 560448
rect 3972 560408 313960 560436
rect 3972 560396 3978 560408
rect 313954 560396 313960 560408
rect 314012 560396 314018 560448
rect 1600 560272 583316 560368
rect 1600 559728 583316 559824
rect 1600 559184 583316 559280
rect 1600 558640 583316 558736
rect 1600 558096 583316 558192
rect 1600 557552 583316 557648
rect 1600 557008 583316 557104
rect 1600 556464 583316 556560
rect 1600 555920 583316 556016
rect 1600 555376 583316 555472
rect 1600 554832 583316 554928
rect 266758 554752 266764 554804
rect 266816 554792 266822 554804
rect 580110 554792 580116 554804
rect 266816 554764 580116 554792
rect 266816 554752 266822 554764
rect 580110 554752 580116 554764
rect 580168 554752 580174 554804
rect 1600 554288 583316 554384
rect 1600 553744 583316 553840
rect 443490 553432 443496 553444
rect 443451 553404 443496 553432
rect 443490 553392 443496 553404
rect 443548 553392 443554 553444
rect 573210 553432 573216 553444
rect 573171 553404 573216 553432
rect 573210 553392 573216 553404
rect 573268 553392 573274 553444
rect 1600 553200 583316 553296
rect 1600 552656 583316 552752
rect 313770 552576 313776 552628
rect 313828 552616 313834 552628
rect 314046 552616 314052 552628
rect 313828 552588 314052 552616
rect 313828 552576 313834 552588
rect 314046 552576 314052 552588
rect 314104 552576 314110 552628
rect 1600 552112 583316 552208
rect 1600 551568 583316 551664
rect 1600 551024 583316 551120
rect 378722 550604 378728 550656
rect 378780 550644 378786 550656
rect 378998 550644 379004 550656
rect 378780 550616 379004 550644
rect 378780 550604 378786 550616
rect 378998 550604 379004 550616
rect 379056 550604 379062 550656
rect 443490 550644 443496 550656
rect 443451 550616 443496 550644
rect 443490 550604 443496 550616
rect 443548 550604 443554 550656
rect 508442 550604 508448 550656
rect 508500 550644 508506 550656
rect 508718 550644 508724 550656
rect 508500 550616 508724 550644
rect 508500 550604 508506 550616
rect 508718 550604 508724 550616
rect 508776 550604 508782 550656
rect 573210 550644 573216 550656
rect 573171 550616 573216 550644
rect 573210 550604 573216 550616
rect 573268 550604 573274 550656
rect 1600 550480 583316 550576
rect 1600 549936 583316 550032
rect 1600 549392 583316 549488
rect 1600 548848 583316 548944
rect 1600 548304 583316 548400
rect 1600 547760 583316 547856
rect 1600 547216 583316 547312
rect 1600 546672 583316 546768
rect 1600 546128 583316 546224
rect 1600 545584 583316 545680
rect 1600 545040 583316 545136
rect 1600 544496 583316 544592
rect 1600 543952 583316 544048
rect 378998 543844 379004 543856
rect 378924 543816 379004 543844
rect 3638 543736 3644 543788
rect 3696 543776 3702 543788
rect 315150 543776 315156 543788
rect 3696 543748 315156 543776
rect 3696 543736 3702 543748
rect 315150 543736 315156 543748
rect 315208 543736 315214 543788
rect 378924 543720 378952 543816
rect 378998 543804 379004 543816
rect 379056 543804 379062 543856
rect 508718 543844 508724 543856
rect 508644 543816 508724 543844
rect 443490 543736 443496 543788
rect 443548 543736 443554 543788
rect 378906 543668 378912 543720
rect 378964 543668 378970 543720
rect 443508 543640 443536 543736
rect 508644 543720 508672 543816
rect 508718 543804 508724 543816
rect 508776 543804 508782 543856
rect 573210 543736 573216 543788
rect 573268 543736 573274 543788
rect 508626 543668 508632 543720
rect 508684 543668 508690 543720
rect 443582 543640 443588 543652
rect 443508 543612 443588 543640
rect 443582 543600 443588 543612
rect 443640 543600 443646 543652
rect 573228 543640 573256 543736
rect 573302 543640 573308 543652
rect 573228 543612 573308 543640
rect 573302 543600 573308 543612
rect 573360 543600 573366 543652
rect 1600 543408 583316 543504
rect 1600 542864 583316 542960
rect 1600 542320 583316 542416
rect 1600 541776 583316 541872
rect 1600 541232 583316 541328
rect 1600 540688 583316 540784
rect 1600 540144 583316 540240
rect 268138 539724 268144 539776
rect 268196 539764 268202 539776
rect 580110 539764 580116 539776
rect 268196 539736 580116 539764
rect 268196 539724 268202 539736
rect 580110 539724 580116 539736
rect 580168 539724 580174 539776
rect 1600 539600 583316 539696
rect 1600 539056 583316 539152
rect 1600 538512 583316 538608
rect 313770 538228 313776 538280
rect 313828 538268 313834 538280
rect 314046 538268 314052 538280
rect 313828 538240 314052 538268
rect 313828 538228 313834 538240
rect 314046 538228 314052 538240
rect 314104 538228 314110 538280
rect 1600 537968 583316 538064
rect 1600 537424 583316 537520
rect 1600 536880 583316 536976
rect 1600 536336 583316 536432
rect 1600 535792 583316 535888
rect 1600 535248 583316 535344
rect 1600 534704 583316 534800
rect 1600 534160 583316 534256
rect 378906 534080 378912 534132
rect 378964 534080 378970 534132
rect 443490 534120 443496 534132
rect 443451 534092 443496 534120
rect 443490 534080 443496 534092
rect 443548 534080 443554 534132
rect 508626 534080 508632 534132
rect 508684 534080 508690 534132
rect 573210 534120 573216 534132
rect 573171 534092 573216 534120
rect 573210 534080 573216 534092
rect 573268 534080 573274 534132
rect 378924 533984 378952 534080
rect 378998 533984 379004 533996
rect 378924 533956 379004 533984
rect 378998 533944 379004 533956
rect 379056 533944 379062 533996
rect 508644 533984 508672 534080
rect 508718 533984 508724 533996
rect 508644 533956 508724 533984
rect 508718 533944 508724 533956
rect 508776 533944 508782 533996
rect 1600 533616 583316 533712
rect 1600 533072 583316 533168
rect 1600 532528 583316 532624
rect 1600 531984 583316 532080
rect 1600 531440 583316 531536
rect 443490 531332 443496 531344
rect 443451 531304 443496 531332
rect 443490 531292 443496 531304
rect 443548 531292 443554 531344
rect 573210 531332 573216 531344
rect 573171 531304 573216 531332
rect 573210 531292 573216 531304
rect 573268 531292 573274 531344
rect 443582 531264 443588 531276
rect 443543 531236 443588 531264
rect 443582 531224 443588 531236
rect 443640 531224 443646 531276
rect 573302 531264 573308 531276
rect 573263 531236 573308 531264
rect 573302 531224 573308 531236
rect 573360 531224 573366 531276
rect 1600 530896 583316 530992
rect 1600 530352 583316 530448
rect 1600 529808 583316 529904
rect 1600 529264 583316 529360
rect 1600 528720 583316 528816
rect 313770 528504 313776 528556
rect 313828 528544 313834 528556
rect 314046 528544 314052 528556
rect 313828 528516 314052 528544
rect 313828 528504 313834 528516
rect 314046 528504 314052 528516
rect 314104 528504 314110 528556
rect 1600 528176 583316 528272
rect 1600 527632 583316 527728
rect 3638 527212 3644 527264
rect 3696 527252 3702 527264
rect 317910 527252 317916 527264
rect 3696 527224 317916 527252
rect 3696 527212 3702 527224
rect 317910 527212 317916 527224
rect 317968 527212 317974 527264
rect 1600 527088 583316 527184
rect 1600 526544 583316 526640
rect 1600 526000 583316 526096
rect 1600 525456 583316 525552
rect 1600 524912 583316 525008
rect 1600 524368 583316 524464
rect 443582 524328 443588 524340
rect 443543 524300 443588 524328
rect 443582 524288 443588 524300
rect 443640 524288 443646 524340
rect 573302 524328 573308 524340
rect 573263 524300 573308 524328
rect 573302 524288 573308 524300
rect 573360 524288 573366 524340
rect 1600 523824 583316 523920
rect 1600 523280 583316 523376
rect 266666 522996 266672 523048
rect 266724 523036 266730 523048
rect 580110 523036 580116 523048
rect 266724 523008 580116 523036
rect 266724 522996 266730 523008
rect 580110 522996 580116 523008
rect 580168 522996 580174 523048
rect 1600 522736 583316 522832
rect 1600 522192 583316 522288
rect 1600 521648 583316 521744
rect 1600 521104 583316 521200
rect 1600 520560 583316 520656
rect 1600 520016 583316 520112
rect 1600 519472 583316 519568
rect 1600 518928 583316 519024
rect 1600 518384 583316 518480
rect 1600 517840 583316 517936
rect 1600 517296 583316 517392
rect 1600 516752 583316 516848
rect 1600 516208 583316 516304
rect 1600 515664 583316 515760
rect 1600 515120 583316 515216
rect 1600 514576 583316 514672
rect 378998 514496 379004 514548
rect 379056 514536 379062 514548
rect 379182 514536 379188 514548
rect 379056 514508 379188 514536
rect 379056 514496 379062 514508
rect 379182 514496 379188 514508
rect 379240 514496 379246 514548
rect 508718 514496 508724 514548
rect 508776 514536 508782 514548
rect 508902 514536 508908 514548
rect 508776 514508 508908 514536
rect 508776 514496 508782 514508
rect 508902 514496 508908 514508
rect 508960 514496 508966 514548
rect 1600 514032 583316 514128
rect 313770 513952 313776 514004
rect 313828 513992 313834 514004
rect 314046 513992 314052 514004
rect 313828 513964 314052 513992
rect 313828 513952 313834 513964
rect 314046 513952 314052 513964
rect 314104 513952 314110 514004
rect 1600 513488 583316 513584
rect 1600 512944 583316 513040
rect 1600 512400 583316 512496
rect 1600 511856 583316 511952
rect 1600 511312 583316 511408
rect 1600 510768 583316 510864
rect 4006 510620 4012 510672
rect 4064 510660 4070 510672
rect 316530 510660 316536 510672
rect 4064 510632 316536 510660
rect 4064 510620 4070 510632
rect 316530 510620 316536 510632
rect 316588 510620 316594 510672
rect 1600 510224 583316 510320
rect 1600 509680 583316 509776
rect 1600 509136 583316 509232
rect 1600 508592 583316 508688
rect 1600 508048 583316 508144
rect 263998 507832 264004 507884
rect 264056 507872 264062 507884
rect 580110 507872 580116 507884
rect 264056 507844 580116 507872
rect 264056 507832 264062 507844
rect 580110 507832 580116 507844
rect 580168 507832 580174 507884
rect 1600 507504 583316 507600
rect 1600 506960 583316 507056
rect 1600 506416 583316 506512
rect 1600 505872 583316 505968
rect 1600 505328 583316 505424
rect 1600 504784 583316 504880
rect 1600 504240 583316 504336
rect 1600 503696 583316 503792
rect 1600 503152 583316 503248
rect 1600 502608 583316 502704
rect 378814 502324 378820 502376
rect 378872 502364 378878 502376
rect 378998 502364 379004 502376
rect 378872 502336 379004 502364
rect 378872 502324 378878 502336
rect 378998 502324 379004 502336
rect 379056 502324 379062 502376
rect 443490 502324 443496 502376
rect 443548 502364 443554 502376
rect 443766 502364 443772 502376
rect 443548 502336 443772 502364
rect 443548 502324 443554 502336
rect 443766 502324 443772 502336
rect 443824 502324 443830 502376
rect 508534 502324 508540 502376
rect 508592 502364 508598 502376
rect 508718 502364 508724 502376
rect 508592 502336 508724 502364
rect 508592 502324 508598 502336
rect 508718 502324 508724 502336
rect 508776 502324 508782 502376
rect 573210 502324 573216 502376
rect 573268 502364 573274 502376
rect 573486 502364 573492 502376
rect 573268 502336 573492 502364
rect 573268 502324 573274 502336
rect 573486 502324 573492 502336
rect 573544 502324 573550 502376
rect 1600 502064 583316 502160
rect 1600 501520 583316 501616
rect 1600 500976 583316 501072
rect 1600 500432 583316 500528
rect 1600 499888 583316 499984
rect 313770 499536 313776 499588
rect 313828 499576 313834 499588
rect 314046 499576 314052 499588
rect 313828 499548 314052 499576
rect 313828 499536 313834 499548
rect 314046 499536 314052 499548
rect 314104 499536 314110 499588
rect 1600 499344 583316 499440
rect 1600 498800 583316 498896
rect 1600 498256 583316 498352
rect 1600 497712 583316 497808
rect 1600 497168 583316 497264
rect 1600 496624 583316 496720
rect 1600 496080 583316 496176
rect 1600 495536 583316 495632
rect 1600 494992 583316 495088
rect 1600 494448 583316 494544
rect 3730 494028 3736 494080
rect 3788 494068 3794 494080
rect 318002 494068 318008 494080
rect 3788 494040 318008 494068
rect 3788 494028 3794 494040
rect 318002 494028 318008 494040
rect 318060 494028 318066 494080
rect 1600 493904 583316 494000
rect 1600 493360 583316 493456
rect 1600 492816 583316 492912
rect 265378 492668 265384 492720
rect 265436 492708 265442 492720
rect 580110 492708 580116 492720
rect 265436 492680 580116 492708
rect 265436 492668 265442 492680
rect 580110 492668 580116 492680
rect 580168 492668 580174 492720
rect 1600 492272 583316 492368
rect 1600 491728 583316 491824
rect 1600 491184 583316 491280
rect 1600 490640 583316 490736
rect 1600 490096 583316 490192
rect 313770 489812 313776 489864
rect 313828 489852 313834 489864
rect 314046 489852 314052 489864
rect 313828 489824 314052 489852
rect 313828 489812 313834 489824
rect 314046 489812 314052 489824
rect 314104 489812 314110 489864
rect 1600 489552 583316 489648
rect 1600 489008 583316 489104
rect 1600 488464 583316 488560
rect 1600 487920 583316 488016
rect 1600 487376 583316 487472
rect 1600 486832 583316 486928
rect 1600 486288 583316 486384
rect 443493 485911 443551 485917
rect 443493 485877 443505 485911
rect 443539 485908 443551 485911
rect 443766 485908 443772 485920
rect 443539 485880 443772 485908
rect 443539 485877 443551 485880
rect 443493 485871 443551 485877
rect 443766 485868 443772 485880
rect 443824 485868 443830 485920
rect 573213 485911 573271 485917
rect 573213 485877 573225 485911
rect 573259 485908 573271 485911
rect 573486 485908 573492 485920
rect 573259 485880 573492 485908
rect 573259 485877 573271 485880
rect 573213 485871 573271 485877
rect 573486 485868 573492 485880
rect 573544 485868 573550 485920
rect 1600 485744 583316 485840
rect 443490 485704 443496 485716
rect 443451 485676 443496 485704
rect 443490 485664 443496 485676
rect 443548 485664 443554 485716
rect 573210 485704 573216 485716
rect 573171 485676 573216 485704
rect 573210 485664 573216 485676
rect 573268 485664 573274 485716
rect 1600 485200 583316 485296
rect 1600 484656 583316 484752
rect 1600 484112 583316 484208
rect 1600 483568 583316 483664
rect 1600 483024 583316 483120
rect 1600 482480 583316 482576
rect 1600 481936 583316 482032
rect 1600 481392 583316 481488
rect 1600 480848 583316 480944
rect 1600 480304 583316 480400
rect 313770 480224 313776 480276
rect 313828 480264 313834 480276
rect 314046 480264 314052 480276
rect 313828 480236 314052 480264
rect 313828 480224 313834 480236
rect 314046 480224 314052 480236
rect 314104 480224 314110 480276
rect 378630 480224 378636 480276
rect 378688 480264 378694 480276
rect 378814 480264 378820 480276
rect 378688 480236 378820 480264
rect 378688 480224 378694 480236
rect 378814 480224 378820 480236
rect 378872 480224 378878 480276
rect 508350 480224 508356 480276
rect 508408 480264 508414 480276
rect 508534 480264 508540 480276
rect 508408 480236 508540 480264
rect 508408 480224 508414 480236
rect 508534 480224 508540 480236
rect 508592 480224 508598 480276
rect 1600 479760 583316 479856
rect 1600 479216 583316 479312
rect 1600 478672 583316 478768
rect 1600 478128 583316 478224
rect 1600 477584 583316 477680
rect 3914 477504 3920 477556
rect 3972 477544 3978 477556
rect 320670 477544 320676 477556
rect 3972 477516 320676 477544
rect 3972 477504 3978 477516
rect 320670 477504 320676 477516
rect 320728 477504 320734 477556
rect 1600 477040 583316 477136
rect 1600 476496 583316 476592
rect 262618 476076 262624 476128
rect 262676 476116 262682 476128
rect 580110 476116 580116 476128
rect 262676 476088 580116 476116
rect 262676 476076 262682 476088
rect 580110 476076 580116 476088
rect 580168 476076 580174 476128
rect 1600 475952 583316 476048
rect 1600 475408 583316 475504
rect 313770 475328 313776 475380
rect 313828 475368 313834 475380
rect 314046 475368 314052 475380
rect 313828 475340 314052 475368
rect 313828 475328 313834 475340
rect 314046 475328 314052 475340
rect 314104 475328 314110 475380
rect 1600 474864 583316 474960
rect 1600 474320 583316 474416
rect 1600 473776 583316 473872
rect 1600 473232 583316 473328
rect 1600 472688 583316 472784
rect 1600 472144 583316 472240
rect 443582 471968 443588 471980
rect 443543 471940 443588 471968
rect 443582 471928 443588 471940
rect 443640 471928 443646 471980
rect 573302 471968 573308 471980
rect 573263 471940 573308 471968
rect 573302 471928 573308 471940
rect 573360 471928 573366 471980
rect 1600 471600 583316 471696
rect 1600 471056 583316 471152
rect 1600 470512 583316 470608
rect 1600 469968 583316 470064
rect 1600 469424 583316 469520
rect 1600 468880 583316 468976
rect 1600 468336 583316 468432
rect 1600 467792 583316 467888
rect 1600 467248 583316 467344
rect 1600 466704 583316 466800
rect 1600 466160 583316 466256
rect 1600 465616 583316 465712
rect 1600 465072 583316 465168
rect 1600 464528 583316 464624
rect 1600 463984 583316 464080
rect 302917 463743 302975 463749
rect 302917 463709 302929 463743
rect 302963 463740 302975 463743
rect 314046 463740 314052 463752
rect 302963 463712 314052 463740
rect 302963 463709 302975 463712
rect 302917 463703 302975 463709
rect 314046 463700 314052 463712
rect 314104 463700 314110 463752
rect 268877 463675 268935 463681
rect 268877 463641 268889 463675
rect 268923 463672 268935 463675
rect 359954 463672 359960 463684
rect 268923 463644 359960 463672
rect 268923 463641 268935 463644
rect 268877 463635 268935 463641
rect 359954 463632 359960 463644
rect 360012 463632 360018 463684
rect 257098 463564 257104 463616
rect 257156 463604 257162 463616
rect 355906 463604 355912 463616
rect 257156 463576 355912 463604
rect 257156 463564 257162 463576
rect 355906 463564 355912 463576
rect 355964 463564 355970 463616
rect 1600 463440 583316 463536
rect 258202 463360 258208 463412
rect 258260 463400 258266 463412
rect 358666 463400 358672 463412
rect 258260 463372 358672 463400
rect 258260 463360 258266 463372
rect 358666 463360 358672 463372
rect 358724 463360 358730 463412
rect 253970 463292 253976 463344
rect 254028 463332 254034 463344
rect 354526 463332 354532 463344
rect 254028 463304 354532 463332
rect 254028 463292 254034 463304
rect 354526 463292 354532 463304
rect 354584 463292 354590 463344
rect 185338 463224 185344 463276
rect 185396 463264 185402 463276
rect 283594 463264 283600 463276
rect 185396 463236 283600 463264
rect 185396 463224 185402 463236
rect 283594 463224 283600 463236
rect 283652 463224 283658 463276
rect 283689 463267 283747 463273
rect 283689 463233 283701 463267
rect 283735 463264 283747 463267
rect 284885 463267 284943 463273
rect 283735 463236 284836 463264
rect 283735 463233 283747 463236
rect 283689 463227 283747 463233
rect 250198 463156 250204 463208
rect 250256 463196 250262 463208
rect 284701 463199 284759 463205
rect 284701 463196 284713 463199
rect 250256 463168 284713 463196
rect 250256 463156 250262 463168
rect 284701 463165 284713 463168
rect 284747 463165 284759 463199
rect 284808 463196 284836 463236
rect 284885 463233 284897 463267
rect 284931 463264 284943 463267
rect 293070 463264 293076 463276
rect 284931 463236 293076 463264
rect 284931 463233 284943 463236
rect 284885 463227 284943 463233
rect 293070 463224 293076 463236
rect 293128 463224 293134 463276
rect 293162 463224 293168 463276
rect 293220 463264 293226 463276
rect 378814 463264 378820 463276
rect 293220 463236 378820 463264
rect 293220 463224 293226 463236
rect 378814 463224 378820 463236
rect 378872 463224 378878 463276
rect 302273 463199 302331 463205
rect 284808 463168 302224 463196
rect 284701 463159 284759 463165
rect 261330 463088 261336 463140
rect 261388 463128 261394 463140
rect 268877 463131 268935 463137
rect 268877 463128 268889 463131
rect 261388 463100 268889 463128
rect 261388 463088 261394 463100
rect 268877 463097 268889 463100
rect 268923 463097 268935 463131
rect 268877 463091 268935 463097
rect 278166 463088 278172 463140
rect 278224 463128 278230 463140
rect 282306 463128 282312 463140
rect 278224 463100 282312 463128
rect 278224 463088 278230 463100
rect 282306 463088 282312 463100
rect 282364 463088 282370 463140
rect 282398 463088 282404 463140
rect 282456 463128 282462 463140
rect 283318 463128 283324 463140
rect 282456 463100 283324 463128
rect 282456 463088 282462 463100
rect 283318 463088 283324 463100
rect 283376 463088 283382 463140
rect 283410 463088 283416 463140
rect 283468 463128 283474 463140
rect 283468 463100 288148 463128
rect 283468 463088 283474 463100
rect 264550 463020 264556 463072
rect 264608 463060 264614 463072
rect 265378 463060 265384 463072
rect 264608 463032 265384 463060
rect 264608 463020 264614 463032
rect 265378 463020 265384 463032
rect 265436 463020 265442 463072
rect 265562 463020 265568 463072
rect 265620 463060 265626 463072
rect 266666 463060 266672 463072
rect 265620 463032 266672 463060
rect 265620 463020 265626 463032
rect 266666 463020 266672 463032
rect 266724 463020 266730 463072
rect 268690 463020 268696 463072
rect 268748 463060 268754 463072
rect 269518 463060 269524 463072
rect 268748 463032 269524 463060
rect 268748 463020 268754 463032
rect 269518 463020 269524 463032
rect 269576 463020 269582 463072
rect 269794 463020 269800 463072
rect 269852 463060 269858 463072
rect 270898 463060 270904 463072
rect 269852 463032 270904 463060
rect 269852 463020 269858 463032
rect 270898 463020 270904 463032
rect 270956 463020 270962 463072
rect 272922 463020 272928 463072
rect 272980 463060 272986 463072
rect 273658 463060 273664 463072
rect 272980 463032 273664 463060
rect 272980 463020 272986 463032
rect 273658 463020 273664 463032
rect 273716 463020 273722 463072
rect 273934 463020 273940 463072
rect 273992 463060 273998 463072
rect 274946 463060 274952 463072
rect 273992 463032 274952 463060
rect 273992 463020 273998 463032
rect 274946 463020 274952 463032
rect 275004 463020 275010 463072
rect 279270 463020 279276 463072
rect 279328 463060 279334 463072
rect 280558 463060 280564 463072
rect 279328 463032 280564 463060
rect 279328 463020 279334 463032
rect 280558 463020 280564 463032
rect 280616 463020 280622 463072
rect 281386 463020 281392 463072
rect 281444 463060 281450 463072
rect 283689 463063 283747 463069
rect 283689 463060 283701 463063
rect 281444 463032 283701 463060
rect 281444 463020 281450 463032
rect 283689 463029 283701 463032
rect 283735 463029 283747 463063
rect 283689 463023 283747 463029
rect 283778 463020 283784 463072
rect 283836 463060 283842 463072
rect 284698 463060 284704 463072
rect 283836 463032 284704 463060
rect 283836 463020 283842 463032
rect 284698 463020 284704 463032
rect 284756 463020 284762 463072
rect 286630 463020 286636 463072
rect 286688 463060 286694 463072
rect 287458 463060 287464 463072
rect 286688 463032 287464 463060
rect 286688 463020 286694 463032
rect 287458 463020 287464 463032
rect 287516 463020 287522 463072
rect 288120 463060 288148 463100
rect 288194 463088 288200 463140
rect 288252 463128 288258 463140
rect 291601 463131 291659 463137
rect 291601 463128 291613 463131
rect 288252 463100 291613 463128
rect 288252 463088 288258 463100
rect 291601 463097 291613 463100
rect 291647 463097 291659 463131
rect 291601 463091 291659 463097
rect 291690 463088 291696 463140
rect 291748 463128 291754 463140
rect 292518 463128 292524 463140
rect 291748 463100 292524 463128
rect 291748 463088 291754 463100
rect 292518 463088 292524 463100
rect 292576 463088 292582 463140
rect 292613 463131 292671 463137
rect 292613 463097 292625 463131
rect 292659 463128 292671 463131
rect 301261 463131 301319 463137
rect 301261 463128 301273 463131
rect 292659 463100 301273 463128
rect 292659 463097 292671 463100
rect 292613 463091 292671 463097
rect 301261 463097 301273 463100
rect 301307 463097 301319 463131
rect 301261 463091 301319 463097
rect 301350 463088 301356 463140
rect 301408 463128 301414 463140
rect 302086 463128 302092 463140
rect 301408 463100 302092 463128
rect 301408 463088 301414 463100
rect 302086 463088 302092 463100
rect 302144 463088 302150 463140
rect 302196 463128 302224 463168
rect 302273 463165 302285 463199
rect 302319 463196 302331 463199
rect 443585 463199 443643 463205
rect 443585 463196 443597 463199
rect 302319 463168 443597 463196
rect 302319 463165 302331 463168
rect 302273 463159 302331 463165
rect 443585 463165 443597 463168
rect 443631 463165 443643 463199
rect 443585 463159 443643 463165
rect 508534 463128 508540 463140
rect 302196 463100 508540 463128
rect 508534 463088 508540 463100
rect 508592 463088 508598 463140
rect 573305 463063 573363 463069
rect 573305 463060 573317 463063
rect 288120 463032 573317 463060
rect 573305 463029 573317 463032
rect 573351 463029 573363 463063
rect 573305 463023 573363 463029
rect 1600 462896 583316 462992
rect 255074 462816 255080 462868
rect 255132 462856 255138 462868
rect 357194 462856 357200 462868
rect 255132 462828 357200 462856
rect 255132 462816 255138 462828
rect 357194 462816 357200 462828
rect 357252 462816 357258 462868
rect 4374 462748 4380 462800
rect 4432 462788 4438 462800
rect 330790 462788 330796 462800
rect 4432 462760 330796 462788
rect 4432 462748 4438 462760
rect 330790 462748 330796 462760
rect 330848 462748 330854 462800
rect 4282 462680 4288 462732
rect 4340 462720 4346 462732
rect 333918 462720 333924 462732
rect 4340 462692 333924 462720
rect 4340 462680 4346 462692
rect 333918 462680 333924 462692
rect 333976 462680 333982 462732
rect 4190 462612 4196 462664
rect 4248 462652 4254 462664
rect 337138 462652 337144 462664
rect 4248 462624 337144 462652
rect 4248 462612 4254 462624
rect 337138 462612 337144 462624
rect 337196 462612 337202 462664
rect 4006 462544 4012 462596
rect 4064 462584 4070 462596
rect 339254 462584 339260 462596
rect 4064 462556 339260 462584
rect 4064 462544 4070 462556
rect 339254 462544 339260 462556
rect 339312 462544 339318 462596
rect 4098 462476 4104 462528
rect 4156 462516 4162 462528
rect 340266 462516 340272 462528
rect 4156 462488 340272 462516
rect 4156 462476 4162 462488
rect 340266 462476 340272 462488
rect 340324 462476 340330 462528
rect 1600 462352 583316 462448
rect 291138 462272 291144 462324
rect 291196 462312 291202 462324
rect 292613 462315 292671 462321
rect 292613 462312 292625 462315
rect 291196 462284 292625 462312
rect 291196 462272 291202 462284
rect 292613 462281 292625 462284
rect 292659 462281 292671 462315
rect 292613 462275 292671 462281
rect 313862 462272 313868 462324
rect 313920 462312 313926 462324
rect 314782 462312 314788 462324
rect 313920 462284 314788 462312
rect 313920 462272 313926 462284
rect 314782 462272 314788 462284
rect 314840 462272 314846 462324
rect 284698 462204 284704 462256
rect 284756 462244 284762 462256
rect 302273 462247 302331 462253
rect 302273 462244 302285 462247
rect 284756 462216 302285 462244
rect 284756 462204 284762 462216
rect 302273 462213 302285 462216
rect 302319 462213 302331 462247
rect 302273 462207 302331 462213
rect 291601 462179 291659 462185
rect 291601 462145 291613 462179
rect 291647 462176 291659 462179
rect 296750 462176 296756 462188
rect 291647 462148 296756 462176
rect 291647 462145 291659 462148
rect 291601 462139 291659 462145
rect 296750 462136 296756 462148
rect 296808 462136 296814 462188
rect 301261 462179 301319 462185
rect 301261 462145 301273 462179
rect 301307 462176 301319 462179
rect 302917 462179 302975 462185
rect 302917 462176 302929 462179
rect 301307 462148 302929 462176
rect 301307 462145 301319 462148
rect 301261 462139 301319 462145
rect 302917 462145 302929 462148
rect 302963 462145 302975 462179
rect 302917 462139 302975 462145
rect 1600 461808 583316 461904
rect 228946 461524 228952 461576
rect 229004 461564 229010 461576
rect 328674 461564 328680 461576
rect 229004 461536 328680 461564
rect 229004 461524 229010 461536
rect 328674 461524 328680 461536
rect 328732 461524 328738 461576
rect 220574 461456 220580 461508
rect 220632 461496 220638 461508
rect 324534 461496 324540 461508
rect 220632 461468 324540 461496
rect 220632 461456 220638 461468
rect 324534 461456 324540 461468
rect 324592 461456 324598 461508
rect 240262 461388 240268 461440
rect 240320 461428 240326 461440
rect 351674 461428 351680 461440
rect 240320 461400 351680 461428
rect 240320 461388 240326 461400
rect 351674 461388 351680 461400
rect 351732 461388 351738 461440
rect 1600 461264 583316 461360
rect 235018 461184 235024 461236
rect 235076 461224 235082 461236
rect 361334 461224 361340 461236
rect 235076 461196 361340 461224
rect 235076 461184 235082 461196
rect 361334 461184 361340 461196
rect 361392 461184 361398 461236
rect 259214 461116 259220 461168
rect 259272 461156 259278 461168
rect 411014 461156 411020 461168
rect 259272 461128 411020 461156
rect 259272 461116 259278 461128
rect 411014 461116 411020 461128
rect 411072 461116 411078 461168
rect 179174 461048 179180 461100
rect 179232 461088 179238 461100
rect 332906 461088 332912 461100
rect 179232 461060 332912 461088
rect 179232 461048 179238 461060
rect 332906 461048 332912 461060
rect 332964 461048 332970 461100
rect 6766 460980 6772 461032
rect 6824 461020 6830 461032
rect 322418 461020 322424 461032
rect 6824 460992 322424 461020
rect 6824 460980 6830 460992
rect 322418 460980 322424 460992
rect 322476 460980 322482 461032
rect 260318 460912 260324 460964
rect 260376 460952 260382 460964
rect 580662 460952 580668 460964
rect 260376 460924 580668 460952
rect 260376 460912 260382 460924
rect 580662 460912 580668 460924
rect 580720 460912 580726 460964
rect 1600 460720 583316 460816
rect 228854 460300 228860 460352
rect 228912 460340 228918 460352
rect 335022 460340 335028 460352
rect 228912 460312 335028 460340
rect 228912 460300 228918 460312
rect 335022 460300 335028 460312
rect 335080 460300 335086 460352
rect 1600 460176 583316 460272
rect 243482 460096 243488 460148
rect 243540 460136 243546 460148
rect 353054 460136 353060 460148
rect 243540 460108 353060 460136
rect 243540 460096 243546 460108
rect 353054 460096 353060 460108
rect 353112 460096 353118 460148
rect 225361 460071 225419 460077
rect 225361 460068 225373 460071
rect 215808 460040 225373 460068
rect 3638 459756 3644 459808
rect 3696 459796 3702 459808
rect 7321 459799 7379 459805
rect 7321 459796 7333 459799
rect 3696 459768 7333 459796
rect 3696 459756 3702 459768
rect 7321 459765 7333 459768
rect 7367 459765 7379 459799
rect 7321 459759 7379 459765
rect 7413 459799 7471 459805
rect 7413 459765 7425 459799
rect 7459 459796 7471 459799
rect 16981 459799 17039 459805
rect 16981 459796 16993 459799
rect 7459 459768 16993 459796
rect 7459 459765 7471 459768
rect 7413 459759 7471 459765
rect 16981 459765 16993 459768
rect 17027 459765 17039 459799
rect 16981 459759 17039 459765
rect 17073 459799 17131 459805
rect 17073 459765 17085 459799
rect 17119 459796 17131 459799
rect 26641 459799 26699 459805
rect 26641 459796 26653 459799
rect 17119 459768 26653 459796
rect 17119 459765 17131 459768
rect 17073 459759 17131 459765
rect 26641 459765 26653 459768
rect 26687 459765 26699 459799
rect 26641 459759 26699 459765
rect 26733 459799 26791 459805
rect 26733 459765 26745 459799
rect 26779 459796 26791 459799
rect 36301 459799 36359 459805
rect 36301 459796 36313 459799
rect 26779 459768 36313 459796
rect 26779 459765 26791 459768
rect 26733 459759 26791 459765
rect 36301 459765 36313 459768
rect 36347 459765 36359 459799
rect 36301 459759 36359 459765
rect 36393 459799 36451 459805
rect 36393 459765 36405 459799
rect 36439 459796 36451 459799
rect 45961 459799 46019 459805
rect 45961 459796 45973 459799
rect 36439 459768 45973 459796
rect 36439 459765 36451 459768
rect 36393 459759 36451 459765
rect 45961 459765 45973 459768
rect 46007 459765 46019 459799
rect 45961 459759 46019 459765
rect 46053 459799 46111 459805
rect 46053 459765 46065 459799
rect 46099 459796 46111 459799
rect 55621 459799 55679 459805
rect 55621 459796 55633 459799
rect 46099 459768 55633 459796
rect 46099 459765 46111 459768
rect 46053 459759 46111 459765
rect 55621 459765 55633 459768
rect 55667 459765 55679 459799
rect 55621 459759 55679 459765
rect 55713 459799 55771 459805
rect 55713 459765 55725 459799
rect 55759 459796 55771 459799
rect 65281 459799 65339 459805
rect 65281 459796 65293 459799
rect 55759 459768 65293 459796
rect 55759 459765 55771 459768
rect 55713 459759 55771 459765
rect 65281 459765 65293 459768
rect 65327 459765 65339 459799
rect 65281 459759 65339 459765
rect 65373 459799 65431 459805
rect 65373 459765 65385 459799
rect 65419 459796 65431 459799
rect 74941 459799 74999 459805
rect 74941 459796 74953 459799
rect 65419 459768 74953 459796
rect 65419 459765 65431 459768
rect 65373 459759 65431 459765
rect 74941 459765 74953 459768
rect 74987 459765 74999 459799
rect 74941 459759 74999 459765
rect 75033 459799 75091 459805
rect 75033 459765 75045 459799
rect 75079 459796 75091 459799
rect 84601 459799 84659 459805
rect 84601 459796 84613 459799
rect 75079 459768 84613 459796
rect 75079 459765 75091 459768
rect 75033 459759 75091 459765
rect 84601 459765 84613 459768
rect 84647 459765 84659 459799
rect 84601 459759 84659 459765
rect 84693 459799 84751 459805
rect 84693 459765 84705 459799
rect 84739 459796 84751 459799
rect 94261 459799 94319 459805
rect 94261 459796 94273 459799
rect 84739 459768 94273 459796
rect 84739 459765 84751 459768
rect 84693 459759 84751 459765
rect 94261 459765 94273 459768
rect 94307 459765 94319 459799
rect 94261 459759 94319 459765
rect 94353 459799 94411 459805
rect 94353 459765 94365 459799
rect 94399 459796 94411 459799
rect 103921 459799 103979 459805
rect 103921 459796 103933 459799
rect 94399 459768 103933 459796
rect 94399 459765 94411 459768
rect 94353 459759 94411 459765
rect 103921 459765 103933 459768
rect 103967 459765 103979 459799
rect 103921 459759 103979 459765
rect 104013 459799 104071 459805
rect 104013 459765 104025 459799
rect 104059 459796 104071 459799
rect 113581 459799 113639 459805
rect 113581 459796 113593 459799
rect 104059 459768 113593 459796
rect 104059 459765 104071 459768
rect 104013 459759 104071 459765
rect 113581 459765 113593 459768
rect 113627 459765 113639 459799
rect 113581 459759 113639 459765
rect 113673 459799 113731 459805
rect 113673 459765 113685 459799
rect 113719 459796 113731 459799
rect 123241 459799 123299 459805
rect 123241 459796 123253 459799
rect 113719 459768 123253 459796
rect 113719 459765 113731 459768
rect 113673 459759 113731 459765
rect 123241 459765 123253 459768
rect 123287 459765 123299 459799
rect 123241 459759 123299 459765
rect 123333 459799 123391 459805
rect 123333 459765 123345 459799
rect 123379 459796 123391 459799
rect 132901 459799 132959 459805
rect 132901 459796 132913 459799
rect 123379 459768 132913 459796
rect 123379 459765 123391 459768
rect 123333 459759 123391 459765
rect 132901 459765 132913 459768
rect 132947 459765 132959 459799
rect 132901 459759 132959 459765
rect 132993 459799 133051 459805
rect 132993 459765 133005 459799
rect 133039 459796 133051 459799
rect 142561 459799 142619 459805
rect 142561 459796 142573 459799
rect 133039 459768 142573 459796
rect 133039 459765 133051 459768
rect 132993 459759 133051 459765
rect 142561 459765 142573 459768
rect 142607 459765 142619 459799
rect 142561 459759 142619 459765
rect 142653 459799 142711 459805
rect 142653 459765 142665 459799
rect 142699 459796 142711 459799
rect 152221 459799 152279 459805
rect 152221 459796 152233 459799
rect 142699 459768 152233 459796
rect 142699 459765 142711 459768
rect 142653 459759 142711 459765
rect 152221 459765 152233 459768
rect 152267 459765 152279 459799
rect 152221 459759 152279 459765
rect 152313 459799 152371 459805
rect 152313 459765 152325 459799
rect 152359 459796 152371 459799
rect 161881 459799 161939 459805
rect 161881 459796 161893 459799
rect 152359 459768 161893 459796
rect 152359 459765 152371 459768
rect 152313 459759 152371 459765
rect 161881 459765 161893 459768
rect 161927 459765 161939 459799
rect 161881 459759 161939 459765
rect 161973 459799 162031 459805
rect 161973 459765 161985 459799
rect 162019 459796 162031 459799
rect 171541 459799 171599 459805
rect 171541 459796 171553 459799
rect 162019 459768 171553 459796
rect 162019 459765 162031 459768
rect 161973 459759 162031 459765
rect 171541 459765 171553 459768
rect 171587 459765 171599 459799
rect 171541 459759 171599 459765
rect 171633 459799 171691 459805
rect 171633 459765 171645 459799
rect 171679 459796 171691 459799
rect 181201 459799 181259 459805
rect 181201 459796 181213 459799
rect 171679 459768 181213 459796
rect 171679 459765 171691 459768
rect 171633 459759 171691 459765
rect 181201 459765 181213 459768
rect 181247 459765 181259 459799
rect 181201 459759 181259 459765
rect 181293 459799 181351 459805
rect 181293 459765 181305 459799
rect 181339 459796 181351 459799
rect 190861 459799 190919 459805
rect 190861 459796 190873 459799
rect 181339 459768 190873 459796
rect 181339 459765 181351 459768
rect 181293 459759 181351 459765
rect 190861 459765 190873 459768
rect 190907 459765 190919 459799
rect 190861 459759 190919 459765
rect 190953 459799 191011 459805
rect 190953 459765 190965 459799
rect 190999 459796 191011 459799
rect 200521 459799 200579 459805
rect 200521 459796 200533 459799
rect 190999 459768 200533 459796
rect 190999 459765 191011 459768
rect 190953 459759 191011 459765
rect 200521 459765 200533 459768
rect 200567 459765 200579 459799
rect 200521 459759 200579 459765
rect 200613 459799 200671 459805
rect 200613 459765 200625 459799
rect 200659 459796 200671 459799
rect 210181 459799 210239 459805
rect 210181 459796 210193 459799
rect 200659 459768 210193 459796
rect 200659 459765 200671 459768
rect 200613 459759 200671 459765
rect 210181 459765 210193 459768
rect 210227 459765 210239 459799
rect 210181 459759 210239 459765
rect 210273 459799 210331 459805
rect 210273 459765 210285 459799
rect 210319 459796 210331 459799
rect 215808 459796 215836 460040
rect 225361 460037 225373 460040
rect 225407 460037 225419 460071
rect 225361 460031 225419 460037
rect 227566 460028 227572 460080
rect 227624 460068 227630 460080
rect 325270 460068 325276 460080
rect 227624 460040 325276 460068
rect 227624 460028 227630 460040
rect 325270 460028 325276 460040
rect 325328 460028 325334 460080
rect 223334 459960 223340 460012
rect 223392 460000 223398 460012
rect 326374 460000 326380 460012
rect 223392 459972 326380 460000
rect 223392 459960 223398 459972
rect 326374 459960 326380 459972
rect 326432 459960 326438 460012
rect 252774 459892 252780 459944
rect 252832 459932 252838 459944
rect 355814 459932 355820 459944
rect 252832 459904 355820 459932
rect 252832 459892 252838 459904
rect 355814 459892 355820 459904
rect 355872 459892 355878 459944
rect 225361 459867 225419 459873
rect 225361 459833 225373 459867
rect 225407 459864 225419 459867
rect 229501 459867 229559 459873
rect 229501 459864 229513 459867
rect 225407 459836 229513 459864
rect 225407 459833 225419 459836
rect 225361 459827 225419 459833
rect 229501 459833 229513 459836
rect 229547 459833 229559 459867
rect 229501 459827 229559 459833
rect 248082 459824 248088 459876
rect 248140 459864 248146 459876
rect 358574 459864 358580 459876
rect 248140 459836 358580 459864
rect 248140 459824 248146 459836
rect 358574 459824 358580 459836
rect 358632 459824 358638 459876
rect 210319 459768 215836 459796
rect 210319 459765 210331 459768
rect 210273 459759 210331 459765
rect 224714 459756 224720 459808
rect 224772 459796 224778 459808
rect 335850 459796 335856 459808
rect 224772 459768 335856 459796
rect 224772 459756 224778 459768
rect 335850 459756 335856 459768
rect 335908 459756 335914 459808
rect 261333 459731 261391 459737
rect 261333 459728 261345 459731
rect 1600 459632 230496 459728
rect 261256 459700 261345 459728
rect 234282 459660 234288 459672
rect 234243 459632 234288 459660
rect 234282 459620 234288 459632
rect 234340 459620 234346 459672
rect 242013 459663 242071 459669
rect 242013 459660 242025 459663
rect 235864 459632 242025 459660
rect 7413 459595 7471 459601
rect 7413 459561 7425 459595
rect 7459 459561 7471 459595
rect 7413 459555 7471 459561
rect 16981 459595 17039 459601
rect 16981 459561 16993 459595
rect 17027 459592 17039 459595
rect 17073 459595 17131 459601
rect 17073 459592 17085 459595
rect 17027 459564 17085 459592
rect 17027 459561 17039 459564
rect 16981 459555 17039 459561
rect 17073 459561 17085 459564
rect 17119 459561 17131 459595
rect 17073 459555 17131 459561
rect 26733 459595 26791 459601
rect 26733 459561 26745 459595
rect 26779 459561 26791 459595
rect 26733 459555 26791 459561
rect 36301 459595 36359 459601
rect 36301 459561 36313 459595
rect 36347 459592 36359 459595
rect 36393 459595 36451 459601
rect 36393 459592 36405 459595
rect 36347 459564 36405 459592
rect 36347 459561 36359 459564
rect 36301 459555 36359 459561
rect 36393 459561 36405 459564
rect 36439 459561 36451 459595
rect 36393 459555 36451 459561
rect 46053 459595 46111 459601
rect 46053 459561 46065 459595
rect 46099 459561 46111 459595
rect 46053 459555 46111 459561
rect 55621 459595 55679 459601
rect 55621 459561 55633 459595
rect 55667 459592 55679 459595
rect 55713 459595 55771 459601
rect 55713 459592 55725 459595
rect 55667 459564 55725 459592
rect 55667 459561 55679 459564
rect 55621 459555 55679 459561
rect 55713 459561 55725 459564
rect 55759 459561 55771 459595
rect 55713 459555 55771 459561
rect 65373 459595 65431 459601
rect 65373 459561 65385 459595
rect 65419 459561 65431 459595
rect 65373 459555 65431 459561
rect 74941 459595 74999 459601
rect 74941 459561 74953 459595
rect 74987 459592 74999 459595
rect 75033 459595 75091 459601
rect 75033 459592 75045 459595
rect 74987 459564 75045 459592
rect 74987 459561 74999 459564
rect 74941 459555 74999 459561
rect 75033 459561 75045 459564
rect 75079 459561 75091 459595
rect 75033 459555 75091 459561
rect 84693 459595 84751 459601
rect 84693 459561 84705 459595
rect 84739 459561 84751 459595
rect 84693 459555 84751 459561
rect 94261 459595 94319 459601
rect 94261 459561 94273 459595
rect 94307 459592 94319 459595
rect 94353 459595 94411 459601
rect 94353 459592 94365 459595
rect 94307 459564 94365 459592
rect 94307 459561 94319 459564
rect 94261 459555 94319 459561
rect 94353 459561 94365 459564
rect 94399 459561 94411 459595
rect 94353 459555 94411 459561
rect 104013 459595 104071 459601
rect 104013 459561 104025 459595
rect 104059 459561 104071 459595
rect 104013 459555 104071 459561
rect 113581 459595 113639 459601
rect 113581 459561 113593 459595
rect 113627 459592 113639 459595
rect 113673 459595 113731 459601
rect 113673 459592 113685 459595
rect 113627 459564 113685 459592
rect 113627 459561 113639 459564
rect 113581 459555 113639 459561
rect 113673 459561 113685 459564
rect 113719 459561 113731 459595
rect 113673 459555 113731 459561
rect 123333 459595 123391 459601
rect 123333 459561 123345 459595
rect 123379 459561 123391 459595
rect 123333 459555 123391 459561
rect 132901 459595 132959 459601
rect 132901 459561 132913 459595
rect 132947 459592 132959 459595
rect 132993 459595 133051 459601
rect 132993 459592 133005 459595
rect 132947 459564 133005 459592
rect 132947 459561 132959 459564
rect 132901 459555 132959 459561
rect 132993 459561 133005 459564
rect 133039 459561 133051 459595
rect 132993 459555 133051 459561
rect 142653 459595 142711 459601
rect 142653 459561 142665 459595
rect 142699 459561 142711 459595
rect 142653 459555 142711 459561
rect 152221 459595 152279 459601
rect 152221 459561 152233 459595
rect 152267 459592 152279 459595
rect 152313 459595 152371 459601
rect 152313 459592 152325 459595
rect 152267 459564 152325 459592
rect 152267 459561 152279 459564
rect 152221 459555 152279 459561
rect 152313 459561 152325 459564
rect 152359 459561 152371 459595
rect 152313 459555 152371 459561
rect 161973 459595 162031 459601
rect 161973 459561 161985 459595
rect 162019 459561 162031 459595
rect 161973 459555 162031 459561
rect 171541 459595 171599 459601
rect 171541 459561 171553 459595
rect 171587 459592 171599 459595
rect 171633 459595 171691 459601
rect 171633 459592 171645 459595
rect 171587 459564 171645 459592
rect 171587 459561 171599 459564
rect 171541 459555 171599 459561
rect 171633 459561 171645 459564
rect 171679 459561 171691 459595
rect 171633 459555 171691 459561
rect 181293 459595 181351 459601
rect 181293 459561 181305 459595
rect 181339 459561 181351 459595
rect 181293 459555 181351 459561
rect 190861 459595 190919 459601
rect 190861 459561 190873 459595
rect 190907 459592 190919 459595
rect 190953 459595 191011 459601
rect 190953 459592 190965 459595
rect 190907 459564 190965 459592
rect 190907 459561 190919 459564
rect 190861 459555 190919 459561
rect 190953 459561 190965 459564
rect 190999 459561 191011 459595
rect 190953 459555 191011 459561
rect 200613 459595 200671 459601
rect 200613 459561 200625 459595
rect 200659 459561 200671 459595
rect 200613 459555 200671 459561
rect 210181 459595 210239 459601
rect 210181 459561 210193 459595
rect 210227 459592 210239 459595
rect 210273 459595 210331 459601
rect 210273 459592 210285 459595
rect 210227 459564 210285 459592
rect 210227 459561 210239 459564
rect 210181 459555 210239 459561
rect 210273 459561 210285 459564
rect 210319 459561 210331 459595
rect 210273 459555 210331 459561
rect 229501 459595 229559 459601
rect 229501 459561 229513 459595
rect 229547 459592 229559 459595
rect 235021 459595 235079 459601
rect 235021 459592 235033 459595
rect 229547 459564 235033 459592
rect 229547 459561 229559 459564
rect 229501 459555 229559 459561
rect 235021 459561 235033 459564
rect 235067 459561 235079 459595
rect 235021 459555 235079 459561
rect 235113 459595 235171 459601
rect 235113 459561 235125 459595
rect 235159 459592 235171 459595
rect 235864 459592 235892 459632
rect 242013 459629 242025 459632
rect 242059 459629 242071 459663
rect 250106 459660 250112 459672
rect 250067 459632 250112 459660
rect 242013 459623 242071 459629
rect 250106 459620 250112 459632
rect 250164 459620 250170 459672
rect 256362 459660 256368 459672
rect 256323 459632 256368 459660
rect 256362 459620 256368 459632
rect 256420 459620 256426 459672
rect 261256 459669 261284 459700
rect 261333 459697 261345 459700
rect 261379 459697 261391 459731
rect 280653 459731 280711 459737
rect 280653 459728 280665 459731
rect 261333 459691 261391 459697
rect 275792 459700 280665 459728
rect 261241 459663 261299 459669
rect 261241 459629 261253 459663
rect 261287 459629 261299 459663
rect 261241 459623 261299 459629
rect 235159 459564 235892 459592
rect 251581 459595 251639 459601
rect 235159 459561 235171 459564
rect 235113 459555 235171 459561
rect 251581 459561 251593 459595
rect 251627 459592 251639 459595
rect 270901 459595 270959 459601
rect 251627 459564 251716 459592
rect 251627 459561 251639 459564
rect 251581 459555 251639 459561
rect 7321 459527 7379 459533
rect 7321 459493 7333 459527
rect 7367 459524 7379 459527
rect 7428 459524 7456 459555
rect 7367 459496 7456 459524
rect 26641 459527 26699 459533
rect 7367 459493 7379 459496
rect 7321 459487 7379 459493
rect 26641 459493 26653 459527
rect 26687 459524 26699 459527
rect 26748 459524 26776 459555
rect 26687 459496 26776 459524
rect 45961 459527 46019 459533
rect 26687 459493 26699 459496
rect 26641 459487 26699 459493
rect 45961 459493 45973 459527
rect 46007 459524 46019 459527
rect 46068 459524 46096 459555
rect 46007 459496 46096 459524
rect 65281 459527 65339 459533
rect 46007 459493 46019 459496
rect 45961 459487 46019 459493
rect 65281 459493 65293 459527
rect 65327 459524 65339 459527
rect 65388 459524 65416 459555
rect 65327 459496 65416 459524
rect 84601 459527 84659 459533
rect 65327 459493 65339 459496
rect 65281 459487 65339 459493
rect 84601 459493 84613 459527
rect 84647 459524 84659 459527
rect 84708 459524 84736 459555
rect 84647 459496 84736 459524
rect 103921 459527 103979 459533
rect 84647 459493 84659 459496
rect 84601 459487 84659 459493
rect 103921 459493 103933 459527
rect 103967 459524 103979 459527
rect 104028 459524 104056 459555
rect 103967 459496 104056 459524
rect 123241 459527 123299 459533
rect 103967 459493 103979 459496
rect 103921 459487 103979 459493
rect 123241 459493 123253 459527
rect 123287 459524 123299 459527
rect 123348 459524 123376 459555
rect 123287 459496 123376 459524
rect 142561 459527 142619 459533
rect 123287 459493 123299 459496
rect 123241 459487 123299 459493
rect 142561 459493 142573 459527
rect 142607 459524 142619 459527
rect 142668 459524 142696 459555
rect 142607 459496 142696 459524
rect 161881 459527 161939 459533
rect 142607 459493 142619 459496
rect 142561 459487 142619 459493
rect 161881 459493 161893 459527
rect 161927 459524 161939 459527
rect 161988 459524 162016 459555
rect 161927 459496 162016 459524
rect 181201 459527 181259 459533
rect 161927 459493 161939 459496
rect 161881 459487 161939 459493
rect 181201 459493 181213 459527
rect 181247 459524 181259 459527
rect 181308 459524 181336 459555
rect 181247 459496 181336 459524
rect 200521 459527 200579 459533
rect 181247 459493 181259 459496
rect 181201 459487 181259 459493
rect 200521 459493 200533 459527
rect 200567 459524 200579 459527
rect 200628 459524 200656 459555
rect 251688 459533 251716 459564
rect 270901 459561 270913 459595
rect 270947 459592 270959 459595
rect 275792 459592 275820 459700
rect 280653 459697 280665 459700
rect 280699 459697 280711 459731
rect 319934 459728 319940 459740
rect 280653 459691 280711 459697
rect 313604 459700 319940 459728
rect 290221 459663 290279 459669
rect 290221 459629 290233 459663
rect 290267 459660 290279 459663
rect 292981 459663 293039 459669
rect 292981 459660 292993 459663
rect 290267 459632 292993 459660
rect 290267 459629 290279 459632
rect 290221 459623 290279 459629
rect 292981 459629 292993 459632
rect 293027 459629 293039 459663
rect 292981 459623 293039 459629
rect 309541 459663 309599 459669
rect 309541 459629 309553 459663
rect 309587 459660 309599 459663
rect 312301 459663 312359 459669
rect 312301 459660 312313 459663
rect 309587 459632 312313 459660
rect 309587 459629 309599 459632
rect 309541 459623 309599 459629
rect 312301 459629 312313 459632
rect 312347 459629 312359 459663
rect 312301 459623 312359 459629
rect 312393 459663 312451 459669
rect 312393 459629 312405 459663
rect 312439 459660 312451 459663
rect 313604 459660 313632 459700
rect 319934 459688 319940 459700
rect 319992 459688 319998 459740
rect 323522 459660 323528 459672
rect 312439 459632 313632 459660
rect 323483 459632 323528 459660
rect 312439 459629 312451 459632
rect 312393 459623 312451 459629
rect 323522 459620 323528 459632
rect 323580 459620 323586 459672
rect 327478 459660 327484 459672
rect 327439 459632 327484 459660
rect 327478 459620 327484 459632
rect 327536 459620 327542 459672
rect 329502 459660 329508 459672
rect 329463 459632 329508 459660
rect 329502 459620 329508 459632
rect 329560 459620 329566 459672
rect 331710 459660 331716 459672
rect 331671 459632 331716 459660
rect 331710 459620 331716 459632
rect 331768 459620 331774 459672
rect 337782 459660 337788 459672
rect 337743 459632 337788 459660
rect 337782 459620 337788 459632
rect 337840 459620 337846 459672
rect 341186 459620 341192 459672
rect 341244 459620 341250 459672
rect 345602 459660 345608 459672
rect 345563 459632 345608 459660
rect 345602 459620 345608 459632
rect 345660 459620 345666 459672
rect 350248 459632 583316 459728
rect 270947 459564 275820 459592
rect 293165 459595 293223 459601
rect 270947 459561 270959 459564
rect 270901 459555 270959 459561
rect 293165 459561 293177 459595
rect 293211 459592 293223 459595
rect 299973 459595 300031 459601
rect 299973 459592 299985 459595
rect 293211 459564 299985 459592
rect 293211 459561 293223 459564
rect 293165 459555 293223 459561
rect 299973 459561 299985 459564
rect 300019 459561 300031 459595
rect 299973 459555 300031 459561
rect 200567 459496 200656 459524
rect 251673 459527 251731 459533
rect 200567 459493 200579 459496
rect 200521 459487 200579 459493
rect 251673 459493 251685 459527
rect 251719 459493 251731 459527
rect 251673 459487 251731 459493
rect 280653 459527 280711 459533
rect 280653 459493 280665 459527
rect 280699 459524 280711 459527
rect 290221 459527 290279 459533
rect 290221 459524 290233 459527
rect 280699 459496 290233 459524
rect 280699 459493 280711 459496
rect 280653 459487 280711 459493
rect 290221 459493 290233 459496
rect 290267 459493 290279 459527
rect 290221 459487 290279 459493
rect 242013 459459 242071 459465
rect 242013 459425 242025 459459
rect 242059 459456 242071 459459
rect 251581 459459 251639 459465
rect 251581 459456 251593 459459
rect 242059 459428 251593 459456
rect 242059 459425 242071 459428
rect 242013 459419 242071 459425
rect 251581 459425 251593 459428
rect 251627 459425 251639 459459
rect 251581 459419 251639 459425
rect 261333 459459 261391 459465
rect 261333 459425 261345 459459
rect 261379 459456 261391 459459
rect 270901 459459 270959 459465
rect 270901 459456 270913 459459
rect 261379 459428 270913 459456
rect 261379 459425 261391 459428
rect 261333 459419 261391 459425
rect 270901 459425 270913 459428
rect 270947 459425 270959 459459
rect 270901 459419 270959 459425
rect 299973 459459 300031 459465
rect 299973 459425 299985 459459
rect 300019 459456 300031 459459
rect 309541 459459 309599 459465
rect 309541 459456 309553 459459
rect 300019 459428 309553 459456
rect 300019 459425 300031 459428
rect 299973 459419 300031 459425
rect 309541 459425 309553 459428
rect 309587 459425 309599 459459
rect 309541 459419 309599 459425
rect 251673 459391 251731 459397
rect 251673 459357 251685 459391
rect 251719 459388 251731 459391
rect 261241 459391 261299 459397
rect 261241 459388 261253 459391
rect 251719 459360 261253 459388
rect 251719 459357 251731 459360
rect 251673 459351 251731 459357
rect 261241 459357 261253 459360
rect 261287 459357 261299 459391
rect 261241 459351 261299 459357
rect 1600 459088 230496 459184
rect 227474 458940 227480 458992
rect 227532 458980 227538 458992
rect 341204 458980 341232 459620
rect 350248 459088 583316 459184
rect 227532 458952 341232 458980
rect 227532 458940 227538 458952
rect 250109 458915 250167 458921
rect 250109 458881 250121 458915
rect 250155 458912 250167 458915
rect 354434 458912 354440 458924
rect 250155 458884 354440 458912
rect 250155 458881 250167 458884
rect 250109 458875 250167 458881
rect 354434 458872 354440 458884
rect 354492 458872 354498 458924
rect 226186 458804 226192 458856
rect 226244 458844 226250 458856
rect 323525 458847 323583 458853
rect 323525 458844 323537 458847
rect 226244 458816 323537 458844
rect 226244 458804 226250 458816
rect 323525 458813 323537 458816
rect 323571 458813 323583 458847
rect 323525 458807 323583 458813
rect 226094 458736 226100 458788
rect 226152 458776 226158 458788
rect 329505 458779 329563 458785
rect 329505 458776 329517 458779
rect 226152 458748 329517 458776
rect 226152 458736 226158 458748
rect 329505 458745 329517 458748
rect 329551 458745 329563 458779
rect 329505 458739 329563 458745
rect 221954 458668 221960 458720
rect 222012 458708 222018 458720
rect 327481 458711 327539 458717
rect 327481 458708 327493 458711
rect 222012 458680 327493 458708
rect 222012 458668 222018 458680
rect 327481 458677 327493 458680
rect 327527 458677 327539 458711
rect 327481 458671 327539 458677
rect 1600 458544 230496 458640
rect 350248 458544 583316 458640
rect 219194 458464 219200 458516
rect 219252 458504 219258 458516
rect 345605 458507 345663 458513
rect 345605 458504 345617 458507
rect 219252 458476 345617 458504
rect 219252 458464 219258 458476
rect 345605 458473 345617 458476
rect 345651 458473 345663 458507
rect 345605 458467 345663 458473
rect 256365 458439 256423 458445
rect 256365 458405 256377 458439
rect 256411 458436 256423 458439
rect 406874 458436 406880 458448
rect 256411 458408 406880 458436
rect 256411 458405 256423 458408
rect 256365 458399 256423 458405
rect 406874 458396 406880 458408
rect 406932 458396 406938 458448
rect 6674 458328 6680 458380
rect 6732 458368 6738 458380
rect 331713 458371 331771 458377
rect 331713 458368 331725 458371
rect 6732 458340 331725 458368
rect 6732 458328 6738 458340
rect 331713 458337 331725 458340
rect 331759 458337 331771 458371
rect 331713 458331 331771 458337
rect 9434 458260 9440 458312
rect 9492 458300 9498 458312
rect 337785 458303 337843 458309
rect 337785 458300 337797 458303
rect 9492 458272 337797 458300
rect 9492 458260 9498 458272
rect 337785 458269 337797 458272
rect 337831 458269 337843 458303
rect 337785 458263 337843 458269
rect 234285 458235 234343 458241
rect 234285 458201 234297 458235
rect 234331 458232 234343 458235
rect 580754 458232 580760 458244
rect 234331 458204 580760 458232
rect 234331 458201 234343 458204
rect 234285 458195 234343 458201
rect 580754 458192 580760 458204
rect 580812 458192 580818 458244
rect 1600 458000 230496 458096
rect 350248 458000 583316 458096
rect 1600 457456 230496 457552
rect 350248 457456 583316 457552
rect 1600 456912 230496 457008
rect 350248 456912 583316 457008
rect 1600 456368 230496 456464
rect 350248 456368 583316 456464
rect 1600 455824 230496 455920
rect 350248 455824 583316 455920
rect 1600 455280 230496 455376
rect 350248 455280 583316 455376
rect 1600 454736 230496 454832
rect 350248 454736 583316 454832
rect 1600 454192 230496 454288
rect 350248 454192 583316 454288
rect 1600 453648 230496 453744
rect 350248 453648 583316 453744
rect 1600 453104 230496 453200
rect 350248 453104 583316 453200
rect 1600 452560 230496 452656
rect 350248 452560 583316 452656
rect 1600 452016 230496 452112
rect 350248 452016 583316 452112
rect 1600 451472 230496 451568
rect 350248 451472 583316 451568
rect 1600 450928 230496 451024
rect 350248 450928 583316 451024
rect 1600 450384 230496 450480
rect 350248 450384 583316 450480
rect 1600 449840 230496 449936
rect 350248 449840 583316 449936
rect 1600 449296 230496 449392
rect 350248 449296 583316 449392
rect 1600 448752 230496 448848
rect 350248 448752 583316 448848
rect 1600 448208 230496 448304
rect 350248 448208 583316 448304
rect 1600 447664 230496 447760
rect 350248 447664 583316 447760
rect 1600 447120 230496 447216
rect 350248 447120 583316 447216
rect 359954 447040 359960 447092
rect 360012 447080 360018 447092
rect 580662 447080 580668 447092
rect 360012 447052 580668 447080
rect 360012 447040 360018 447052
rect 580662 447040 580668 447052
rect 580720 447040 580726 447092
rect 1600 446576 230496 446672
rect 350248 446576 583316 446672
rect 1600 446032 230496 446128
rect 350248 446032 583316 446128
rect 1600 445488 230496 445584
rect 350248 445488 583316 445584
rect 1600 444944 230496 445040
rect 350248 444944 583316 445040
rect 1600 444400 230496 444496
rect 350248 444400 583316 444496
rect 3638 444116 3644 444168
rect 3696 444156 3702 444168
rect 6766 444156 6772 444168
rect 3696 444128 6772 444156
rect 3696 444116 3702 444128
rect 6766 444116 6772 444128
rect 6824 444116 6830 444168
rect 1600 443856 230496 443952
rect 350248 443856 583316 443952
rect 1600 443312 230496 443408
rect 350248 443312 583316 443408
rect 1600 442768 230496 442864
rect 350248 442768 583316 442864
rect 1600 442224 230496 442320
rect 350248 442224 583316 442320
rect 1600 441680 230496 441776
rect 350248 441680 583316 441776
rect 1600 441136 230496 441232
rect 350248 441136 583316 441232
rect 1600 440592 230496 440688
rect 350248 440592 583316 440688
rect 1600 440048 230496 440144
rect 350248 440048 583316 440144
rect 1600 439504 230496 439600
rect 350248 439504 583316 439600
rect 1600 438960 230496 439056
rect 350248 438960 583316 439056
rect 1600 438416 230496 438512
rect 350248 438416 583316 438512
rect 1600 437872 230496 437968
rect 350248 437872 583316 437968
rect 1600 437328 230496 437424
rect 350248 437328 583316 437424
rect 1600 436784 230496 436880
rect 350248 436784 583316 436880
rect 1600 436240 230496 436336
rect 350248 436240 583316 436336
rect 1600 435696 230496 435792
rect 350248 435696 583316 435792
rect 1600 435152 230496 435248
rect 350248 435152 583316 435248
rect 1600 434608 230496 434704
rect 350248 434608 583316 434704
rect 1600 434064 230496 434160
rect 350248 434064 583316 434160
rect 1600 433520 230496 433616
rect 350248 433520 583316 433616
rect 1600 432976 230496 433072
rect 350248 432976 583316 433072
rect 1600 432432 230496 432528
rect 350248 432432 583316 432528
rect 1600 431888 230496 431984
rect 350248 431888 583316 431984
rect 1600 431344 230496 431440
rect 350248 431344 583316 431440
rect 1600 430800 230496 430896
rect 350248 430800 583316 430896
rect 411014 430516 411020 430568
rect 411072 430556 411078 430568
rect 580662 430556 580668 430568
rect 411072 430528 580668 430556
rect 411072 430516 411078 430528
rect 580662 430516 580668 430528
rect 580720 430516 580726 430568
rect 1600 430256 230496 430352
rect 350248 430256 583316 430352
rect 1600 429712 230496 429808
rect 350248 429712 583316 429808
rect 1600 429168 230496 429264
rect 350248 429168 583316 429264
rect 1600 428624 230496 428720
rect 350248 428624 583316 428720
rect 1600 428080 230496 428176
rect 350248 428080 583316 428176
rect 3638 427728 3644 427780
rect 3696 427768 3702 427780
rect 220574 427768 220580 427780
rect 3696 427740 220580 427768
rect 3696 427728 3702 427740
rect 220574 427728 220580 427740
rect 220632 427728 220638 427780
rect 1600 427536 230496 427632
rect 350248 427536 583316 427632
rect 1600 426992 230496 427088
rect 350248 426992 583316 427088
rect 1600 426448 230496 426544
rect 350248 426448 583316 426544
rect 1600 425904 230496 426000
rect 350248 425904 583316 426000
rect 1600 425360 230496 425456
rect 350248 425360 583316 425456
rect 1600 424816 230496 424912
rect 350248 424816 583316 424912
rect 1600 424272 230496 424368
rect 350248 424272 583316 424368
rect 1600 423728 230496 423824
rect 350248 423728 583316 423824
rect 1600 423184 230496 423280
rect 350248 423184 583316 423280
rect 1600 422640 230496 422736
rect 350248 422640 583316 422736
rect 1600 422096 230496 422192
rect 350248 422096 583316 422192
rect 1600 421552 230496 421648
rect 350248 421552 583316 421648
rect 1600 421008 230496 421104
rect 350248 421008 583316 421104
rect 1600 420464 230496 420560
rect 350248 420464 583316 420560
rect 1600 419920 230496 420016
rect 350248 419920 583316 420016
rect 1600 419376 230496 419472
rect 350248 419376 583316 419472
rect 1600 418832 230496 418928
rect 350248 418832 583316 418928
rect 1600 418288 230496 418384
rect 350248 418288 583316 418384
rect 1600 417744 230496 417840
rect 350248 417744 583316 417840
rect 1600 417200 230496 417296
rect 350248 417200 583316 417296
rect 1600 416656 230496 416752
rect 350248 416656 583316 416752
rect 1600 416112 230496 416208
rect 350248 416112 583316 416208
rect 1600 415568 230496 415664
rect 350248 415568 583316 415664
rect 355906 415352 355912 415404
rect 355964 415392 355970 415404
rect 580662 415392 580668 415404
rect 355964 415364 580668 415392
rect 355964 415352 355970 415364
rect 580662 415352 580668 415364
rect 580720 415352 580726 415404
rect 1600 415024 230496 415120
rect 350248 415024 583316 415120
rect 1600 414480 230496 414576
rect 350248 414480 583316 414576
rect 1600 413936 230496 414032
rect 350248 413936 583316 414032
rect 1600 413392 230496 413488
rect 350248 413392 583316 413488
rect 1600 412848 230496 412944
rect 350248 412848 583316 412944
rect 1600 412304 230496 412400
rect 350248 412304 583316 412400
rect 1600 411760 230496 411856
rect 350248 411760 583316 411856
rect 1600 411216 230496 411312
rect 350248 411216 583316 411312
rect 3822 411136 3828 411188
rect 3880 411176 3886 411188
rect 226186 411176 226192 411188
rect 3880 411148 226192 411176
rect 3880 411136 3886 411148
rect 226186 411136 226192 411148
rect 226244 411136 226250 411188
rect 1600 410672 230496 410768
rect 350248 410672 583316 410768
rect 1600 410128 230496 410224
rect 350248 410128 583316 410224
rect 1600 409584 230496 409680
rect 350248 409584 583316 409680
rect 1600 409040 230496 409136
rect 350248 409040 583316 409136
rect 1600 408496 230496 408592
rect 350248 408496 583316 408592
rect 1600 407952 230496 408048
rect 350248 407952 583316 408048
rect 1600 407408 230496 407504
rect 350248 407408 583316 407504
rect 1600 406864 230496 406960
rect 350248 406864 583316 406960
rect 1600 406320 230496 406416
rect 350248 406320 583316 406416
rect 1600 405776 230496 405872
rect 350248 405776 583316 405872
rect 1600 405232 230496 405328
rect 350248 405232 583316 405328
rect 1600 404688 230496 404784
rect 350248 404688 583316 404784
rect 1600 404144 230496 404240
rect 350248 404144 583316 404240
rect 1600 403600 230496 403696
rect 350248 403600 583316 403696
rect 1600 403056 230496 403152
rect 350248 403056 583316 403152
rect 1600 402512 230496 402608
rect 350248 402512 583316 402608
rect 1600 401968 230496 402064
rect 350248 401968 583316 402064
rect 1600 401424 230496 401520
rect 350248 401424 583316 401520
rect 1600 400880 230496 400976
rect 350248 400880 583316 400976
rect 1600 400336 230496 400432
rect 350248 400336 583316 400432
rect 358666 400120 358672 400172
rect 358724 400160 358730 400172
rect 580662 400160 580668 400172
rect 358724 400132 580668 400160
rect 358724 400120 358730 400132
rect 580662 400120 580668 400132
rect 580720 400120 580726 400172
rect 1600 399792 230496 399888
rect 350248 399792 583316 399888
rect 1600 399248 230496 399344
rect 350248 399248 583316 399344
rect 1600 398704 230496 398800
rect 350248 398704 583316 398800
rect 1600 398160 230496 398256
rect 350248 398160 583316 398256
rect 1600 397616 230496 397712
rect 350248 397616 583316 397712
rect 1600 397072 230496 397168
rect 350248 397072 583316 397168
rect 1600 396528 230496 396624
rect 350248 396528 583316 396624
rect 1600 395984 230496 396080
rect 350248 395984 583316 396080
rect 1600 395440 230496 395536
rect 350248 395440 583316 395536
rect 1600 394896 230496 394992
rect 350248 394896 583316 394992
rect 3822 394612 3828 394664
rect 3880 394652 3886 394664
rect 227566 394652 227572 394664
rect 3880 394624 227572 394652
rect 3880 394612 3886 394624
rect 227566 394612 227572 394624
rect 227624 394612 227630 394664
rect 1600 394352 230496 394448
rect 350248 394352 583316 394448
rect 1600 393808 230496 393904
rect 350248 393808 583316 393904
rect 1600 393264 230496 393360
rect 350248 393264 583316 393360
rect 1600 392720 230496 392816
rect 350248 392720 583316 392816
rect 1600 392176 230496 392272
rect 350248 392176 583316 392272
rect 1600 391632 230496 391728
rect 350248 391632 583316 391728
rect 1600 391088 230496 391184
rect 350248 391088 583316 391184
rect 1600 390544 230496 390640
rect 350248 390544 583316 390640
rect 1600 390000 230496 390096
rect 350248 390000 583316 390096
rect 1600 389456 230496 389552
rect 350248 389456 583316 389552
rect 1600 388912 230496 389008
rect 350248 388912 583316 389008
rect 1600 388368 230496 388464
rect 350248 388368 583316 388464
rect 1600 387824 230496 387920
rect 350248 387824 583316 387920
rect 1600 387280 230496 387376
rect 350248 387280 583316 387376
rect 1600 386736 230496 386832
rect 350248 386736 583316 386832
rect 1600 386192 230496 386288
rect 350248 386192 583316 386288
rect 1600 385648 230496 385744
rect 350248 385648 583316 385744
rect 1600 385104 230496 385200
rect 350248 385104 583316 385200
rect 1600 384560 230496 384656
rect 350248 384560 583316 384656
rect 1600 384016 230496 384112
rect 350248 384016 583316 384112
rect 406874 383596 406880 383648
rect 406932 383636 406938 383648
rect 580662 383636 580668 383648
rect 406932 383608 580668 383636
rect 406932 383596 406938 383608
rect 580662 383596 580668 383608
rect 580720 383596 580726 383648
rect 1600 383472 230496 383568
rect 350248 383472 583316 383568
rect 1600 382928 230496 383024
rect 350248 382928 583316 383024
rect 1600 382384 230496 382480
rect 350248 382384 583316 382480
rect 1600 381840 230496 381936
rect 350248 381840 583316 381936
rect 1600 381296 230496 381392
rect 350248 381296 583316 381392
rect 1600 380752 230496 380848
rect 350248 380752 583316 380848
rect 1600 380208 230496 380304
rect 350248 380208 583316 380304
rect 1600 379664 230496 379760
rect 350248 379664 583316 379760
rect 1600 379120 230496 379216
rect 350248 379120 583316 379216
rect 1600 378576 230496 378672
rect 350248 378576 583316 378672
rect 1600 378032 230496 378128
rect 350248 378032 583316 378128
rect 3546 377952 3552 378004
rect 3604 377992 3610 378004
rect 221954 377992 221960 378004
rect 3604 377964 221960 377992
rect 3604 377952 3610 377964
rect 221954 377952 221960 377964
rect 222012 377952 222018 378004
rect 1600 377488 230496 377584
rect 350248 377488 583316 377584
rect 1600 376944 230496 377040
rect 350248 376944 583316 377040
rect 1600 376400 230496 376496
rect 350248 376400 583316 376496
rect 1600 375856 230496 375952
rect 350248 375856 583316 375952
rect 1600 375312 230496 375408
rect 350248 375312 583316 375408
rect 1600 374768 230496 374864
rect 350248 374768 583316 374864
rect 1600 374224 230496 374320
rect 350248 374224 583316 374320
rect 1600 373680 230496 373776
rect 350248 373680 583316 373776
rect 1600 373136 230496 373232
rect 350248 373136 583316 373232
rect 1600 372592 230496 372688
rect 350248 372592 583316 372688
rect 1600 372048 230496 372144
rect 350248 372048 583316 372144
rect 1600 371504 230496 371600
rect 350248 371504 583316 371600
rect 1600 370960 230496 371056
rect 350248 370960 583316 371056
rect 1600 370416 230496 370512
rect 350248 370416 583316 370512
rect 1600 369872 230496 369968
rect 350248 369872 583316 369968
rect 1600 369328 230496 369424
rect 350248 369328 583316 369424
rect 1600 368784 230496 368880
rect 350248 368784 583316 368880
rect 354526 368432 354532 368484
rect 354584 368472 354590 368484
rect 580662 368472 580668 368484
rect 354584 368444 580668 368472
rect 354584 368432 354590 368444
rect 580662 368432 580668 368444
rect 580720 368432 580726 368484
rect 1600 368240 230496 368336
rect 350248 368240 583316 368336
rect 1600 367696 230496 367792
rect 350248 367696 583316 367792
rect 1600 367152 230496 367248
rect 350248 367152 583316 367248
rect 1600 366608 230496 366704
rect 350248 366608 583316 366704
rect 1600 366064 230496 366160
rect 350248 366064 583316 366160
rect 1600 365520 230496 365616
rect 350248 365520 583316 365616
rect 1600 364976 230496 365072
rect 350248 364976 583316 365072
rect 1600 364432 230496 364528
rect 350248 364432 583316 364528
rect 1600 363888 230496 363984
rect 350248 363888 583316 363984
rect 1600 363344 230496 363440
rect 350248 363344 583316 363440
rect 1600 362800 230496 362896
rect 350248 362800 583316 362896
rect 1600 362256 230496 362352
rect 350248 362256 583316 362352
rect 1600 361712 230496 361808
rect 350248 361712 583316 361808
rect 3822 361496 3828 361548
rect 3880 361536 3886 361548
rect 223334 361536 223340 361548
rect 3880 361508 223340 361536
rect 3880 361496 3886 361508
rect 223334 361496 223340 361508
rect 223392 361496 223398 361548
rect 1600 361168 230496 361264
rect 350248 361168 583316 361264
rect 1600 360624 230496 360720
rect 350248 360624 583316 360720
rect 1600 360080 230496 360176
rect 350248 360080 583316 360176
rect 1600 359536 230496 359632
rect 350248 359536 583316 359632
rect 1600 358992 230496 359088
rect 350248 358992 583316 359088
rect 1600 358448 230496 358544
rect 350248 358448 583316 358544
rect 1600 357904 230496 358000
rect 350248 357904 583316 358000
rect 1600 357360 230496 357456
rect 350248 357360 583316 357456
rect 1600 356816 230496 356912
rect 350248 356816 583316 356912
rect 1600 356272 230496 356368
rect 350248 356272 583316 356368
rect 1600 355728 230496 355824
rect 350248 355728 583316 355824
rect 1600 355184 230496 355280
rect 350248 355184 583316 355280
rect 1600 354640 230496 354736
rect 350248 354640 583316 354736
rect 1600 354096 230496 354192
rect 350248 354096 583316 354192
rect 1600 353552 230496 353648
rect 350248 353552 583316 353648
rect 357194 353200 357200 353252
rect 357252 353240 357258 353252
rect 580662 353240 580668 353252
rect 357252 353212 580668 353240
rect 357252 353200 357258 353212
rect 580662 353200 580668 353212
rect 580720 353200 580726 353252
rect 1600 353008 230496 353104
rect 350248 353008 583316 353104
rect 1600 352464 230496 352560
rect 350248 352464 583316 352560
rect 1600 351920 230496 352016
rect 350248 351920 583316 352016
rect 1600 351376 230496 351472
rect 350248 351376 583316 351472
rect 1600 350832 230496 350928
rect 350248 350832 583316 350928
rect 1600 350288 230496 350384
rect 350248 350288 583316 350384
rect 1600 349744 230496 349840
rect 350248 349744 583316 349840
rect 1600 349200 230496 349296
rect 350248 349200 583316 349296
rect 1600 348656 230496 348752
rect 350248 348656 583316 348752
rect 1600 348112 230496 348208
rect 350248 348112 583316 348208
rect 1600 347568 230496 347664
rect 350248 347568 583316 347664
rect 1600 347024 230496 347120
rect 350248 347024 583316 347120
rect 1600 346480 230496 346576
rect 350248 346480 583316 346576
rect 1600 345936 230496 346032
rect 350248 345936 583316 346032
rect 1600 345392 230496 345488
rect 350248 345392 583316 345488
rect 1600 344848 230496 344944
rect 350248 344848 583316 344944
rect 1600 344304 230496 344400
rect 350248 344304 583316 344400
rect 1600 343760 230496 343856
rect 350248 343760 583316 343856
rect 3822 343544 3828 343596
rect 3880 343584 3886 343596
rect 228946 343584 228952 343596
rect 3880 343556 228952 343584
rect 3880 343544 3886 343556
rect 228946 343544 228952 343556
rect 229004 343544 229010 343596
rect 1600 343216 230496 343312
rect 350248 343216 583316 343312
rect 1600 342672 230496 342768
rect 350248 342672 583316 342768
rect 1600 342128 230496 342224
rect 350248 342128 583316 342224
rect 1600 341584 230496 341680
rect 350248 341584 583316 341680
rect 1600 341040 230496 341136
rect 350248 341040 583316 341136
rect 1600 340496 230496 340592
rect 350248 340496 583316 340592
rect 1600 339952 583316 340048
rect 1600 339408 583316 339504
rect 240906 339056 240912 339108
rect 240964 339096 240970 339108
rect 241274 339096 241280 339108
rect 240964 339068 241280 339096
rect 240964 339056 240970 339068
rect 241274 339056 241280 339068
rect 241332 339056 241338 339108
rect 242102 339056 242108 339108
rect 242160 339096 242166 339108
rect 242470 339096 242476 339108
rect 242160 339068 242476 339096
rect 242160 339056 242166 339068
rect 242470 339056 242476 339068
rect 242528 339056 242534 339108
rect 268230 339056 268236 339108
rect 268288 339096 268294 339108
rect 268690 339096 268696 339108
rect 268288 339068 268696 339096
rect 268288 339056 268294 339068
rect 268690 339056 268696 339068
rect 268748 339056 268754 339108
rect 1600 338864 583316 338960
rect 254798 338512 254804 338564
rect 254856 338552 254862 338564
rect 255166 338552 255172 338564
rect 254856 338524 255172 338552
rect 254856 338512 254862 338524
rect 255166 338512 255172 338524
rect 255224 338512 255230 338564
rect 272646 338444 272652 338496
rect 272704 338484 272710 338496
rect 273106 338484 273112 338496
rect 272704 338456 273112 338484
rect 272704 338444 272710 338456
rect 273106 338444 273112 338456
rect 273164 338444 273170 338496
rect 278902 338444 278908 338496
rect 278960 338484 278966 338496
rect 279178 338484 279184 338496
rect 278960 338456 279184 338484
rect 278960 338444 278966 338456
rect 279178 338444 279184 338456
rect 279236 338444 279242 338496
rect 1600 338320 583316 338416
rect 119193 338283 119251 338289
rect 119193 338249 119205 338283
rect 119239 338280 119251 338283
rect 230145 338283 230203 338289
rect 119239 338252 128804 338280
rect 119239 338249 119251 338252
rect 119193 338243 119251 338249
rect 113673 338147 113731 338153
rect 113673 338113 113685 338147
rect 113719 338144 113731 338147
rect 119285 338147 119343 338153
rect 119285 338144 119297 338147
rect 113719 338116 119297 338144
rect 113719 338113 113731 338116
rect 113673 338107 113731 338113
rect 119285 338113 119297 338116
rect 119331 338113 119343 338147
rect 128776 338144 128804 338252
rect 230145 338249 230157 338283
rect 230191 338280 230203 338283
rect 234745 338283 234803 338289
rect 234745 338280 234757 338283
rect 230191 338252 234757 338280
rect 230191 338249 230203 338252
rect 230145 338243 230203 338249
rect 234745 338249 234757 338252
rect 234791 338249 234803 338283
rect 234745 338243 234803 338249
rect 128945 338215 129003 338221
rect 128945 338181 128957 338215
rect 128991 338212 129003 338215
rect 138329 338215 138387 338221
rect 138329 338212 138341 338215
rect 128991 338184 138341 338212
rect 128991 338181 129003 338184
rect 128945 338175 129003 338181
rect 138329 338181 138341 338184
rect 138375 338181 138387 338215
rect 138329 338175 138387 338181
rect 225453 338215 225511 338221
rect 225453 338181 225465 338215
rect 225499 338212 225511 338215
rect 234190 338212 234196 338224
rect 225499 338184 234196 338212
rect 225499 338181 225511 338184
rect 225453 338175 225511 338181
rect 234190 338172 234196 338184
rect 234248 338172 234254 338224
rect 129218 338144 129224 338156
rect 128776 338116 129224 338144
rect 119285 338107 119343 338113
rect 129218 338104 129224 338116
rect 129276 338104 129282 338156
rect 129405 338147 129463 338153
rect 129405 338113 129417 338147
rect 129451 338144 129463 338147
rect 142558 338144 142564 338156
rect 129451 338116 142564 338144
rect 129451 338113 129463 338116
rect 129405 338107 129463 338113
rect 142558 338104 142564 338116
rect 142616 338104 142622 338156
rect 142653 338147 142711 338153
rect 142653 338113 142665 338147
rect 142699 338144 142711 338147
rect 152218 338144 152224 338156
rect 142699 338116 152224 338144
rect 142699 338113 142711 338116
rect 142653 338107 142711 338113
rect 152218 338104 152224 338116
rect 152276 338104 152282 338156
rect 152313 338147 152371 338153
rect 152313 338113 152325 338147
rect 152359 338144 152371 338147
rect 161878 338144 161884 338156
rect 152359 338116 161884 338144
rect 152359 338113 152371 338116
rect 152313 338107 152371 338113
rect 161878 338104 161884 338116
rect 161936 338104 161942 338156
rect 161973 338147 162031 338153
rect 161973 338113 161985 338147
rect 162019 338144 162031 338147
rect 171538 338144 171544 338156
rect 162019 338116 171544 338144
rect 162019 338113 162031 338116
rect 161973 338107 162031 338113
rect 171538 338104 171544 338116
rect 171596 338104 171602 338156
rect 171633 338147 171691 338153
rect 171633 338113 171645 338147
rect 171679 338144 171691 338147
rect 181198 338144 181204 338156
rect 171679 338116 181204 338144
rect 171679 338113 171691 338116
rect 171633 338107 171691 338113
rect 181198 338104 181204 338116
rect 181256 338104 181262 338156
rect 181293 338147 181351 338153
rect 181293 338113 181305 338147
rect 181339 338144 181351 338147
rect 190858 338144 190864 338156
rect 181339 338116 190864 338144
rect 181339 338113 181351 338116
rect 181293 338107 181351 338113
rect 190858 338104 190864 338116
rect 190916 338104 190922 338156
rect 190953 338147 191011 338153
rect 190953 338113 190965 338147
rect 190999 338144 191011 338147
rect 200518 338144 200524 338156
rect 190999 338116 200524 338144
rect 190999 338113 191011 338116
rect 190953 338107 191011 338113
rect 200518 338104 200524 338116
rect 200576 338104 200582 338156
rect 200613 338147 200671 338153
rect 200613 338113 200625 338147
rect 200659 338144 200671 338147
rect 210178 338144 210184 338156
rect 200659 338116 210184 338144
rect 200659 338113 200671 338116
rect 200613 338107 200671 338113
rect 210178 338104 210184 338116
rect 210236 338104 210242 338156
rect 210273 338147 210331 338153
rect 210273 338113 210285 338147
rect 210319 338144 210331 338147
rect 219838 338144 219844 338156
rect 210319 338116 219844 338144
rect 210319 338113 210331 338116
rect 210273 338107 210331 338113
rect 219838 338104 219844 338116
rect 219896 338104 219902 338156
rect 219933 338147 219991 338153
rect 219933 338113 219945 338147
rect 219979 338144 219991 338147
rect 225545 338147 225603 338153
rect 225545 338144 225557 338147
rect 219979 338116 225557 338144
rect 219979 338113 219991 338116
rect 219933 338107 219991 338113
rect 225545 338113 225557 338116
rect 225591 338113 225603 338147
rect 225545 338107 225603 338113
rect 226741 338147 226799 338153
rect 226741 338113 226753 338147
rect 226787 338144 226799 338147
rect 232350 338144 232356 338156
rect 226787 338116 232356 338144
rect 226787 338113 226799 338116
rect 226741 338107 226799 338113
rect 232350 338104 232356 338116
rect 232408 338104 232414 338156
rect 308894 338104 308900 338156
rect 308952 338144 308958 338156
rect 309538 338144 309544 338156
rect 308952 338116 309544 338144
rect 308952 338104 308958 338116
rect 309538 338104 309544 338116
rect 309596 338104 309602 338156
rect 62518 338036 62524 338088
rect 62576 338076 62582 338088
rect 242930 338076 242936 338088
rect 62576 338048 242936 338076
rect 62576 338036 62582 338048
rect 242930 338036 242936 338048
rect 242988 338036 242994 338088
rect 259125 338079 259183 338085
rect 259125 338045 259137 338079
rect 259171 338076 259183 338079
rect 259214 338076 259220 338088
rect 259171 338048 259220 338076
rect 259171 338045 259183 338048
rect 259125 338039 259183 338045
rect 259214 338036 259220 338048
rect 259272 338036 259278 338088
rect 278537 338079 278595 338085
rect 278537 338045 278549 338079
rect 278583 338076 278595 338079
rect 283870 338076 283876 338088
rect 278583 338048 283876 338076
rect 278583 338045 278595 338048
rect 278537 338039 278595 338045
rect 283870 338036 283876 338048
rect 283928 338036 283934 338088
rect 303926 338036 303932 338088
rect 303984 338076 303990 338088
rect 356550 338076 356556 338088
rect 303984 338048 356556 338076
rect 303984 338036 303990 338048
rect 356550 338036 356556 338048
rect 356608 338036 356614 338088
rect 36393 338011 36451 338017
rect 36393 337977 36405 338011
rect 36439 338008 36451 338011
rect 45958 338008 45964 338020
rect 36439 337980 45964 338008
rect 36439 337977 36451 337980
rect 36393 337971 36451 337977
rect 45958 337968 45964 337980
rect 46016 337968 46022 338020
rect 55618 337968 55624 338020
rect 55676 338008 55682 338020
rect 230145 338011 230203 338017
rect 230145 338008 230157 338011
rect 55676 337980 230157 338008
rect 55676 337968 55682 337980
rect 230145 337977 230157 337980
rect 230191 337977 230203 338011
rect 230145 337971 230203 337977
rect 230237 338011 230295 338017
rect 230237 337977 230249 338011
rect 230283 338008 230295 338011
rect 236306 338008 236312 338020
rect 230283 337980 236312 338008
rect 230283 337977 230295 337980
rect 230237 337971 230295 337977
rect 236306 337968 236312 337980
rect 236364 337968 236370 338020
rect 280653 338011 280711 338017
rect 280653 338008 280665 338011
rect 270916 337980 280665 338008
rect 26733 337943 26791 337949
rect 26733 337909 26745 337943
rect 26779 337940 26791 337943
rect 36301 337943 36359 337949
rect 36301 337940 36313 337943
rect 26779 337912 36313 337940
rect 26779 337909 26791 337912
rect 26733 337903 26791 337909
rect 36301 337909 36313 337912
rect 36347 337909 36359 337943
rect 36301 337903 36359 337909
rect 44578 337900 44584 337952
rect 44636 337940 44642 337952
rect 129405 337943 129463 337949
rect 129405 337940 129417 337943
rect 44636 337912 129417 337940
rect 44636 337900 44642 337912
rect 129405 337909 129417 337912
rect 129451 337909 129463 337943
rect 129405 337903 129463 337909
rect 129497 337943 129555 337949
rect 129497 337909 129509 337943
rect 129543 337940 129555 337943
rect 142469 337943 142527 337949
rect 142469 337940 142481 337943
rect 129543 337912 142481 337940
rect 129543 337909 129555 337912
rect 129497 337903 129555 337909
rect 142469 337909 142481 337912
rect 142515 337909 142527 337943
rect 142469 337903 142527 337909
rect 142558 337900 142564 337952
rect 142616 337940 142622 337952
rect 142653 337943 142711 337949
rect 142653 337940 142665 337943
rect 142616 337912 142665 337940
rect 142616 337900 142622 337912
rect 142653 337909 142665 337912
rect 142699 337909 142711 337943
rect 142653 337903 142711 337909
rect 142745 337943 142803 337949
rect 142745 337909 142757 337943
rect 142791 337940 142803 337943
rect 152129 337943 152187 337949
rect 152129 337940 152141 337943
rect 142791 337912 152141 337940
rect 142791 337909 142803 337912
rect 142745 337903 142803 337909
rect 152129 337909 152141 337912
rect 152175 337909 152187 337943
rect 152129 337903 152187 337909
rect 152218 337900 152224 337952
rect 152276 337940 152282 337952
rect 152313 337943 152371 337949
rect 152313 337940 152325 337943
rect 152276 337912 152325 337940
rect 152276 337900 152282 337912
rect 152313 337909 152325 337912
rect 152359 337909 152371 337943
rect 152313 337903 152371 337909
rect 152405 337943 152463 337949
rect 152405 337909 152417 337943
rect 152451 337940 152463 337943
rect 161789 337943 161847 337949
rect 161789 337940 161801 337943
rect 152451 337912 161801 337940
rect 152451 337909 152463 337912
rect 152405 337903 152463 337909
rect 161789 337909 161801 337912
rect 161835 337909 161847 337943
rect 161789 337903 161847 337909
rect 161878 337900 161884 337952
rect 161936 337940 161942 337952
rect 161973 337943 162031 337949
rect 161973 337940 161985 337943
rect 161936 337912 161985 337940
rect 161936 337900 161942 337912
rect 161973 337909 161985 337912
rect 162019 337909 162031 337943
rect 161973 337903 162031 337909
rect 162065 337943 162123 337949
rect 162065 337909 162077 337943
rect 162111 337940 162123 337943
rect 171449 337943 171507 337949
rect 171449 337940 171461 337943
rect 162111 337912 171461 337940
rect 162111 337909 162123 337912
rect 162065 337903 162123 337909
rect 171449 337909 171461 337912
rect 171495 337909 171507 337943
rect 171449 337903 171507 337909
rect 171538 337900 171544 337952
rect 171596 337940 171602 337952
rect 171633 337943 171691 337949
rect 171633 337940 171645 337943
rect 171596 337912 171645 337940
rect 171596 337900 171602 337912
rect 171633 337909 171645 337912
rect 171679 337909 171691 337943
rect 171633 337903 171691 337909
rect 171725 337943 171783 337949
rect 171725 337909 171737 337943
rect 171771 337940 171783 337943
rect 181109 337943 181167 337949
rect 181109 337940 181121 337943
rect 171771 337912 181121 337940
rect 171771 337909 171783 337912
rect 171725 337903 171783 337909
rect 181109 337909 181121 337912
rect 181155 337909 181167 337943
rect 181109 337903 181167 337909
rect 181198 337900 181204 337952
rect 181256 337940 181262 337952
rect 181293 337943 181351 337949
rect 181293 337940 181305 337943
rect 181256 337912 181305 337940
rect 181256 337900 181262 337912
rect 181293 337909 181305 337912
rect 181339 337909 181351 337943
rect 181293 337903 181351 337909
rect 181385 337943 181443 337949
rect 181385 337909 181397 337943
rect 181431 337940 181443 337943
rect 190769 337943 190827 337949
rect 190769 337940 190781 337943
rect 181431 337912 190781 337940
rect 181431 337909 181443 337912
rect 181385 337903 181443 337909
rect 190769 337909 190781 337912
rect 190815 337909 190827 337943
rect 190769 337903 190827 337909
rect 190858 337900 190864 337952
rect 190916 337940 190922 337952
rect 190953 337943 191011 337949
rect 190953 337940 190965 337943
rect 190916 337912 190965 337940
rect 190916 337900 190922 337912
rect 190953 337909 190965 337912
rect 190999 337909 191011 337943
rect 190953 337903 191011 337909
rect 191045 337943 191103 337949
rect 191045 337909 191057 337943
rect 191091 337940 191103 337943
rect 200429 337943 200487 337949
rect 200429 337940 200441 337943
rect 191091 337912 200441 337940
rect 191091 337909 191103 337912
rect 191045 337903 191103 337909
rect 200429 337909 200441 337912
rect 200475 337909 200487 337943
rect 200429 337903 200487 337909
rect 200518 337900 200524 337952
rect 200576 337940 200582 337952
rect 200613 337943 200671 337949
rect 200613 337940 200625 337943
rect 200576 337912 200625 337940
rect 200576 337900 200582 337912
rect 200613 337909 200625 337912
rect 200659 337909 200671 337943
rect 200613 337903 200671 337909
rect 200705 337943 200763 337949
rect 200705 337909 200717 337943
rect 200751 337940 200763 337943
rect 210089 337943 210147 337949
rect 210089 337940 210101 337943
rect 200751 337912 210101 337940
rect 200751 337909 200763 337912
rect 200705 337903 200763 337909
rect 210089 337909 210101 337912
rect 210135 337909 210147 337943
rect 210089 337903 210147 337909
rect 210178 337900 210184 337952
rect 210236 337940 210242 337952
rect 210273 337943 210331 337949
rect 210273 337940 210285 337943
rect 210236 337912 210285 337940
rect 210236 337900 210242 337912
rect 210273 337909 210285 337912
rect 210319 337909 210331 337943
rect 210273 337903 210331 337909
rect 210365 337943 210423 337949
rect 210365 337909 210377 337943
rect 210411 337940 210423 337943
rect 219749 337943 219807 337949
rect 219749 337940 219761 337943
rect 210411 337912 219761 337940
rect 210411 337909 210423 337912
rect 210365 337903 210423 337909
rect 219749 337909 219761 337912
rect 219795 337909 219807 337943
rect 219749 337903 219807 337909
rect 219838 337900 219844 337952
rect 219896 337940 219902 337952
rect 219933 337943 219991 337949
rect 219933 337940 219945 337943
rect 219896 337912 219945 337940
rect 219896 337900 219902 337912
rect 219933 337909 219945 337912
rect 219979 337909 219991 337943
rect 219933 337903 219991 337909
rect 220025 337943 220083 337949
rect 220025 337909 220037 337943
rect 220071 337940 220083 337943
rect 237778 337940 237784 337952
rect 220071 337912 237784 337940
rect 220071 337909 220083 337912
rect 220025 337903 220083 337909
rect 237778 337900 237784 337912
rect 237836 337900 237842 337952
rect 270916 337949 270944 337980
rect 280653 337977 280665 337980
rect 280699 337977 280711 338011
rect 280653 337971 280711 337977
rect 292610 337968 292616 338020
rect 292668 338008 292674 338020
rect 293806 338008 293812 338020
rect 292668 337980 293812 338008
rect 292668 337968 292674 337980
rect 293806 337968 293812 337980
rect 293864 337968 293870 338020
rect 297302 337968 297308 338020
rect 297360 338008 297366 338020
rect 304754 338008 304760 338020
rect 297360 337980 304760 338008
rect 297360 337968 297366 337980
rect 304754 337968 304760 337980
rect 304812 337968 304818 338020
rect 305398 337968 305404 338020
rect 305456 338008 305462 338020
rect 364830 338008 364836 338020
rect 305456 337980 364836 338008
rect 305456 337968 305462 337980
rect 364830 337968 364836 337980
rect 364888 337968 364894 338020
rect 270901 337943 270959 337949
rect 270901 337909 270913 337943
rect 270947 337909 270959 337943
rect 270901 337903 270959 337909
rect 298222 337900 298228 337952
rect 298280 337940 298286 337952
rect 298498 337940 298504 337952
rect 298280 337912 298504 337940
rect 298280 337900 298286 337912
rect 298498 337900 298504 337912
rect 298556 337900 298562 337952
rect 300246 337900 300252 337952
rect 300304 337940 300310 337952
rect 303466 337940 303472 337952
rect 300304 337912 303472 337940
rect 300304 337900 300310 337912
rect 303466 337900 303472 337912
rect 303524 337900 303530 337952
rect 304938 337900 304944 337952
rect 304996 337940 305002 337952
rect 305122 337940 305128 337952
rect 304996 337912 305128 337940
rect 304996 337900 305002 337912
rect 305122 337900 305128 337912
rect 305180 337900 305186 337952
rect 309078 337900 309084 337952
rect 309136 337940 309142 337952
rect 309538 337940 309544 337952
rect 309136 337912 309544 337940
rect 309136 337900 309142 337912
rect 309538 337900 309544 337912
rect 309596 337900 309602 337952
rect 317177 337943 317235 337949
rect 317177 337909 317189 337943
rect 317223 337940 317235 337943
rect 371917 337943 371975 337949
rect 371917 337940 371929 337943
rect 317223 337912 371929 337940
rect 317223 337909 317235 337912
rect 317177 337903 317235 337909
rect 371917 337909 371929 337912
rect 371963 337909 371975 337943
rect 371917 337903 371975 337909
rect 1600 337776 583316 337872
rect 22498 337696 22504 337748
rect 22556 337736 22562 337748
rect 26733 337739 26791 337745
rect 26733 337736 26745 337739
rect 22556 337708 26745 337736
rect 22556 337696 22562 337708
rect 26733 337705 26745 337708
rect 26779 337705 26791 337739
rect 26733 337699 26791 337705
rect 37678 337696 37684 337748
rect 37736 337736 37742 337748
rect 129497 337739 129555 337745
rect 129497 337736 129509 337739
rect 37736 337708 129509 337736
rect 37736 337696 37742 337708
rect 129497 337705 129509 337708
rect 129543 337705 129555 337739
rect 142561 337739 142619 337745
rect 129497 337699 129555 337705
rect 130248 337708 142512 337736
rect 30778 337628 30784 337680
rect 30836 337668 30842 337680
rect 130248 337668 130276 337708
rect 138326 337668 138332 337680
rect 30836 337640 130276 337668
rect 130340 337640 138332 337668
rect 30836 337628 30842 337640
rect 36301 337603 36359 337609
rect 36301 337569 36313 337603
rect 36347 337600 36359 337603
rect 36393 337603 36451 337609
rect 36393 337600 36405 337603
rect 36347 337572 36405 337600
rect 36347 337569 36359 337572
rect 36301 337563 36359 337569
rect 36393 337569 36405 337572
rect 36439 337569 36451 337603
rect 36393 337563 36451 337569
rect 45958 337560 45964 337612
rect 46016 337600 46022 337612
rect 55713 337603 55771 337609
rect 55713 337600 55725 337603
rect 46016 337572 55725 337600
rect 46016 337560 46022 337572
rect 55713 337569 55725 337572
rect 55759 337569 55771 337603
rect 55713 337563 55771 337569
rect 65278 337560 65284 337612
rect 65336 337600 65342 337612
rect 75033 337603 75091 337609
rect 75033 337600 75045 337603
rect 65336 337572 75045 337600
rect 65336 337560 65342 337572
rect 75033 337569 75045 337572
rect 75079 337569 75091 337603
rect 75033 337563 75091 337569
rect 84598 337560 84604 337612
rect 84656 337600 84662 337612
rect 94353 337603 94411 337609
rect 94353 337600 94365 337603
rect 84656 337572 94365 337600
rect 84656 337560 84662 337572
rect 94353 337569 94365 337572
rect 94399 337569 94411 337603
rect 94353 337563 94411 337569
rect 103829 337603 103887 337609
rect 103829 337569 103841 337603
rect 103875 337600 103887 337603
rect 113673 337603 113731 337609
rect 113673 337600 113685 337603
rect 103875 337572 113685 337600
rect 103875 337569 103887 337572
rect 103829 337563 103887 337569
rect 113673 337569 113685 337572
rect 113719 337569 113731 337603
rect 113673 337563 113731 337569
rect 113765 337603 113823 337609
rect 113765 337569 113777 337603
rect 113811 337600 113823 337603
rect 123977 337603 124035 337609
rect 123977 337600 123989 337603
rect 113811 337572 123989 337600
rect 113811 337569 113823 337572
rect 113765 337563 113823 337569
rect 123977 337569 123989 337572
rect 124023 337569 124035 337603
rect 123977 337563 124035 337569
rect 125998 337560 126004 337612
rect 126056 337600 126062 337612
rect 126056 337572 128712 337600
rect 126056 337560 126062 337572
rect 12838 337492 12844 337544
rect 12896 337532 12902 337544
rect 116249 337535 116307 337541
rect 116249 337532 116261 337535
rect 12896 337504 116261 337532
rect 12896 337492 12902 337504
rect 116249 337501 116261 337504
rect 116295 337501 116307 337535
rect 116249 337495 116307 337501
rect 116338 337492 116344 337544
rect 116396 337532 116402 337544
rect 128574 337532 128580 337544
rect 116396 337504 128580 337532
rect 116396 337492 116402 337504
rect 128574 337492 128580 337504
rect 128632 337492 128638 337544
rect 128684 337532 128712 337572
rect 128758 337560 128764 337612
rect 128816 337600 128822 337612
rect 128945 337603 129003 337609
rect 128945 337600 128957 337603
rect 128816 337572 128957 337600
rect 128816 337560 128822 337572
rect 128945 337569 128957 337572
rect 128991 337569 129003 337603
rect 128945 337563 129003 337569
rect 129034 337560 129040 337612
rect 129092 337600 129098 337612
rect 130340 337600 130368 337640
rect 138326 337628 138332 337640
rect 138384 337628 138390 337680
rect 138418 337628 138424 337680
rect 138476 337668 138482 337680
rect 142377 337671 142435 337677
rect 142377 337668 142389 337671
rect 138476 337640 142389 337668
rect 138476 337628 138482 337640
rect 142377 337637 142389 337640
rect 142423 337637 142435 337671
rect 142484 337668 142512 337708
rect 142561 337705 142573 337739
rect 142607 337736 142619 337739
rect 142653 337739 142711 337745
rect 142653 337736 142665 337739
rect 142607 337708 142665 337736
rect 142607 337705 142619 337708
rect 142561 337699 142619 337705
rect 142653 337705 142665 337708
rect 142699 337705 142711 337739
rect 152221 337739 152279 337745
rect 142653 337699 142711 337705
rect 142760 337708 152172 337736
rect 142760 337668 142788 337708
rect 142484 337640 142788 337668
rect 142837 337671 142895 337677
rect 142377 337631 142435 337637
rect 142837 337637 142849 337671
rect 142883 337668 142895 337671
rect 152037 337671 152095 337677
rect 152037 337668 152049 337671
rect 142883 337640 152049 337668
rect 142883 337637 142895 337640
rect 142837 337631 142895 337637
rect 152037 337637 152049 337640
rect 152083 337637 152095 337671
rect 152144 337668 152172 337708
rect 152221 337705 152233 337739
rect 152267 337736 152279 337739
rect 152313 337739 152371 337745
rect 152313 337736 152325 337739
rect 152267 337708 152325 337736
rect 152267 337705 152279 337708
rect 152221 337699 152279 337705
rect 152313 337705 152325 337708
rect 152359 337705 152371 337739
rect 161881 337739 161939 337745
rect 152313 337699 152371 337705
rect 152420 337708 161832 337736
rect 152420 337668 152448 337708
rect 152144 337640 152448 337668
rect 152497 337671 152555 337677
rect 152037 337631 152095 337637
rect 152497 337637 152509 337671
rect 152543 337668 152555 337671
rect 161697 337671 161755 337677
rect 161697 337668 161709 337671
rect 152543 337640 161709 337668
rect 152543 337637 152555 337640
rect 152497 337631 152555 337637
rect 161697 337637 161709 337640
rect 161743 337637 161755 337671
rect 161804 337668 161832 337708
rect 161881 337705 161893 337739
rect 161927 337736 161939 337739
rect 161973 337739 162031 337745
rect 161973 337736 161985 337739
rect 161927 337708 161985 337736
rect 161927 337705 161939 337708
rect 161881 337699 161939 337705
rect 161973 337705 161985 337708
rect 162019 337705 162031 337739
rect 171541 337739 171599 337745
rect 161973 337699 162031 337705
rect 162080 337708 171492 337736
rect 162080 337668 162108 337708
rect 161804 337640 162108 337668
rect 162157 337671 162215 337677
rect 161697 337631 161755 337637
rect 162157 337637 162169 337671
rect 162203 337668 162215 337671
rect 171357 337671 171415 337677
rect 171357 337668 171369 337671
rect 162203 337640 171369 337668
rect 162203 337637 162215 337640
rect 162157 337631 162215 337637
rect 171357 337637 171369 337640
rect 171403 337637 171415 337671
rect 171464 337668 171492 337708
rect 171541 337705 171553 337739
rect 171587 337736 171599 337739
rect 171633 337739 171691 337745
rect 171633 337736 171645 337739
rect 171587 337708 171645 337736
rect 171587 337705 171599 337708
rect 171541 337699 171599 337705
rect 171633 337705 171645 337708
rect 171679 337705 171691 337739
rect 181201 337739 181259 337745
rect 171633 337699 171691 337705
rect 171740 337708 181152 337736
rect 171740 337668 171768 337708
rect 171464 337640 171768 337668
rect 171817 337671 171875 337677
rect 171357 337631 171415 337637
rect 171817 337637 171829 337671
rect 171863 337668 171875 337671
rect 181017 337671 181075 337677
rect 181017 337668 181029 337671
rect 171863 337640 181029 337668
rect 171863 337637 171875 337640
rect 171817 337631 171875 337637
rect 181017 337637 181029 337640
rect 181063 337637 181075 337671
rect 181124 337668 181152 337708
rect 181201 337705 181213 337739
rect 181247 337736 181259 337739
rect 181293 337739 181351 337745
rect 181293 337736 181305 337739
rect 181247 337708 181305 337736
rect 181247 337705 181259 337708
rect 181201 337699 181259 337705
rect 181293 337705 181305 337708
rect 181339 337705 181351 337739
rect 190861 337739 190919 337745
rect 181293 337699 181351 337705
rect 181400 337708 190812 337736
rect 181400 337668 181428 337708
rect 181124 337640 181428 337668
rect 181477 337671 181535 337677
rect 181017 337631 181075 337637
rect 181477 337637 181489 337671
rect 181523 337668 181535 337671
rect 190677 337671 190735 337677
rect 190677 337668 190689 337671
rect 181523 337640 190689 337668
rect 181523 337637 181535 337640
rect 181477 337631 181535 337637
rect 190677 337637 190689 337640
rect 190723 337637 190735 337671
rect 190784 337668 190812 337708
rect 190861 337705 190873 337739
rect 190907 337736 190919 337739
rect 190953 337739 191011 337745
rect 190953 337736 190965 337739
rect 190907 337708 190965 337736
rect 190907 337705 190919 337708
rect 190861 337699 190919 337705
rect 190953 337705 190965 337708
rect 190999 337705 191011 337739
rect 200521 337739 200579 337745
rect 190953 337699 191011 337705
rect 191060 337708 200472 337736
rect 191060 337668 191088 337708
rect 190784 337640 191088 337668
rect 191137 337671 191195 337677
rect 190677 337631 190735 337637
rect 191137 337637 191149 337671
rect 191183 337668 191195 337671
rect 200337 337671 200395 337677
rect 200337 337668 200349 337671
rect 191183 337640 200349 337668
rect 191183 337637 191195 337640
rect 191137 337631 191195 337637
rect 200337 337637 200349 337640
rect 200383 337637 200395 337671
rect 200444 337668 200472 337708
rect 200521 337705 200533 337739
rect 200567 337736 200579 337739
rect 200613 337739 200671 337745
rect 200613 337736 200625 337739
rect 200567 337708 200625 337736
rect 200567 337705 200579 337708
rect 200521 337699 200579 337705
rect 200613 337705 200625 337708
rect 200659 337705 200671 337739
rect 210181 337739 210239 337745
rect 200613 337699 200671 337705
rect 200720 337708 210132 337736
rect 200720 337668 200748 337708
rect 200444 337640 200748 337668
rect 200797 337671 200855 337677
rect 200337 337631 200395 337637
rect 200797 337637 200809 337671
rect 200843 337668 200855 337671
rect 209997 337671 210055 337677
rect 209997 337668 210009 337671
rect 200843 337640 210009 337668
rect 200843 337637 200855 337640
rect 200797 337631 200855 337637
rect 209997 337637 210009 337640
rect 210043 337637 210055 337671
rect 210104 337668 210132 337708
rect 210181 337705 210193 337739
rect 210227 337736 210239 337739
rect 210273 337739 210331 337745
rect 210273 337736 210285 337739
rect 210227 337708 210285 337736
rect 210227 337705 210239 337708
rect 210181 337699 210239 337705
rect 210273 337705 210285 337708
rect 210319 337705 210331 337739
rect 219841 337739 219899 337745
rect 210273 337699 210331 337705
rect 210380 337708 219792 337736
rect 210380 337668 210408 337708
rect 210104 337640 210408 337668
rect 210457 337671 210515 337677
rect 209997 337631 210055 337637
rect 210457 337637 210469 337671
rect 210503 337668 210515 337671
rect 219657 337671 219715 337677
rect 219657 337668 219669 337671
rect 210503 337640 219669 337668
rect 210503 337637 210515 337640
rect 210457 337631 210515 337637
rect 219657 337637 219669 337640
rect 219703 337637 219715 337671
rect 219764 337668 219792 337708
rect 219841 337705 219853 337739
rect 219887 337736 219899 337739
rect 219933 337739 219991 337745
rect 219933 337736 219945 337739
rect 219887 337708 219945 337736
rect 219887 337705 219899 337708
rect 219841 337699 219899 337705
rect 219933 337705 219945 337708
rect 219979 337705 219991 337739
rect 230237 337739 230295 337745
rect 230237 337736 230249 337739
rect 219933 337699 219991 337705
rect 220040 337708 230249 337736
rect 220040 337668 220068 337708
rect 230237 337705 230249 337708
rect 230283 337705 230295 337739
rect 230237 337699 230295 337705
rect 230329 337739 230387 337745
rect 230329 337705 230341 337739
rect 230375 337736 230387 337739
rect 232626 337736 232632 337748
rect 230375 337708 232632 337736
rect 230375 337705 230387 337708
rect 230329 337699 230387 337705
rect 232626 337696 232632 337708
rect 232684 337696 232690 337748
rect 232810 337696 232816 337748
rect 232868 337736 232874 337748
rect 234650 337736 234656 337748
rect 232868 337708 234656 337736
rect 232868 337696 232874 337708
rect 234650 337696 234656 337708
rect 234708 337696 234714 337748
rect 234745 337739 234803 337745
rect 234745 337705 234757 337739
rect 234791 337736 234803 337739
rect 241458 337736 241464 337748
rect 234791 337708 241464 337736
rect 234791 337705 234803 337708
rect 234745 337699 234803 337705
rect 241458 337696 241464 337708
rect 241516 337696 241522 337748
rect 264734 337696 264740 337748
rect 264792 337736 264798 337748
rect 280650 337736 280656 337748
rect 264792 337708 280656 337736
rect 264792 337696 264798 337708
rect 280650 337696 280656 337708
rect 280708 337696 280714 337748
rect 280745 337739 280803 337745
rect 280745 337705 280757 337739
rect 280791 337736 280803 337739
rect 284054 337736 284060 337748
rect 280791 337708 284060 337736
rect 280791 337705 280803 337708
rect 280745 337699 280803 337705
rect 284054 337696 284060 337708
rect 284112 337696 284118 337748
rect 293346 337696 293352 337748
rect 293404 337736 293410 337748
rect 294174 337736 294180 337748
rect 293404 337708 294180 337736
rect 293404 337696 293410 337708
rect 294174 337696 294180 337708
rect 294232 337696 294238 337748
rect 294818 337696 294824 337748
rect 294876 337736 294882 337748
rect 295738 337736 295744 337748
rect 294876 337708 295744 337736
rect 294876 337696 294882 337708
rect 295738 337696 295744 337708
rect 295796 337696 295802 337748
rect 296290 337696 296296 337748
rect 296348 337736 296354 337748
rect 296750 337736 296756 337748
rect 296348 337708 296756 337736
rect 296348 337696 296354 337708
rect 296750 337696 296756 337708
rect 296808 337696 296814 337748
rect 296842 337696 296848 337748
rect 296900 337736 296906 337748
rect 297026 337736 297032 337748
rect 296900 337708 297032 337736
rect 296900 337696 296906 337708
rect 297026 337696 297032 337708
rect 297084 337696 297090 337748
rect 297578 337696 297584 337748
rect 297636 337736 297642 337748
rect 298314 337736 298320 337748
rect 297636 337708 298320 337736
rect 297636 337696 297642 337708
rect 298314 337696 298320 337708
rect 298372 337696 298378 337748
rect 298774 337696 298780 337748
rect 298832 337736 298838 337748
rect 299510 337736 299516 337748
rect 298832 337708 299516 337736
rect 298832 337696 298838 337708
rect 299510 337696 299516 337708
rect 299568 337696 299574 337748
rect 300706 337696 300712 337748
rect 300764 337736 300770 337748
rect 301166 337736 301172 337748
rect 300764 337708 301172 337736
rect 300764 337696 300770 337708
rect 301166 337696 301172 337708
rect 301224 337696 301230 337748
rect 302178 337696 302184 337748
rect 302236 337736 302242 337748
rect 302454 337736 302460 337748
rect 302236 337708 302460 337736
rect 302236 337696 302242 337708
rect 302454 337696 302460 337708
rect 302512 337696 302518 337748
rect 302914 337696 302920 337748
rect 302972 337736 302978 337748
rect 303926 337736 303932 337748
rect 302972 337708 303932 337736
rect 302972 337696 302978 337708
rect 303926 337696 303932 337708
rect 303984 337696 303990 337748
rect 304662 337696 304668 337748
rect 304720 337736 304726 337748
rect 305214 337736 305220 337748
rect 304720 337708 305220 337736
rect 304720 337696 304726 337708
rect 305214 337696 305220 337708
rect 305272 337696 305278 337748
rect 306410 337696 306416 337748
rect 306468 337736 306474 337748
rect 306594 337736 306600 337748
rect 306468 337708 306600 337736
rect 306468 337696 306474 337708
rect 306594 337696 306600 337708
rect 306652 337696 306658 337748
rect 307330 337696 307336 337748
rect 307388 337736 307394 337748
rect 307974 337736 307980 337748
rect 307388 337708 307980 337736
rect 307388 337696 307394 337708
rect 307974 337696 307980 337708
rect 308032 337696 308038 337748
rect 309998 337696 310004 337748
rect 310056 337736 310062 337748
rect 310826 337736 310832 337748
rect 310056 337708 310832 337736
rect 310056 337696 310062 337708
rect 310826 337696 310832 337708
rect 310884 337696 310890 337748
rect 312022 337696 312028 337748
rect 312080 337736 312086 337748
rect 312298 337736 312304 337748
rect 312080 337708 312304 337736
rect 312080 337696 312086 337708
rect 312298 337696 312304 337708
rect 312356 337696 312362 337748
rect 315061 337739 315119 337745
rect 315061 337705 315073 337739
rect 315107 337736 315119 337739
rect 378630 337736 378636 337748
rect 315107 337708 378636 337736
rect 315107 337705 315119 337708
rect 315061 337699 315119 337705
rect 378630 337696 378636 337708
rect 378688 337696 378694 337748
rect 219764 337640 220068 337668
rect 220117 337671 220175 337677
rect 219657 337631 219715 337637
rect 220117 337637 220129 337671
rect 220163 337668 220175 337671
rect 230050 337668 230056 337680
rect 220163 337640 230056 337668
rect 220163 337637 220175 337640
rect 220117 337631 220175 337637
rect 230050 337628 230056 337640
rect 230108 337628 230114 337680
rect 266761 337671 266819 337677
rect 266761 337637 266773 337671
rect 266807 337668 266819 337671
rect 278537 337671 278595 337677
rect 278537 337668 278549 337671
rect 266807 337640 278549 337668
rect 266807 337637 266819 337640
rect 266761 337631 266819 337637
rect 278537 337637 278549 337640
rect 278583 337637 278595 337671
rect 278537 337631 278595 337637
rect 292886 337628 292892 337680
rect 292944 337668 292950 337680
rect 293714 337668 293720 337680
rect 292944 337640 293720 337668
rect 292944 337628 292950 337640
rect 293714 337628 293720 337640
rect 293772 337628 293778 337680
rect 293898 337628 293904 337680
rect 293956 337668 293962 337680
rect 295186 337668 295192 337680
rect 293956 337640 295192 337668
rect 293956 337628 293962 337640
rect 295186 337628 295192 337640
rect 295244 337628 295250 337680
rect 295370 337628 295376 337680
rect 295428 337668 295434 337680
rect 295554 337668 295560 337680
rect 295428 337640 295560 337668
rect 295428 337628 295434 337640
rect 295554 337628 295560 337640
rect 295612 337628 295618 337680
rect 296566 337628 296572 337680
rect 296624 337668 296630 337680
rect 296624 337640 299004 337668
rect 296624 337628 296630 337640
rect 129092 337572 130368 337600
rect 133177 337603 133235 337609
rect 129092 337560 129098 337572
rect 133177 337569 133189 337603
rect 133223 337600 133235 337603
rect 142466 337600 142472 337612
rect 133223 337572 142472 337600
rect 133223 337569 133235 337572
rect 133177 337563 133235 337569
rect 142466 337560 142472 337572
rect 142524 337560 142530 337612
rect 142561 337603 142619 337609
rect 142561 337569 142573 337603
rect 142607 337600 142619 337603
rect 142650 337600 142656 337612
rect 142607 337572 142656 337600
rect 142607 337569 142619 337572
rect 142561 337563 142619 337569
rect 142650 337560 142656 337572
rect 142708 337560 142714 337612
rect 142742 337560 142748 337612
rect 142800 337600 142806 337612
rect 152126 337600 152132 337612
rect 142800 337572 152132 337600
rect 142800 337560 142806 337572
rect 152126 337560 152132 337572
rect 152184 337560 152190 337612
rect 152218 337560 152224 337612
rect 152276 337600 152282 337612
rect 152313 337603 152371 337609
rect 152313 337600 152325 337603
rect 152276 337572 152325 337600
rect 152276 337560 152282 337572
rect 152313 337569 152325 337572
rect 152359 337569 152371 337603
rect 152313 337563 152371 337569
rect 152402 337560 152408 337612
rect 152460 337600 152466 337612
rect 161786 337600 161792 337612
rect 152460 337572 161792 337600
rect 152460 337560 152466 337572
rect 161786 337560 161792 337572
rect 161844 337560 161850 337612
rect 161881 337603 161939 337609
rect 161881 337569 161893 337603
rect 161927 337600 161939 337603
rect 161970 337600 161976 337612
rect 161927 337572 161976 337600
rect 161927 337569 161939 337572
rect 161881 337563 161939 337569
rect 161970 337560 161976 337572
rect 162028 337560 162034 337612
rect 162062 337560 162068 337612
rect 162120 337600 162126 337612
rect 171446 337600 171452 337612
rect 162120 337572 171452 337600
rect 162120 337560 162126 337572
rect 171446 337560 171452 337572
rect 171504 337560 171510 337612
rect 171538 337560 171544 337612
rect 171596 337600 171602 337612
rect 171633 337603 171691 337609
rect 171633 337600 171645 337603
rect 171596 337572 171645 337600
rect 171596 337560 171602 337572
rect 171633 337569 171645 337572
rect 171679 337569 171691 337603
rect 171633 337563 171691 337569
rect 171722 337560 171728 337612
rect 171780 337600 171786 337612
rect 181106 337600 181112 337612
rect 171780 337572 181112 337600
rect 171780 337560 171786 337572
rect 181106 337560 181112 337572
rect 181164 337560 181170 337612
rect 181201 337603 181259 337609
rect 181201 337569 181213 337603
rect 181247 337600 181259 337603
rect 181290 337600 181296 337612
rect 181247 337572 181296 337600
rect 181247 337569 181259 337572
rect 181201 337563 181259 337569
rect 181290 337560 181296 337572
rect 181348 337560 181354 337612
rect 181382 337560 181388 337612
rect 181440 337600 181446 337612
rect 190766 337600 190772 337612
rect 181440 337572 190772 337600
rect 181440 337560 181446 337572
rect 190766 337560 190772 337572
rect 190824 337560 190830 337612
rect 190858 337560 190864 337612
rect 190916 337600 190922 337612
rect 190953 337603 191011 337609
rect 190953 337600 190965 337603
rect 190916 337572 190965 337600
rect 190916 337560 190922 337572
rect 190953 337569 190965 337572
rect 190999 337569 191011 337603
rect 190953 337563 191011 337569
rect 191042 337560 191048 337612
rect 191100 337600 191106 337612
rect 200426 337600 200432 337612
rect 191100 337572 200432 337600
rect 191100 337560 191106 337572
rect 200426 337560 200432 337572
rect 200484 337560 200490 337612
rect 200521 337603 200579 337609
rect 200521 337569 200533 337603
rect 200567 337600 200579 337603
rect 200610 337600 200616 337612
rect 200567 337572 200616 337600
rect 200567 337569 200579 337572
rect 200521 337563 200579 337569
rect 200610 337560 200616 337572
rect 200668 337560 200674 337612
rect 200702 337560 200708 337612
rect 200760 337600 200766 337612
rect 210086 337600 210092 337612
rect 200760 337572 210092 337600
rect 200760 337560 200766 337572
rect 210086 337560 210092 337572
rect 210144 337560 210150 337612
rect 210178 337560 210184 337612
rect 210236 337600 210242 337612
rect 210273 337603 210331 337609
rect 210273 337600 210285 337603
rect 210236 337572 210285 337600
rect 210236 337560 210242 337572
rect 210273 337569 210285 337572
rect 210319 337569 210331 337603
rect 210273 337563 210331 337569
rect 210362 337560 210368 337612
rect 210420 337600 210426 337612
rect 219746 337600 219752 337612
rect 210420 337572 219752 337600
rect 210420 337560 210426 337572
rect 219746 337560 219752 337572
rect 219804 337560 219810 337612
rect 219841 337603 219899 337609
rect 219841 337569 219853 337603
rect 219887 337600 219899 337603
rect 219930 337600 219936 337612
rect 219887 337572 219936 337600
rect 219887 337569 219899 337572
rect 219841 337563 219899 337569
rect 219930 337560 219936 337572
rect 219988 337560 219994 337612
rect 220022 337560 220028 337612
rect 220080 337600 220086 337612
rect 225453 337603 225511 337609
rect 225453 337600 225465 337603
rect 220080 337572 225465 337600
rect 220080 337560 220086 337572
rect 225453 337569 225465 337572
rect 225499 337569 225511 337603
rect 225453 337563 225511 337569
rect 225545 337603 225603 337609
rect 225545 337569 225557 337603
rect 225591 337600 225603 337603
rect 239250 337600 239256 337612
rect 225591 337572 239256 337600
rect 225591 337569 225603 337572
rect 225545 337563 225603 337569
rect 239250 337560 239256 337572
rect 239308 337560 239314 337612
rect 251578 337560 251584 337612
rect 251636 337600 251642 337612
rect 281846 337600 281852 337612
rect 251636 337572 281852 337600
rect 251636 337560 251642 337572
rect 281846 337560 281852 337572
rect 281904 337560 281910 337612
rect 293622 337560 293628 337612
rect 293680 337600 293686 337612
rect 294358 337600 294364 337612
rect 293680 337572 294364 337600
rect 293680 337560 293686 337572
rect 294358 337560 294364 337572
rect 294416 337560 294422 337612
rect 296106 337560 296112 337612
rect 296164 337600 296170 337612
rect 297026 337600 297032 337612
rect 296164 337572 297032 337600
rect 296164 337560 296170 337572
rect 297026 337560 297032 337572
rect 297084 337560 297090 337612
rect 297762 337560 297768 337612
rect 297820 337600 297826 337612
rect 298406 337600 298412 337612
rect 297820 337572 298412 337600
rect 297820 337560 297826 337572
rect 298406 337560 298412 337572
rect 298464 337560 298470 337612
rect 128850 337532 128856 337544
rect 128684 337504 128856 337532
rect 128850 337492 128856 337504
rect 128908 337492 128914 337544
rect 129126 337492 129132 337544
rect 129184 337532 129190 337544
rect 253970 337532 253976 337544
rect 129184 337504 253976 337532
rect 129184 337492 129190 337504
rect 253970 337492 253976 337504
rect 254028 337492 254034 337544
rect 254338 337492 254344 337544
rect 254396 337532 254402 337544
rect 282582 337532 282588 337544
rect 254396 337504 282588 337532
rect 254396 337492 254402 337504
rect 282582 337492 282588 337504
rect 282640 337492 282646 337544
rect 295830 337492 295836 337544
rect 295888 337532 295894 337544
rect 297118 337532 297124 337544
rect 295888 337504 297124 337532
rect 295888 337492 295894 337504
rect 297118 337492 297124 337504
rect 297176 337492 297182 337544
rect 298976 337532 299004 337640
rect 299234 337628 299240 337680
rect 299292 337668 299298 337680
rect 299878 337668 299884 337680
rect 299292 337640 299884 337668
rect 299292 337628 299298 337640
rect 299878 337628 299884 337640
rect 299936 337628 299942 337680
rect 299970 337628 299976 337680
rect 300028 337668 300034 337680
rect 301258 337668 301264 337680
rect 300028 337640 301264 337668
rect 300028 337628 300034 337640
rect 301258 337628 301264 337640
rect 301316 337628 301322 337680
rect 301994 337628 302000 337680
rect 302052 337668 302058 337680
rect 302546 337668 302552 337680
rect 302052 337640 302552 337668
rect 302052 337628 302058 337640
rect 302546 337628 302552 337640
rect 302604 337628 302610 337680
rect 304386 337628 304392 337680
rect 304444 337668 304450 337680
rect 305306 337668 305312 337680
rect 304444 337640 305312 337668
rect 304444 337628 304450 337640
rect 305306 337628 305312 337640
rect 305364 337628 305370 337680
rect 305858 337628 305864 337680
rect 305916 337668 305922 337680
rect 306686 337668 306692 337680
rect 305916 337640 306692 337668
rect 305916 337628 305922 337640
rect 306686 337628 306692 337640
rect 306744 337628 306750 337680
rect 310274 337628 310280 337680
rect 310332 337668 310338 337680
rect 310642 337668 310648 337680
rect 310332 337640 310648 337668
rect 310332 337628 310338 337640
rect 310642 337628 310648 337640
rect 310700 337628 310706 337680
rect 311470 337628 311476 337680
rect 311528 337668 311534 337680
rect 312114 337668 312120 337680
rect 311528 337640 312120 337668
rect 311528 337628 311534 337640
rect 312114 337628 312120 337640
rect 312172 337628 312178 337680
rect 317085 337671 317143 337677
rect 317085 337637 317097 337671
rect 317131 337668 317143 337671
rect 385530 337668 385536 337680
rect 317131 337640 385536 337668
rect 317131 337637 317143 337640
rect 317085 337631 317143 337637
rect 385530 337628 385536 337640
rect 385588 337628 385594 337680
rect 299050 337560 299056 337612
rect 299108 337600 299114 337612
rect 299786 337600 299792 337612
rect 299108 337572 299792 337600
rect 299108 337560 299114 337572
rect 299786 337560 299792 337572
rect 299844 337560 299850 337612
rect 301442 337560 301448 337612
rect 301500 337600 301506 337612
rect 302638 337600 302644 337612
rect 301500 337572 302644 337600
rect 301500 337560 301506 337572
rect 302638 337560 302644 337572
rect 302696 337560 302702 337612
rect 306134 337560 306140 337612
rect 306192 337600 306198 337612
rect 306594 337600 306600 337612
rect 306192 337572 306600 337600
rect 306192 337560 306198 337572
rect 306594 337560 306600 337572
rect 306652 337560 306658 337612
rect 311010 337560 311016 337612
rect 311068 337600 311074 337612
rect 312022 337600 312028 337612
rect 311068 337572 312028 337600
rect 311068 337560 311074 337572
rect 312022 337560 312028 337572
rect 312080 337560 312086 337612
rect 321961 337603 322019 337609
rect 321961 337569 321973 337603
rect 322007 337600 322019 337603
rect 392430 337600 392436 337612
rect 322007 337572 392436 337600
rect 322007 337569 322019 337572
rect 321961 337563 322019 337569
rect 392430 337560 392436 337572
rect 392488 337560 392494 337612
rect 303374 337532 303380 337544
rect 298976 337504 303380 337532
rect 303374 337492 303380 337504
rect 303432 337492 303438 337544
rect 306870 337492 306876 337544
rect 306928 337532 306934 337544
rect 306928 337504 310504 337532
rect 306928 337492 306934 337504
rect 21118 337424 21124 337476
rect 21176 337464 21182 337476
rect 133177 337467 133235 337473
rect 133177 337464 133189 337467
rect 21176 337436 133189 337464
rect 21176 337424 21182 337436
rect 133177 337433 133189 337436
rect 133223 337433 133235 337467
rect 133177 337427 133235 337433
rect 142374 337424 142380 337476
rect 142432 337464 142438 337476
rect 152494 337464 152500 337476
rect 142432 337436 152500 337464
rect 142432 337424 142438 337436
rect 152494 337424 152500 337436
rect 152552 337424 152558 337476
rect 161694 337424 161700 337476
rect 161752 337464 161758 337476
rect 171814 337464 171820 337476
rect 161752 337436 171820 337464
rect 161752 337424 161758 337436
rect 171814 337424 171820 337436
rect 171872 337424 171878 337476
rect 181014 337424 181020 337476
rect 181072 337464 181078 337476
rect 191134 337464 191140 337476
rect 181072 337436 191140 337464
rect 181072 337424 181078 337436
rect 191134 337424 191140 337436
rect 191192 337424 191198 337476
rect 200334 337424 200340 337476
rect 200392 337464 200398 337476
rect 210454 337464 210460 337476
rect 200392 337436 210460 337464
rect 200392 337424 200398 337436
rect 210454 337424 210460 337436
rect 210512 337424 210518 337476
rect 219654 337424 219660 337476
rect 219712 337464 219718 337476
rect 219712 337436 226876 337464
rect 219712 337424 219718 337436
rect 11458 337356 11464 337408
rect 11516 337396 11522 337408
rect 17073 337399 17131 337405
rect 17073 337396 17085 337399
rect 11516 337368 17085 337396
rect 11516 337356 11522 337368
rect 17073 337365 17085 337368
rect 17119 337365 17131 337399
rect 17073 337359 17131 337365
rect 26638 337356 26644 337408
rect 26696 337396 26702 337408
rect 36390 337396 36396 337408
rect 26696 337368 36396 337396
rect 26696 337356 26702 337368
rect 36390 337356 36396 337368
rect 36448 337356 36454 337408
rect 45958 337356 45964 337408
rect 46016 337396 46022 337408
rect 55710 337396 55716 337408
rect 46016 337368 55716 337396
rect 46016 337356 46022 337368
rect 55710 337356 55716 337368
rect 55768 337356 55774 337408
rect 65278 337356 65284 337408
rect 65336 337396 65342 337408
rect 75030 337396 75036 337408
rect 65336 337368 75036 337396
rect 65336 337356 65342 337368
rect 75030 337356 75036 337368
rect 75088 337356 75094 337408
rect 84598 337356 84604 337408
rect 84656 337396 84662 337408
rect 94350 337396 94356 337408
rect 84656 337368 94356 337396
rect 84656 337356 84662 337368
rect 94350 337356 94356 337368
rect 94408 337356 94414 337408
rect 103918 337356 103924 337408
rect 103976 337396 103982 337408
rect 113673 337399 113731 337405
rect 113673 337396 113685 337399
rect 103976 337368 113685 337396
rect 103976 337356 103982 337368
rect 113673 337365 113685 337368
rect 113719 337365 113731 337399
rect 113673 337359 113731 337365
rect 113857 337399 113915 337405
rect 113857 337365 113869 337399
rect 113903 337396 113915 337399
rect 119193 337399 119251 337405
rect 119193 337396 119205 337399
rect 113903 337368 119205 337396
rect 113903 337365 113915 337368
rect 113857 337359 113915 337365
rect 119193 337365 119205 337368
rect 119239 337365 119251 337399
rect 119193 337359 119251 337365
rect 119285 337399 119343 337405
rect 119285 337365 119297 337399
rect 119331 337396 119343 337399
rect 123882 337396 123888 337408
rect 119331 337368 123888 337396
rect 119331 337365 119343 337368
rect 119285 337359 119343 337365
rect 123882 337356 123888 337368
rect 123940 337356 123946 337408
rect 123977 337399 124035 337405
rect 123977 337365 123989 337399
rect 124023 337396 124035 337399
rect 138326 337396 138332 337408
rect 124023 337368 138332 337396
rect 124023 337365 124035 337368
rect 123977 337359 124035 337365
rect 138326 337356 138332 337368
rect 138384 337356 138390 337408
rect 138421 337399 138479 337405
rect 138421 337365 138433 337399
rect 138467 337396 138479 337399
rect 142469 337399 142527 337405
rect 142469 337396 142481 337399
rect 138467 337368 142481 337396
rect 138467 337365 138479 337368
rect 138421 337359 138479 337365
rect 142469 337365 142481 337368
rect 142515 337365 142527 337399
rect 142469 337359 142527 337365
rect 142558 337356 142564 337408
rect 142616 337396 142622 337408
rect 152310 337396 152316 337408
rect 142616 337368 152316 337396
rect 142616 337356 142622 337368
rect 152310 337356 152316 337368
rect 152368 337356 152374 337408
rect 152405 337399 152463 337405
rect 152405 337365 152417 337399
rect 152451 337396 152463 337399
rect 161789 337399 161847 337405
rect 161789 337396 161801 337399
rect 152451 337368 161801 337396
rect 152451 337365 152463 337368
rect 152405 337359 152463 337365
rect 161789 337365 161801 337368
rect 161835 337365 161847 337399
rect 161789 337359 161847 337365
rect 161878 337356 161884 337408
rect 161936 337396 161942 337408
rect 171630 337396 171636 337408
rect 161936 337368 171636 337396
rect 161936 337356 161942 337368
rect 171630 337356 171636 337368
rect 171688 337356 171694 337408
rect 171725 337399 171783 337405
rect 171725 337365 171737 337399
rect 171771 337396 171783 337399
rect 181109 337399 181167 337405
rect 181109 337396 181121 337399
rect 171771 337368 181121 337396
rect 171771 337365 171783 337368
rect 171725 337359 171783 337365
rect 181109 337365 181121 337368
rect 181155 337365 181167 337399
rect 181109 337359 181167 337365
rect 181198 337356 181204 337408
rect 181256 337396 181262 337408
rect 190950 337396 190956 337408
rect 181256 337368 190956 337396
rect 181256 337356 181262 337368
rect 190950 337356 190956 337368
rect 191008 337356 191014 337408
rect 191045 337399 191103 337405
rect 191045 337365 191057 337399
rect 191091 337396 191103 337399
rect 200429 337399 200487 337405
rect 200429 337396 200441 337399
rect 191091 337368 200441 337396
rect 191091 337365 191103 337368
rect 191045 337359 191103 337365
rect 200429 337365 200441 337368
rect 200475 337365 200487 337399
rect 200429 337359 200487 337365
rect 200518 337356 200524 337408
rect 200576 337396 200582 337408
rect 210270 337396 210276 337408
rect 200576 337368 210276 337396
rect 200576 337356 200582 337368
rect 210270 337356 210276 337368
rect 210328 337356 210334 337408
rect 210365 337399 210423 337405
rect 210365 337365 210377 337399
rect 210411 337396 210423 337399
rect 219749 337399 219807 337405
rect 219749 337396 219761 337399
rect 210411 337368 219761 337396
rect 210411 337365 210423 337368
rect 210365 337359 210423 337365
rect 219749 337365 219761 337368
rect 219795 337365 219807 337399
rect 219749 337359 219807 337365
rect 219838 337356 219844 337408
rect 219896 337396 219902 337408
rect 226741 337399 226799 337405
rect 226741 337396 226753 337399
rect 219896 337368 226753 337396
rect 219896 337356 219902 337368
rect 226741 337365 226753 337368
rect 226787 337365 226799 337399
rect 226848 337396 226876 337436
rect 226922 337424 226928 337476
rect 226980 337464 226986 337476
rect 229961 337467 230019 337473
rect 229961 337464 229973 337467
rect 226980 337436 229973 337464
rect 226980 337424 226986 337436
rect 229961 337433 229973 337436
rect 230007 337433 230019 337467
rect 229961 337427 230019 337433
rect 230050 337424 230056 337476
rect 230108 337464 230114 337476
rect 256178 337464 256184 337476
rect 230108 337436 256184 337464
rect 230108 337424 230114 337436
rect 256178 337424 256184 337436
rect 256236 337424 256242 337476
rect 257098 337424 257104 337476
rect 257156 337464 257162 337476
rect 283134 337464 283140 337476
rect 257156 337436 283140 337464
rect 257156 337424 257162 337436
rect 283134 337424 283140 337436
rect 283192 337424 283198 337476
rect 294634 337424 294640 337476
rect 294692 337464 294698 337476
rect 310274 337464 310280 337476
rect 294692 337436 310280 337464
rect 294692 337424 294698 337436
rect 310274 337424 310280 337436
rect 310332 337424 310338 337476
rect 310476 337464 310504 337504
rect 310550 337492 310556 337544
rect 310608 337532 310614 337544
rect 310918 337532 310924 337544
rect 310608 337504 310924 337532
rect 310608 337492 310614 337504
rect 310918 337492 310924 337504
rect 310976 337492 310982 337544
rect 311286 337492 311292 337544
rect 311344 337532 311350 337544
rect 314141 337535 314199 337541
rect 314141 337532 314153 337535
rect 311344 337504 314153 337532
rect 311344 337492 311350 337504
rect 314141 337501 314153 337504
rect 314187 337501 314199 337535
rect 314141 337495 314199 337501
rect 314230 337492 314236 337544
rect 314288 337532 314294 337544
rect 318189 337535 318247 337541
rect 314288 337504 318140 337532
rect 314288 337492 314294 337504
rect 317177 337467 317235 337473
rect 317177 337464 317189 337467
rect 310476 337436 317189 337464
rect 317177 337433 317189 337436
rect 317223 337433 317235 337467
rect 318112 337464 318140 337504
rect 318189 337501 318201 337535
rect 318235 337532 318247 337535
rect 400710 337532 400716 337544
rect 318235 337504 400716 337532
rect 318235 337501 318247 337504
rect 318189 337495 318247 337501
rect 400710 337492 400716 337504
rect 400768 337492 400774 337544
rect 407610 337464 407616 337476
rect 318112 337436 407616 337464
rect 317177 337427 317235 337433
rect 407610 337424 407616 337436
rect 407668 337424 407674 337476
rect 252498 337396 252504 337408
rect 226848 337368 252504 337396
rect 226741 337359 226799 337365
rect 252498 337356 252504 337368
rect 252556 337356 252562 337408
rect 254246 337356 254252 337408
rect 254304 337396 254310 337408
rect 282398 337396 282404 337408
rect 254304 337368 282404 337396
rect 254304 337356 254310 337368
rect 282398 337356 282404 337368
rect 282456 337356 282462 337408
rect 295094 337356 295100 337408
rect 295152 337396 295158 337408
rect 308437 337399 308495 337405
rect 308437 337396 308449 337399
rect 295152 337368 308449 337396
rect 295152 337356 295158 337368
rect 308437 337365 308449 337368
rect 308483 337365 308495 337399
rect 308437 337359 308495 337365
rect 308526 337356 308532 337408
rect 308584 337396 308590 337408
rect 309354 337396 309360 337408
rect 308584 337368 309360 337396
rect 308584 337356 308590 337368
rect 309354 337356 309360 337368
rect 309412 337356 309418 337408
rect 312758 337356 312764 337408
rect 312816 337396 312822 337408
rect 313678 337396 313684 337408
rect 312816 337368 313684 337396
rect 312816 337356 312822 337368
rect 313678 337356 313684 337368
rect 313736 337356 313742 337408
rect 315702 337356 315708 337408
rect 315760 337396 315766 337408
rect 414510 337396 414516 337408
rect 315760 337368 414516 337396
rect 315760 337356 315766 337368
rect 414510 337356 414516 337368
rect 414568 337356 414574 337408
rect 1600 337232 583316 337328
rect 17073 337195 17131 337201
rect 17073 337161 17085 337195
rect 17119 337192 17131 337195
rect 26638 337192 26644 337204
rect 17119 337164 26644 337192
rect 17119 337161 17131 337164
rect 17073 337155 17131 337161
rect 26638 337152 26644 337164
rect 26696 337152 26702 337204
rect 55713 337195 55771 337201
rect 55713 337161 55725 337195
rect 55759 337192 55771 337195
rect 65186 337192 65192 337204
rect 55759 337164 65192 337192
rect 55759 337161 55771 337164
rect 55713 337155 55771 337161
rect 65186 337152 65192 337164
rect 65244 337152 65250 337204
rect 69418 337152 69424 337204
rect 69476 337192 69482 337204
rect 244402 337192 244408 337204
rect 69476 337164 244408 337192
rect 69476 337152 69482 337164
rect 244402 337152 244408 337164
rect 244460 337152 244466 337204
rect 245325 337195 245383 337201
rect 245325 337161 245337 337195
rect 245371 337192 245383 337195
rect 251026 337192 251032 337204
rect 245371 337164 251032 337192
rect 245371 337161 245383 337164
rect 245325 337155 245383 337161
rect 251026 337152 251032 337164
rect 251084 337152 251090 337204
rect 280098 337152 280104 337204
rect 280156 337192 280162 337204
rect 287274 337192 287280 337204
rect 280156 337164 287280 337192
rect 280156 337152 280162 337164
rect 287274 337152 287280 337164
rect 287332 337152 287338 337204
rect 293162 337152 293168 337204
rect 293220 337192 293226 337204
rect 295094 337192 295100 337204
rect 293220 337164 295100 337192
rect 293220 337152 293226 337164
rect 295094 337152 295100 337164
rect 295152 337152 295158 337204
rect 301718 337152 301724 337204
rect 301776 337192 301782 337204
rect 313034 337192 313040 337204
rect 301776 337164 313040 337192
rect 301776 337152 301782 337164
rect 313034 337152 313040 337164
rect 313092 337152 313098 337204
rect 313678 337152 313684 337204
rect 313736 337192 313742 337204
rect 318189 337195 318247 337201
rect 318189 337192 318201 337195
rect 313736 337164 318201 337192
rect 313736 337152 313742 337164
rect 318189 337161 318201 337164
rect 318235 337161 318247 337195
rect 318189 337155 318247 337161
rect 342382 337152 342388 337204
rect 342440 337192 342446 337204
rect 342658 337192 342664 337204
rect 342440 337164 342664 337192
rect 342440 337152 342446 337164
rect 342658 337152 342664 337164
rect 342716 337152 342722 337204
rect 342842 337152 342848 337204
rect 342900 337192 342906 337204
rect 343762 337192 343768 337204
rect 342900 337164 343768 337192
rect 342900 337152 342906 337164
rect 343762 337152 343768 337164
rect 343820 337152 343826 337204
rect 344590 337152 344596 337204
rect 344648 337192 344654 337204
rect 345418 337192 345424 337204
rect 344648 337164 345424 337192
rect 344648 337152 344654 337164
rect 345418 337152 345424 337164
rect 345476 337152 345482 337204
rect 346246 337152 346252 337204
rect 346304 337192 346310 337204
rect 346522 337192 346528 337204
rect 346304 337164 346528 337192
rect 346304 337152 346310 337164
rect 346522 337152 346528 337164
rect 346580 337152 346586 337204
rect 347534 337152 347540 337204
rect 347592 337192 347598 337204
rect 348178 337192 348184 337204
rect 347592 337164 348184 337192
rect 347592 337152 347598 337164
rect 348178 337152 348184 337164
rect 348236 337152 348242 337204
rect 348270 337152 348276 337204
rect 348328 337192 348334 337204
rect 349190 337192 349196 337204
rect 348328 337164 349196 337192
rect 348328 337152 348334 337164
rect 349190 337152 349196 337164
rect 349248 337152 349254 337204
rect 349282 337152 349288 337204
rect 349340 337192 349346 337204
rect 349466 337192 349472 337204
rect 349340 337164 349472 337192
rect 349340 337152 349346 337164
rect 349466 337152 349472 337164
rect 349524 337152 349530 337204
rect 349926 337152 349932 337204
rect 349984 337192 349990 337204
rect 350938 337192 350944 337204
rect 349984 337164 350944 337192
rect 349984 337152 349990 337164
rect 350938 337152 350944 337164
rect 350996 337152 351002 337204
rect 76318 337084 76324 337136
rect 76376 337124 76382 337136
rect 245874 337124 245880 337136
rect 76376 337096 245880 337124
rect 76376 337084 76382 337096
rect 245874 337084 245880 337096
rect 245932 337084 245938 337136
rect 278534 337084 278540 337136
rect 278592 337124 278598 337136
rect 286538 337124 286544 337136
rect 278592 337096 286544 337124
rect 278592 337084 278598 337096
rect 286538 337084 286544 337096
rect 286596 337084 286602 337136
rect 291414 337084 291420 337136
rect 291472 337124 291478 337136
rect 293898 337124 293904 337136
rect 291472 337096 293904 337124
rect 291472 337084 291478 337096
rect 293898 337084 293904 337096
rect 293956 337084 293962 337136
rect 308437 337127 308495 337133
rect 308437 337093 308449 337127
rect 308483 337124 308495 337127
rect 314138 337124 314144 337136
rect 308483 337096 314144 337124
rect 308483 337093 308495 337096
rect 308437 337087 308495 337093
rect 314138 337084 314144 337096
rect 314196 337084 314202 337136
rect 314233 337127 314291 337133
rect 314233 337093 314245 337127
rect 314279 337124 314291 337127
rect 321961 337127 322019 337133
rect 321961 337124 321973 337127
rect 314279 337096 321973 337124
rect 314279 337093 314291 337096
rect 314233 337087 314291 337093
rect 321961 337093 321973 337096
rect 322007 337093 322019 337127
rect 321961 337087 322019 337093
rect 341370 337084 341376 337136
rect 341428 337124 341434 337136
rect 342474 337124 342480 337136
rect 341428 337096 342480 337124
rect 341428 337084 341434 337096
rect 342474 337084 342480 337096
rect 342532 337084 342538 337136
rect 344314 337084 344320 337136
rect 344372 337124 344378 337136
rect 345050 337124 345056 337136
rect 344372 337096 345056 337124
rect 344372 337084 344378 337096
rect 345050 337084 345056 337096
rect 345108 337084 345114 337136
rect 346062 337084 346068 337136
rect 346120 337124 346126 337136
rect 346798 337124 346804 337136
rect 346120 337096 346804 337124
rect 346120 337084 346126 337096
rect 346798 337084 346804 337096
rect 346856 337084 346862 337136
rect 346982 337084 346988 337136
rect 347040 337124 347046 337136
rect 347994 337124 348000 337136
rect 347040 337096 348000 337124
rect 347040 337084 347046 337096
rect 347994 337084 348000 337096
rect 348052 337084 348058 337136
rect 348730 337084 348736 337136
rect 348788 337124 348794 337136
rect 351766 337124 351772 337136
rect 348788 337096 351772 337124
rect 348788 337084 348794 337096
rect 351766 337084 351772 337096
rect 351824 337084 351830 337136
rect 36390 337016 36396 337068
rect 36448 337056 36454 337068
rect 45958 337056 45964 337068
rect 36448 337028 45964 337056
rect 36448 337016 36454 337028
rect 45958 337016 45964 337028
rect 46016 337016 46022 337068
rect 55710 337016 55716 337068
rect 55768 337056 55774 337068
rect 65278 337056 65284 337068
rect 55768 337028 65284 337056
rect 55768 337016 55774 337028
rect 65278 337016 65284 337028
rect 65336 337016 65342 337068
rect 83218 337016 83224 337068
rect 83276 337056 83282 337068
rect 247346 337056 247352 337068
rect 83276 337028 247352 337056
rect 83276 337016 83282 337028
rect 247346 337016 247352 337028
rect 247404 337016 247410 337068
rect 261238 337016 261244 337068
rect 261296 337056 261302 337068
rect 266761 337059 266819 337065
rect 266761 337056 266773 337059
rect 261296 337028 266773 337056
rect 261296 337016 261302 337028
rect 266761 337025 266773 337028
rect 266807 337025 266819 337059
rect 266761 337019 266819 337025
rect 283502 337016 283508 337068
rect 283560 337056 283566 337068
rect 284146 337056 284152 337068
rect 283560 337028 284152 337056
rect 283560 337016 283566 337028
rect 284146 337016 284152 337028
rect 284204 337016 284210 337068
rect 291138 337016 291144 337068
rect 291196 337056 291202 337068
rect 292242 337056 292248 337068
rect 291196 337028 292248 337056
rect 291196 337016 291202 337028
rect 292242 337016 292248 337028
rect 292300 337016 292306 337068
rect 300522 337016 300528 337068
rect 300580 337056 300586 337068
rect 300982 337056 300988 337068
rect 300580 337028 300988 337056
rect 300580 337016 300586 337028
rect 300982 337016 300988 337028
rect 301040 337016 301046 337068
rect 309814 337016 309820 337068
rect 309872 337056 309878 337068
rect 317085 337059 317143 337065
rect 317085 337056 317097 337059
rect 309872 337028 317097 337056
rect 309872 337016 309878 337028
rect 317085 337025 317097 337028
rect 317131 337025 317143 337059
rect 317085 337019 317143 337025
rect 318370 337016 318376 337068
rect 318428 337056 318434 337068
rect 318830 337056 318836 337068
rect 318428 337028 318836 337056
rect 318428 337016 318434 337028
rect 318830 337016 318836 337028
rect 318888 337016 318894 337068
rect 321038 337016 321044 337068
rect 321096 337056 321102 337068
rect 321590 337056 321596 337068
rect 321096 337028 321596 337056
rect 321096 337016 321102 337028
rect 321590 337016 321596 337028
rect 321648 337016 321654 337068
rect 326650 337016 326656 337068
rect 326708 337056 326714 337068
rect 327386 337056 327392 337068
rect 326708 337028 327392 337056
rect 326708 337016 326714 337028
rect 327386 337016 327392 337028
rect 327444 337016 327450 337068
rect 332078 337016 332084 337068
rect 332136 337056 332142 337068
rect 332630 337056 332636 337068
rect 332136 337028 332636 337056
rect 332136 337016 332142 337028
rect 332630 337016 332636 337028
rect 332688 337016 332694 337068
rect 336218 337016 336224 337068
rect 336276 337056 336282 337068
rect 336770 337056 336776 337068
rect 336276 337028 336776 337056
rect 336276 337016 336282 337028
rect 336770 337016 336776 337028
rect 336828 337016 336834 337068
rect 341646 337016 341652 337068
rect 341704 337056 341710 337068
rect 342658 337056 342664 337068
rect 341704 337028 342664 337056
rect 341704 337016 341710 337028
rect 342658 337016 342664 337028
rect 342716 337016 342722 337068
rect 343118 337016 343124 337068
rect 343176 337056 343182 337068
rect 343578 337056 343584 337068
rect 343176 337028 343584 337056
rect 343176 337016 343182 337028
rect 343578 337016 343584 337028
rect 343636 337016 343642 337068
rect 343670 337016 343676 337068
rect 343728 337056 343734 337068
rect 344038 337056 344044 337068
rect 343728 337028 344044 337056
rect 343728 337016 343734 337028
rect 344038 337016 344044 337028
rect 344096 337016 344102 337068
rect 345510 337016 345516 337068
rect 345568 337056 345574 337068
rect 346614 337056 346620 337068
rect 345568 337028 346620 337056
rect 345568 337016 345574 337028
rect 346614 337016 346620 337028
rect 346672 337016 346678 337068
rect 347258 337016 347264 337068
rect 347316 337056 347322 337068
rect 347810 337056 347816 337068
rect 347316 337028 347816 337056
rect 347316 337016 347322 337028
rect 347810 337016 347816 337028
rect 347868 337016 347874 337068
rect 348454 337016 348460 337068
rect 348512 337056 348518 337068
rect 349466 337056 349472 337068
rect 348512 337028 349472 337056
rect 348512 337016 348518 337028
rect 349466 337016 349472 337028
rect 349524 337016 349530 337068
rect 75033 336991 75091 336997
rect 75033 336957 75045 336991
rect 75079 336988 75091 336991
rect 84506 336988 84512 337000
rect 75079 336960 84512 336988
rect 75079 336957 75091 336960
rect 75033 336951 75091 336957
rect 84506 336948 84512 336960
rect 84564 336948 84570 337000
rect 87358 336948 87364 337000
rect 87416 336988 87422 337000
rect 248082 336988 248088 337000
rect 87416 336960 248088 336988
rect 87416 336948 87422 336960
rect 248082 336948 248088 336960
rect 248140 336948 248146 337000
rect 288010 336988 288016 337000
rect 284072 336960 288016 336988
rect 94258 336880 94264 336932
rect 94316 336920 94322 336932
rect 249554 336920 249560 336932
rect 94316 336892 249560 336920
rect 94316 336880 94322 336892
rect 249554 336880 249560 336892
rect 249612 336880 249618 336932
rect 284072 336864 284100 336960
rect 288010 336948 288016 336960
rect 288068 336948 288074 337000
rect 290494 336948 290500 337000
rect 290552 336988 290558 337000
rect 291506 336988 291512 337000
rect 290552 336960 291512 336988
rect 290552 336948 290558 336960
rect 291506 336948 291512 336960
rect 291564 336948 291570 337000
rect 291874 336948 291880 337000
rect 291932 336988 291938 337000
rect 292886 336988 292892 337000
rect 291932 336960 292892 336988
rect 291932 336948 291938 336960
rect 292886 336948 292892 336960
rect 292944 336948 292950 337000
rect 298038 336948 298044 337000
rect 298096 336988 298102 337000
rect 306134 336988 306140 337000
rect 298096 336960 306140 336988
rect 298096 336948 298102 336960
rect 306134 336948 306140 336960
rect 306192 336948 306198 337000
rect 308342 336948 308348 337000
rect 308400 336988 308406 337000
rect 315061 336991 315119 336997
rect 315061 336988 315073 336991
rect 308400 336960 315073 336988
rect 308400 336948 308406 336960
rect 315061 336957 315073 336960
rect 315107 336957 315119 336991
rect 315061 336951 315119 336957
rect 315150 336948 315156 337000
rect 315208 336988 315214 337000
rect 316346 336988 316352 337000
rect 315208 336960 316352 336988
rect 315208 336948 315214 336960
rect 316346 336948 316352 336960
rect 316404 336948 316410 337000
rect 316622 336948 316628 337000
rect 316680 336988 316686 337000
rect 317634 336988 317640 337000
rect 316680 336960 317640 336988
rect 316680 336948 316686 336960
rect 317634 336948 317640 336960
rect 317692 336948 317698 337000
rect 318646 336948 318652 337000
rect 318704 336988 318710 337000
rect 319198 336988 319204 337000
rect 318704 336960 319204 336988
rect 318704 336948 318710 336960
rect 319198 336948 319204 336960
rect 319256 336948 319262 337000
rect 320118 336948 320124 337000
rect 320176 336988 320182 337000
rect 320486 336988 320492 337000
rect 320176 336960 320492 336988
rect 320176 336948 320182 336960
rect 320486 336948 320492 336960
rect 320544 336948 320550 337000
rect 320762 336948 320768 337000
rect 320820 336988 320826 337000
rect 321958 336988 321964 337000
rect 320820 336960 321964 336988
rect 320820 336948 320826 336960
rect 321958 336948 321964 336960
rect 322016 336948 322022 337000
rect 326466 336948 326472 337000
rect 326524 336988 326530 337000
rect 327202 336988 327208 337000
rect 326524 336960 327208 336988
rect 326524 336948 326530 336960
rect 327202 336948 327208 336960
rect 327260 336948 327266 337000
rect 328122 336948 328128 337000
rect 328180 336988 328186 337000
rect 328766 336988 328772 337000
rect 328180 336960 328772 336988
rect 328180 336948 328186 336960
rect 328766 336948 328772 336960
rect 328824 336948 328830 337000
rect 330882 336948 330888 337000
rect 330940 336988 330946 337000
rect 331158 336988 331164 337000
rect 330940 336960 331164 336988
rect 330940 336948 330946 336960
rect 331158 336948 331164 336960
rect 331216 336948 331222 337000
rect 331802 336948 331808 337000
rect 331860 336988 331866 337000
rect 332906 336988 332912 337000
rect 331860 336960 332912 336988
rect 331860 336948 331866 336960
rect 332906 336948 332912 336960
rect 332964 336948 332970 337000
rect 333826 336948 333832 337000
rect 333884 336988 333890 337000
rect 334378 336988 334384 337000
rect 333884 336960 334384 336988
rect 333884 336948 333890 336960
rect 334378 336948 334384 336960
rect 334436 336948 334442 337000
rect 334562 336948 334568 337000
rect 334620 336988 334626 337000
rect 335666 336988 335672 337000
rect 334620 336960 335672 336988
rect 334620 336948 334626 336960
rect 335666 336948 335672 336960
rect 335724 336948 335730 337000
rect 335942 336948 335948 337000
rect 336000 336988 336006 337000
rect 336954 336988 336960 337000
rect 336000 336960 336960 336988
rect 336000 336948 336006 336960
rect 336954 336948 336960 336960
rect 337012 336948 337018 337000
rect 338886 336948 338892 337000
rect 338944 336988 338950 337000
rect 339806 336988 339812 337000
rect 338944 336960 339812 336988
rect 338944 336948 338950 336960
rect 339806 336948 339812 336960
rect 339864 336948 339870 337000
rect 340174 336948 340180 337000
rect 340232 336988 340238 337000
rect 341278 336988 341284 337000
rect 340232 336960 341284 336988
rect 340232 336948 340238 336960
rect 341278 336948 341284 336960
rect 341336 336948 341342 337000
rect 345786 336948 345792 337000
rect 345844 336988 345850 337000
rect 346338 336988 346344 337000
rect 345844 336960 346344 336988
rect 345844 336948 345850 336960
rect 346338 336948 346344 336960
rect 346396 336948 346402 337000
rect 347718 336948 347724 337000
rect 347776 336988 347782 337000
rect 348086 336988 348092 337000
rect 347776 336960 348092 336988
rect 347776 336948 347782 336960
rect 348086 336948 348092 336960
rect 348144 336948 348150 337000
rect 349742 336948 349748 337000
rect 349800 336988 349806 337000
rect 350754 336988 350760 337000
rect 349800 336960 350760 336988
rect 349800 336948 349806 336960
rect 350754 336948 350760 336960
rect 350812 336948 350818 337000
rect 290954 336880 290960 336932
rect 291012 336920 291018 336932
rect 291598 336920 291604 336932
rect 291012 336892 291604 336920
rect 291012 336880 291018 336892
rect 291598 336880 291604 336892
rect 291656 336880 291662 336932
rect 291690 336880 291696 336932
rect 291748 336920 291754 336932
rect 292794 336920 292800 336932
rect 291748 336892 292800 336920
rect 291748 336880 291754 336892
rect 292794 336880 292800 336892
rect 292852 336880 292858 336932
rect 307606 336880 307612 336932
rect 307664 336920 307670 336932
rect 307882 336920 307888 336932
rect 307664 336892 307888 336920
rect 307664 336880 307670 336892
rect 307882 336880 307888 336892
rect 307940 336880 307946 336932
rect 313954 336880 313960 336932
rect 314012 336920 314018 336932
rect 314782 336920 314788 336932
rect 314012 336892 314788 336920
rect 314012 336880 314018 336892
rect 314782 336880 314788 336892
rect 314840 336880 314846 336932
rect 315886 336880 315892 336932
rect 315944 336920 315950 336932
rect 316254 336920 316260 336932
rect 315944 336892 316260 336920
rect 315944 336880 315950 336892
rect 316254 336880 316260 336892
rect 316312 336880 316318 336932
rect 317174 336880 317180 336932
rect 317232 336920 317238 336932
rect 317818 336920 317824 336932
rect 317232 336892 317824 336920
rect 317232 336880 317238 336892
rect 317818 336880 317824 336892
rect 317876 336880 317882 336932
rect 319566 336880 319572 336932
rect 319624 336920 319630 336932
rect 320302 336920 320308 336932
rect 319624 336892 320308 336920
rect 319624 336880 319630 336892
rect 320302 336880 320308 336892
rect 320360 336880 320366 336932
rect 321314 336880 321320 336932
rect 321372 336920 321378 336932
rect 321774 336920 321780 336932
rect 321372 336892 321780 336920
rect 321372 336880 321378 336892
rect 321774 336880 321780 336892
rect 321832 336880 321838 336932
rect 322786 336880 322792 336932
rect 322844 336920 322850 336932
rect 323154 336920 323160 336932
rect 322844 336892 323160 336920
rect 322844 336880 322850 336892
rect 323154 336880 323160 336892
rect 323212 336880 323218 336932
rect 323522 336880 323528 336932
rect 323580 336920 323586 336932
rect 324442 336920 324448 336932
rect 323580 336892 324448 336920
rect 323580 336880 323586 336892
rect 324442 336880 324448 336892
rect 324500 336880 324506 336932
rect 325178 336880 325184 336932
rect 325236 336920 325242 336932
rect 326098 336920 326104 336932
rect 325236 336892 326104 336920
rect 325236 336880 325242 336892
rect 326098 336880 326104 336892
rect 326156 336880 326162 336932
rect 326926 336880 326932 336932
rect 326984 336920 326990 336932
rect 327294 336920 327300 336932
rect 326984 336892 327300 336920
rect 326984 336880 326990 336892
rect 327294 336880 327300 336892
rect 327352 336880 327358 336932
rect 329134 336880 329140 336932
rect 329192 336920 329198 336932
rect 330054 336920 330060 336932
rect 329192 336892 330060 336920
rect 329192 336880 329198 336892
rect 330054 336880 330060 336892
rect 330112 336880 330118 336932
rect 330330 336880 330336 336932
rect 330388 336920 330394 336932
rect 331434 336920 331440 336932
rect 330388 336892 331440 336920
rect 330388 336880 330394 336892
rect 331434 336880 331440 336892
rect 331492 336880 331498 336932
rect 332354 336880 332360 336932
rect 332412 336920 332418 336932
rect 332998 336920 333004 336932
rect 332412 336892 333004 336920
rect 332412 336880 332418 336892
rect 332998 336880 333004 336892
rect 333056 336880 333062 336932
rect 333274 336880 333280 336932
rect 333332 336920 333338 336932
rect 334194 336920 334200 336932
rect 333332 336892 334200 336920
rect 333332 336880 333338 336892
rect 334194 336880 334200 336892
rect 334252 336880 334258 336932
rect 335298 336880 335304 336932
rect 335356 336920 335362 336932
rect 335574 336920 335580 336932
rect 335356 336892 335580 336920
rect 335356 336880 335362 336892
rect 335574 336880 335580 336892
rect 335632 336880 335638 336932
rect 336494 336880 336500 336932
rect 336552 336920 336558 336932
rect 337138 336920 337144 336932
rect 336552 336892 337144 336920
rect 336552 336880 336558 336892
rect 337138 336880 337144 336892
rect 337196 336880 337202 336932
rect 337414 336880 337420 336932
rect 337472 336920 337478 336932
rect 338242 336920 338248 336932
rect 337472 336892 338248 336920
rect 337472 336880 337478 336892
rect 338242 336880 338248 336892
rect 338300 336880 338306 336932
rect 339346 336880 339352 336932
rect 339404 336920 339410 336932
rect 339622 336920 339628 336932
rect 339404 336892 339628 336920
rect 339404 336880 339410 336892
rect 339622 336880 339628 336892
rect 339680 336880 339686 336932
rect 340634 336880 340640 336932
rect 340692 336920 340698 336932
rect 341094 336920 341100 336932
rect 340692 336892 341100 336920
rect 340692 336880 340698 336892
rect 341094 336880 341100 336892
rect 341152 336880 341158 336932
rect 342750 336880 342756 336932
rect 342808 336920 342814 336932
rect 343302 336920 343308 336932
rect 342808 336892 343308 336920
rect 342808 336880 342814 336892
rect 343302 336880 343308 336892
rect 343360 336880 343366 336932
rect 75030 336812 75036 336864
rect 75088 336852 75094 336864
rect 84598 336852 84604 336864
rect 75088 336824 84604 336852
rect 75088 336812 75094 336824
rect 84598 336812 84604 336824
rect 84656 336812 84662 336864
rect 94353 336855 94411 336861
rect 94353 336821 94365 336855
rect 94399 336852 94411 336855
rect 101069 336855 101127 336861
rect 101069 336852 101081 336855
rect 94399 336824 101081 336852
rect 94399 336821 94411 336824
rect 94353 336815 94411 336821
rect 101069 336821 101081 336824
rect 101115 336821 101127 336855
rect 101069 336815 101127 336821
rect 101158 336812 101164 336864
rect 101216 336852 101222 336864
rect 245325 336855 245383 336861
rect 245325 336852 245337 336855
rect 101216 336824 245337 336852
rect 101216 336812 101222 336824
rect 245325 336821 245337 336824
rect 245371 336821 245383 336855
rect 245325 336815 245383 336821
rect 245414 336812 245420 336864
rect 245472 336852 245478 336864
rect 247622 336852 247628 336864
rect 245472 336824 247628 336852
rect 245472 336812 245478 336824
rect 247622 336812 247628 336824
rect 247680 336812 247686 336864
rect 249738 336812 249744 336864
rect 249796 336852 249802 336864
rect 250566 336852 250572 336864
rect 249796 336824 250572 336852
rect 249796 336812 249802 336824
rect 250566 336812 250572 336824
rect 250624 336812 250630 336864
rect 256822 336812 256828 336864
rect 256880 336852 256886 336864
rect 258662 336852 258668 336864
rect 256880 336824 258668 336852
rect 256880 336812 256886 336824
rect 258662 336812 258668 336824
rect 258720 336812 258726 336864
rect 276142 336812 276148 336864
rect 276200 336852 276206 336864
rect 278718 336852 278724 336864
rect 276200 336824 278724 336852
rect 276200 336812 276206 336824
rect 278718 336812 278724 336824
rect 278776 336812 278782 336864
rect 284054 336812 284060 336864
rect 284112 336812 284118 336864
rect 284146 336812 284152 336864
rect 284204 336852 284210 336864
rect 285066 336852 285072 336864
rect 284204 336824 285072 336852
rect 284204 336812 284210 336824
rect 285066 336812 285072 336824
rect 285124 336812 285130 336864
rect 287090 336812 287096 336864
rect 287148 336852 287154 336864
rect 287550 336852 287556 336864
rect 287148 336824 287556 336852
rect 287148 336812 287154 336824
rect 287550 336812 287556 336824
rect 287608 336812 287614 336864
rect 288838 336812 288844 336864
rect 288896 336852 288902 336864
rect 289482 336852 289488 336864
rect 288896 336824 289488 336852
rect 288896 336812 288902 336824
rect 289482 336812 289488 336824
rect 289540 336812 289546 336864
rect 290678 336812 290684 336864
rect 290736 336852 290742 336864
rect 291414 336852 291420 336864
rect 290736 336824 291420 336852
rect 290736 336812 290742 336824
rect 291414 336812 291420 336824
rect 291472 336812 291478 336864
rect 292426 336812 292432 336864
rect 292484 336852 292490 336864
rect 292978 336852 292984 336864
rect 292484 336824 292984 336852
rect 292484 336812 292490 336824
rect 292978 336812 292984 336824
rect 293036 336812 293042 336864
rect 312482 336812 312488 336864
rect 312540 336852 312546 336864
rect 313310 336852 313316 336864
rect 312540 336824 313316 336852
rect 312540 336812 312546 336824
rect 313310 336812 313316 336824
rect 313368 336812 313374 336864
rect 313494 336812 313500 336864
rect 313552 336852 313558 336864
rect 313678 336852 313684 336864
rect 313552 336824 313684 336852
rect 313552 336812 313558 336824
rect 313678 336812 313684 336824
rect 313736 336812 313742 336864
rect 314414 336812 314420 336864
rect 314472 336852 314478 336864
rect 314966 336852 314972 336864
rect 314472 336824 314972 336852
rect 314472 336812 314478 336824
rect 314966 336812 314972 336824
rect 315024 336812 315030 336864
rect 315426 336812 315432 336864
rect 315484 336852 315490 336864
rect 316070 336852 316076 336864
rect 315484 336824 316076 336852
rect 315484 336812 315490 336824
rect 316070 336812 316076 336824
rect 316128 336812 316134 336864
rect 316898 336812 316904 336864
rect 316956 336852 316962 336864
rect 317266 336852 317272 336864
rect 316956 336824 317272 336852
rect 316956 336812 316962 336824
rect 317266 336812 317272 336824
rect 317324 336812 317330 336864
rect 317358 336812 317364 336864
rect 317416 336852 317422 336864
rect 317726 336852 317732 336864
rect 317416 336824 317732 336852
rect 317416 336812 317422 336824
rect 317726 336812 317732 336824
rect 317784 336812 317790 336864
rect 318094 336812 318100 336864
rect 318152 336852 318158 336864
rect 318922 336852 318928 336864
rect 318152 336824 318928 336852
rect 318152 336812 318158 336824
rect 318922 336812 318928 336824
rect 318980 336812 318986 336864
rect 319658 336812 319664 336864
rect 319716 336852 319722 336864
rect 320026 336852 320032 336864
rect 319716 336824 320032 336852
rect 319716 336812 319722 336824
rect 320026 336812 320032 336824
rect 320084 336812 320090 336864
rect 320210 336812 320216 336864
rect 320268 336852 320274 336864
rect 320578 336852 320584 336864
rect 320268 336824 320584 336852
rect 320268 336812 320274 336824
rect 320578 336812 320584 336824
rect 320636 336812 320642 336864
rect 321498 336812 321504 336864
rect 321556 336852 321562 336864
rect 321866 336852 321872 336864
rect 321556 336824 321872 336852
rect 321556 336812 321562 336824
rect 321866 336812 321872 336824
rect 321924 336812 321930 336864
rect 322234 336812 322240 336864
rect 322292 336852 322298 336864
rect 322878 336852 322884 336864
rect 322292 336824 322884 336852
rect 322292 336812 322298 336824
rect 322878 336812 322884 336824
rect 322936 336812 322942 336864
rect 322970 336812 322976 336864
rect 323028 336852 323034 336864
rect 323246 336852 323252 336864
rect 323028 336824 323252 336852
rect 323028 336812 323034 336824
rect 323246 336812 323252 336824
rect 323304 336812 323310 336864
rect 323706 336812 323712 336864
rect 323764 336852 323770 336864
rect 324166 336852 324172 336864
rect 323764 336824 324172 336852
rect 323764 336812 323770 336824
rect 324166 336812 324172 336824
rect 324224 336812 324230 336864
rect 324258 336812 324264 336864
rect 324316 336852 324322 336864
rect 324718 336852 324724 336864
rect 324316 336824 324724 336852
rect 324316 336812 324322 336824
rect 324718 336812 324724 336824
rect 324776 336812 324782 336864
rect 324994 336812 325000 336864
rect 325052 336852 325058 336864
rect 325730 336852 325736 336864
rect 325052 336824 325736 336852
rect 325052 336812 325058 336824
rect 325730 336812 325736 336824
rect 325788 336812 325794 336864
rect 326190 336812 326196 336864
rect 326248 336852 326254 336864
rect 327018 336852 327024 336864
rect 326248 336824 327024 336852
rect 326248 336812 326254 336824
rect 327018 336812 327024 336824
rect 327076 336812 327082 336864
rect 327938 336812 327944 336864
rect 327996 336852 328002 336864
rect 328490 336852 328496 336864
rect 327996 336824 328496 336852
rect 327996 336812 328002 336824
rect 328490 336812 328496 336824
rect 328548 336812 328554 336864
rect 329410 336812 329416 336864
rect 329468 336852 329474 336864
rect 329962 336852 329968 336864
rect 329468 336824 329968 336852
rect 329468 336812 329474 336824
rect 329962 336812 329968 336824
rect 330020 336812 330026 336864
rect 331066 336812 331072 336864
rect 331124 336852 331130 336864
rect 331342 336852 331348 336864
rect 331124 336824 331348 336852
rect 331124 336812 331130 336824
rect 331342 336812 331348 336824
rect 331400 336812 331406 336864
rect 332538 336812 332544 336864
rect 332596 336852 332602 336864
rect 332814 336852 332820 336864
rect 332596 336824 332820 336852
rect 332596 336812 332602 336824
rect 332814 336812 332820 336824
rect 332872 336812 332878 336864
rect 334010 336812 334016 336864
rect 334068 336852 334074 336864
rect 334286 336852 334292 336864
rect 334068 336824 334292 336852
rect 334068 336812 334074 336824
rect 334286 336812 334292 336824
rect 334344 336812 334350 336864
rect 334746 336812 334752 336864
rect 334804 336852 334810 336864
rect 335390 336852 335396 336864
rect 334804 336824 335396 336852
rect 334804 336812 334810 336824
rect 335390 336812 335396 336824
rect 335448 336812 335454 336864
rect 336678 336812 336684 336864
rect 336736 336852 336742 336864
rect 337046 336852 337052 336864
rect 336736 336824 337052 336852
rect 336736 336812 336742 336824
rect 337046 336812 337052 336824
rect 337104 336812 337110 336864
rect 337230 336812 337236 336864
rect 337288 336852 337294 336864
rect 338058 336852 338064 336864
rect 337288 336824 338064 336852
rect 337288 336812 337294 336824
rect 338058 336812 338064 336824
rect 338116 336812 338122 336864
rect 338150 336812 338156 336864
rect 338208 336852 338214 336864
rect 338426 336852 338432 336864
rect 338208 336824 338432 336852
rect 338208 336812 338214 336824
rect 338426 336812 338432 336824
rect 338484 336812 338490 336864
rect 339162 336812 339168 336864
rect 339220 336852 339226 336864
rect 339530 336852 339536 336864
rect 339220 336824 339536 336852
rect 339220 336812 339226 336824
rect 339530 336812 339536 336824
rect 339588 336812 339594 336864
rect 340910 336812 340916 336864
rect 340968 336852 340974 336864
rect 341186 336852 341192 336864
rect 340968 336824 341192 336852
rect 340968 336812 340974 336824
rect 341186 336812 341192 336824
rect 341244 336812 341250 336864
rect 1600 336688 583316 336784
rect 101069 336651 101127 336657
rect 101069 336617 101081 336651
rect 101115 336648 101127 336651
rect 103829 336651 103887 336657
rect 103829 336648 103841 336651
rect 101115 336620 103841 336648
rect 101115 336617 101127 336620
rect 101069 336611 101127 336617
rect 103829 336617 103841 336620
rect 103875 336617 103887 336651
rect 103829 336611 103887 336617
rect 108058 336608 108064 336660
rect 108116 336648 108122 336660
rect 113857 336651 113915 336657
rect 113857 336648 113869 336651
rect 108116 336620 113869 336648
rect 108116 336608 108122 336620
rect 113857 336617 113869 336620
rect 113903 336617 113915 336651
rect 113857 336611 113915 336617
rect 142377 336651 142435 336657
rect 142377 336617 142389 336651
rect 142423 336648 142435 336651
rect 142837 336651 142895 336657
rect 142837 336648 142849 336651
rect 142423 336620 142849 336648
rect 142423 336617 142435 336620
rect 142377 336611 142435 336617
rect 142837 336617 142849 336620
rect 142883 336617 142895 336651
rect 142837 336611 142895 336617
rect 152037 336651 152095 336657
rect 152037 336617 152049 336651
rect 152083 336648 152095 336651
rect 152497 336651 152555 336657
rect 152497 336648 152509 336651
rect 152083 336620 152509 336648
rect 152083 336617 152095 336620
rect 152037 336611 152095 336617
rect 152497 336617 152509 336620
rect 152543 336617 152555 336651
rect 152497 336611 152555 336617
rect 161697 336651 161755 336657
rect 161697 336617 161709 336651
rect 161743 336648 161755 336651
rect 162157 336651 162215 336657
rect 162157 336648 162169 336651
rect 161743 336620 162169 336648
rect 161743 336617 161755 336620
rect 161697 336611 161755 336617
rect 162157 336617 162169 336620
rect 162203 336617 162215 336651
rect 162157 336611 162215 336617
rect 171357 336651 171415 336657
rect 171357 336617 171369 336651
rect 171403 336648 171415 336651
rect 171817 336651 171875 336657
rect 171817 336648 171829 336651
rect 171403 336620 171829 336648
rect 171403 336617 171415 336620
rect 171357 336611 171415 336617
rect 171817 336617 171829 336620
rect 171863 336617 171875 336651
rect 171817 336611 171875 336617
rect 181017 336651 181075 336657
rect 181017 336617 181029 336651
rect 181063 336648 181075 336651
rect 181477 336651 181535 336657
rect 181477 336648 181489 336651
rect 181063 336620 181489 336648
rect 181063 336617 181075 336620
rect 181017 336611 181075 336617
rect 181477 336617 181489 336620
rect 181523 336617 181535 336651
rect 181477 336611 181535 336617
rect 190677 336651 190735 336657
rect 190677 336617 190689 336651
rect 190723 336648 190735 336651
rect 191137 336651 191195 336657
rect 191137 336648 191149 336651
rect 190723 336620 191149 336648
rect 190723 336617 190735 336620
rect 190677 336611 190735 336617
rect 191137 336617 191149 336620
rect 191183 336617 191195 336651
rect 191137 336611 191195 336617
rect 200337 336651 200395 336657
rect 200337 336617 200349 336651
rect 200383 336648 200395 336651
rect 200797 336651 200855 336657
rect 200797 336648 200809 336651
rect 200383 336620 200809 336648
rect 200383 336617 200395 336620
rect 200337 336611 200395 336617
rect 200797 336617 200809 336620
rect 200843 336617 200855 336651
rect 200797 336611 200855 336617
rect 209997 336651 210055 336657
rect 209997 336617 210009 336651
rect 210043 336648 210055 336651
rect 210457 336651 210515 336657
rect 210457 336648 210469 336651
rect 210043 336620 210469 336648
rect 210043 336617 210055 336620
rect 209997 336611 210055 336617
rect 210457 336617 210469 336620
rect 210503 336617 210515 336651
rect 210457 336611 210515 336617
rect 219657 336651 219715 336657
rect 219657 336617 219669 336651
rect 219703 336648 219715 336651
rect 220117 336651 220175 336657
rect 220117 336648 220129 336651
rect 219703 336620 220129 336648
rect 219703 336617 219715 336620
rect 219657 336611 219715 336617
rect 220117 336617 220129 336620
rect 220163 336617 220175 336651
rect 220117 336611 220175 336617
rect 355814 336608 355820 336660
rect 355872 336648 355878 336660
rect 580386 336648 580392 336660
rect 355872 336620 580392 336648
rect 355872 336608 355878 336620
rect 580386 336608 580392 336620
rect 580444 336608 580450 336660
rect 116249 336447 116307 336453
rect 116249 336413 116261 336447
rect 116295 336444 116307 336447
rect 119282 336444 119288 336456
rect 116295 336416 119288 336444
rect 116295 336413 116307 336416
rect 116249 336407 116307 336413
rect 119282 336404 119288 336416
rect 119340 336404 119346 336456
rect 284974 336444 284980 336456
rect 284935 336416 284980 336444
rect 284974 336404 284980 336416
rect 285032 336404 285038 336456
rect 225358 336268 225364 336320
rect 225416 336308 225422 336320
rect 276510 336308 276516 336320
rect 225416 336280 276516 336308
rect 225416 336268 225422 336280
rect 276510 336268 276516 336280
rect 276568 336268 276574 336320
rect 302730 336268 302736 336320
rect 302788 336308 302794 336320
rect 351030 336308 351036 336320
rect 302788 336280 351036 336308
rect 302788 336268 302794 336280
rect 351030 336268 351036 336280
rect 351088 336268 351094 336320
rect 1600 336144 583316 336240
rect 181198 336064 181204 336116
rect 181256 336104 181262 336116
rect 267402 336104 267408 336116
rect 181256 336076 267408 336104
rect 181256 336064 181262 336076
rect 267402 336064 267408 336076
rect 267460 336064 267466 336116
rect 304202 336064 304208 336116
rect 304260 336104 304266 336116
rect 357930 336104 357936 336116
rect 304260 336076 357936 336104
rect 304260 336064 304266 336076
rect 357930 336064 357936 336076
rect 357988 336064 357994 336116
rect 127378 335996 127384 336048
rect 127436 336036 127442 336048
rect 256454 336036 256460 336048
rect 127436 336008 256460 336036
rect 127436 335996 127442 336008
rect 256454 335996 256460 336008
rect 256512 335996 256518 336048
rect 323982 335996 323988 336048
rect 324040 336036 324046 336048
rect 454530 336036 454536 336048
rect 324040 336008 454536 336036
rect 324040 335996 324046 336008
rect 454530 335996 454536 336008
rect 454588 335996 454594 336048
rect 275222 335860 275228 335912
rect 275280 335900 275286 335912
rect 275406 335900 275412 335912
rect 275280 335872 275412 335900
rect 275280 335860 275286 335872
rect 275406 335860 275412 335872
rect 275464 335860 275470 335912
rect 275130 335792 275136 335844
rect 275188 335832 275194 335844
rect 275590 335832 275596 335844
rect 275188 335804 275596 335832
rect 275188 335792 275194 335804
rect 275590 335792 275596 335804
rect 275648 335792 275654 335844
rect 231062 335724 231068 335776
rect 231120 335764 231126 335776
rect 231614 335764 231620 335776
rect 231120 335736 231620 335764
rect 231120 335724 231126 335736
rect 231614 335724 231620 335736
rect 231672 335724 231678 335776
rect 235202 335724 235208 335776
rect 235260 335764 235266 335776
rect 235478 335764 235484 335776
rect 235260 335736 235484 335764
rect 235260 335724 235266 335736
rect 235478 335724 235484 335736
rect 235536 335724 235542 335776
rect 237962 335724 237968 335776
rect 238020 335764 238026 335776
rect 238422 335764 238428 335776
rect 238020 335736 238428 335764
rect 238020 335724 238026 335736
rect 238422 335724 238428 335736
rect 238480 335724 238486 335776
rect 239342 335724 239348 335776
rect 239400 335764 239406 335776
rect 239894 335764 239900 335776
rect 239400 335736 239900 335764
rect 239400 335724 239406 335736
rect 239894 335724 239900 335736
rect 239952 335724 239958 335776
rect 245046 335724 245052 335776
rect 245104 335764 245110 335776
rect 245230 335764 245236 335776
rect 245104 335736 245236 335764
rect 245104 335724 245110 335736
rect 245230 335724 245236 335736
rect 245288 335724 245294 335776
rect 247898 335724 247904 335776
rect 247956 335764 247962 335776
rect 248634 335764 248640 335776
rect 247956 335736 248640 335764
rect 247956 335724 247962 335736
rect 248634 335724 248640 335736
rect 248692 335724 248698 335776
rect 253142 335724 253148 335776
rect 253200 335764 253206 335776
rect 254062 335764 254068 335776
rect 253200 335736 254068 335764
rect 253200 335724 253206 335736
rect 254062 335724 254068 335736
rect 254120 335724 254126 335776
rect 254614 335724 254620 335776
rect 254672 335764 254678 335776
rect 255534 335764 255540 335776
rect 254672 335736 255540 335764
rect 254672 335724 254678 335736
rect 255534 335724 255540 335736
rect 255592 335724 255598 335776
rect 260042 335724 260048 335776
rect 260100 335764 260106 335776
rect 260870 335764 260876 335776
rect 260100 335736 260876 335764
rect 260100 335724 260106 335736
rect 260870 335724 260876 335736
rect 260928 335724 260934 335776
rect 264182 335724 264188 335776
rect 264240 335764 264246 335776
rect 264826 335764 264832 335776
rect 264240 335736 264832 335764
rect 264240 335724 264246 335736
rect 264826 335724 264832 335736
rect 264884 335724 264890 335776
rect 265654 335724 265660 335776
rect 265712 335764 265718 335776
rect 266298 335764 266304 335776
rect 265712 335736 266304 335764
rect 265712 335724 265718 335736
rect 266298 335724 266304 335736
rect 266356 335724 266362 335776
rect 268322 335724 268328 335776
rect 268380 335764 268386 335776
rect 268966 335764 268972 335776
rect 268380 335736 268972 335764
rect 268380 335724 268386 335736
rect 268966 335724 268972 335736
rect 269024 335724 269030 335776
rect 269794 335724 269800 335776
rect 269852 335764 269858 335776
rect 270438 335764 270444 335776
rect 269852 335736 270444 335764
rect 269852 335724 269858 335736
rect 270438 335724 270444 335736
rect 270496 335724 270502 335776
rect 271174 335724 271180 335776
rect 271232 335764 271238 335776
rect 271910 335764 271916 335776
rect 271232 335736 271916 335764
rect 271232 335724 271238 335736
rect 271910 335724 271916 335736
rect 271968 335724 271974 335776
rect 273750 335724 273756 335776
rect 273808 335764 273814 335776
rect 274854 335764 274860 335776
rect 273808 335736 274860 335764
rect 273808 335724 273814 335736
rect 274854 335724 274860 335736
rect 274912 335724 274918 335776
rect 276510 335724 276516 335776
rect 276568 335764 276574 335776
rect 276786 335764 276792 335776
rect 276568 335736 276792 335764
rect 276568 335724 276574 335736
rect 276786 335724 276792 335736
rect 276844 335724 276850 335776
rect 328214 335724 328220 335776
rect 328272 335764 328278 335776
rect 328674 335764 328680 335776
rect 328272 335736 328680 335764
rect 328272 335724 328278 335736
rect 328674 335724 328680 335736
rect 328732 335724 328738 335776
rect 1600 335600 583316 335696
rect 229958 335520 229964 335572
rect 230016 335560 230022 335572
rect 230694 335560 230700 335572
rect 230016 335532 230700 335560
rect 230016 335520 230022 335532
rect 230694 335520 230700 335532
rect 230752 335520 230758 335572
rect 231338 335520 231344 335572
rect 231396 335560 231402 335572
rect 231982 335560 231988 335572
rect 231396 335532 231988 335560
rect 231396 335520 231402 335532
rect 231982 335520 231988 335532
rect 232040 335520 232046 335572
rect 232994 335520 233000 335572
rect 233052 335560 233058 335572
rect 233454 335560 233460 335572
rect 233052 335532 233460 335560
rect 233052 335520 233058 335532
rect 233454 335520 233460 335532
rect 233512 335520 233518 335572
rect 233822 335520 233828 335572
rect 233880 335560 233886 335572
rect 234742 335560 234748 335572
rect 233880 335532 234748 335560
rect 233880 335520 233886 335532
rect 234742 335520 234748 335532
rect 234800 335520 234806 335572
rect 235294 335520 235300 335572
rect 235352 335560 235358 335572
rect 235662 335560 235668 335572
rect 235352 335532 235668 335560
rect 235352 335520 235358 335532
rect 235662 335520 235668 335532
rect 235720 335520 235726 335572
rect 236766 335520 236772 335572
rect 236824 335560 236830 335572
rect 237134 335560 237140 335572
rect 236824 335532 237140 335560
rect 236824 335520 236830 335532
rect 237134 335520 237140 335532
rect 237192 335520 237198 335572
rect 238146 335520 238152 335572
rect 238204 335560 238210 335572
rect 238606 335560 238612 335572
rect 238204 335532 238612 335560
rect 238204 335520 238210 335532
rect 238606 335520 238612 335532
rect 238664 335520 238670 335572
rect 239618 335520 239624 335572
rect 239676 335560 239682 335572
rect 240354 335560 240360 335572
rect 239676 335532 240360 335560
rect 239676 335520 239682 335532
rect 240354 335520 240360 335532
rect 240412 335520 240418 335572
rect 240814 335520 240820 335572
rect 240872 335560 240878 335572
rect 241090 335560 241096 335572
rect 240872 335532 241096 335560
rect 240872 335520 240878 335532
rect 241090 335520 241096 335532
rect 241148 335520 241154 335572
rect 242378 335520 242384 335572
rect 242436 335560 242442 335572
rect 242562 335560 242568 335572
rect 242436 335532 242568 335560
rect 242436 335520 242442 335532
rect 242562 335520 242568 335532
rect 242620 335520 242626 335572
rect 244034 335520 244040 335572
rect 244092 335560 244098 335572
rect 244494 335560 244500 335572
rect 244092 335532 244500 335560
rect 244092 335520 244098 335532
rect 244494 335520 244500 335532
rect 244552 335520 244558 335572
rect 244862 335520 244868 335572
rect 244920 335560 244926 335572
rect 245506 335560 245512 335572
rect 244920 335532 245512 335560
rect 244920 335520 244926 335532
rect 245506 335520 245512 335532
rect 245564 335520 245570 335572
rect 247714 335520 247720 335572
rect 247772 335560 247778 335572
rect 248450 335560 248456 335572
rect 247772 335532 248456 335560
rect 247772 335520 247778 335532
rect 248450 335520 248456 335532
rect 248508 335520 248514 335572
rect 249002 335520 249008 335572
rect 249060 335560 249066 335572
rect 249922 335560 249928 335572
rect 249060 335532 249928 335560
rect 249060 335520 249066 335532
rect 249922 335520 249928 335532
rect 249980 335520 249986 335572
rect 253326 335520 253332 335572
rect 253384 335560 253390 335572
rect 253602 335560 253608 335572
rect 253384 335532 253608 335560
rect 253384 335520 253390 335532
rect 253602 335520 253608 335532
rect 253660 335520 253666 335572
rect 254706 335520 254712 335572
rect 254764 335560 254770 335572
rect 255258 335560 255264 335572
rect 254764 335532 255264 335560
rect 254764 335520 254770 335532
rect 255258 335520 255264 335532
rect 255316 335520 255322 335572
rect 257466 335520 257472 335572
rect 257524 335560 257530 335572
rect 258202 335560 258208 335572
rect 257524 335532 258208 335560
rect 257524 335520 257530 335532
rect 258202 335520 258208 335532
rect 258260 335520 258266 335572
rect 258754 335520 258760 335572
rect 258812 335560 258818 335572
rect 259490 335560 259496 335572
rect 258812 335532 259496 335560
rect 258812 335520 258818 335532
rect 259490 335520 259496 335532
rect 259548 335520 259554 335572
rect 260226 335520 260232 335572
rect 260284 335560 260290 335572
rect 260686 335560 260692 335572
rect 260284 335532 260692 335560
rect 260284 335520 260290 335532
rect 260686 335520 260692 335532
rect 260744 335520 260750 335572
rect 261698 335520 261704 335572
rect 261756 335560 261762 335572
rect 262342 335560 262348 335572
rect 261756 335532 262348 335560
rect 261756 335520 261762 335532
rect 262342 335520 262348 335532
rect 262400 335520 262406 335572
rect 262894 335520 262900 335572
rect 262952 335560 262958 335572
rect 263354 335560 263360 335572
rect 262952 335532 263360 335560
rect 262952 335520 262958 335532
rect 263354 335520 263360 335532
rect 263412 335520 263418 335572
rect 264090 335520 264096 335572
rect 264148 335560 264154 335572
rect 264366 335560 264372 335572
rect 264148 335532 264372 335560
rect 264148 335520 264154 335532
rect 264366 335520 264372 335532
rect 264424 335520 264430 335572
rect 265838 335520 265844 335572
rect 265896 335560 265902 335572
rect 266574 335560 266580 335572
rect 265896 335532 266580 335560
rect 265896 335520 265902 335532
rect 266574 335520 266580 335532
rect 266632 335520 266638 335572
rect 267126 335520 267132 335572
rect 267184 335560 267190 335572
rect 267770 335560 267776 335572
rect 267184 335532 267776 335560
rect 267184 335520 267190 335532
rect 267770 335520 267776 335532
rect 267828 335520 267834 335572
rect 268506 335520 268512 335572
rect 268564 335560 268570 335572
rect 269242 335560 269248 335572
rect 268564 335532 269248 335560
rect 268564 335520 268570 335532
rect 269242 335520 269248 335532
rect 269300 335520 269306 335572
rect 269978 335520 269984 335572
rect 270036 335560 270042 335572
rect 270714 335560 270720 335572
rect 270036 335532 270720 335560
rect 270036 335520 270042 335532
rect 270714 335520 270720 335532
rect 270772 335520 270778 335572
rect 274118 335520 274124 335572
rect 274176 335560 274182 335572
rect 274670 335560 274676 335572
rect 274176 335532 274676 335560
rect 274176 335520 274182 335532
rect 274670 335520 274676 335532
rect 274728 335520 274734 335572
rect 276786 335520 276792 335572
rect 276844 335560 276850 335572
rect 277338 335560 277344 335572
rect 276844 335532 277344 335560
rect 276844 335520 276850 335532
rect 277338 335520 277344 335532
rect 277396 335520 277402 335572
rect 278074 335520 278080 335572
rect 278132 335560 278138 335572
rect 278810 335560 278816 335572
rect 278132 335532 278816 335560
rect 278132 335520 278138 335532
rect 278810 335520 278816 335532
rect 278868 335520 278874 335572
rect 279270 335520 279276 335572
rect 279328 335560 279334 335572
rect 280282 335560 280288 335572
rect 279328 335532 280288 335560
rect 279328 335520 279334 335532
rect 280282 335520 280288 335532
rect 280340 335520 280346 335572
rect 280742 335520 280748 335572
rect 280800 335560 280806 335572
rect 281478 335560 281484 335572
rect 280800 335532 281484 335560
rect 280800 335520 280806 335532
rect 281478 335520 281484 335532
rect 281536 335520 281542 335572
rect 327846 335520 327852 335572
rect 327904 335560 327910 335572
rect 328674 335560 328680 335572
rect 327904 335532 328680 335560
rect 327904 335520 327910 335532
rect 328674 335520 328680 335532
rect 328732 335520 328738 335572
rect 333182 335520 333188 335572
rect 333240 335560 333246 335572
rect 334286 335560 334292 335572
rect 333240 335532 334292 335560
rect 333240 335520 333246 335532
rect 334286 335520 334292 335532
rect 334344 335520 334350 335572
rect 337966 335520 337972 335572
rect 338024 335560 338030 335572
rect 338426 335560 338432 335572
rect 338024 335532 338432 335560
rect 338024 335520 338030 335532
rect 338426 335520 338432 335532
rect 338484 335520 338490 335572
rect 231062 335452 231068 335504
rect 231120 335492 231126 335504
rect 231798 335492 231804 335504
rect 231120 335464 231804 335492
rect 231120 335452 231126 335464
rect 231798 335452 231804 335464
rect 231856 335452 231862 335504
rect 232718 335452 232724 335504
rect 232776 335492 232782 335504
rect 233270 335492 233276 335504
rect 232776 335464 233276 335492
rect 232776 335452 232782 335464
rect 233270 335452 233276 335464
rect 233328 335452 233334 335504
rect 237870 335452 237876 335504
rect 237928 335492 237934 335504
rect 238882 335492 238888 335504
rect 237928 335464 238888 335492
rect 237928 335452 237934 335464
rect 238882 335452 238888 335464
rect 238940 335452 238946 335504
rect 239434 335452 239440 335504
rect 239492 335492 239498 335504
rect 240078 335492 240084 335504
rect 239492 335464 240084 335492
rect 239492 335452 239498 335464
rect 240078 335452 240084 335464
rect 240136 335452 240142 335504
rect 242010 335452 242016 335504
rect 242068 335492 242074 335504
rect 242286 335492 242292 335504
rect 242068 335464 242292 335492
rect 242068 335452 242074 335464
rect 242286 335452 242292 335464
rect 242344 335452 242350 335504
rect 243574 335452 243580 335504
rect 243632 335492 243638 335504
rect 243942 335492 243948 335504
rect 243632 335464 243948 335492
rect 243632 335452 243638 335464
rect 243942 335452 243948 335464
rect 244000 335452 244006 335504
rect 270070 335452 270076 335504
rect 270128 335492 270134 335504
rect 270254 335492 270260 335504
rect 270128 335464 270260 335492
rect 270128 335452 270134 335464
rect 270254 335452 270260 335464
rect 270312 335452 270318 335504
rect 272646 335452 272652 335504
rect 272704 335492 272710 335504
rect 273382 335492 273388 335504
rect 272704 335464 273388 335492
rect 272704 335452 272710 335464
rect 273382 335452 273388 335464
rect 273440 335452 273446 335504
rect 284974 335452 284980 335504
rect 285032 335492 285038 335504
rect 285618 335492 285624 335504
rect 285032 335464 285624 335492
rect 285032 335452 285038 335464
rect 285618 335452 285624 335464
rect 285676 335452 285682 335504
rect 289022 335452 289028 335504
rect 289080 335492 289086 335504
rect 289666 335492 289672 335504
rect 289080 335464 289672 335492
rect 289080 335452 289086 335464
rect 289666 335452 289672 335464
rect 289724 335452 289730 335504
rect 313126 335452 313132 335504
rect 313184 335492 313190 335504
rect 313586 335492 313592 335504
rect 313184 335464 313592 335492
rect 313184 335452 313190 335464
rect 313586 335452 313592 335464
rect 313644 335452 313650 335504
rect 318002 335452 318008 335504
rect 318060 335492 318066 335504
rect 319198 335492 319204 335504
rect 318060 335464 319204 335492
rect 318060 335452 318066 335464
rect 319198 335452 319204 335464
rect 319256 335452 319262 335504
rect 319474 335452 319480 335504
rect 319532 335492 319538 335504
rect 320486 335492 320492 335504
rect 319532 335464 320492 335492
rect 319532 335452 319538 335464
rect 320486 335452 320492 335464
rect 320544 335452 320550 335504
rect 322142 335452 322148 335504
rect 322200 335492 322206 335504
rect 323062 335492 323068 335504
rect 322200 335464 323068 335492
rect 322200 335452 322206 335464
rect 323062 335452 323068 335464
rect 323120 335452 323126 335504
rect 240814 335384 240820 335436
rect 240872 335424 240878 335436
rect 241550 335424 241556 335436
rect 240872 335396 241556 335424
rect 240872 335384 240878 335396
rect 241550 335384 241556 335396
rect 241608 335384 241614 335436
rect 264366 335384 264372 335436
rect 264424 335424 264430 335436
rect 265102 335424 265108 335436
rect 264424 335396 265108 335424
rect 264424 335384 264430 335396
rect 265102 335384 265108 335396
rect 265160 335384 265166 335436
rect 250382 335316 250388 335368
rect 250440 335356 250446 335368
rect 251118 335356 251124 335368
rect 250440 335328 251124 335356
rect 250440 335316 250446 335328
rect 251118 335316 251124 335328
rect 251176 335316 251182 335368
rect 251854 335316 251860 335368
rect 251912 335356 251918 335368
rect 252590 335356 252596 335368
rect 251912 335328 252596 335356
rect 251912 335316 251918 335328
rect 252590 335316 252596 335328
rect 252648 335316 252654 335368
rect 338794 335316 338800 335368
rect 338852 335356 338858 335368
rect 339806 335356 339812 335368
rect 338852 335328 339812 335356
rect 338852 335316 338858 335328
rect 339806 335316 339812 335328
rect 339864 335316 339870 335368
rect 250474 335248 250480 335300
rect 250532 335288 250538 335300
rect 250750 335288 250756 335300
rect 250532 335260 250756 335288
rect 250532 335248 250538 335260
rect 250750 335248 250756 335260
rect 250808 335248 250814 335300
rect 251946 335248 251952 335300
rect 252004 335288 252010 335300
rect 252406 335288 252412 335300
rect 252004 335260 252412 335288
rect 252004 335248 252010 335260
rect 252406 335248 252412 335260
rect 252464 335248 252470 335300
rect 277062 335248 277068 335300
rect 277120 335288 277126 335300
rect 277522 335288 277528 335300
rect 277120 335260 277528 335288
rect 277120 335248 277126 335260
rect 277522 335248 277528 335260
rect 277580 335248 277586 335300
rect 319934 335288 319940 335300
rect 319895 335260 319940 335288
rect 319934 335248 319940 335260
rect 319992 335248 319998 335300
rect 1600 335056 583316 335152
rect 263170 334908 263176 334960
rect 263228 334948 263234 334960
rect 263814 334948 263820 334960
rect 263228 334920 263820 334948
rect 263228 334908 263234 334920
rect 263814 334908 263820 334920
rect 263872 334908 263878 334960
rect 305582 334704 305588 334756
rect 305640 334744 305646 334756
rect 366210 334744 366216 334756
rect 305640 334716 366216 334744
rect 305640 334704 305646 334716
rect 366210 334704 366216 334716
rect 366268 334704 366274 334756
rect 152221 334679 152279 334685
rect 152221 334645 152233 334679
rect 152267 334676 152279 334679
rect 261514 334676 261520 334688
rect 152267 334648 261520 334676
rect 152267 334645 152279 334648
rect 152221 334639 152279 334645
rect 261514 334636 261520 334648
rect 261572 334636 261578 334688
rect 342750 334636 342756 334688
rect 342808 334676 342814 334688
rect 548370 334676 548376 334688
rect 342808 334648 548376 334676
rect 342808 334636 342814 334648
rect 548370 334636 548376 334648
rect 548428 334636 548434 334688
rect 1600 334512 583316 334608
rect 279825 334339 279883 334345
rect 279825 334305 279837 334339
rect 279871 334336 279883 334339
rect 280006 334336 280012 334348
rect 279871 334308 280012 334336
rect 279871 334305 279883 334308
rect 279825 334299 279883 334305
rect 280006 334296 280012 334308
rect 280064 334296 280070 334348
rect 1600 333968 583316 334064
rect 276510 333888 276516 333940
rect 276568 333928 276574 333940
rect 276568 333900 276613 333928
rect 276568 333888 276574 333900
rect 236674 333548 236680 333600
rect 236732 333588 236738 333600
rect 237410 333588 237416 333600
rect 236732 333560 237416 333588
rect 236732 333548 236738 333560
rect 237410 333548 237416 333560
rect 237468 333548 237474 333600
rect 1600 333424 583316 333520
rect 204658 333344 204664 333396
rect 204716 333384 204722 333396
rect 272370 333384 272376 333396
rect 204716 333356 272376 333384
rect 204716 333344 204722 333356
rect 272370 333344 272376 333356
rect 272428 333344 272434 333396
rect 303098 333344 303104 333396
rect 303156 333384 303162 333396
rect 353790 333384 353796 333396
rect 303156 333356 353796 333384
rect 303156 333344 303162 333356
rect 353790 333344 353796 333356
rect 353848 333344 353854 333396
rect 163258 333276 163264 333328
rect 163316 333316 163322 333328
rect 263722 333316 263728 333328
rect 163316 333288 263728 333316
rect 163316 333276 163322 333288
rect 263722 333276 263728 333288
rect 263780 333276 263786 333328
rect 284882 333276 284888 333328
rect 284940 333316 284946 333328
rect 285158 333316 285164 333328
rect 284940 333288 285164 333316
rect 284940 333276 284946 333288
rect 285158 333276 285164 333288
rect 285216 333276 285222 333328
rect 329870 333276 329876 333328
rect 329928 333316 329934 333328
rect 483510 333316 483516 333328
rect 329928 333288 483516 333316
rect 329928 333276 329934 333288
rect 483510 333276 483516 333288
rect 483568 333276 483574 333328
rect 145318 333208 145324 333260
rect 145376 333248 145382 333260
rect 260134 333248 260140 333260
rect 145376 333220 260140 333248
rect 145376 333208 145382 333220
rect 260134 333208 260140 333220
rect 260192 333208 260198 333260
rect 262618 333208 262624 333260
rect 262676 333248 262682 333260
rect 270901 333251 270959 333257
rect 270901 333248 270913 333251
rect 262676 333220 270913 333248
rect 262676 333208 262682 333220
rect 270901 333217 270913 333220
rect 270947 333217 270959 333251
rect 270901 333211 270959 333217
rect 348822 333208 348828 333260
rect 348880 333248 348886 333260
rect 575970 333248 575976 333260
rect 348880 333220 575976 333248
rect 348880 333208 348886 333220
rect 575970 333208 575976 333220
rect 576028 333208 576034 333260
rect 1600 332880 583316 332976
rect 279362 332800 279368 332852
rect 279420 332840 279426 332852
rect 279730 332840 279736 332852
rect 279420 332812 279736 332840
rect 279420 332800 279426 332812
rect 279730 332800 279736 332812
rect 279788 332800 279794 332852
rect 1600 332336 583316 332432
rect 214321 332027 214379 332033
rect 214321 331993 214333 332027
rect 214367 332024 214379 332027
rect 274302 332024 274308 332036
rect 214367 331996 274308 332024
rect 214367 331993 214379 331996
rect 214321 331987 214379 331993
rect 274302 331984 274308 331996
rect 274360 331984 274366 332036
rect 287918 331984 287924 332036
rect 287976 332024 287982 332036
rect 288378 332024 288384 332036
rect 287976 331996 288384 332024
rect 287976 331984 287982 331996
rect 288378 331984 288384 331996
rect 288436 331984 288442 332036
rect 307054 331984 307060 332036
rect 307112 332024 307118 332036
rect 373018 332024 373024 332036
rect 307112 331996 373024 332024
rect 307112 331984 307118 331996
rect 373018 331984 373024 331996
rect 373076 331984 373082 332036
rect 117718 331916 117724 331968
rect 117776 331956 117782 331968
rect 254430 331956 254436 331968
rect 117776 331928 254436 331956
rect 117776 331916 117782 331928
rect 254430 331916 254436 331928
rect 254488 331916 254494 331968
rect 278721 331959 278779 331965
rect 278721 331925 278733 331959
rect 278767 331956 278779 331959
rect 278810 331956 278816 331968
rect 278767 331928 278816 331956
rect 278767 331925 278779 331928
rect 278721 331919 278779 331925
rect 278810 331916 278816 331928
rect 278868 331916 278874 331968
rect 337690 331916 337696 331968
rect 337748 331956 337754 331968
rect 520770 331956 520776 331968
rect 337748 331928 520776 331956
rect 337748 331916 337754 331928
rect 520770 331916 520776 331928
rect 520828 331916 520834 331968
rect 1600 331792 583316 331888
rect 282306 331576 282312 331628
rect 282364 331616 282370 331628
rect 283226 331616 283232 331628
rect 282364 331588 283232 331616
rect 282364 331576 282370 331588
rect 283226 331576 283232 331588
rect 283284 331576 283290 331628
rect 285345 331483 285403 331489
rect 285345 331449 285357 331483
rect 285391 331480 285403 331483
rect 285434 331480 285440 331492
rect 285391 331452 285440 331480
rect 285391 331449 285403 331452
rect 285345 331443 285403 331449
rect 285434 331440 285440 331452
rect 285492 331440 285498 331492
rect 259033 331415 259091 331421
rect 259033 331381 259045 331415
rect 259079 331412 259091 331415
rect 259122 331412 259128 331424
rect 259079 331384 259128 331412
rect 259079 331381 259091 331384
rect 259033 331375 259091 331381
rect 259122 331372 259128 331384
rect 259180 331372 259186 331424
rect 1600 331248 583316 331344
rect 254706 331168 254712 331220
rect 254764 331208 254770 331220
rect 254890 331208 254896 331220
rect 254764 331180 254896 331208
rect 254764 331168 254770 331180
rect 254890 331168 254896 331180
rect 254948 331168 254954 331220
rect 259030 331208 259036 331220
rect 258991 331180 259036 331208
rect 259030 331168 259036 331180
rect 259088 331168 259094 331220
rect 340818 331168 340824 331220
rect 340876 331208 340882 331220
rect 341186 331208 341192 331220
rect 340876 331180 341192 331208
rect 340876 331168 340882 331180
rect 341186 331168 341192 331180
rect 341244 331168 341250 331220
rect 259122 331140 259128 331152
rect 259083 331112 259128 331140
rect 259122 331100 259128 331112
rect 259180 331100 259186 331152
rect 284977 331143 285035 331149
rect 284977 331109 284989 331143
rect 285023 331140 285035 331143
rect 285158 331140 285164 331152
rect 285023 331112 285164 331140
rect 285023 331109 285035 331112
rect 284977 331103 285035 331109
rect 285158 331100 285164 331112
rect 285216 331100 285222 331152
rect 285434 331100 285440 331152
rect 285492 331140 285498 331152
rect 288746 331140 288752 331152
rect 285492 331112 288752 331140
rect 285492 331100 285498 331112
rect 288746 331100 288752 331112
rect 288804 331100 288810 331152
rect 371914 331140 371920 331152
rect 371875 331112 371920 331140
rect 371914 331100 371920 331112
rect 371972 331100 371978 331152
rect 246426 331032 246432 331084
rect 246484 331072 246490 331084
rect 246702 331072 246708 331084
rect 246484 331044 246708 331072
rect 246484 331032 246490 331044
rect 246702 331032 246708 331044
rect 246760 331032 246766 331084
rect 271358 331032 271364 331084
rect 271416 331072 271422 331084
rect 271726 331072 271732 331084
rect 271416 331044 271732 331072
rect 271416 331032 271422 331044
rect 271726 331032 271732 331044
rect 271784 331032 271790 331084
rect 1600 330704 583316 330800
rect 167398 330624 167404 330676
rect 167456 330664 167462 330676
rect 264090 330664 264096 330676
rect 167456 330636 264096 330664
rect 167456 330624 167462 330636
rect 264090 330624 264096 330636
rect 264148 330624 264154 330676
rect 303558 330624 303564 330676
rect 303616 330664 303622 330676
rect 355170 330664 355176 330676
rect 303616 330636 355176 330664
rect 303616 330624 303622 330636
rect 355170 330624 355176 330636
rect 355228 330624 355234 330676
rect 156358 330556 156364 330608
rect 156416 330596 156422 330608
rect 262066 330596 262072 330608
rect 156416 330568 262072 330596
rect 156416 330556 156422 330568
rect 262066 330556 262072 330568
rect 262124 330556 262130 330608
rect 330514 330556 330520 330608
rect 330572 330596 330578 330608
rect 486270 330596 486276 330608
rect 330572 330568 486276 330596
rect 330572 330556 330578 330568
rect 486270 330556 486276 330568
rect 486328 330556 486334 330608
rect 23878 330488 23884 330540
rect 23936 330528 23942 330540
rect 235110 330528 235116 330540
rect 23936 330500 235116 330528
rect 23936 330488 23942 330500
rect 235110 330488 235116 330500
rect 235168 330488 235174 330540
rect 342014 330488 342020 330540
rect 342072 330528 342078 330540
rect 342382 330528 342388 330540
rect 342072 330500 342388 330528
rect 342072 330488 342078 330500
rect 342382 330488 342388 330500
rect 342440 330488 342446 330540
rect 530430 330528 530436 330540
rect 342492 330500 530436 330528
rect 339346 330420 339352 330472
rect 339404 330460 339410 330472
rect 342492 330460 342520 330500
rect 530430 330488 530436 330500
rect 530488 330488 530494 330540
rect 339404 330432 342520 330460
rect 339404 330420 339410 330432
rect 1600 330160 583316 330256
rect 1600 329616 583316 329712
rect 221218 329196 221224 329248
rect 221276 329236 221282 329248
rect 275130 329236 275136 329248
rect 221276 329208 275136 329236
rect 221276 329196 221282 329208
rect 275130 329196 275136 329208
rect 275188 329196 275194 329248
rect 322510 329196 322516 329248
rect 322568 329236 322574 329248
rect 447630 329236 447636 329248
rect 322568 329208 447636 329236
rect 322568 329196 322574 329208
rect 447630 329196 447636 329208
rect 447688 329196 447694 329248
rect 1600 329072 583316 329168
rect 1600 328528 583316 328624
rect 252498 328448 252504 328500
rect 252556 328488 252562 328500
rect 252866 328488 252872 328500
rect 252556 328460 252872 328488
rect 252556 328448 252562 328460
rect 252866 328448 252872 328460
rect 252924 328448 252930 328500
rect 259306 328448 259312 328500
rect 259364 328488 259370 328500
rect 259766 328488 259772 328500
rect 259364 328460 259772 328488
rect 259364 328448 259370 328460
rect 259766 328448 259772 328460
rect 259824 328448 259830 328500
rect 285342 328488 285348 328500
rect 285303 328460 285348 328488
rect 285342 328448 285348 328460
rect 285400 328448 285406 328500
rect 285710 328448 285716 328500
rect 285768 328488 285774 328500
rect 285986 328488 285992 328500
rect 285768 328460 285992 328488
rect 285768 328448 285774 328460
rect 285986 328448 285992 328460
rect 286044 328448 286050 328500
rect 333366 328448 333372 328500
rect 333424 328488 333430 328500
rect 333918 328488 333924 328500
rect 333424 328460 333924 328488
rect 333424 328448 333430 328460
rect 333918 328448 333924 328460
rect 333976 328448 333982 328500
rect 229869 328423 229927 328429
rect 229869 328389 229881 328423
rect 229915 328420 229927 328423
rect 229958 328420 229964 328432
rect 229915 328392 229964 328420
rect 229915 328389 229927 328392
rect 229869 328383 229927 328389
rect 229958 328380 229964 328392
rect 230016 328380 230022 328432
rect 235481 328423 235539 328429
rect 235481 328389 235493 328423
rect 235527 328420 235539 328423
rect 235570 328420 235576 328432
rect 235527 328392 235576 328420
rect 235527 328389 235539 328392
rect 235481 328383 235539 328389
rect 235570 328380 235576 328392
rect 235628 328380 235634 328432
rect 268598 328420 268604 328432
rect 268559 328392 268604 328420
rect 268598 328380 268604 328392
rect 268656 328380 268662 328432
rect 318646 328420 318652 328432
rect 318607 328392 318652 328420
rect 318646 328380 318652 328392
rect 318704 328380 318710 328432
rect 328122 328380 328128 328432
rect 328180 328420 328186 328432
rect 328214 328420 328220 328432
rect 328180 328392 328220 328420
rect 328180 328380 328186 328392
rect 328214 328380 328220 328392
rect 328272 328380 328278 328432
rect 371914 328420 371920 328432
rect 371875 328392 371920 328420
rect 371914 328380 371920 328392
rect 371972 328380 371978 328432
rect 1600 327984 583316 328080
rect 218458 327836 218464 327888
rect 218516 327876 218522 327888
rect 273750 327876 273756 327888
rect 218516 327848 273756 327876
rect 218516 327836 218522 327848
rect 273750 327836 273756 327848
rect 273808 327836 273814 327888
rect 305122 327836 305128 327888
rect 305180 327876 305186 327888
rect 362070 327876 362076 327888
rect 305180 327848 362076 327876
rect 305180 327836 305186 327848
rect 362070 327836 362076 327848
rect 362128 327836 362134 327888
rect 170161 327811 170219 327817
rect 170161 327777 170173 327811
rect 170207 327808 170219 327811
rect 264366 327808 264372 327820
rect 170207 327780 264372 327808
rect 170207 327777 170219 327780
rect 170161 327771 170219 327777
rect 264366 327768 264372 327780
rect 264424 327768 264430 327820
rect 331250 327768 331256 327820
rect 331308 327808 331314 327820
rect 490410 327808 490416 327820
rect 331308 327780 490416 327808
rect 331308 327768 331314 327780
rect 490410 327768 490416 327780
rect 490468 327768 490474 327820
rect 77698 327700 77704 327752
rect 77756 327740 77762 327752
rect 246150 327740 246156 327752
rect 77756 327712 246156 327740
rect 77756 327700 77762 327712
rect 246150 327700 246156 327712
rect 246208 327700 246214 327752
rect 341830 327700 341836 327752
rect 341888 327740 341894 327752
rect 541470 327740 541476 327752
rect 341888 327712 541476 327740
rect 341888 327700 341894 327712
rect 541470 327700 541476 327712
rect 541528 327700 541534 327752
rect 1600 327440 583316 327536
rect 152218 327128 152224 327140
rect 152179 327100 152224 327128
rect 152218 327088 152224 327100
rect 152276 327088 152282 327140
rect 170158 327128 170164 327140
rect 170119 327100 170164 327128
rect 170158 327088 170164 327100
rect 170216 327088 170222 327140
rect 214318 327128 214324 327140
rect 214279 327100 214324 327128
rect 214318 327088 214324 327100
rect 214376 327088 214382 327140
rect 246518 327088 246524 327140
rect 246576 327128 246582 327140
rect 246702 327128 246708 327140
rect 246576 327100 246708 327128
rect 246576 327088 246582 327100
rect 246702 327088 246708 327100
rect 246760 327088 246766 327140
rect 279822 327128 279828 327140
rect 279783 327100 279828 327128
rect 279822 327088 279828 327100
rect 279880 327088 279886 327140
rect 392246 327088 392252 327140
rect 392304 327128 392310 327140
rect 392430 327128 392436 327140
rect 392304 327100 392436 327128
rect 392304 327088 392310 327100
rect 392430 327088 392436 327100
rect 392488 327088 392494 327140
rect 328122 327060 328128 327072
rect 328083 327032 328128 327060
rect 328122 327020 328128 327032
rect 328180 327020 328186 327072
rect 373018 327060 373024 327072
rect 372979 327032 373024 327060
rect 373018 327020 373024 327032
rect 373076 327020 373082 327072
rect 1600 326896 583316 326992
rect 278718 326856 278724 326868
rect 278679 326828 278724 326856
rect 278718 326816 278724 326828
rect 278776 326816 278782 326868
rect 186718 326476 186724 326528
rect 186776 326516 186782 326528
rect 268230 326516 268236 326528
rect 186776 326488 268236 326516
rect 186776 326476 186782 326488
rect 268230 326476 268236 326488
rect 268288 326476 268294 326528
rect 327018 326476 327024 326528
rect 327076 326516 327082 326528
rect 465570 326516 465576 326528
rect 327076 326488 465576 326516
rect 327076 326476 327082 326488
rect 465570 326476 465576 326488
rect 465628 326476 465634 326528
rect 1600 326352 583316 326448
rect 1600 325808 583316 325904
rect 1600 325264 583316 325360
rect 229498 325048 229504 325100
rect 229556 325088 229562 325100
rect 276878 325088 276884 325100
rect 229556 325060 276884 325088
rect 229556 325048 229562 325060
rect 276878 325048 276884 325060
rect 276936 325048 276942 325100
rect 306502 325048 306508 325100
rect 306560 325088 306566 325100
rect 368970 325088 368976 325100
rect 306560 325060 368976 325088
rect 306560 325048 306566 325060
rect 368970 325048 368976 325060
rect 369028 325048 369034 325100
rect 174298 324980 174304 325032
rect 174356 325020 174362 325032
rect 265930 325020 265936 325032
rect 174356 324992 265936 325020
rect 174356 324980 174362 324992
rect 265930 324980 265936 324992
rect 265988 324980 265994 325032
rect 332630 324980 332636 325032
rect 332688 325020 332694 325032
rect 494550 325020 494556 325032
rect 332688 324992 494556 325020
rect 332688 324980 332694 324992
rect 494550 324980 494556 324992
rect 494608 324980 494614 325032
rect 73558 324912 73564 324964
rect 73616 324952 73622 324964
rect 245046 324952 245052 324964
rect 73616 324924 245052 324952
rect 73616 324912 73622 324924
rect 245046 324912 245052 324924
rect 245104 324912 245110 324964
rect 345050 324912 345056 324964
rect 345108 324952 345114 324964
rect 553890 324952 553896 324964
rect 345108 324924 553896 324952
rect 345108 324912 345114 324924
rect 553890 324912 553896 324924
rect 553948 324912 553954 324964
rect 1600 324720 583316 324816
rect 275774 324368 275780 324420
rect 275832 324408 275838 324420
rect 276142 324408 276148 324420
rect 275832 324380 276148 324408
rect 275832 324368 275838 324380
rect 276142 324368 276148 324380
rect 276200 324368 276206 324420
rect 276513 324411 276571 324417
rect 276513 324377 276525 324411
rect 276559 324408 276571 324411
rect 276602 324408 276608 324420
rect 276559 324380 276608 324408
rect 276559 324377 276571 324380
rect 276513 324371 276571 324377
rect 276602 324368 276608 324380
rect 276660 324368 276666 324420
rect 272922 324300 272928 324352
rect 272980 324340 272986 324352
rect 273014 324340 273020 324352
rect 272980 324312 273020 324340
rect 272980 324300 272986 324312
rect 273014 324300 273020 324312
rect 273072 324300 273078 324352
rect 275682 324300 275688 324352
rect 275740 324340 275746 324352
rect 275958 324340 275964 324352
rect 275740 324312 275964 324340
rect 275740 324300 275746 324312
rect 275958 324300 275964 324312
rect 276016 324300 276022 324352
rect 1600 324176 583316 324272
rect 1600 323632 583316 323728
rect 194906 323552 194912 323604
rect 194964 323592 194970 323604
rect 270162 323592 270168 323604
rect 194964 323564 270168 323592
rect 194964 323552 194970 323564
rect 270162 323552 270168 323564
rect 270220 323552 270226 323604
rect 313310 323552 313316 323604
rect 313368 323592 313374 323604
rect 399330 323592 399336 323604
rect 313368 323564 399336 323592
rect 313368 323552 313374 323564
rect 399330 323552 399336 323564
rect 399388 323552 399394 323604
rect 1600 323088 583316 323184
rect 1600 322544 583316 322640
rect 177058 322260 177064 322312
rect 177116 322300 177122 322312
rect 265838 322300 265844 322312
rect 177116 322272 265844 322300
rect 177116 322260 177122 322272
rect 265838 322260 265844 322272
rect 265896 322260 265902 322312
rect 332722 322260 332728 322312
rect 332780 322300 332786 322312
rect 497310 322300 497316 322312
rect 332780 322272 497316 322300
rect 332780 322260 332786 322272
rect 497310 322260 497316 322272
rect 497368 322260 497374 322312
rect 135658 322192 135664 322244
rect 135716 322232 135722 322244
rect 257926 322232 257932 322244
rect 135716 322204 257932 322232
rect 135716 322192 135722 322204
rect 257926 322192 257932 322204
rect 257984 322192 257990 322244
rect 299510 322192 299516 322244
rect 299568 322232 299574 322244
rect 331710 322232 331716 322244
rect 299568 322204 331716 322232
rect 299568 322192 299574 322204
rect 331710 322192 331716 322204
rect 331768 322192 331774 322244
rect 343670 322192 343676 322244
rect 343728 322232 343734 322244
rect 552510 322232 552516 322244
rect 343728 322204 552516 322232
rect 343728 322192 343734 322204
rect 552510 322192 552516 322204
rect 552568 322192 552574 322244
rect 1600 322000 583316 322096
rect 235665 321963 235723 321969
rect 235665 321929 235677 321963
rect 235711 321960 235723 321963
rect 235754 321960 235760 321972
rect 235711 321932 235760 321960
rect 235711 321929 235723 321932
rect 235665 321923 235723 321929
rect 235754 321920 235760 321932
rect 235812 321920 235818 321972
rect 239250 321580 239256 321632
rect 239308 321620 239314 321632
rect 239434 321620 239440 321632
rect 239308 321592 239440 321620
rect 239308 321580 239314 321592
rect 239434 321580 239440 321592
rect 239492 321580 239498 321632
rect 258938 321580 258944 321632
rect 258996 321620 259002 321632
rect 259122 321620 259128 321632
rect 258996 321592 259128 321620
rect 258996 321580 259002 321592
rect 259122 321580 259128 321592
rect 259180 321580 259186 321632
rect 272554 321580 272560 321632
rect 272612 321620 272618 321632
rect 272738 321620 272744 321632
rect 272612 321592 272744 321620
rect 272612 321580 272618 321592
rect 272738 321580 272744 321592
rect 272796 321580 272802 321632
rect 340818 321580 340824 321632
rect 340876 321620 340882 321632
rect 341186 321620 341192 321632
rect 340876 321592 341192 321620
rect 340876 321580 340882 321592
rect 341186 321580 341192 321592
rect 341244 321580 341250 321632
rect 1600 321456 583316 321552
rect 229866 321416 229872 321428
rect 229827 321388 229872 321416
rect 229866 321376 229872 321388
rect 229924 321376 229930 321428
rect 268601 321419 268659 321425
rect 268601 321385 268613 321419
rect 268647 321416 268659 321419
rect 268690 321416 268696 321428
rect 268647 321388 268696 321416
rect 268647 321385 268659 321388
rect 268601 321379 268659 321385
rect 268690 321376 268696 321388
rect 268748 321376 268754 321428
rect 318646 321416 318652 321428
rect 318607 321388 318652 321416
rect 318646 321376 318652 321388
rect 318704 321376 318710 321428
rect 340818 321376 340824 321428
rect 340876 321416 340882 321428
rect 341186 321416 341192 321428
rect 340876 321388 341192 321416
rect 340876 321376 340882 321388
rect 341186 321376 341192 321388
rect 341244 321376 341250 321428
rect 371914 321416 371920 321428
rect 371875 321388 371920 321416
rect 371914 321376 371920 321388
rect 371972 321376 371978 321428
rect 1600 320912 583316 321008
rect 110818 320832 110824 320884
rect 110876 320872 110882 320884
rect 252498 320872 252504 320884
rect 110876 320844 252504 320872
rect 110876 320832 110882 320844
rect 252498 320832 252504 320844
rect 252556 320832 252562 320884
rect 261238 320668 261244 320680
rect 261199 320640 261244 320668
rect 261238 320628 261244 320640
rect 261296 320628 261302 320680
rect 254154 320492 254160 320544
rect 254212 320532 254218 320544
rect 261146 320532 261152 320544
rect 254212 320504 261152 320532
rect 254212 320492 254218 320504
rect 261146 320492 261152 320504
rect 261204 320492 261210 320544
rect 488294 320492 488300 320544
rect 488352 320532 488358 320544
rect 493078 320532 493084 320544
rect 488352 320504 493084 320532
rect 488352 320492 488358 320504
rect 493078 320492 493084 320504
rect 493136 320492 493142 320544
rect 1600 320368 583316 320464
rect 418558 320288 418564 320340
rect 418616 320328 418622 320340
rect 425458 320328 425464 320340
rect 418616 320300 425464 320328
rect 418616 320288 418622 320300
rect 425458 320288 425464 320300
rect 425516 320288 425522 320340
rect 437878 320288 437884 320340
rect 437936 320328 437942 320340
rect 444778 320328 444784 320340
rect 437936 320300 444784 320328
rect 437936 320288 437942 320300
rect 444778 320288 444784 320300
rect 444836 320288 444842 320340
rect 457198 320288 457204 320340
rect 457256 320328 457262 320340
rect 464098 320328 464104 320340
rect 457256 320300 464104 320328
rect 457256 320288 457262 320300
rect 464098 320288 464104 320300
rect 464156 320288 464162 320340
rect 476518 320288 476524 320340
rect 476576 320328 476582 320340
rect 483418 320328 483424 320340
rect 476576 320300 483424 320328
rect 476576 320288 476582 320300
rect 483418 320288 483424 320300
rect 483476 320288 483482 320340
rect 541562 320288 541568 320340
rect 541620 320328 541626 320340
rect 544322 320328 544328 320340
rect 541620 320300 544328 320328
rect 541620 320288 541626 320300
rect 544322 320288 544328 320300
rect 544380 320288 544386 320340
rect 261238 320260 261244 320272
rect 261199 320232 261244 320260
rect 261238 320220 261244 320232
rect 261296 320220 261302 320272
rect 290310 320220 290316 320272
rect 290368 320260 290374 320272
rect 294634 320260 294640 320272
rect 290368 320232 294640 320260
rect 290368 320220 290374 320232
rect 294634 320220 294640 320232
rect 294692 320220 294698 320272
rect 1600 319824 583316 319920
rect 311930 319540 311936 319592
rect 311988 319580 311994 319592
rect 395190 319580 395196 319592
rect 311988 319552 395196 319580
rect 311988 319540 311994 319552
rect 395190 319540 395196 319552
rect 395248 319540 395254 319592
rect 185338 319472 185344 319524
rect 185396 319512 185402 319524
rect 267586 319512 267592 319524
rect 185396 319484 267592 319512
rect 185396 319472 185402 319484
rect 267586 319472 267592 319484
rect 267644 319472 267650 319524
rect 333918 319472 333924 319524
rect 333976 319512 333982 319524
rect 501450 319512 501456 319524
rect 333976 319484 501456 319512
rect 333976 319472 333982 319484
rect 501450 319472 501456 319484
rect 501508 319472 501514 319524
rect 134186 319404 134192 319456
rect 134244 319444 134250 319456
rect 257558 319444 257564 319456
rect 134244 319416 257564 319444
rect 134244 319404 134250 319416
rect 257558 319404 257564 319416
rect 257616 319404 257622 319456
rect 346338 319404 346344 319456
rect 346396 319444 346402 319456
rect 560790 319444 560796 319456
rect 346396 319416 560796 319444
rect 346396 319404 346402 319416
rect 560790 319404 560796 319416
rect 560848 319404 560854 319456
rect 1600 319280 583316 319376
rect 235478 318900 235484 318912
rect 235439 318872 235484 318900
rect 235478 318860 235484 318872
rect 235536 318860 235542 318912
rect 235662 318900 235668 318912
rect 235623 318872 235668 318900
rect 235662 318860 235668 318872
rect 235720 318860 235726 318912
rect 276973 318903 277031 318909
rect 276973 318869 276985 318903
rect 277019 318900 277031 318903
rect 277062 318900 277068 318912
rect 277019 318872 277068 318900
rect 277019 318869 277031 318872
rect 276973 318863 277031 318869
rect 277062 318860 277068 318872
rect 277120 318860 277126 318912
rect 1600 318736 583316 318832
rect 235478 318696 235484 318708
rect 235439 318668 235484 318696
rect 235478 318656 235484 318668
rect 235536 318656 235542 318708
rect 235662 318656 235668 318708
rect 235720 318696 235726 318708
rect 235938 318696 235944 318708
rect 235720 318668 235944 318696
rect 235720 318656 235726 318668
rect 235938 318656 235944 318668
rect 235996 318656 236002 318708
rect 276970 318696 276976 318708
rect 276931 318668 276976 318696
rect 276970 318656 276976 318668
rect 277028 318656 277034 318708
rect 285250 318696 285256 318708
rect 285211 318668 285256 318696
rect 285250 318656 285256 318668
rect 285308 318656 285314 318708
rect 285618 318696 285624 318708
rect 285579 318668 285624 318696
rect 285618 318656 285624 318668
rect 285676 318656 285682 318708
rect 318922 318696 318928 318708
rect 318883 318668 318928 318696
rect 318922 318656 318928 318668
rect 318980 318656 318986 318708
rect 319106 318696 319112 318708
rect 319067 318668 319112 318696
rect 319106 318656 319112 318668
rect 319164 318656 319170 318708
rect 373021 318699 373079 318705
rect 373021 318665 373033 318699
rect 373067 318696 373079 318699
rect 373110 318696 373116 318708
rect 373067 318668 373116 318696
rect 373067 318665 373079 318668
rect 373021 318659 373079 318665
rect 373110 318656 373116 318668
rect 373168 318656 373174 318708
rect 319198 318588 319204 318640
rect 319256 318588 319262 318640
rect 319216 318504 319244 318588
rect 319198 318452 319204 318504
rect 319256 318452 319262 318504
rect 1600 318192 583316 318288
rect 197758 318112 197764 318164
rect 197816 318152 197822 318164
rect 269978 318152 269984 318164
rect 197816 318124 269984 318152
rect 197816 318112 197822 318124
rect 269978 318112 269984 318124
rect 270036 318112 270042 318164
rect 314782 318112 314788 318164
rect 314840 318152 314846 318164
rect 406230 318152 406236 318164
rect 314840 318124 406236 318152
rect 314840 318112 314846 318124
rect 406230 318112 406236 318124
rect 406288 318112 406294 318164
rect 138418 318044 138424 318096
rect 138476 318084 138482 318096
rect 256454 318084 256460 318096
rect 138476 318056 256460 318084
rect 138476 318044 138482 318056
rect 256454 318044 256460 318056
rect 256512 318044 256518 318096
rect 334010 318044 334016 318096
rect 334068 318084 334074 318096
rect 504210 318084 504216 318096
rect 334068 318056 504216 318084
rect 334068 318044 334074 318056
rect 504210 318044 504216 318056
rect 504268 318044 504274 318096
rect 1600 317648 583316 317744
rect 319937 317475 319995 317481
rect 319937 317441 319949 317475
rect 319983 317472 319995 317475
rect 320118 317472 320124 317484
rect 319983 317444 320124 317472
rect 319983 317441 319995 317444
rect 319937 317435 319995 317441
rect 320118 317432 320124 317444
rect 320176 317432 320182 317484
rect 328125 317475 328183 317481
rect 328125 317441 328137 317475
rect 328171 317472 328183 317475
rect 328398 317472 328404 317484
rect 328171 317444 328404 317472
rect 328171 317441 328183 317444
rect 328125 317435 328183 317441
rect 328398 317432 328404 317444
rect 328456 317432 328462 317484
rect 135658 317404 135664 317416
rect 135619 317376 135664 317404
rect 135658 317364 135664 317376
rect 135716 317364 135722 317416
rect 152218 317404 152224 317416
rect 152179 317376 152224 317404
rect 152218 317364 152224 317376
rect 152276 317364 152282 317416
rect 170158 317404 170164 317416
rect 170119 317376 170164 317404
rect 170158 317364 170164 317376
rect 170216 317364 170222 317416
rect 214318 317404 214324 317416
rect 214279 317376 214324 317404
rect 214318 317364 214324 317376
rect 214376 317364 214382 317416
rect 385530 317364 385536 317416
rect 385588 317404 385594 317416
rect 392430 317404 392436 317416
rect 385588 317376 385633 317404
rect 392391 317376 392436 317404
rect 385588 317364 385594 317376
rect 392430 317364 392436 317376
rect 392488 317364 392494 317416
rect 1600 317104 583316 317200
rect 342198 316752 342204 316804
rect 342256 316792 342262 316804
rect 342382 316792 342388 316804
rect 342256 316764 342388 316792
rect 342256 316752 342262 316764
rect 342382 316752 342388 316764
rect 342440 316752 342446 316804
rect 121858 316684 121864 316736
rect 121916 316724 121922 316736
rect 254798 316724 254804 316736
rect 121916 316696 254804 316724
rect 121916 316684 121922 316696
rect 254798 316684 254804 316696
rect 254856 316684 254862 316736
rect 317450 316684 317456 316736
rect 317508 316724 317514 316736
rect 420030 316724 420036 316736
rect 317508 316696 420036 316724
rect 317508 316684 317514 316696
rect 420030 316684 420036 316696
rect 420088 316684 420094 316736
rect 1600 316560 583316 316656
rect 1600 316016 583316 316112
rect 1600 315472 583316 315568
rect 201898 315324 201904 315376
rect 201956 315364 201962 315376
rect 271634 315364 271640 315376
rect 201956 315336 271640 315364
rect 201956 315324 201962 315336
rect 271634 315324 271640 315336
rect 271692 315324 271698 315376
rect 316070 315324 316076 315376
rect 316128 315364 316134 315376
rect 413130 315364 413136 315376
rect 316128 315336 413136 315364
rect 316128 315324 316134 315336
rect 413130 315324 413136 315336
rect 413188 315324 413194 315376
rect 142558 315256 142564 315308
rect 142616 315296 142622 315308
rect 258938 315296 258944 315308
rect 142616 315268 258944 315296
rect 142616 315256 142622 315268
rect 258938 315256 258944 315268
rect 258996 315256 259002 315308
rect 335298 315256 335304 315308
rect 335356 315296 335362 315308
rect 508350 315296 508356 315308
rect 335356 315268 508356 315296
rect 335356 315256 335362 315268
rect 508350 315256 508356 315268
rect 508408 315256 508414 315308
rect 1600 314928 583316 315024
rect 275498 314644 275504 314696
rect 275556 314684 275562 314696
rect 275682 314684 275688 314696
rect 275556 314656 275688 314684
rect 275556 314644 275562 314656
rect 275682 314644 275688 314656
rect 275740 314644 275746 314696
rect 1600 314384 583316 314480
rect 318922 314072 318928 314084
rect 318883 314044 318928 314072
rect 318922 314032 318928 314044
rect 318980 314032 318986 314084
rect 242654 313964 242660 314016
rect 242712 314004 242718 314016
rect 242838 314004 242844 314016
rect 242712 313976 242844 314004
rect 242712 313964 242718 313976
rect 242838 313964 242844 313976
rect 242896 313964 242902 314016
rect 305214 313964 305220 314016
rect 305272 314004 305278 314016
rect 360690 314004 360696 314016
rect 305272 313976 360696 314004
rect 305272 313964 305278 313976
rect 360690 313964 360696 313976
rect 360748 313964 360754 314016
rect 1600 313840 583316 313936
rect 1600 313296 583316 313392
rect 1600 312752 583316 312848
rect 149458 312604 149464 312656
rect 149516 312644 149522 312656
rect 260226 312644 260232 312656
rect 149516 312616 260232 312644
rect 149516 312604 149522 312616
rect 260226 312604 260232 312616
rect 260284 312604 260290 312656
rect 313402 312604 313408 312656
rect 313460 312644 313466 312656
rect 402090 312644 402096 312656
rect 313460 312616 402096 312644
rect 313460 312604 313466 312616
rect 402090 312604 402096 312616
rect 402148 312604 402154 312656
rect 14218 312536 14224 312588
rect 14276 312576 14282 312588
rect 233086 312576 233092 312588
rect 14276 312548 233092 312576
rect 14276 312536 14282 312548
rect 233086 312536 233092 312548
rect 233144 312536 233150 312588
rect 350754 312536 350760 312588
rect 350812 312576 350818 312588
rect 579374 312576 579380 312588
rect 350812 312548 579380 312576
rect 350812 312536 350818 312548
rect 579374 312536 579380 312548
rect 579432 312536 579438 312588
rect 1600 312208 583316 312304
rect 268690 311964 268696 311976
rect 268651 311936 268696 311964
rect 268690 311924 268696 311936
rect 268748 311924 268754 311976
rect 318738 311924 318744 311976
rect 318796 311924 318802 311976
rect 331158 311964 331164 311976
rect 331119 311936 331164 311964
rect 331158 311924 331164 311936
rect 331216 311924 331222 311976
rect 372006 311964 372012 311976
rect 371932 311936 372012 311964
rect 318756 311840 318784 311924
rect 371932 311840 371960 311936
rect 372006 311924 372012 311936
rect 372064 311924 372070 311976
rect 235481 311831 235539 311837
rect 235481 311797 235493 311831
rect 235527 311828 235539 311831
rect 235570 311828 235576 311840
rect 235527 311800 235576 311828
rect 235527 311797 235539 311800
rect 235481 311791 235539 311797
rect 235570 311788 235576 311800
rect 235628 311788 235634 311840
rect 249462 311788 249468 311840
rect 249520 311828 249526 311840
rect 249646 311828 249652 311840
rect 249520 311800 249652 311828
rect 249520 311788 249526 311800
rect 249646 311788 249652 311800
rect 249704 311788 249710 311840
rect 309170 311828 309176 311840
rect 309131 311800 309176 311828
rect 309170 311788 309176 311800
rect 309228 311788 309234 311840
rect 318738 311788 318744 311840
rect 318796 311788 318802 311840
rect 371914 311788 371920 311840
rect 371972 311788 371978 311840
rect 1600 311664 583316 311760
rect 268690 311624 268696 311636
rect 268651 311596 268696 311624
rect 268690 311584 268696 311596
rect 268748 311584 268754 311636
rect 306594 311244 306600 311296
rect 306652 311284 306658 311296
rect 367590 311284 367596 311296
rect 306652 311256 367596 311284
rect 306652 311244 306658 311256
rect 367590 311244 367596 311256
rect 367648 311244 367654 311296
rect 1600 311120 583316 311216
rect 1600 310576 583316 310672
rect 3638 310428 3644 310480
rect 3696 310468 3702 310480
rect 226094 310468 226100 310480
rect 3696 310440 226100 310468
rect 3696 310428 3702 310440
rect 226094 310428 226100 310440
rect 226152 310428 226158 310480
rect 1600 310032 583316 310128
rect 319106 309856 319112 309868
rect 319067 309828 319112 309856
rect 319106 309816 319112 309828
rect 319164 309816 319170 309868
rect 321590 309816 321596 309868
rect 321648 309856 321654 309868
rect 440730 309856 440736 309868
rect 321648 309828 440736 309856
rect 321648 309816 321654 309828
rect 440730 309816 440736 309828
rect 440788 309816 440794 309868
rect 190861 309791 190919 309797
rect 190861 309757 190873 309791
rect 190907 309788 190919 309791
rect 268506 309788 268512 309800
rect 190907 309760 268512 309788
rect 190907 309757 190919 309760
rect 190861 309751 190919 309757
rect 268506 309748 268512 309760
rect 268564 309748 268570 309800
rect 345142 309748 345148 309800
rect 345200 309788 345206 309800
rect 555270 309788 555276 309800
rect 345200 309760 555276 309788
rect 345200 309748 345206 309760
rect 555270 309748 555276 309760
rect 555328 309748 555334 309800
rect 1600 309488 583316 309584
rect 285434 309272 285440 309324
rect 285492 309272 285498 309324
rect 285452 309188 285480 309272
rect 331161 309247 331219 309253
rect 331161 309213 331173 309247
rect 331207 309244 331219 309247
rect 331250 309244 331256 309256
rect 331207 309216 331256 309244
rect 331207 309213 331219 309216
rect 331161 309207 331219 309213
rect 331250 309204 331256 309216
rect 331308 309204 331314 309256
rect 242470 309136 242476 309188
rect 242528 309176 242534 309188
rect 242562 309176 242568 309188
rect 242528 309148 242568 309176
rect 242528 309136 242534 309148
rect 242562 309136 242568 309148
rect 242620 309136 242626 309188
rect 285253 309179 285311 309185
rect 285253 309145 285265 309179
rect 285299 309176 285311 309179
rect 285342 309176 285348 309188
rect 285299 309148 285348 309176
rect 285299 309145 285311 309148
rect 285253 309139 285311 309145
rect 285342 309136 285348 309148
rect 285400 309136 285406 309188
rect 285434 309136 285440 309188
rect 285492 309136 285498 309188
rect 285621 309179 285679 309185
rect 285621 309145 285633 309179
rect 285667 309176 285679 309179
rect 285710 309176 285716 309188
rect 285667 309148 285716 309176
rect 285667 309145 285679 309148
rect 285621 309139 285679 309145
rect 285710 309136 285716 309148
rect 285768 309136 285774 309188
rect 309170 309176 309176 309188
rect 309131 309148 309176 309176
rect 309170 309136 309176 309148
rect 309228 309136 309234 309188
rect 340818 309136 340824 309188
rect 340876 309176 340882 309188
rect 341186 309176 341192 309188
rect 340876 309148 341192 309176
rect 340876 309136 340882 309148
rect 341186 309136 341192 309148
rect 341244 309136 341250 309188
rect 225358 309108 225364 309120
rect 225319 309080 225364 309108
rect 225358 309068 225364 309080
rect 225416 309068 225422 309120
rect 259306 309108 259312 309120
rect 259267 309080 259312 309108
rect 259306 309068 259312 309080
rect 259364 309068 259370 309120
rect 357930 309068 357936 309120
rect 357988 309108 357994 309120
rect 371825 309111 371883 309117
rect 357988 309080 358033 309108
rect 357988 309068 357994 309080
rect 371825 309077 371837 309111
rect 371871 309108 371883 309111
rect 371914 309108 371920 309120
rect 371871 309080 371920 309108
rect 371871 309077 371883 309080
rect 371825 309071 371883 309077
rect 371914 309068 371920 309080
rect 371972 309068 371978 309120
rect 373110 309068 373116 309120
rect 373168 309108 373174 309120
rect 373202 309108 373208 309120
rect 373168 309080 373208 309108
rect 373168 309068 373174 309080
rect 373202 309068 373208 309080
rect 373260 309068 373266 309120
rect 552510 309068 552516 309120
rect 552568 309108 552574 309120
rect 552602 309108 552608 309120
rect 552568 309080 552608 309108
rect 552568 309068 552574 309080
rect 552602 309068 552608 309080
rect 552660 309068 552666 309120
rect 1600 308944 583316 309040
rect 1600 308400 583316 308496
rect 1600 307856 583316 307952
rect 135658 307816 135664 307828
rect 135619 307788 135664 307816
rect 135658 307776 135664 307788
rect 135716 307776 135722 307828
rect 152218 307816 152224 307828
rect 152179 307788 152224 307816
rect 152218 307776 152224 307788
rect 152276 307776 152282 307828
rect 170158 307816 170164 307828
rect 170119 307788 170164 307816
rect 170158 307776 170164 307788
rect 170216 307776 170222 307828
rect 190858 307816 190864 307828
rect 190819 307788 190864 307816
rect 190858 307776 190864 307788
rect 190916 307776 190922 307828
rect 214318 307816 214324 307828
rect 214279 307788 214324 307816
rect 214318 307776 214324 307788
rect 214376 307776 214382 307828
rect 319934 307776 319940 307828
rect 319992 307816 319998 307828
rect 320118 307816 320124 307828
rect 319992 307788 320124 307816
rect 319992 307776 319998 307788
rect 320118 307776 320124 307788
rect 320176 307776 320182 307828
rect 385530 307776 385536 307828
rect 385588 307816 385594 307828
rect 392430 307816 392436 307828
rect 385588 307788 385633 307816
rect 392391 307788 392436 307816
rect 385588 307776 385594 307788
rect 392430 307776 392436 307788
rect 392488 307776 392494 307828
rect 229866 307708 229872 307760
rect 229924 307748 229930 307760
rect 229958 307748 229964 307760
rect 229924 307720 229964 307748
rect 229924 307708 229930 307720
rect 229958 307708 229964 307720
rect 230016 307708 230022 307760
rect 372926 307708 372932 307760
rect 372984 307748 372990 307760
rect 373202 307748 373208 307760
rect 372984 307720 373208 307748
rect 372984 307708 372990 307720
rect 373202 307708 373208 307720
rect 373260 307708 373266 307760
rect 1600 307312 583316 307408
rect 247732 307176 247944 307204
rect 160498 307096 160504 307148
rect 160556 307136 160562 307148
rect 247732 307136 247760 307176
rect 160556 307108 247760 307136
rect 247916 307136 247944 307176
rect 263078 307136 263084 307148
rect 247916 307108 263084 307136
rect 160556 307096 160562 307108
rect 263078 307096 263084 307108
rect 263136 307096 263142 307148
rect 321682 307096 321688 307148
rect 321740 307136 321746 307148
rect 443582 307136 443588 307148
rect 321740 307108 443588 307136
rect 321740 307096 321746 307108
rect 443582 307096 443588 307108
rect 443640 307096 443646 307148
rect 103918 307028 103924 307080
rect 103976 307068 103982 307080
rect 250934 307068 250940 307080
rect 103976 307040 250940 307068
rect 103976 307028 103982 307040
rect 250934 307028 250940 307040
rect 250992 307028 250998 307080
rect 339530 307028 339536 307080
rect 339588 307068 339594 307080
rect 529050 307068 529056 307080
rect 339588 307040 529056 307068
rect 339588 307028 339594 307040
rect 529050 307028 529056 307040
rect 529108 307028 529114 307080
rect 1600 306768 583316 306864
rect 342198 306348 342204 306400
rect 342256 306388 342262 306400
rect 342382 306388 342388 306400
rect 342256 306360 342388 306388
rect 342256 306348 342262 306360
rect 342382 306348 342388 306360
rect 342440 306348 342446 306400
rect 1600 306224 583316 306320
rect 1600 305680 583316 305776
rect 1600 305136 583316 305232
rect 272554 304920 272560 304972
rect 272612 304960 272618 304972
rect 272830 304960 272836 304972
rect 272612 304932 272836 304960
rect 272612 304920 272618 304932
rect 272830 304920 272836 304932
rect 272888 304920 272894 304972
rect 273014 304920 273020 304972
rect 273072 304960 273078 304972
rect 273198 304960 273204 304972
rect 273072 304932 273204 304960
rect 273072 304920 273078 304932
rect 273198 304920 273204 304932
rect 273256 304920 273262 304972
rect 276602 304920 276608 304972
rect 276660 304920 276666 304972
rect 276694 304920 276700 304972
rect 276752 304960 276758 304972
rect 276970 304960 276976 304972
rect 276752 304932 276976 304960
rect 276752 304920 276758 304932
rect 276970 304920 276976 304932
rect 277028 304920 277034 304972
rect 276620 304892 276648 304920
rect 277246 304892 277252 304904
rect 276620 304864 277252 304892
rect 277246 304852 277252 304864
rect 277304 304852 277310 304904
rect 1600 304592 583316 304688
rect 322970 304308 322976 304360
rect 323028 304348 323034 304360
rect 451770 304348 451776 304360
rect 323028 304320 451776 304348
rect 323028 304308 323034 304320
rect 451770 304308 451776 304320
rect 451828 304308 451834 304360
rect 128758 304240 128764 304292
rect 128816 304280 128822 304292
rect 255994 304280 256000 304292
rect 128816 304252 256000 304280
rect 128816 304240 128822 304252
rect 255994 304240 256000 304252
rect 256052 304240 256058 304292
rect 343762 304240 343768 304292
rect 343820 304280 343826 304292
rect 546990 304280 546996 304292
rect 343820 304252 546996 304280
rect 343820 304240 343826 304252
rect 546990 304240 546996 304252
rect 547048 304240 547054 304292
rect 1600 304048 583316 304144
rect 1600 303504 583316 303600
rect 1600 302960 583316 303056
rect 1600 302416 583316 302512
rect 235754 302308 235760 302320
rect 235680 302280 235760 302308
rect 235680 302184 235708 302280
rect 235754 302268 235760 302280
rect 235812 302268 235818 302320
rect 239250 302268 239256 302320
rect 239308 302268 239314 302320
rect 239342 302268 239348 302320
rect 239400 302268 239406 302320
rect 285342 302308 285348 302320
rect 285268 302280 285348 302308
rect 239268 302184 239296 302268
rect 239360 302184 239388 302268
rect 285268 302184 285296 302280
rect 285342 302268 285348 302280
rect 285400 302268 285406 302320
rect 285710 302268 285716 302320
rect 285768 302268 285774 302320
rect 235662 302132 235668 302184
rect 235720 302132 235726 302184
rect 239250 302132 239256 302184
rect 239308 302132 239314 302184
rect 239342 302132 239348 302184
rect 239400 302132 239406 302184
rect 285250 302132 285256 302184
rect 285308 302132 285314 302184
rect 285728 302104 285756 302268
rect 331158 302200 331164 302252
rect 331216 302200 331222 302252
rect 331176 302172 331204 302200
rect 331250 302172 331256 302184
rect 331176 302144 331256 302172
rect 331250 302132 331256 302144
rect 331308 302132 331314 302184
rect 340818 302132 340824 302184
rect 340876 302172 340882 302184
rect 341186 302172 341192 302184
rect 340876 302144 341192 302172
rect 340876 302132 340882 302144
rect 341186 302132 341192 302144
rect 341244 302132 341250 302184
rect 371822 302172 371828 302184
rect 371783 302144 371828 302172
rect 371822 302132 371828 302144
rect 371880 302132 371886 302184
rect 285802 302104 285808 302116
rect 285728 302076 285808 302104
rect 285802 302064 285808 302076
rect 285860 302064 285866 302116
rect 1600 301872 583316 301968
rect 324350 301520 324356 301572
rect 324408 301560 324414 301572
rect 458670 301560 458676 301572
rect 324408 301532 458676 301560
rect 324408 301520 324414 301532
rect 458670 301520 458676 301532
rect 458728 301520 458734 301572
rect 139798 301452 139804 301504
rect 139856 301492 139862 301504
rect 258846 301492 258852 301504
rect 139856 301464 258852 301492
rect 139856 301452 139862 301464
rect 258846 301452 258852 301464
rect 258904 301452 258910 301504
rect 346430 301452 346436 301504
rect 346488 301492 346494 301504
rect 563550 301492 563556 301504
rect 346488 301464 563556 301492
rect 346488 301452 346494 301464
rect 563550 301452 563556 301464
rect 563608 301452 563614 301504
rect 1600 301328 583316 301424
rect 1600 300784 583316 300880
rect 1600 300240 583316 300336
rect 325730 300160 325736 300212
rect 325788 300200 325794 300212
rect 461430 300200 461436 300212
rect 325788 300172 461436 300200
rect 325788 300160 325794 300172
rect 461430 300160 461436 300172
rect 461488 300160 461494 300212
rect 142466 300092 142472 300144
rect 142524 300132 142530 300144
rect 258754 300132 258760 300144
rect 142524 300104 258760 300132
rect 142524 300092 142530 300104
rect 258754 300092 258760 300104
rect 258812 300092 258818 300144
rect 347810 300092 347816 300144
rect 347868 300132 347874 300144
rect 567690 300132 567696 300144
rect 347868 300104 567696 300132
rect 347868 300092 347874 300104
rect 567690 300092 567696 300104
rect 567748 300092 567754 300144
rect 1600 299696 583316 299792
rect 225358 299520 225364 299532
rect 225319 299492 225364 299520
rect 225358 299480 225364 299492
rect 225416 299480 225422 299532
rect 242470 299480 242476 299532
rect 242528 299520 242534 299532
rect 242562 299520 242568 299532
rect 242528 299492 242568 299520
rect 242528 299480 242534 299492
rect 242562 299480 242568 299492
rect 242620 299480 242626 299532
rect 259309 299523 259367 299529
rect 259309 299489 259321 299523
rect 259355 299520 259367 299523
rect 259398 299520 259404 299532
rect 259355 299492 259404 299520
rect 259355 299489 259367 299492
rect 259309 299483 259367 299489
rect 259398 299480 259404 299492
rect 259456 299480 259462 299532
rect 271358 299480 271364 299532
rect 271416 299480 271422 299532
rect 275501 299523 275559 299529
rect 275501 299489 275513 299523
rect 275547 299520 275559 299523
rect 275682 299520 275688 299532
rect 275547 299492 275688 299520
rect 275547 299489 275559 299492
rect 275501 299483 275559 299489
rect 275682 299480 275688 299492
rect 275740 299480 275746 299532
rect 357930 299480 357936 299532
rect 357988 299520 357994 299532
rect 357988 299492 358033 299520
rect 357988 299480 357994 299492
rect 235662 299452 235668 299464
rect 235623 299424 235668 299452
rect 235662 299412 235668 299424
rect 235720 299412 235726 299464
rect 239250 299412 239256 299464
rect 239308 299452 239314 299464
rect 239434 299452 239440 299464
rect 239308 299424 239440 299452
rect 239308 299412 239314 299424
rect 239434 299412 239440 299424
rect 239492 299412 239498 299464
rect 271376 299384 271404 299480
rect 309170 299452 309176 299464
rect 309131 299424 309176 299452
rect 309170 299412 309176 299424
rect 309228 299412 309234 299464
rect 553798 299412 553804 299464
rect 553856 299452 553862 299464
rect 553890 299452 553896 299464
rect 553856 299424 553896 299452
rect 553856 299412 553862 299424
rect 553890 299412 553896 299424
rect 553948 299412 553954 299464
rect 271450 299384 271456 299396
rect 271376 299356 271456 299384
rect 271450 299344 271456 299356
rect 271508 299344 271514 299396
rect 1600 299152 583316 299248
rect 272554 298732 272560 298784
rect 272612 298772 272618 298784
rect 272922 298772 272928 298784
rect 272612 298744 272928 298772
rect 272612 298732 272618 298744
rect 272922 298732 272928 298744
rect 272980 298732 272986 298784
rect 1600 298608 583316 298704
rect 1600 298064 583316 298160
rect 229866 297984 229872 298036
rect 229924 298024 229930 298036
rect 230234 298024 230240 298036
rect 229924 297996 230240 298024
rect 229924 297984 229930 297996
rect 230234 297984 230240 297996
rect 230292 297984 230298 298036
rect 319934 298024 319940 298036
rect 319895 297996 319940 298024
rect 319934 297984 319940 297996
rect 319992 297984 319998 298036
rect 1600 297520 583316 297616
rect 183958 297440 183964 297492
rect 184016 297480 184022 297492
rect 267126 297480 267132 297492
rect 184016 297452 267132 297480
rect 184016 297440 184022 297452
rect 267126 297440 267132 297452
rect 267184 297440 267190 297492
rect 307882 297440 307888 297492
rect 307940 297480 307946 297492
rect 374490 297480 374496 297492
rect 307940 297452 374496 297480
rect 307940 297440 307946 297452
rect 374490 297440 374496 297452
rect 374548 297440 374554 297492
rect 29398 297372 29404 297424
rect 29456 297412 29462 297424
rect 235665 297415 235723 297421
rect 235665 297412 235677 297415
rect 29456 297384 235677 297412
rect 29456 297372 29462 297384
rect 235665 297381 235677 297384
rect 235711 297381 235723 297415
rect 235665 297375 235723 297381
rect 340910 297372 340916 297424
rect 340968 297412 340974 297424
rect 534570 297412 534576 297424
rect 340968 297384 534576 297412
rect 340968 297372 340974 297384
rect 534570 297372 534576 297384
rect 534628 297372 534634 297424
rect 1600 296976 583316 297072
rect 275498 296936 275504 296948
rect 275459 296908 275504 296936
rect 275498 296896 275504 296908
rect 275556 296896 275562 296948
rect 278718 296692 278724 296744
rect 278776 296732 278782 296744
rect 278902 296732 278908 296744
rect 278776 296704 278908 296732
rect 278776 296692 278782 296704
rect 278902 296692 278908 296704
rect 278960 296692 278966 296744
rect 342198 296692 342204 296744
rect 342256 296732 342262 296744
rect 342382 296732 342388 296744
rect 342256 296704 342388 296732
rect 342256 296692 342262 296704
rect 342382 296692 342388 296704
rect 342440 296692 342446 296744
rect 1600 296432 583316 296528
rect 1600 295888 583316 295984
rect 272646 295576 272652 295588
rect 272607 295548 272652 295576
rect 272646 295536 272652 295548
rect 272704 295536 272710 295588
rect 272738 295508 272744 295520
rect 272699 295480 272744 295508
rect 272738 295468 272744 295480
rect 272796 295468 272802 295520
rect 1600 295344 583316 295440
rect 249370 295264 249376 295316
rect 249428 295304 249434 295316
rect 249646 295304 249652 295316
rect 249428 295276 249652 295304
rect 249428 295264 249434 295276
rect 249646 295264 249652 295276
rect 249704 295264 249710 295316
rect 272738 295304 272744 295316
rect 272699 295276 272744 295304
rect 272738 295264 272744 295276
rect 272796 295264 272802 295316
rect 276694 295304 276700 295316
rect 276655 295276 276700 295304
rect 276694 295264 276700 295276
rect 276752 295264 276758 295316
rect 278442 295264 278448 295316
rect 278500 295304 278506 295316
rect 278718 295304 278724 295316
rect 278500 295276 278724 295304
rect 278500 295264 278506 295276
rect 278718 295264 278724 295276
rect 278776 295264 278782 295316
rect 272646 295236 272652 295248
rect 272607 295208 272652 295236
rect 272646 295196 272652 295208
rect 272704 295196 272710 295248
rect 276602 295236 276608 295248
rect 276563 295208 276608 295236
rect 276602 295196 276608 295208
rect 276660 295196 276666 295248
rect 340818 294924 340824 294976
rect 340876 294964 340882 294976
rect 341186 294964 341192 294976
rect 340876 294936 341192 294964
rect 340876 294924 340882 294936
rect 341186 294924 341192 294936
rect 341244 294924 341250 294976
rect 1600 294800 583316 294896
rect 81838 294584 81844 294636
rect 81896 294624 81902 294636
rect 246426 294624 246432 294636
rect 81896 294596 246432 294624
rect 81896 294584 81902 294596
rect 246426 294584 246432 294596
rect 246484 294584 246490 294636
rect 303466 294584 303472 294636
rect 303524 294624 303530 294636
rect 339990 294624 339996 294636
rect 303524 294596 339996 294624
rect 303524 294584 303530 294596
rect 339990 294584 339996 294596
rect 340048 294584 340054 294636
rect 341002 294584 341008 294636
rect 341060 294624 341066 294636
rect 537330 294624 537336 294636
rect 341060 294596 537336 294624
rect 341060 294584 341066 294596
rect 537330 294584 537336 294596
rect 537388 294584 537394 294636
rect 1600 294256 583316 294352
rect 3546 293836 3552 293888
rect 3604 293876 3610 293888
rect 6674 293876 6680 293888
rect 3604 293848 6680 293876
rect 3604 293836 3610 293848
rect 6674 293836 6680 293848
rect 6732 293836 6738 293888
rect 1600 293712 583316 293808
rect 1600 293168 583316 293264
rect 1600 292624 583316 292720
rect 331158 292544 331164 292596
rect 331216 292584 331222 292596
rect 331216 292556 331296 292584
rect 331216 292544 331222 292556
rect 331268 292528 331296 292556
rect 268690 292476 268696 292528
rect 268748 292476 268754 292528
rect 331250 292476 331256 292528
rect 331308 292476 331314 292528
rect 268708 292392 268736 292476
rect 319937 292451 319995 292457
rect 319937 292417 319949 292451
rect 319983 292448 319995 292451
rect 320118 292448 320124 292460
rect 319983 292420 320124 292448
rect 319983 292417 319995 292420
rect 319937 292411 319995 292417
rect 320118 292408 320124 292420
rect 320176 292408 320182 292460
rect 268690 292340 268696 292392
rect 268748 292340 268754 292392
rect 1600 292080 583316 292176
rect 84598 291796 84604 291848
rect 84656 291836 84662 291848
rect 245414 291836 245420 291848
rect 84656 291808 245420 291836
rect 84656 291796 84662 291808
rect 245414 291796 245420 291808
rect 245472 291796 245478 291848
rect 342290 291796 342296 291848
rect 342348 291836 342354 291848
rect 545610 291836 545616 291848
rect 342348 291808 545616 291836
rect 342348 291796 342354 291808
rect 545610 291796 545616 291808
rect 545668 291796 545674 291848
rect 1600 291536 583316 291632
rect 1600 290992 583316 291088
rect 1600 290448 583316 290544
rect 1600 289904 583316 290000
rect 235478 289824 235484 289876
rect 235536 289864 235542 289876
rect 235570 289864 235576 289876
rect 235536 289836 235576 289864
rect 235536 289824 235542 289836
rect 235570 289824 235576 289836
rect 235628 289824 235634 289876
rect 309170 289864 309176 289876
rect 309131 289836 309176 289864
rect 309170 289824 309176 289836
rect 309228 289824 309234 289876
rect 259398 289796 259404 289808
rect 259359 289768 259404 289796
rect 259398 289756 259404 289768
rect 259456 289756 259462 289808
rect 340913 289799 340971 289805
rect 340913 289765 340925 289799
rect 340959 289796 340971 289799
rect 341186 289796 341192 289808
rect 340959 289768 341192 289796
rect 340959 289765 340971 289768
rect 340913 289759 340971 289765
rect 341186 289756 341192 289768
rect 341244 289756 341250 289808
rect 354434 289756 354440 289808
rect 354492 289796 354498 289808
rect 580662 289796 580668 289808
rect 354492 289768 580668 289796
rect 354492 289756 354498 289768
rect 580662 289756 580668 289768
rect 580720 289756 580726 289808
rect 357930 289688 357936 289740
rect 357988 289728 357994 289740
rect 358025 289731 358083 289737
rect 358025 289728 358037 289731
rect 357988 289700 358037 289728
rect 357988 289688 357994 289700
rect 358025 289697 358037 289700
rect 358071 289697 358083 289731
rect 371914 289728 371920 289740
rect 371875 289700 371920 289728
rect 358025 289691 358083 289697
rect 371914 289688 371920 289700
rect 371972 289688 371978 289740
rect 553890 289728 553896 289740
rect 553851 289700 553896 289728
rect 553890 289688 553896 289700
rect 553948 289688 553954 289740
rect 1600 289360 583316 289456
rect 88738 289076 88744 289128
rect 88796 289116 88802 289128
rect 248266 289116 248272 289128
rect 88796 289088 248272 289116
rect 88796 289076 88802 289088
rect 248266 289076 248272 289088
rect 248324 289076 248330 289128
rect 1600 288816 583316 288912
rect 135474 288396 135480 288448
rect 135532 288436 135538 288448
rect 135658 288436 135664 288448
rect 135532 288408 135664 288436
rect 135532 288396 135538 288408
rect 135658 288396 135664 288408
rect 135716 288396 135722 288448
rect 152034 288396 152040 288448
rect 152092 288436 152098 288448
rect 152218 288436 152224 288448
rect 152092 288408 152224 288436
rect 152092 288396 152098 288408
rect 152218 288396 152224 288408
rect 152276 288396 152282 288448
rect 170158 288396 170164 288448
rect 170216 288436 170222 288448
rect 170342 288436 170348 288448
rect 170216 288408 170348 288436
rect 170216 288396 170222 288408
rect 170342 288396 170348 288408
rect 170400 288396 170406 288448
rect 190674 288396 190680 288448
rect 190732 288436 190738 288448
rect 190858 288436 190864 288448
rect 190732 288408 190864 288436
rect 190732 288396 190738 288408
rect 190858 288396 190864 288408
rect 190916 288396 190922 288448
rect 214318 288396 214324 288448
rect 214376 288436 214382 288448
rect 214502 288436 214508 288448
rect 214376 288408 214508 288436
rect 214376 288396 214382 288408
rect 214502 288396 214508 288408
rect 214560 288396 214566 288448
rect 385530 288396 385536 288448
rect 385588 288436 385594 288448
rect 385714 288436 385720 288448
rect 385588 288408 385720 288436
rect 385588 288396 385594 288408
rect 385714 288396 385720 288408
rect 385772 288396 385778 288448
rect 392430 288396 392436 288448
rect 392488 288436 392494 288448
rect 392614 288436 392620 288448
rect 392488 288408 392620 288436
rect 392488 288396 392494 288408
rect 392614 288396 392620 288408
rect 392672 288396 392678 288448
rect 528866 288396 528872 288448
rect 528924 288436 528930 288448
rect 529050 288436 529056 288448
rect 528924 288408 529056 288436
rect 528924 288396 528930 288408
rect 529050 288396 529056 288408
rect 529108 288396 529114 288448
rect 1600 288272 583316 288368
rect 372834 288192 372840 288244
rect 372892 288232 372898 288244
rect 373110 288232 373116 288244
rect 372892 288204 373116 288232
rect 372892 288192 372898 288204
rect 373110 288192 373116 288204
rect 373168 288192 373174 288244
rect 1600 287728 583316 287824
rect 1600 287184 583316 287280
rect 229958 287036 229964 287088
rect 230016 287076 230022 287088
rect 230142 287076 230148 287088
rect 230016 287048 230148 287076
rect 230016 287036 230022 287048
rect 230142 287036 230148 287048
rect 230200 287036 230206 287088
rect 1600 286640 583316 286736
rect 314874 286356 314880 286408
rect 314932 286396 314938 286408
rect 408990 286396 408996 286408
rect 314932 286368 408996 286396
rect 314932 286356 314938 286368
rect 408990 286356 408996 286368
rect 409048 286356 409054 286408
rect 91501 286331 91559 286337
rect 91501 286297 91513 286331
rect 91547 286328 91559 286331
rect 249186 286328 249192 286340
rect 91547 286300 249192 286328
rect 91547 286297 91559 286300
rect 91501 286291 91559 286297
rect 249186 286288 249192 286300
rect 249244 286288 249250 286340
rect 347902 286288 347908 286340
rect 347960 286328 347966 286340
rect 571830 286328 571836 286340
rect 347960 286300 571836 286328
rect 347960 286288 347966 286300
rect 571830 286288 571836 286300
rect 571888 286288 571894 286340
rect 1600 286096 583316 286192
rect 276602 285716 276608 285728
rect 276563 285688 276608 285716
rect 276602 285676 276608 285688
rect 276660 285676 276666 285728
rect 276697 285719 276755 285725
rect 276697 285685 276709 285719
rect 276743 285716 276755 285719
rect 276970 285716 276976 285728
rect 276743 285688 276976 285716
rect 276743 285685 276755 285688
rect 276697 285679 276755 285685
rect 276970 285676 276976 285688
rect 277028 285676 277034 285728
rect 1600 285552 583316 285648
rect 235478 285308 235484 285320
rect 235439 285280 235484 285308
rect 235478 285268 235484 285280
rect 235536 285268 235542 285320
rect 276697 285175 276755 285181
rect 276697 285141 276709 285175
rect 276743 285172 276755 285175
rect 276970 285172 276976 285184
rect 276743 285144 276976 285172
rect 276743 285141 276755 285144
rect 276697 285135 276755 285141
rect 276970 285132 276976 285144
rect 277028 285132 277034 285184
rect 1600 285008 583316 285104
rect 268690 284968 268696 284980
rect 268651 284940 268696 284968
rect 268690 284928 268696 284940
rect 268748 284928 268754 284980
rect 1600 284464 583316 284560
rect 272830 284248 272836 284300
rect 272888 284288 272894 284300
rect 272922 284288 272928 284300
rect 272888 284260 272928 284288
rect 272888 284248 272894 284260
rect 272922 284248 272928 284260
rect 272980 284248 272986 284300
rect 1600 283920 583316 284016
rect 316162 283636 316168 283688
rect 316220 283676 316226 283688
rect 417362 283676 417368 283688
rect 316220 283648 417368 283676
rect 316220 283636 316226 283648
rect 417362 283636 417368 283648
rect 417420 283636 417426 283688
rect 95638 283568 95644 283620
rect 95696 283608 95702 283620
rect 249370 283608 249376 283620
rect 95696 283580 249376 283608
rect 95696 283568 95702 283580
rect 249370 283568 249376 283580
rect 249428 283568 249434 283620
rect 349282 283568 349288 283620
rect 349340 283608 349346 283620
rect 577994 283608 578000 283620
rect 349340 283580 578000 283608
rect 349340 283568 349346 283580
rect 577994 283568 578000 283580
rect 578052 283568 578058 283620
rect 1600 283376 583316 283472
rect 271450 283064 271456 283076
rect 271411 283036 271456 283064
rect 271450 283024 271456 283036
rect 271508 283024 271514 283076
rect 341094 282996 341100 283008
rect 341055 282968 341100 282996
rect 341094 282956 341100 282968
rect 341152 282956 341158 283008
rect 1600 282832 583316 282928
rect 235481 282795 235539 282801
rect 235481 282761 235493 282795
rect 235527 282792 235539 282795
rect 235570 282792 235576 282804
rect 235527 282764 235576 282792
rect 235527 282761 235539 282764
rect 235481 282755 235539 282761
rect 235570 282752 235576 282764
rect 235628 282752 235634 282804
rect 268693 282795 268751 282801
rect 268693 282761 268705 282795
rect 268739 282792 268751 282795
rect 268782 282792 268788 282804
rect 268739 282764 268788 282792
rect 268739 282761 268751 282764
rect 268693 282755 268751 282761
rect 268782 282752 268788 282764
rect 268840 282752 268846 282804
rect 271450 282792 271456 282804
rect 271411 282764 271456 282792
rect 271450 282752 271456 282764
rect 271508 282752 271514 282804
rect 341094 282792 341100 282804
rect 341055 282764 341100 282792
rect 341094 282752 341100 282764
rect 341152 282752 341158 282804
rect 371914 282792 371920 282804
rect 371875 282764 371920 282792
rect 371914 282752 371920 282764
rect 371972 282752 371978 282804
rect 1600 282288 583316 282384
rect 1600 281744 583316 281840
rect 1600 281200 583316 281296
rect 1600 280656 583316 280752
rect 276786 280480 276792 280492
rect 276747 280452 276792 280480
rect 276786 280440 276792 280452
rect 276844 280440 276850 280492
rect 357930 280304 357936 280356
rect 357988 280344 357994 280356
rect 358025 280347 358083 280353
rect 358025 280344 358037 280347
rect 357988 280316 358037 280344
rect 357988 280304 357994 280316
rect 358025 280313 358037 280316
rect 358071 280313 358083 280347
rect 358025 280307 358083 280313
rect 91498 280276 91504 280288
rect 91459 280248 91504 280276
rect 91498 280236 91504 280248
rect 91556 280236 91562 280288
rect 259398 280276 259404 280288
rect 259359 280248 259404 280276
rect 259398 280236 259404 280248
rect 259456 280236 259462 280288
rect 340910 280276 340916 280288
rect 340871 280248 340916 280276
rect 340910 280236 340916 280248
rect 340968 280236 340974 280288
rect 372929 280279 372987 280285
rect 372929 280245 372941 280279
rect 372975 280276 372987 280279
rect 373110 280276 373116 280288
rect 372975 280248 373116 280276
rect 372975 280245 372987 280248
rect 372929 280239 372987 280245
rect 373110 280236 373116 280248
rect 373168 280236 373174 280288
rect 553890 280276 553896 280288
rect 553851 280248 553896 280276
rect 553890 280236 553896 280248
rect 553948 280236 553954 280288
rect 1600 280112 583316 280208
rect 276786 280072 276792 280084
rect 276747 280044 276792 280072
rect 276786 280032 276792 280044
rect 276844 280032 276850 280084
rect 309170 280072 309176 280084
rect 309131 280044 309176 280072
rect 309170 280032 309176 280044
rect 309228 280032 309234 280084
rect 331250 280072 331256 280084
rect 331211 280044 331256 280072
rect 331250 280032 331256 280044
rect 331308 280032 331314 280084
rect 276694 280004 276700 280016
rect 276655 279976 276700 280004
rect 276694 279964 276700 279976
rect 276752 279964 276758 280016
rect 285158 279868 285164 279880
rect 285119 279840 285164 279868
rect 285158 279828 285164 279840
rect 285216 279828 285222 279880
rect 285250 279828 285256 279880
rect 285308 279868 285314 279880
rect 285308 279840 285353 279868
rect 285308 279828 285314 279840
rect 1600 279568 583316 279664
rect 99778 279420 99784 279472
rect 99836 279460 99842 279472
rect 249554 279460 249560 279472
rect 99836 279432 249560 279460
rect 99836 279420 99842 279432
rect 249554 279420 249560 279432
rect 249612 279420 249618 279472
rect 335390 279420 335396 279472
rect 335448 279460 335454 279472
rect 506970 279460 506976 279472
rect 335448 279432 506976 279460
rect 335448 279420 335454 279432
rect 506970 279420 506976 279432
rect 507028 279420 507034 279472
rect 1600 279024 583316 279120
rect 242102 278848 242108 278860
rect 242063 278820 242108 278848
rect 242102 278808 242108 278820
rect 242160 278808 242166 278860
rect 246610 278848 246616 278860
rect 246571 278820 246616 278848
rect 246610 278808 246616 278820
rect 246668 278808 246674 278860
rect 229958 278740 229964 278792
rect 230016 278780 230022 278792
rect 230050 278780 230056 278792
rect 230016 278752 230056 278780
rect 230016 278740 230022 278752
rect 230050 278740 230056 278752
rect 230108 278740 230114 278792
rect 372926 278780 372932 278792
rect 372887 278752 372932 278780
rect 372926 278740 372932 278752
rect 372984 278740 372990 278792
rect 552510 278740 552516 278792
rect 552568 278780 552574 278792
rect 552602 278780 552608 278792
rect 552568 278752 552608 278780
rect 552568 278740 552574 278752
rect 552602 278740 552608 278752
rect 552660 278740 552666 278792
rect 285710 278672 285716 278724
rect 285768 278712 285774 278724
rect 285802 278712 285808 278724
rect 285768 278684 285808 278712
rect 285768 278672 285774 278684
rect 285802 278672 285808 278684
rect 285860 278672 285866 278724
rect 1600 278480 583316 278576
rect 1600 277936 583316 278032
rect 1600 277392 583316 277488
rect 242102 277352 242108 277364
rect 242063 277324 242108 277352
rect 242102 277312 242108 277324
rect 242160 277312 242166 277364
rect 246610 277352 246616 277364
rect 246571 277324 246616 277352
rect 246610 277312 246616 277324
rect 246668 277312 246674 277364
rect 1600 276848 583316 276944
rect 90118 276632 90124 276684
rect 90176 276672 90182 276684
rect 247714 276672 247720 276684
rect 90176 276644 247720 276672
rect 90176 276632 90182 276644
rect 247714 276632 247720 276644
rect 247772 276632 247778 276684
rect 336770 276632 336776 276684
rect 336828 276672 336834 276684
rect 513870 276672 513876 276684
rect 336828 276644 513876 276672
rect 336828 276632 336834 276644
rect 513870 276632 513876 276644
rect 513928 276632 513934 276684
rect 1600 276304 583316 276400
rect 273014 275952 273020 276004
rect 273072 275992 273078 276004
rect 273106 275992 273112 276004
rect 273072 275964 273112 275992
rect 273072 275952 273078 275964
rect 273106 275952 273112 275964
rect 273164 275952 273170 276004
rect 328214 275952 328220 276004
rect 328272 275992 328278 276004
rect 328398 275992 328404 276004
rect 328272 275964 328404 275992
rect 328272 275952 328278 275964
rect 328398 275952 328404 275964
rect 328456 275952 328462 276004
rect 1600 275760 583316 275856
rect 1600 275216 583316 275312
rect 1600 274672 583316 274768
rect 272830 274592 272836 274644
rect 272888 274632 272894 274644
rect 273014 274632 273020 274644
rect 272888 274604 273020 274632
rect 272888 274592 272894 274604
rect 273014 274592 273020 274604
rect 273072 274592 273078 274644
rect 358574 274592 358580 274644
rect 358632 274632 358638 274644
rect 580662 274632 580668 274644
rect 358632 274604 580668 274632
rect 358632 274592 358638 274604
rect 580662 274592 580668 274604
rect 580720 274592 580726 274644
rect 1600 274128 583316 274224
rect 19738 273912 19744 273964
rect 19796 273952 19802 273964
rect 234098 273952 234104 273964
rect 19796 273924 234104 273952
rect 19796 273912 19802 273924
rect 234098 273912 234104 273924
rect 234156 273912 234162 273964
rect 1600 273584 583316 273680
rect 246794 273340 246800 273352
rect 246720 273312 246800 273340
rect 239250 273232 239256 273284
rect 239308 273272 239314 273284
rect 239434 273272 239440 273284
rect 239308 273244 239440 273272
rect 239308 273232 239314 273244
rect 239434 273232 239440 273244
rect 239492 273232 239498 273284
rect 246720 273216 246748 273312
rect 246794 273300 246800 273312
rect 246852 273300 246858 273352
rect 259309 273343 259367 273349
rect 259309 273309 259321 273343
rect 259355 273340 259367 273343
rect 259398 273340 259404 273352
rect 259355 273312 259404 273340
rect 259355 273309 259367 273312
rect 259309 273303 259367 273309
rect 259398 273300 259404 273312
rect 259456 273300 259462 273352
rect 372006 273340 372012 273352
rect 371932 273312 372012 273340
rect 371932 273216 371960 273312
rect 372006 273300 372012 273312
rect 372064 273300 372070 273352
rect 246702 273164 246708 273216
rect 246760 273164 246766 273216
rect 371914 273164 371920 273216
rect 371972 273164 371978 273216
rect 1600 273040 583316 273136
rect 1600 272496 583316 272592
rect 1600 271952 583316 272048
rect 1600 271408 583316 271504
rect 125906 271124 125912 271176
rect 125964 271164 125970 271176
rect 255902 271164 255908 271176
rect 125964 271136 255908 271164
rect 125964 271124 125970 271136
rect 255902 271124 255908 271136
rect 255960 271124 255966 271176
rect 341094 271124 341100 271176
rect 341152 271164 341158 271176
rect 535953 271167 536011 271173
rect 535953 271164 535965 271167
rect 341152 271136 535965 271164
rect 341152 271124 341158 271136
rect 535953 271133 535965 271136
rect 535999 271133 536011 271167
rect 535953 271127 536011 271133
rect 1600 270864 583316 270960
rect 259306 270552 259312 270564
rect 259267 270524 259312 270552
rect 259306 270512 259312 270524
rect 259364 270512 259370 270564
rect 285253 270555 285311 270561
rect 285253 270521 285265 270555
rect 285299 270552 285311 270555
rect 285342 270552 285348 270564
rect 285299 270524 285348 270552
rect 285299 270521 285311 270524
rect 285253 270515 285311 270521
rect 285342 270512 285348 270524
rect 285400 270512 285406 270564
rect 309170 270552 309176 270564
rect 309131 270524 309176 270552
rect 309170 270512 309176 270524
rect 309228 270512 309234 270564
rect 331250 270552 331256 270564
rect 331211 270524 331256 270552
rect 331250 270512 331256 270524
rect 331308 270512 331314 270564
rect 91498 270484 91504 270496
rect 91459 270456 91504 270484
rect 91498 270444 91504 270456
rect 91556 270444 91562 270496
rect 225358 270484 225364 270496
rect 225319 270456 225364 270484
rect 225358 270444 225364 270456
rect 225416 270444 225422 270496
rect 357930 270444 357936 270496
rect 357988 270484 357994 270496
rect 553890 270484 553896 270496
rect 357988 270456 358033 270484
rect 553851 270456 553896 270484
rect 357988 270444 357994 270456
rect 553890 270444 553896 270456
rect 553948 270444 553954 270496
rect 1600 270320 583316 270416
rect 278442 270240 278448 270292
rect 278500 270280 278506 270292
rect 278810 270280 278816 270292
rect 278500 270252 278816 270280
rect 278500 270240 278506 270252
rect 278810 270240 278816 270252
rect 278868 270240 278874 270292
rect 1600 269776 583316 269872
rect 242746 269736 242752 269748
rect 242707 269708 242752 269736
rect 242746 269696 242752 269708
rect 242804 269696 242810 269748
rect 1600 269232 583316 269328
rect 135474 269084 135480 269136
rect 135532 269124 135538 269136
rect 135658 269124 135664 269136
rect 135532 269096 135664 269124
rect 135532 269084 135538 269096
rect 135658 269084 135664 269096
rect 135716 269084 135722 269136
rect 152034 269084 152040 269136
rect 152092 269124 152098 269136
rect 152218 269124 152224 269136
rect 152092 269096 152224 269124
rect 152092 269084 152098 269096
rect 152218 269084 152224 269096
rect 152276 269084 152282 269136
rect 170158 269084 170164 269136
rect 170216 269124 170222 269136
rect 170342 269124 170348 269136
rect 170216 269096 170348 269124
rect 170216 269084 170222 269096
rect 170342 269084 170348 269096
rect 170400 269084 170406 269136
rect 190674 269084 190680 269136
rect 190732 269124 190738 269136
rect 190858 269124 190864 269136
rect 190732 269096 190864 269124
rect 190732 269084 190738 269096
rect 190858 269084 190864 269096
rect 190916 269084 190922 269136
rect 214318 269084 214324 269136
rect 214376 269124 214382 269136
rect 214502 269124 214508 269136
rect 214376 269096 214508 269124
rect 214376 269084 214382 269096
rect 214502 269084 214508 269096
rect 214560 269084 214566 269136
rect 229774 269084 229780 269136
rect 229832 269124 229838 269136
rect 229866 269124 229872 269136
rect 229832 269096 229872 269124
rect 229832 269084 229838 269096
rect 229866 269084 229872 269096
rect 229924 269084 229930 269136
rect 235386 269084 235392 269136
rect 235444 269124 235450 269136
rect 235570 269124 235576 269136
rect 235444 269096 235576 269124
rect 235444 269084 235450 269096
rect 235570 269084 235576 269096
rect 235628 269084 235634 269136
rect 268598 269084 268604 269136
rect 268656 269124 268662 269136
rect 268690 269124 268696 269136
rect 268656 269096 268696 269124
rect 268656 269084 268662 269096
rect 268690 269084 268696 269096
rect 268748 269084 268754 269136
rect 279822 269084 279828 269136
rect 279880 269124 279886 269136
rect 280006 269124 280012 269136
rect 279880 269096 280012 269124
rect 279880 269084 279886 269096
rect 280006 269084 280012 269096
rect 280064 269084 280070 269136
rect 285158 269124 285164 269136
rect 285119 269096 285164 269124
rect 285158 269084 285164 269096
rect 285216 269084 285222 269136
rect 372926 269084 372932 269136
rect 372984 269124 372990 269136
rect 373110 269124 373116 269136
rect 372984 269096 373116 269124
rect 372984 269084 372990 269096
rect 373110 269084 373116 269096
rect 373168 269084 373174 269136
rect 385530 269084 385536 269136
rect 385588 269124 385594 269136
rect 385714 269124 385720 269136
rect 385588 269096 385720 269124
rect 385588 269084 385594 269096
rect 385714 269084 385720 269096
rect 385772 269084 385778 269136
rect 392430 269084 392436 269136
rect 392488 269124 392494 269136
rect 392614 269124 392620 269136
rect 392488 269096 392620 269124
rect 392488 269084 392494 269096
rect 392614 269084 392620 269096
rect 392672 269084 392678 269136
rect 528866 269084 528872 269136
rect 528924 269124 528930 269136
rect 529050 269124 529056 269136
rect 528924 269096 529056 269124
rect 528924 269084 528930 269096
rect 529050 269084 529056 269096
rect 529108 269084 529114 269136
rect 535950 269124 535956 269136
rect 535911 269096 535956 269124
rect 535950 269084 535956 269096
rect 536008 269084 536014 269136
rect 552602 269084 552608 269136
rect 552660 269124 552666 269136
rect 552786 269124 552792 269136
rect 552660 269096 552792 269124
rect 552660 269084 552666 269096
rect 552786 269084 552792 269096
rect 552844 269084 552850 269136
rect 571830 269084 571836 269136
rect 571888 269124 571894 269136
rect 572014 269124 572020 269136
rect 571888 269096 572020 269124
rect 571888 269084 571894 269096
rect 572014 269084 572020 269096
rect 572072 269084 572078 269136
rect 1600 268688 583316 268784
rect 342382 268336 342388 268388
rect 342440 268376 342446 268388
rect 542850 268376 542856 268388
rect 342440 268348 542856 268376
rect 342440 268336 342446 268348
rect 542850 268336 542856 268348
rect 542908 268336 542914 268388
rect 1600 268144 583316 268240
rect 242562 267832 242568 267844
rect 242488 267804 242568 267832
rect 242488 267776 242516 267804
rect 242562 267792 242568 267804
rect 242620 267792 242626 267844
rect 242470 267724 242476 267776
rect 242528 267724 242534 267776
rect 1600 267600 583316 267696
rect 242749 267563 242807 267569
rect 242749 267529 242761 267563
rect 242795 267560 242807 267563
rect 242930 267560 242936 267572
rect 242795 267532 242936 267560
rect 242795 267529 242807 267532
rect 242749 267523 242807 267529
rect 242930 267520 242936 267532
rect 242988 267520 242994 267572
rect 1600 267056 583316 267152
rect 1600 266512 583316 266608
rect 1600 265968 583316 266064
rect 300890 265616 300896 265668
rect 300948 265656 300954 265668
rect 342750 265656 342756 265668
rect 300948 265628 342756 265656
rect 300948 265616 300954 265628
rect 342750 265616 342756 265628
rect 342808 265616 342814 265668
rect 343854 265616 343860 265668
rect 343912 265656 343918 265668
rect 549750 265656 549756 265668
rect 343912 265628 549756 265656
rect 343912 265616 343918 265628
rect 549750 265616 549756 265628
rect 549808 265616 549814 265668
rect 1600 265424 583316 265520
rect 1600 264880 583316 264976
rect 242841 264843 242899 264849
rect 242841 264809 242853 264843
rect 242887 264840 242899 264843
rect 242930 264840 242936 264852
rect 242887 264812 242936 264840
rect 242887 264809 242899 264812
rect 242841 264803 242899 264809
rect 242930 264800 242936 264812
rect 242988 264800 242994 264852
rect 1600 264336 583316 264432
rect 1600 263792 583316 263888
rect 235570 263644 235576 263696
rect 235628 263644 235634 263696
rect 285342 263684 285348 263696
rect 285268 263656 285348 263684
rect 235588 263492 235616 263644
rect 239250 263576 239256 263628
rect 239308 263616 239314 263628
rect 239434 263616 239440 263628
rect 239308 263588 239440 263616
rect 239308 263576 239314 263588
rect 239434 263576 239440 263588
rect 239492 263576 239498 263628
rect 285268 263560 285296 263656
rect 285342 263644 285348 263656
rect 285400 263644 285406 263696
rect 328398 263684 328404 263696
rect 328324 263656 328404 263684
rect 320026 263616 320032 263628
rect 319987 263588 320032 263616
rect 320026 263576 320032 263588
rect 320084 263576 320090 263628
rect 328324 263560 328352 263656
rect 328398 263644 328404 263656
rect 328456 263644 328462 263696
rect 341186 263684 341192 263696
rect 341112 263656 341192 263684
rect 341112 263560 341140 263656
rect 341186 263644 341192 263656
rect 341244 263644 341250 263696
rect 285250 263508 285256 263560
rect 285308 263508 285314 263560
rect 328306 263508 328312 263560
rect 328364 263508 328370 263560
rect 341094 263508 341100 263560
rect 341152 263508 341158 263560
rect 235570 263440 235576 263492
rect 235628 263440 235634 263492
rect 1600 263248 583316 263344
rect 345234 262828 345240 262880
rect 345292 262868 345298 262880
rect 556650 262868 556656 262880
rect 345292 262840 556656 262868
rect 345292 262828 345298 262840
rect 556650 262828 556656 262840
rect 556708 262828 556714 262880
rect 1600 262704 583316 262800
rect 1600 262160 583316 262256
rect 1600 261616 583316 261712
rect 351766 261468 351772 261520
rect 351824 261508 351830 261520
rect 574590 261508 574596 261520
rect 351824 261480 574596 261508
rect 351824 261468 351830 261480
rect 574590 261468 574596 261480
rect 574648 261468 574654 261520
rect 1600 261072 583316 261168
rect 553890 260964 553896 260976
rect 553851 260936 553896 260964
rect 553890 260924 553896 260936
rect 553948 260924 553954 260976
rect 91498 260896 91504 260908
rect 91459 260868 91504 260896
rect 91498 260856 91504 260868
rect 91556 260856 91562 260908
rect 225358 260896 225364 260908
rect 225319 260868 225364 260896
rect 225358 260856 225364 260868
rect 225416 260856 225422 260908
rect 279730 260856 279736 260908
rect 279788 260896 279794 260908
rect 279822 260896 279828 260908
rect 279788 260868 279828 260896
rect 279788 260856 279794 260868
rect 279822 260856 279828 260868
rect 279880 260856 279886 260908
rect 357930 260856 357936 260908
rect 357988 260896 357994 260908
rect 357988 260868 358033 260896
rect 357988 260856 357994 260868
rect 3822 260788 3828 260840
rect 3880 260828 3886 260840
rect 179174 260828 179180 260840
rect 3880 260800 179180 260828
rect 3880 260788 3886 260800
rect 179174 260788 179180 260800
rect 179232 260788 179238 260840
rect 235570 260828 235576 260840
rect 235531 260800 235576 260828
rect 235570 260788 235576 260800
rect 235628 260788 235634 260840
rect 285618 260828 285624 260840
rect 285579 260800 285624 260828
rect 285618 260788 285624 260800
rect 285676 260788 285682 260840
rect 331250 260828 331256 260840
rect 331211 260800 331256 260828
rect 331250 260788 331256 260800
rect 331308 260788 331314 260840
rect 341094 260828 341100 260840
rect 341055 260800 341100 260828
rect 341094 260788 341100 260800
rect 341152 260788 341158 260840
rect 553890 260788 553896 260840
rect 553948 260788 553954 260840
rect 285250 260760 285256 260772
rect 285211 260732 285256 260760
rect 285250 260720 285256 260732
rect 285308 260720 285314 260772
rect 553798 260720 553804 260772
rect 553856 260760 553862 260772
rect 553908 260760 553936 260788
rect 553856 260732 553936 260760
rect 553856 260720 553862 260732
rect 1600 260528 583316 260624
rect 1600 259984 583316 260080
rect 1600 259440 583316 259536
rect 305030 259400 305036 259412
rect 304991 259372 305036 259400
rect 305030 259360 305036 259372
rect 305088 259360 305094 259412
rect 1600 258896 583316 258992
rect 1600 258352 583316 258448
rect 320026 258108 320032 258120
rect 319987 258080 320032 258108
rect 320026 258068 320032 258080
rect 320084 258068 320090 258120
rect 1600 257808 583316 257904
rect 1600 257264 583316 257360
rect 273014 256884 273020 256896
rect 272975 256856 273020 256884
rect 273014 256844 273020 256856
rect 273072 256844 273078 256896
rect 1600 256720 583316 256816
rect 328306 256680 328312 256692
rect 328267 256652 328312 256680
rect 328306 256640 328312 256652
rect 328364 256640 328370 256692
rect 1600 256176 583316 256272
rect 279730 256028 279736 256080
rect 279788 256028 279794 256080
rect 279748 256000 279776 256028
rect 279822 256000 279828 256012
rect 279748 255972 279828 256000
rect 279822 255960 279828 255972
rect 279880 255960 279886 256012
rect 1600 255632 583316 255728
rect 242838 255320 242844 255332
rect 242799 255292 242844 255320
rect 242838 255280 242844 255292
rect 242896 255280 242902 255332
rect 273014 255320 273020 255332
rect 272975 255292 273020 255320
rect 273014 255280 273020 255292
rect 273072 255280 273078 255332
rect 242562 255252 242568 255264
rect 242523 255224 242568 255252
rect 242562 255212 242568 255224
rect 242620 255212 242626 255264
rect 275593 255255 275651 255261
rect 275593 255221 275605 255255
rect 275639 255252 275651 255255
rect 275682 255252 275688 255264
rect 275639 255224 275688 255252
rect 275639 255221 275651 255224
rect 275593 255215 275651 255221
rect 275682 255212 275688 255224
rect 275740 255212 275746 255264
rect 1600 255088 583316 255184
rect 1600 254544 583316 254640
rect 246521 254167 246579 254173
rect 246521 254133 246533 254167
rect 246567 254164 246579 254167
rect 246610 254164 246616 254176
rect 246567 254136 246616 254164
rect 246567 254133 246579 254136
rect 246521 254127 246579 254133
rect 246610 254124 246616 254136
rect 246668 254124 246674 254176
rect 1600 254000 583316 254096
rect 308986 253920 308992 253972
rect 309044 253960 309050 253972
rect 309044 253932 309124 253960
rect 309044 253920 309050 253932
rect 309096 253904 309124 253932
rect 371914 253920 371920 253972
rect 371972 253960 371978 253972
rect 372098 253960 372104 253972
rect 371972 253932 372104 253960
rect 371972 253920 371978 253932
rect 372098 253920 372104 253932
rect 372156 253920 372162 253972
rect 273014 253892 273020 253904
rect 272975 253864 273020 253892
rect 273014 253852 273020 253864
rect 273072 253852 273078 253904
rect 309078 253852 309084 253904
rect 309136 253852 309142 253904
rect 328306 253892 328312 253904
rect 328267 253864 328312 253892
rect 328306 253852 328312 253864
rect 328364 253852 328370 253904
rect 235570 253824 235576 253836
rect 235531 253796 235576 253824
rect 235570 253784 235576 253796
rect 235628 253784 235634 253836
rect 1600 253456 583316 253552
rect 302362 253172 302368 253224
rect 302420 253212 302426 253224
rect 349650 253212 349656 253224
rect 302420 253184 349656 253212
rect 302420 253172 302426 253184
rect 349650 253172 349656 253184
rect 349708 253172 349714 253224
rect 350846 253172 350852 253224
rect 350904 253212 350910 253224
rect 581490 253212 581496 253224
rect 350904 253184 581496 253212
rect 350904 253172 350910 253184
rect 581490 253172 581496 253184
rect 581548 253172 581554 253224
rect 1600 252912 583316 253008
rect 1600 252368 583316 252464
rect 1600 251824 583316 251920
rect 1600 251280 583316 251376
rect 278810 251200 278816 251252
rect 278868 251200 278874 251252
rect 285253 251243 285311 251249
rect 285253 251209 285265 251243
rect 285299 251240 285311 251243
rect 285342 251240 285348 251252
rect 285299 251212 285348 251240
rect 285299 251209 285311 251212
rect 285253 251203 285311 251209
rect 285342 251200 285348 251212
rect 285400 251200 285406 251252
rect 285621 251243 285679 251249
rect 285621 251209 285633 251243
rect 285667 251240 285679 251243
rect 285710 251240 285716 251252
rect 285667 251212 285716 251240
rect 285667 251209 285679 251212
rect 285621 251203 285679 251209
rect 285710 251200 285716 251212
rect 285768 251200 285774 251252
rect 331250 251240 331256 251252
rect 331211 251212 331256 251240
rect 331250 251200 331256 251212
rect 331308 251200 331314 251252
rect 341097 251243 341155 251249
rect 341097 251209 341109 251243
rect 341143 251240 341155 251243
rect 341186 251240 341192 251252
rect 341143 251212 341192 251240
rect 341143 251209 341155 251212
rect 341097 251203 341155 251209
rect 341186 251200 341192 251212
rect 341244 251200 341250 251252
rect 91498 251172 91504 251184
rect 91459 251144 91504 251172
rect 91498 251132 91504 251144
rect 91556 251132 91562 251184
rect 225358 251172 225364 251184
rect 225319 251144 225364 251172
rect 225358 251132 225364 251144
rect 225416 251132 225422 251184
rect 229958 251172 229964 251184
rect 229919 251144 229964 251172
rect 229958 251132 229964 251144
rect 230016 251132 230022 251184
rect 278828 251116 278856 251200
rect 357930 251132 357936 251184
rect 357988 251172 357994 251184
rect 553890 251172 553896 251184
rect 357988 251144 358033 251172
rect 553851 251144 553896 251172
rect 357988 251132 357994 251144
rect 553890 251132 553896 251144
rect 553948 251132 553954 251184
rect 278810 251064 278816 251116
rect 278868 251064 278874 251116
rect 1600 250736 583316 250832
rect 1600 250192 583316 250288
rect 135474 249772 135480 249824
rect 135532 249812 135538 249824
rect 135658 249812 135664 249824
rect 135532 249784 135664 249812
rect 135532 249772 135538 249784
rect 135658 249772 135664 249784
rect 135716 249772 135722 249824
rect 152034 249772 152040 249824
rect 152092 249812 152098 249824
rect 152218 249812 152224 249824
rect 152092 249784 152224 249812
rect 152092 249772 152098 249784
rect 152218 249772 152224 249784
rect 152276 249772 152282 249824
rect 170158 249772 170164 249824
rect 170216 249812 170222 249824
rect 170342 249812 170348 249824
rect 170216 249784 170348 249812
rect 170216 249772 170222 249784
rect 170342 249772 170348 249784
rect 170400 249772 170406 249824
rect 190674 249772 190680 249824
rect 190732 249812 190738 249824
rect 190858 249812 190864 249824
rect 190732 249784 190864 249812
rect 190732 249772 190738 249784
rect 190858 249772 190864 249784
rect 190916 249772 190922 249824
rect 214318 249772 214324 249824
rect 214376 249812 214382 249824
rect 214502 249812 214508 249824
rect 214376 249784 214508 249812
rect 214376 249772 214382 249784
rect 214502 249772 214508 249784
rect 214560 249772 214566 249824
rect 246518 249812 246524 249824
rect 246479 249784 246524 249812
rect 246518 249772 246524 249784
rect 246576 249772 246582 249824
rect 305033 249815 305091 249821
rect 305033 249781 305045 249815
rect 305079 249812 305091 249815
rect 305122 249812 305128 249824
rect 305079 249784 305128 249812
rect 305079 249781 305091 249784
rect 305033 249775 305091 249781
rect 305122 249772 305128 249784
rect 305180 249772 305186 249824
rect 372926 249772 372932 249824
rect 372984 249812 372990 249824
rect 373110 249812 373116 249824
rect 372984 249784 373116 249812
rect 372984 249772 372990 249784
rect 373110 249772 373116 249784
rect 373168 249772 373174 249824
rect 385530 249772 385536 249824
rect 385588 249812 385594 249824
rect 385714 249812 385720 249824
rect 385588 249784 385720 249812
rect 385588 249772 385594 249784
rect 385714 249772 385720 249784
rect 385772 249772 385778 249824
rect 392430 249772 392436 249824
rect 392488 249812 392494 249824
rect 392614 249812 392620 249824
rect 392488 249784 392620 249812
rect 392488 249772 392494 249784
rect 392614 249772 392620 249784
rect 392672 249772 392678 249824
rect 528866 249772 528872 249824
rect 528924 249812 528930 249824
rect 529050 249812 529056 249824
rect 528924 249784 529056 249812
rect 528924 249772 528930 249784
rect 529050 249772 529056 249784
rect 529108 249772 529114 249824
rect 535950 249772 535956 249824
rect 536008 249812 536014 249824
rect 536134 249812 536140 249824
rect 536008 249784 536140 249812
rect 536008 249772 536014 249784
rect 536134 249772 536140 249784
rect 536192 249772 536198 249824
rect 571830 249772 571836 249824
rect 571888 249812 571894 249824
rect 572014 249812 572020 249824
rect 571888 249784 572020 249812
rect 571888 249772 571894 249784
rect 572014 249772 572020 249784
rect 572072 249772 572078 249824
rect 1600 249648 583316 249744
rect 1600 249104 583316 249200
rect 1600 248560 583316 248656
rect 1600 248016 583316 248112
rect 1600 247472 583316 247568
rect 1600 246928 583316 247024
rect 242746 246820 242752 246832
rect 242707 246792 242752 246820
rect 242746 246780 242752 246792
rect 242804 246780 242810 246832
rect 1600 246384 583316 246480
rect 1600 245840 583316 245936
rect 242565 245667 242623 245673
rect 242565 245633 242577 245667
rect 242611 245664 242623 245667
rect 242654 245664 242660 245676
rect 242611 245636 242660 245664
rect 242611 245633 242623 245636
rect 242565 245627 242623 245633
rect 242654 245624 242660 245636
rect 242712 245624 242718 245676
rect 275590 245664 275596 245676
rect 275551 245636 275596 245664
rect 275590 245624 275596 245636
rect 275648 245624 275654 245676
rect 1600 245296 583316 245392
rect 1600 244752 583316 244848
rect 239250 244332 239256 244384
rect 239308 244372 239314 244384
rect 239434 244372 239440 244384
rect 239308 244344 239440 244372
rect 239308 244332 239314 244344
rect 239434 244332 239440 244344
rect 239492 244332 239498 244384
rect 285342 244372 285348 244384
rect 285303 244344 285348 244372
rect 285342 244332 285348 244344
rect 285400 244332 285406 244384
rect 1600 244208 583316 244304
rect 3822 244128 3828 244180
rect 3880 244168 3886 244180
rect 228854 244168 228860 244180
rect 3880 244140 228860 244168
rect 3880 244128 3886 244140
rect 228854 244128 228860 244140
rect 228912 244128 228918 244180
rect 229958 244168 229964 244180
rect 229919 244140 229964 244168
rect 229958 244128 229964 244140
rect 230016 244128 230022 244180
rect 239250 244128 239256 244180
rect 239308 244168 239314 244180
rect 239434 244168 239440 244180
rect 239308 244140 239440 244168
rect 239308 244128 239314 244140
rect 239434 244128 239440 244140
rect 239492 244128 239498 244180
rect 285342 244168 285348 244180
rect 285303 244140 285348 244168
rect 285342 244128 285348 244140
rect 285400 244128 285406 244180
rect 1600 243664 583316 243760
rect 328306 243448 328312 243500
rect 328364 243488 328370 243500
rect 328398 243488 328404 243500
rect 328364 243460 328404 243488
rect 328364 243448 328370 243460
rect 328398 243448 328404 243460
rect 328456 243448 328462 243500
rect 1600 243120 583316 243216
rect 1600 242576 583316 242672
rect 1600 242032 583316 242128
rect 242746 241992 242752 242004
rect 242707 241964 242752 241992
rect 242746 241952 242752 241964
rect 242804 241952 242810 242004
rect 251670 241748 251676 241800
rect 251728 241788 251734 241800
rect 261146 241788 261152 241800
rect 251728 241760 261152 241788
rect 251728 241748 251734 241760
rect 261146 241748 261152 241760
rect 261204 241748 261210 241800
rect 91498 241652 91504 241664
rect 91459 241624 91504 241652
rect 91498 241612 91504 241624
rect 91556 241612 91562 241664
rect 225358 241652 225364 241664
rect 225319 241624 225364 241652
rect 225358 241612 225364 241624
rect 225416 241612 225422 241664
rect 290310 241612 290316 241664
rect 290368 241652 290374 241664
rect 294818 241652 294824 241664
rect 290368 241624 294824 241652
rect 290368 241612 290374 241624
rect 294818 241612 294824 241624
rect 294876 241612 294882 241664
rect 357930 241612 357936 241664
rect 357988 241652 357994 241664
rect 553890 241652 553896 241664
rect 357988 241624 358033 241652
rect 553851 241624 553896 241652
rect 357988 241612 357994 241624
rect 553890 241612 553896 241624
rect 553948 241612 553954 241664
rect 1600 241488 583316 241584
rect 246426 241408 246432 241460
rect 246484 241448 246490 241460
rect 246702 241448 246708 241460
rect 246484 241420 246708 241448
rect 246484 241408 246490 241420
rect 246702 241408 246708 241420
rect 246760 241408 246766 241460
rect 309170 241448 309176 241460
rect 309131 241420 309176 241448
rect 309170 241408 309176 241420
rect 309228 241408 309234 241460
rect 1600 240944 583316 241040
rect 1600 240400 583316 240496
rect 279454 240116 279460 240168
rect 279512 240156 279518 240168
rect 279730 240156 279736 240168
rect 279512 240128 279736 240156
rect 279512 240116 279518 240128
rect 279730 240116 279736 240128
rect 279788 240116 279794 240168
rect 235478 240088 235484 240100
rect 235439 240060 235484 240088
rect 235478 240048 235484 240060
rect 235536 240048 235542 240100
rect 1600 239856 583316 239952
rect 1600 239312 583316 239408
rect 1600 238768 583316 238864
rect 1600 238224 583316 238320
rect 1600 237680 583316 237776
rect 242470 237368 242476 237380
rect 242431 237340 242476 237368
rect 242470 237328 242476 237340
rect 242528 237328 242534 237380
rect 276694 237328 276700 237380
rect 276752 237368 276758 237380
rect 276878 237368 276884 237380
rect 276752 237340 276884 237368
rect 276752 237328 276758 237340
rect 276878 237328 276884 237340
rect 276936 237328 276942 237380
rect 1600 237136 583316 237232
rect 285342 236756 285348 236768
rect 285303 236728 285348 236756
rect 285342 236716 285348 236728
rect 285400 236716 285406 236768
rect 1600 236592 583316 236688
rect 1600 236048 583316 236144
rect 273014 236008 273020 236020
rect 272975 235980 273020 236008
rect 273014 235968 273020 235980
rect 273072 235968 273078 236020
rect 272830 235940 272836 235952
rect 272791 235912 272836 235940
rect 272830 235900 272836 235912
rect 272888 235900 272894 235952
rect 328306 235940 328312 235952
rect 328267 235912 328312 235940
rect 328306 235900 328312 235912
rect 328364 235900 328370 235952
rect 1600 235504 583316 235600
rect 1600 234960 583316 235056
rect 371822 234716 371828 234728
rect 371748 234688 371828 234716
rect 371748 234592 371776 234688
rect 371822 234676 371828 234688
rect 371880 234676 371886 234728
rect 275682 234580 275688 234592
rect 275643 234552 275688 234580
rect 275682 234540 275688 234552
rect 275740 234540 275746 234592
rect 371730 234540 371736 234592
rect 371788 234540 371794 234592
rect 1600 234416 583316 234512
rect 309170 234376 309176 234388
rect 309131 234348 309176 234376
rect 309170 234336 309176 234348
rect 309228 234336 309234 234388
rect 319934 234336 319940 234388
rect 319992 234376 319998 234388
rect 320118 234376 320124 234388
rect 319992 234348 320124 234376
rect 319992 234336 319998 234348
rect 320118 234336 320124 234348
rect 320176 234336 320182 234388
rect 1600 233872 583316 233968
rect 1600 233328 583316 233424
rect 1600 232784 583316 232880
rect 276513 232611 276571 232617
rect 276513 232577 276525 232611
rect 276559 232608 276571 232611
rect 276602 232608 276608 232620
rect 276559 232580 276608 232608
rect 276559 232577 276571 232580
rect 276513 232571 276571 232577
rect 276602 232568 276608 232580
rect 276660 232568 276666 232620
rect 277062 232500 277068 232552
rect 277120 232540 277126 232552
rect 277246 232540 277252 232552
rect 277120 232512 277252 232540
rect 277120 232500 277126 232512
rect 277246 232500 277252 232512
rect 277304 232500 277310 232552
rect 1600 232240 583316 232336
rect 285342 231928 285348 231940
rect 285303 231900 285348 231928
rect 285342 231888 285348 231900
rect 285400 231888 285406 231940
rect 242102 231820 242108 231872
rect 242160 231860 242166 231872
rect 242194 231860 242200 231872
rect 242160 231832 242200 231860
rect 242160 231820 242166 231832
rect 242194 231820 242200 231832
rect 242252 231820 242258 231872
rect 246610 231820 246616 231872
rect 246668 231860 246674 231872
rect 246702 231860 246708 231872
rect 246668 231832 246708 231860
rect 246668 231820 246674 231832
rect 246702 231820 246708 231832
rect 246760 231820 246766 231872
rect 285710 231820 285716 231872
rect 285768 231860 285774 231872
rect 285802 231860 285808 231872
rect 285768 231832 285808 231860
rect 285768 231820 285774 231832
rect 285802 231820 285808 231832
rect 285860 231820 285866 231872
rect 331066 231820 331072 231872
rect 331124 231860 331130 231872
rect 331250 231860 331256 231872
rect 331124 231832 331256 231860
rect 331124 231820 331130 231832
rect 331250 231820 331256 231832
rect 331308 231820 331314 231872
rect 341002 231820 341008 231872
rect 341060 231860 341066 231872
rect 341094 231860 341100 231872
rect 341060 231832 341100 231860
rect 341060 231820 341066 231832
rect 341094 231820 341100 231832
rect 341152 231820 341158 231872
rect 1600 231696 583316 231792
rect 272833 231591 272891 231597
rect 272833 231557 272845 231591
rect 272879 231588 272891 231591
rect 272922 231588 272928 231600
rect 272879 231560 272928 231588
rect 272879 231557 272891 231560
rect 272833 231551 272891 231557
rect 272922 231548 272928 231560
rect 272980 231548 272986 231600
rect 1600 231152 583316 231248
rect 1600 230608 583316 230704
rect 135474 230460 135480 230512
rect 135532 230500 135538 230512
rect 135658 230500 135664 230512
rect 135532 230472 135664 230500
rect 135532 230460 135538 230472
rect 135658 230460 135664 230472
rect 135716 230460 135722 230512
rect 152034 230460 152040 230512
rect 152092 230500 152098 230512
rect 152218 230500 152224 230512
rect 152092 230472 152224 230500
rect 152092 230460 152098 230472
rect 152218 230460 152224 230472
rect 152276 230460 152282 230512
rect 170158 230460 170164 230512
rect 170216 230500 170222 230512
rect 170342 230500 170348 230512
rect 170216 230472 170348 230500
rect 170216 230460 170222 230472
rect 170342 230460 170348 230472
rect 170400 230460 170406 230512
rect 190674 230460 190680 230512
rect 190732 230500 190738 230512
rect 190858 230500 190864 230512
rect 190732 230472 190864 230500
rect 190732 230460 190738 230472
rect 190858 230460 190864 230472
rect 190916 230460 190922 230512
rect 214318 230460 214324 230512
rect 214376 230500 214382 230512
rect 214502 230500 214508 230512
rect 214376 230472 214508 230500
rect 214376 230460 214382 230472
rect 214502 230460 214508 230472
rect 214560 230460 214566 230512
rect 235481 230503 235539 230509
rect 235481 230469 235493 230503
rect 235527 230500 235539 230503
rect 235662 230500 235668 230512
rect 235527 230472 235668 230500
rect 235527 230469 235539 230472
rect 235481 230463 235539 230469
rect 235662 230460 235668 230472
rect 235720 230460 235726 230512
rect 385530 230460 385536 230512
rect 385588 230500 385594 230512
rect 385714 230500 385720 230512
rect 385588 230472 385720 230500
rect 385588 230460 385594 230472
rect 385714 230460 385720 230472
rect 385772 230460 385778 230512
rect 392430 230460 392436 230512
rect 392488 230500 392494 230512
rect 392614 230500 392620 230512
rect 392488 230472 392620 230500
rect 392488 230460 392494 230472
rect 392614 230460 392620 230472
rect 392672 230460 392678 230512
rect 528866 230460 528872 230512
rect 528924 230500 528930 230512
rect 529050 230500 529056 230512
rect 528924 230472 529056 230500
rect 528924 230460 528930 230472
rect 529050 230460 529056 230472
rect 529108 230460 529114 230512
rect 535950 230460 535956 230512
rect 536008 230500 536014 230512
rect 536134 230500 536140 230512
rect 536008 230472 536140 230500
rect 536008 230460 536014 230472
rect 536134 230460 536140 230472
rect 536192 230460 536198 230512
rect 552326 230460 552332 230512
rect 552384 230500 552390 230512
rect 552418 230500 552424 230512
rect 552384 230472 552424 230500
rect 552384 230460 552390 230472
rect 552418 230460 552424 230472
rect 552476 230460 552482 230512
rect 571830 230460 571836 230512
rect 571888 230500 571894 230512
rect 572014 230500 572020 230512
rect 571888 230472 572020 230500
rect 571888 230460 571894 230472
rect 572014 230460 572020 230472
rect 572072 230460 572078 230512
rect 1600 230064 583316 230160
rect 1600 229520 583316 229616
rect 1600 228976 583316 229072
rect 1600 228432 583316 228528
rect 1600 227888 583316 227984
rect 242473 227783 242531 227789
rect 242473 227749 242485 227783
rect 242519 227780 242531 227783
rect 242838 227780 242844 227792
rect 242519 227752 242844 227780
rect 242519 227749 242531 227752
rect 242473 227743 242531 227749
rect 242838 227740 242844 227752
rect 242896 227740 242902 227792
rect 276510 227740 276516 227792
rect 276568 227780 276574 227792
rect 276568 227752 276613 227780
rect 276568 227740 276574 227752
rect 1600 227344 583316 227440
rect 268690 227032 268696 227044
rect 268651 227004 268696 227032
rect 268690 226992 268696 227004
rect 268748 226992 268754 227044
rect 1600 226800 583316 226896
rect 300430 226584 300436 226636
rect 300488 226624 300494 226636
rect 308158 226624 308164 226636
rect 300488 226596 308164 226624
rect 300488 226584 300494 226596
rect 308158 226584 308164 226596
rect 308216 226584 308222 226636
rect 360598 226516 360604 226568
rect 360656 226556 360662 226568
rect 362254 226556 362260 226568
rect 360656 226528 362260 226556
rect 360656 226516 360662 226528
rect 362254 226516 362260 226528
rect 362312 226516 362318 226568
rect 1600 226256 583316 226352
rect 1600 225712 583316 225808
rect 239250 225632 239256 225684
rect 239308 225672 239314 225684
rect 239434 225672 239440 225684
rect 239308 225644 239440 225672
rect 239308 225632 239314 225644
rect 239434 225632 239440 225644
rect 239492 225632 239498 225684
rect 1600 225168 583316 225264
rect 341094 225060 341100 225072
rect 341020 225032 341100 225060
rect 229774 224952 229780 225004
rect 229832 224992 229838 225004
rect 229958 224992 229964 225004
rect 229832 224964 229964 224992
rect 229832 224952 229838 224964
rect 229958 224952 229964 224964
rect 230016 224952 230022 225004
rect 275682 224992 275688 225004
rect 275643 224964 275688 224992
rect 275682 224952 275688 224964
rect 275740 224952 275746 225004
rect 285253 224995 285311 225001
rect 285253 224961 285265 224995
rect 285299 224992 285311 224995
rect 285342 224992 285348 225004
rect 285299 224964 285348 224992
rect 285299 224961 285311 224964
rect 285253 224955 285311 224961
rect 285342 224952 285348 224964
rect 285400 224952 285406 225004
rect 285526 224952 285532 225004
rect 285584 224992 285590 225004
rect 285710 224992 285716 225004
rect 285584 224964 285716 224992
rect 285584 224952 285590 224964
rect 285710 224952 285716 224964
rect 285768 224952 285774 225004
rect 304938 224952 304944 225004
rect 304996 224952 305002 225004
rect 320026 224992 320032 225004
rect 319987 224964 320032 224992
rect 320026 224952 320032 224964
rect 320084 224952 320090 225004
rect 271358 224884 271364 224936
rect 271416 224924 271422 224936
rect 271542 224924 271548 224936
rect 271416 224896 271548 224924
rect 271416 224884 271422 224896
rect 271542 224884 271548 224896
rect 271600 224884 271606 224936
rect 272922 224884 272928 224936
rect 272980 224924 272986 224936
rect 272980 224896 273025 224924
rect 272980 224884 272986 224896
rect 304956 224868 304984 224952
rect 341020 224936 341048 225032
rect 341094 225020 341100 225032
rect 341152 225020 341158 225072
rect 341002 224884 341008 224936
rect 341060 224884 341066 224936
rect 275593 224859 275651 224865
rect 275593 224825 275605 224859
rect 275639 224856 275651 224859
rect 275682 224856 275688 224868
rect 275639 224828 275688 224856
rect 275639 224825 275651 224828
rect 275593 224819 275651 224825
rect 275682 224816 275688 224828
rect 275740 224816 275746 224868
rect 304938 224816 304944 224868
rect 304996 224816 305002 224868
rect 1600 224624 583316 224720
rect 1600 224080 583316 224176
rect 1600 223536 583316 223632
rect 1600 222992 583316 223088
rect 1600 222448 583316 222544
rect 239342 222232 239348 222284
rect 239400 222232 239406 222284
rect 242194 222272 242200 222284
rect 242120 222244 242200 222272
rect 91314 222164 91320 222216
rect 91372 222204 91378 222216
rect 91498 222204 91504 222216
rect 91372 222176 91504 222204
rect 91372 222164 91378 222176
rect 91498 222164 91504 222176
rect 91556 222164 91562 222216
rect 239360 222148 239388 222232
rect 242120 222148 242148 222244
rect 242194 222232 242200 222244
rect 242252 222232 242258 222284
rect 246610 222272 246616 222284
rect 246536 222244 246616 222272
rect 246536 222148 246564 222244
rect 246610 222232 246616 222244
rect 246668 222232 246674 222284
rect 246794 222164 246800 222216
rect 246852 222164 246858 222216
rect 268693 222207 268751 222213
rect 268693 222173 268705 222207
rect 268739 222204 268751 222207
rect 268782 222204 268788 222216
rect 268739 222176 268788 222204
rect 268739 222173 268751 222176
rect 268693 222167 268751 222173
rect 268782 222164 268788 222176
rect 268840 222164 268846 222216
rect 276694 222164 276700 222216
rect 276752 222204 276758 222216
rect 276878 222204 276884 222216
rect 276752 222176 276884 222204
rect 276752 222164 276758 222176
rect 276878 222164 276884 222176
rect 276936 222164 276942 222216
rect 357930 222164 357936 222216
rect 357988 222204 357994 222216
rect 358114 222204 358120 222216
rect 357988 222176 358120 222204
rect 357988 222164 357994 222176
rect 358114 222164 358120 222176
rect 358172 222164 358178 222216
rect 371546 222164 371552 222216
rect 371604 222204 371610 222216
rect 371822 222204 371828 222216
rect 371604 222176 371828 222204
rect 371604 222164 371610 222176
rect 371822 222164 371828 222176
rect 371880 222164 371886 222216
rect 553706 222164 553712 222216
rect 553764 222204 553770 222216
rect 553890 222204 553896 222216
rect 553764 222176 553896 222204
rect 553764 222164 553770 222176
rect 553890 222164 553896 222176
rect 553948 222164 553954 222216
rect 239342 222096 239348 222148
rect 239400 222096 239406 222148
rect 242102 222096 242108 222148
rect 242160 222096 242166 222148
rect 246518 222096 246524 222148
rect 246576 222096 246582 222148
rect 246812 222080 246840 222164
rect 246794 222028 246800 222080
rect 246852 222028 246858 222080
rect 1600 221904 583316 222000
rect 1600 221360 583316 221456
rect 320026 220980 320032 220992
rect 319987 220952 320032 220980
rect 320026 220940 320032 220952
rect 320084 220940 320090 220992
rect 1600 220816 583316 220912
rect 276694 220776 276700 220788
rect 276655 220748 276700 220776
rect 276694 220736 276700 220748
rect 276752 220736 276758 220788
rect 341002 220776 341008 220788
rect 340963 220748 341008 220776
rect 341002 220736 341008 220748
rect 341060 220736 341066 220788
rect 373202 220776 373208 220788
rect 373163 220748 373208 220776
rect 373202 220736 373208 220748
rect 373260 220736 373266 220788
rect 1600 220272 583316 220368
rect 1600 219728 583316 219824
rect 279730 219444 279736 219496
rect 279788 219484 279794 219496
rect 279822 219484 279828 219496
rect 279788 219456 279828 219484
rect 279788 219444 279794 219456
rect 279822 219444 279828 219456
rect 279880 219444 279886 219496
rect 285250 219484 285256 219496
rect 285211 219456 285256 219484
rect 285250 219444 285256 219456
rect 285308 219444 285314 219496
rect 1600 219184 583316 219280
rect 1600 218640 583316 218736
rect 1600 218096 583316 218192
rect 272922 217988 272928 218000
rect 272883 217960 272928 217988
rect 272922 217948 272928 217960
rect 272980 217948 272986 218000
rect 1600 217552 583316 217648
rect 1600 217008 583316 217104
rect 242470 216628 242476 216640
rect 242431 216600 242476 216628
rect 242470 216588 242476 216600
rect 242528 216588 242534 216640
rect 1600 216464 583316 216560
rect 1600 215920 583316 216016
rect 1600 215376 583316 215472
rect 275590 215336 275596 215348
rect 275551 215308 275596 215336
rect 275590 215296 275596 215308
rect 275648 215296 275654 215348
rect 272830 215268 272836 215280
rect 272791 215240 272836 215268
rect 272830 215228 272836 215240
rect 272888 215228 272894 215280
rect 341005 215271 341063 215277
rect 341005 215237 341017 215271
rect 341051 215268 341063 215271
rect 341094 215268 341100 215280
rect 341051 215240 341100 215268
rect 341051 215237 341063 215240
rect 341005 215231 341063 215237
rect 341094 215228 341100 215240
rect 341152 215228 341158 215280
rect 1600 214832 583316 214928
rect 1600 214288 583316 214384
rect 1600 213744 583316 213840
rect 1600 213200 583316 213296
rect 1600 212656 583316 212752
rect 331066 212508 331072 212560
rect 331124 212548 331130 212560
rect 331250 212548 331256 212560
rect 331124 212520 331256 212548
rect 331124 212508 331130 212520
rect 331250 212508 331256 212520
rect 331308 212508 331314 212560
rect 553706 212508 553712 212560
rect 553764 212548 553770 212560
rect 553890 212548 553896 212560
rect 553764 212520 553896 212548
rect 553764 212508 553770 212520
rect 553890 212508 553896 212520
rect 553948 212508 553954 212560
rect 279730 212440 279736 212492
rect 279788 212480 279794 212492
rect 279822 212480 279828 212492
rect 279788 212452 279828 212480
rect 279788 212440 279794 212452
rect 279822 212440 279828 212452
rect 279880 212440 279886 212492
rect 357930 212440 357936 212492
rect 357988 212480 357994 212492
rect 373202 212480 373208 212492
rect 357988 212452 358033 212480
rect 373163 212452 373208 212480
rect 357988 212440 357994 212452
rect 373202 212440 373208 212452
rect 373260 212440 373266 212492
rect 1600 212112 583316 212208
rect 1600 211568 583316 211664
rect 275590 211256 275596 211268
rect 275551 211228 275596 211256
rect 275590 211216 275596 211228
rect 275648 211216 275654 211268
rect 235386 211148 235392 211200
rect 235444 211188 235450 211200
rect 235478 211188 235484 211200
rect 235444 211160 235484 211188
rect 235444 211148 235450 211160
rect 235478 211148 235484 211160
rect 235536 211148 235542 211200
rect 276694 211188 276700 211200
rect 276655 211160 276700 211188
rect 276694 211148 276700 211160
rect 276752 211148 276758 211200
rect 328306 211188 328312 211200
rect 328267 211160 328312 211188
rect 328306 211148 328312 211160
rect 328364 211148 328370 211200
rect 385530 211148 385536 211200
rect 385588 211188 385594 211200
rect 385714 211188 385720 211200
rect 385588 211160 385720 211188
rect 385588 211148 385594 211160
rect 385714 211148 385720 211160
rect 385772 211148 385778 211200
rect 392430 211148 392436 211200
rect 392488 211188 392494 211200
rect 392614 211188 392620 211200
rect 392488 211160 392620 211188
rect 392488 211148 392494 211160
rect 392614 211148 392620 211160
rect 392672 211148 392678 211200
rect 528866 211148 528872 211200
rect 528924 211188 528930 211200
rect 529050 211188 529056 211200
rect 528924 211160 529056 211188
rect 528924 211148 528930 211160
rect 529050 211148 529056 211160
rect 529108 211148 529114 211200
rect 535950 211148 535956 211200
rect 536008 211188 536014 211200
rect 536134 211188 536140 211200
rect 536008 211160 536140 211188
rect 536008 211148 536014 211160
rect 536134 211148 536140 211160
rect 536192 211148 536198 211200
rect 552326 211148 552332 211200
rect 552384 211188 552390 211200
rect 552510 211188 552516 211200
rect 552384 211160 552516 211188
rect 552384 211148 552390 211160
rect 552510 211148 552516 211160
rect 552568 211148 552574 211200
rect 571830 211148 571836 211200
rect 571888 211188 571894 211200
rect 572014 211188 572020 211200
rect 571888 211160 572020 211188
rect 571888 211148 571894 211160
rect 572014 211148 572020 211160
rect 572072 211148 572078 211200
rect 1600 211024 583316 211120
rect 1600 210480 583316 210576
rect 272830 210440 272836 210452
rect 272791 210412 272836 210440
rect 272830 210400 272836 210412
rect 272888 210400 272894 210452
rect 275590 210440 275596 210452
rect 275551 210412 275596 210440
rect 275590 210400 275596 210412
rect 275648 210400 275654 210452
rect 1600 209936 583316 210032
rect 3730 209720 3736 209772
rect 3788 209760 3794 209772
rect 224714 209760 224720 209772
rect 3788 209732 224720 209760
rect 3788 209720 3794 209732
rect 224714 209720 224720 209732
rect 224772 209720 224778 209772
rect 328398 209760 328404 209772
rect 328359 209732 328404 209760
rect 328398 209720 328404 209732
rect 328456 209720 328462 209772
rect 1600 209392 583316 209488
rect 1600 208848 583316 208944
rect 285250 208564 285256 208616
rect 285308 208564 285314 208616
rect 285268 208480 285296 208564
rect 285250 208428 285256 208480
rect 285308 208428 285314 208480
rect 1600 208304 583316 208400
rect 285069 208267 285127 208273
rect 285069 208233 285081 208267
rect 285115 208264 285127 208267
rect 285250 208264 285256 208276
rect 285115 208236 285256 208264
rect 285115 208233 285127 208236
rect 285069 208227 285127 208233
rect 285250 208224 285256 208236
rect 285308 208224 285314 208276
rect 1600 207760 583316 207856
rect 268690 207720 268696 207732
rect 268651 207692 268696 207720
rect 268690 207680 268696 207692
rect 268748 207680 268754 207732
rect 1600 207216 583316 207312
rect 242470 207040 242476 207052
rect 242431 207012 242476 207040
rect 242470 207000 242476 207012
rect 242528 207000 242534 207052
rect 273014 206932 273020 206984
rect 273072 206932 273078 206984
rect 273032 206904 273060 206932
rect 273106 206904 273112 206916
rect 273032 206876 273112 206904
rect 273106 206864 273112 206876
rect 273164 206864 273170 206916
rect 1600 206672 583316 206768
rect 1600 206128 583316 206224
rect 229961 205819 230019 205825
rect 229961 205785 229973 205819
rect 230007 205816 230019 205819
rect 230050 205816 230056 205828
rect 230007 205788 230056 205816
rect 230007 205785 230019 205788
rect 229961 205779 230019 205785
rect 230050 205776 230056 205788
rect 230108 205776 230114 205828
rect 341097 205819 341155 205825
rect 341097 205785 341109 205819
rect 341143 205816 341155 205819
rect 341186 205816 341192 205828
rect 341143 205788 341192 205816
rect 341143 205785 341155 205788
rect 341097 205779 341155 205785
rect 341186 205776 341192 205788
rect 341244 205776 341250 205828
rect 235478 205748 235484 205760
rect 235439 205720 235484 205748
rect 235478 205708 235484 205720
rect 235536 205708 235542 205760
rect 271450 205748 271456 205760
rect 271411 205720 271456 205748
rect 271450 205708 271456 205720
rect 271508 205708 271514 205760
rect 309078 205748 309084 205760
rect 309039 205720 309084 205748
rect 309078 205708 309084 205720
rect 309136 205708 309142 205760
rect 1600 205584 583316 205680
rect 229958 205544 229964 205556
rect 229919 205516 229964 205544
rect 229958 205504 229964 205516
rect 230016 205504 230022 205556
rect 239250 205504 239256 205556
rect 239308 205544 239314 205556
rect 239434 205544 239440 205556
rect 239308 205516 239440 205544
rect 239308 205504 239314 205516
rect 239434 205504 239440 205516
rect 239492 205504 239498 205556
rect 268693 205547 268751 205553
rect 268693 205513 268705 205547
rect 268739 205544 268751 205547
rect 268782 205544 268788 205556
rect 268739 205516 268788 205544
rect 268739 205513 268751 205516
rect 268693 205507 268751 205513
rect 268782 205504 268788 205516
rect 268840 205504 268846 205556
rect 271450 205544 271456 205556
rect 271411 205516 271456 205544
rect 271450 205504 271456 205516
rect 271508 205504 271514 205556
rect 309078 205544 309084 205556
rect 309039 205516 309084 205544
rect 309078 205504 309084 205516
rect 309136 205504 309142 205556
rect 341094 205544 341100 205556
rect 341055 205516 341100 205544
rect 341094 205504 341100 205516
rect 341152 205504 341158 205556
rect 1600 205040 583316 205136
rect 328398 204932 328404 204944
rect 328359 204904 328404 204932
rect 328398 204892 328404 204904
rect 328456 204892 328462 204944
rect 1600 204496 583316 204592
rect 1600 203952 583316 204048
rect 1600 203408 583316 203504
rect 91314 202988 91320 203040
rect 91372 203028 91378 203040
rect 91498 203028 91504 203040
rect 91372 203000 91504 203028
rect 91372 202988 91378 203000
rect 91498 202988 91504 203000
rect 91556 202988 91562 203040
rect 225358 202988 225364 203040
rect 225416 203028 225422 203040
rect 225542 203028 225548 203040
rect 225416 203000 225548 203028
rect 225416 202988 225422 203000
rect 225542 202988 225548 203000
rect 225600 202988 225606 203040
rect 235478 203028 235484 203040
rect 235439 203000 235484 203028
rect 235478 202988 235484 203000
rect 235536 202988 235542 203040
rect 357930 202988 357936 203040
rect 357988 203028 357994 203040
rect 357988 203000 358033 203028
rect 357988 202988 357994 203000
rect 1600 202864 583316 202960
rect 235570 202824 235576 202836
rect 235531 202796 235576 202824
rect 235570 202784 235576 202796
rect 235628 202784 235634 202836
rect 341094 202824 341100 202836
rect 341055 202796 341100 202824
rect 341094 202784 341100 202796
rect 341152 202784 341158 202836
rect 1600 202320 583316 202416
rect 1600 201776 583316 201872
rect 242470 201492 242476 201544
rect 242528 201492 242534 201544
rect 285618 201492 285624 201544
rect 285676 201532 285682 201544
rect 285710 201532 285716 201544
rect 285676 201504 285716 201532
rect 285676 201492 285682 201504
rect 285710 201492 285716 201504
rect 285768 201492 285774 201544
rect 135474 201424 135480 201476
rect 135532 201464 135538 201476
rect 135658 201464 135664 201476
rect 135532 201436 135664 201464
rect 135532 201424 135538 201436
rect 135658 201424 135664 201436
rect 135716 201424 135722 201476
rect 152034 201424 152040 201476
rect 152092 201464 152098 201476
rect 152218 201464 152224 201476
rect 152092 201436 152224 201464
rect 152092 201424 152098 201436
rect 152218 201424 152224 201436
rect 152276 201424 152282 201476
rect 170158 201424 170164 201476
rect 170216 201464 170222 201476
rect 170342 201464 170348 201476
rect 170216 201436 170348 201464
rect 170216 201424 170222 201436
rect 170342 201424 170348 201436
rect 170400 201424 170406 201476
rect 190674 201424 190680 201476
rect 190732 201464 190738 201476
rect 190858 201464 190864 201476
rect 190732 201436 190864 201464
rect 190732 201424 190738 201436
rect 190858 201424 190864 201436
rect 190916 201424 190922 201476
rect 214318 201424 214324 201476
rect 214376 201464 214382 201476
rect 214502 201464 214508 201476
rect 214376 201436 214508 201464
rect 214376 201424 214382 201436
rect 214502 201424 214508 201436
rect 214560 201424 214566 201476
rect 242488 201396 242516 201492
rect 268506 201424 268512 201476
rect 268564 201464 268570 201476
rect 268782 201464 268788 201476
rect 268564 201436 268788 201464
rect 268564 201424 268570 201436
rect 268782 201424 268788 201436
rect 268840 201424 268846 201476
rect 385530 201424 385536 201476
rect 385588 201464 385594 201476
rect 385714 201464 385720 201476
rect 385588 201436 385720 201464
rect 385588 201424 385594 201436
rect 385714 201424 385720 201436
rect 385772 201424 385778 201476
rect 392430 201424 392436 201476
rect 392488 201464 392494 201476
rect 392614 201464 392620 201476
rect 392488 201436 392620 201464
rect 392488 201424 392494 201436
rect 392614 201424 392620 201436
rect 392672 201424 392678 201476
rect 528866 201424 528872 201476
rect 528924 201464 528930 201476
rect 529050 201464 529056 201476
rect 528924 201436 529056 201464
rect 528924 201424 528930 201436
rect 529050 201424 529056 201436
rect 529108 201424 529114 201476
rect 535950 201424 535956 201476
rect 536008 201464 536014 201476
rect 536134 201464 536140 201476
rect 536008 201436 536140 201464
rect 536008 201424 536014 201436
rect 536134 201424 536140 201436
rect 536192 201424 536198 201476
rect 552418 201464 552424 201476
rect 552379 201436 552424 201464
rect 552418 201424 552424 201436
rect 552476 201424 552482 201476
rect 571830 201424 571836 201476
rect 571888 201464 571894 201476
rect 572014 201464 572020 201476
rect 571888 201436 572020 201464
rect 571888 201424 571894 201436
rect 572014 201424 572020 201436
rect 572072 201424 572078 201476
rect 242562 201396 242568 201408
rect 242488 201368 242568 201396
rect 242562 201356 242568 201368
rect 242620 201356 242626 201408
rect 1600 201232 583316 201328
rect 1600 200688 583316 200784
rect 1600 200144 583316 200240
rect 279822 200104 279828 200116
rect 279783 200076 279828 200104
rect 279822 200064 279828 200076
rect 279880 200064 279886 200116
rect 320026 200104 320032 200116
rect 319987 200076 320032 200104
rect 320026 200064 320032 200076
rect 320084 200064 320090 200116
rect 372006 200104 372012 200116
rect 371967 200076 372012 200104
rect 372006 200064 372012 200076
rect 372064 200064 372070 200116
rect 373021 200107 373079 200113
rect 373021 200073 373033 200107
rect 373067 200104 373079 200107
rect 373110 200104 373116 200116
rect 373067 200076 373116 200104
rect 373067 200073 373079 200076
rect 373021 200067 373079 200073
rect 373110 200064 373116 200076
rect 373168 200064 373174 200116
rect 328398 200036 328404 200048
rect 328359 200008 328404 200036
rect 328398 199996 328404 200008
rect 328456 199996 328462 200048
rect 1600 199600 583316 199696
rect 1600 199056 583316 199152
rect 285066 198744 285072 198756
rect 285027 198716 285072 198744
rect 285066 198704 285072 198716
rect 285124 198704 285130 198756
rect 242473 198679 242531 198685
rect 242473 198645 242485 198679
rect 242519 198676 242531 198679
rect 242562 198676 242568 198688
rect 242519 198648 242568 198676
rect 242519 198645 242531 198648
rect 242473 198639 242531 198645
rect 242562 198636 242568 198648
rect 242620 198636 242626 198688
rect 1600 198512 583316 198608
rect 276970 198132 276976 198144
rect 276931 198104 276976 198132
rect 276970 198092 276976 198104
rect 277028 198092 277034 198144
rect 1600 197968 583316 198064
rect 275590 197548 275596 197600
rect 275648 197588 275654 197600
rect 275685 197591 275743 197597
rect 275685 197588 275697 197591
rect 275648 197560 275697 197588
rect 275648 197548 275654 197560
rect 275685 197557 275697 197560
rect 275731 197557 275743 197591
rect 275685 197551 275743 197557
rect 1600 197424 583316 197520
rect 275682 197344 275688 197396
rect 275740 197384 275746 197396
rect 275740 197356 275785 197384
rect 275740 197344 275746 197356
rect 1600 196880 583316 196976
rect 1600 196336 583316 196432
rect 552418 196296 552424 196308
rect 552379 196268 552424 196296
rect 552418 196256 552424 196268
rect 552476 196256 552482 196308
rect 320026 195956 320032 195968
rect 319987 195928 320032 195956
rect 320026 195916 320032 195928
rect 320084 195916 320090 195968
rect 353054 195916 353060 195968
rect 353112 195956 353118 195968
rect 580662 195956 580668 195968
rect 353112 195928 580668 195956
rect 353112 195916 353118 195928
rect 580662 195916 580668 195928
rect 580720 195916 580726 195968
rect 1600 195792 583316 195888
rect 235570 195752 235576 195764
rect 235531 195724 235576 195752
rect 235570 195712 235576 195724
rect 235628 195712 235634 195764
rect 328398 195752 328404 195764
rect 328359 195724 328404 195752
rect 328398 195712 328404 195724
rect 328456 195712 328462 195764
rect 1600 195248 583316 195344
rect 1600 194704 583316 194800
rect 1600 194160 583316 194256
rect 246702 193876 246708 193928
rect 246760 193916 246766 193928
rect 246978 193916 246984 193928
rect 246760 193888 246984 193916
rect 246760 193876 246766 193888
rect 246978 193876 246984 193888
rect 247036 193876 247042 193928
rect 1600 193616 583316 193712
rect 341097 193375 341155 193381
rect 341097 193341 341109 193375
rect 341143 193372 341155 193375
rect 341186 193372 341192 193384
rect 341143 193344 341192 193372
rect 341143 193341 341155 193344
rect 341097 193335 341155 193341
rect 341186 193332 341192 193344
rect 341244 193332 341250 193384
rect 331066 193196 331072 193248
rect 331124 193236 331130 193248
rect 331250 193236 331256 193248
rect 331124 193208 331256 193236
rect 331124 193196 331130 193208
rect 331250 193196 331256 193208
rect 331308 193196 331314 193248
rect 553706 193196 553712 193248
rect 553764 193236 553770 193248
rect 553890 193236 553896 193248
rect 553764 193208 553896 193236
rect 553764 193196 553770 193208
rect 553890 193196 553896 193208
rect 553948 193196 553954 193248
rect 1600 193072 583316 193168
rect 3822 192652 3828 192704
rect 3880 192692 3886 192704
rect 9434 192692 9440 192704
rect 3880 192664 9440 192692
rect 3880 192652 3886 192664
rect 9434 192652 9440 192664
rect 9492 192652 9498 192704
rect 1600 192528 583316 192624
rect 1600 191984 583316 192080
rect 235570 191768 235576 191820
rect 235628 191808 235634 191820
rect 235754 191808 235760 191820
rect 235628 191780 235760 191808
rect 235628 191768 235634 191780
rect 235754 191768 235760 191780
rect 235812 191768 235818 191820
rect 552418 191808 552424 191820
rect 552379 191780 552424 191808
rect 552418 191768 552424 191780
rect 552476 191768 552482 191820
rect 1600 191440 583316 191536
rect 372006 191264 372012 191276
rect 371967 191236 372012 191264
rect 372006 191224 372012 191236
rect 372064 191224 372070 191276
rect 1600 190896 583316 190992
rect 373018 190584 373024 190596
rect 372979 190556 373024 190584
rect 373018 190544 373024 190556
rect 373076 190544 373082 190596
rect 279822 190516 279828 190528
rect 279783 190488 279828 190516
rect 279822 190476 279828 190488
rect 279880 190476 279886 190528
rect 1600 190352 583316 190448
rect 1600 189808 583316 189904
rect 1600 189264 583316 189360
rect 242470 189088 242476 189100
rect 242431 189060 242476 189088
rect 242470 189048 242476 189060
rect 242528 189048 242534 189100
rect 246426 189048 246432 189100
rect 246484 189088 246490 189100
rect 246610 189088 246616 189100
rect 246484 189060 246616 189088
rect 246484 189048 246490 189060
rect 246610 189048 246616 189060
rect 246668 189048 246674 189100
rect 272922 189048 272928 189100
rect 272980 189048 272986 189100
rect 276970 189088 276976 189100
rect 276931 189060 276976 189088
rect 276970 189048 276976 189060
rect 277028 189048 277034 189100
rect 242838 189020 242844 189032
rect 242799 188992 242844 189020
rect 242838 188980 242844 188992
rect 242896 188980 242902 189032
rect 272940 188964 272968 189048
rect 272922 188912 272928 188964
rect 272980 188912 272986 188964
rect 1600 188720 583316 188816
rect 1600 188176 583316 188272
rect 1600 187632 583316 187728
rect 1600 187088 583316 187184
rect 1600 186544 583316 186640
rect 229774 186328 229780 186380
rect 229832 186368 229838 186380
rect 229958 186368 229964 186380
rect 229832 186340 229964 186368
rect 229832 186328 229838 186340
rect 229958 186328 229964 186340
rect 230016 186328 230022 186380
rect 285526 186328 285532 186380
rect 285584 186328 285590 186380
rect 305030 186328 305036 186380
rect 305088 186368 305094 186380
rect 305214 186368 305220 186380
rect 305088 186340 305220 186368
rect 305088 186328 305094 186340
rect 305214 186328 305220 186340
rect 305272 186328 305278 186380
rect 308989 186371 309047 186377
rect 308989 186337 309001 186371
rect 309035 186368 309047 186371
rect 309078 186368 309084 186380
rect 309035 186340 309084 186368
rect 309035 186337 309047 186340
rect 308989 186331 309047 186337
rect 309078 186328 309084 186340
rect 309136 186328 309142 186380
rect 341094 186368 341100 186380
rect 341055 186340 341100 186368
rect 341094 186328 341100 186340
rect 341152 186328 341158 186380
rect 285066 186260 285072 186312
rect 285124 186300 285130 186312
rect 285250 186300 285256 186312
rect 285124 186272 285256 186300
rect 285124 186260 285130 186272
rect 285250 186260 285256 186272
rect 285308 186260 285314 186312
rect 285544 186232 285572 186328
rect 285618 186232 285624 186244
rect 285544 186204 285624 186232
rect 285618 186192 285624 186204
rect 285676 186192 285682 186244
rect 1600 186000 583316 186096
rect 1600 185456 583316 185552
rect 1600 184912 583316 185008
rect 1600 184368 583316 184464
rect 1600 183824 583316 183920
rect 279822 183648 279828 183660
rect 279748 183620 279828 183648
rect 91314 183540 91320 183592
rect 91372 183580 91378 183592
rect 91498 183580 91504 183592
rect 91372 183552 91504 183580
rect 91372 183540 91378 183552
rect 91498 183540 91504 183552
rect 91556 183540 91562 183592
rect 279748 183524 279776 183620
rect 279822 183608 279828 183620
rect 279880 183608 279886 183660
rect 341094 183648 341100 183660
rect 341055 183620 341100 183648
rect 341094 183608 341100 183620
rect 341152 183608 341158 183660
rect 308986 183580 308992 183592
rect 308947 183552 308992 183580
rect 308986 183540 308992 183552
rect 309044 183540 309050 183592
rect 357930 183540 357936 183592
rect 357988 183580 357994 183592
rect 358114 183580 358120 183592
rect 357988 183552 358120 183580
rect 357988 183540 357994 183552
rect 358114 183540 358120 183552
rect 358172 183540 358178 183592
rect 553706 183540 553712 183592
rect 553764 183580 553770 183592
rect 553890 183580 553896 183592
rect 553764 183552 553896 183580
rect 553764 183540 553770 183552
rect 553890 183540 553896 183552
rect 553948 183540 553954 183592
rect 279730 183472 279736 183524
rect 279788 183472 279794 183524
rect 341094 183472 341100 183524
rect 341152 183512 341158 183524
rect 341462 183512 341468 183524
rect 341152 183484 341468 183512
rect 341152 183472 341158 183484
rect 341462 183472 341468 183484
rect 341520 183472 341526 183524
rect 552418 183512 552424 183524
rect 552379 183484 552424 183512
rect 552418 183472 552424 183484
rect 552476 183472 552482 183524
rect 1600 183280 583316 183376
rect 1600 182736 583316 182832
rect 1600 182192 583316 182288
rect 135474 182112 135480 182164
rect 135532 182152 135538 182164
rect 135658 182152 135664 182164
rect 135532 182124 135664 182152
rect 135532 182112 135538 182124
rect 135658 182112 135664 182124
rect 135716 182112 135722 182164
rect 152034 182112 152040 182164
rect 152092 182152 152098 182164
rect 152218 182152 152224 182164
rect 152092 182124 152224 182152
rect 152092 182112 152098 182124
rect 152218 182112 152224 182124
rect 152276 182112 152282 182164
rect 170158 182112 170164 182164
rect 170216 182152 170222 182164
rect 170342 182152 170348 182164
rect 170216 182124 170348 182152
rect 170216 182112 170222 182124
rect 170342 182112 170348 182124
rect 170400 182112 170406 182164
rect 190674 182112 190680 182164
rect 190732 182152 190738 182164
rect 190858 182152 190864 182164
rect 190732 182124 190864 182152
rect 190732 182112 190738 182124
rect 190858 182112 190864 182124
rect 190916 182112 190922 182164
rect 214318 182112 214324 182164
rect 214376 182152 214382 182164
rect 214502 182152 214508 182164
rect 214376 182124 214508 182152
rect 214376 182112 214382 182124
rect 214502 182112 214508 182124
rect 214560 182112 214566 182164
rect 229866 182152 229872 182164
rect 229827 182124 229872 182152
rect 229866 182112 229872 182124
rect 229924 182112 229930 182164
rect 242102 182112 242108 182164
rect 242160 182152 242166 182164
rect 242194 182152 242200 182164
rect 242160 182124 242200 182152
rect 242160 182112 242166 182124
rect 242194 182112 242200 182124
rect 242252 182112 242258 182164
rect 246518 182112 246524 182164
rect 246576 182152 246582 182164
rect 246610 182152 246616 182164
rect 246576 182124 246616 182152
rect 246576 182112 246582 182124
rect 246610 182112 246616 182124
rect 246668 182112 246674 182164
rect 285158 182152 285164 182164
rect 285119 182124 285164 182152
rect 285158 182112 285164 182124
rect 285216 182112 285222 182164
rect 285618 182112 285624 182164
rect 285676 182152 285682 182164
rect 285710 182152 285716 182164
rect 285676 182124 285716 182152
rect 285676 182112 285682 182124
rect 285710 182112 285716 182124
rect 285768 182112 285774 182164
rect 328306 182152 328312 182164
rect 328267 182124 328312 182152
rect 328306 182112 328312 182124
rect 328364 182112 328370 182164
rect 385530 182112 385536 182164
rect 385588 182152 385594 182164
rect 385714 182152 385720 182164
rect 385588 182124 385720 182152
rect 385588 182112 385594 182124
rect 385714 182112 385720 182124
rect 385772 182112 385778 182164
rect 392430 182112 392436 182164
rect 392488 182152 392494 182164
rect 392614 182152 392620 182164
rect 392488 182124 392620 182152
rect 392488 182112 392494 182124
rect 392614 182112 392620 182124
rect 392672 182112 392678 182164
rect 528866 182112 528872 182164
rect 528924 182152 528930 182164
rect 529050 182152 529056 182164
rect 528924 182124 529056 182152
rect 528924 182112 528930 182124
rect 529050 182112 529056 182124
rect 529108 182112 529114 182164
rect 535950 182112 535956 182164
rect 536008 182152 536014 182164
rect 536134 182152 536140 182164
rect 536008 182124 536140 182152
rect 536008 182112 536014 182124
rect 536134 182112 536140 182124
rect 536192 182112 536198 182164
rect 571830 182112 571836 182164
rect 571888 182152 571894 182164
rect 572014 182152 572020 182164
rect 571888 182124 572020 182152
rect 571888 182112 571894 182124
rect 572014 182112 572020 182124
rect 572072 182112 572078 182164
rect 242838 182016 242844 182028
rect 242799 181988 242844 182016
rect 242838 181976 242844 181988
rect 242896 181976 242902 182028
rect 1600 181648 583316 181744
rect 295186 181432 295192 181484
rect 295244 181472 295250 181484
rect 308250 181472 308256 181484
rect 295244 181444 308256 181472
rect 295244 181432 295250 181444
rect 308250 181432 308256 181444
rect 308308 181432 308314 181484
rect 1600 181104 583316 181200
rect 273014 180752 273020 180804
rect 273072 180792 273078 180804
rect 273106 180792 273112 180804
rect 273072 180764 273112 180792
rect 273072 180752 273078 180764
rect 273106 180752 273112 180764
rect 273164 180752 273170 180804
rect 278810 180792 278816 180804
rect 278771 180764 278816 180792
rect 278810 180752 278816 180764
rect 278868 180752 278874 180804
rect 371914 180752 371920 180804
rect 371972 180792 371978 180804
rect 372006 180792 372012 180804
rect 371972 180764 372012 180792
rect 371972 180752 371978 180764
rect 372006 180752 372012 180764
rect 372064 180752 372070 180804
rect 1600 180560 583316 180656
rect 1600 180016 583316 180112
rect 1600 179472 583316 179568
rect 251670 179392 251676 179444
rect 251728 179432 251734 179444
rect 259858 179432 259864 179444
rect 251728 179404 259864 179432
rect 251728 179392 251734 179404
rect 259858 179392 259864 179404
rect 259916 179392 259922 179444
rect 371914 179364 371920 179376
rect 371875 179336 371920 179364
rect 371914 179324 371920 179336
rect 371972 179324 371978 179376
rect 1600 178928 583316 179024
rect 304846 178712 304852 178764
rect 304904 178752 304910 178764
rect 305122 178752 305128 178764
rect 304904 178724 305128 178752
rect 304904 178712 304910 178724
rect 305122 178712 305128 178724
rect 305180 178712 305186 178764
rect 1600 178384 583316 178480
rect 1600 177840 583316 177936
rect 1600 177296 583316 177392
rect 319750 177216 319756 177268
rect 319808 177256 319814 177268
rect 320026 177256 320032 177268
rect 319808 177228 320032 177256
rect 319808 177216 319814 177228
rect 320026 177216 320032 177228
rect 320084 177216 320090 177268
rect 1600 176752 583316 176848
rect 235478 176672 235484 176724
rect 235536 176672 235542 176724
rect 229866 176576 229872 176588
rect 229827 176548 229872 176576
rect 229866 176536 229872 176548
rect 229924 176536 229930 176588
rect 235496 176576 235524 176672
rect 235570 176576 235576 176588
rect 235496 176548 235576 176576
rect 235570 176536 235576 176548
rect 235628 176536 235634 176588
rect 328309 176579 328367 176585
rect 328309 176545 328321 176579
rect 328355 176576 328367 176579
rect 328398 176576 328404 176588
rect 328355 176548 328404 176576
rect 328355 176545 328367 176548
rect 328309 176539 328367 176545
rect 328398 176536 328404 176548
rect 328456 176536 328462 176588
rect 1600 176208 583316 176304
rect 1600 175664 583316 175760
rect 1600 175120 583316 175216
rect 1600 174576 583316 174672
rect 1600 174032 583316 174128
rect 268506 173884 268512 173936
rect 268564 173924 268570 173936
rect 268690 173924 268696 173936
rect 268564 173896 268696 173924
rect 268564 173884 268570 173896
rect 268690 173884 268696 173896
rect 268748 173884 268754 173936
rect 308986 173884 308992 173936
rect 309044 173924 309050 173936
rect 309078 173924 309084 173936
rect 309044 173896 309084 173924
rect 309044 173884 309050 173896
rect 309078 173884 309084 173896
rect 309136 173884 309142 173936
rect 331066 173884 331072 173936
rect 331124 173924 331130 173936
rect 331250 173924 331256 173936
rect 331124 173896 331256 173924
rect 331124 173884 331130 173896
rect 331250 173884 331256 173896
rect 331308 173884 331314 173936
rect 1600 173488 583316 173584
rect 275590 173244 275596 173256
rect 275551 173216 275596 173244
rect 275590 173204 275596 173216
rect 275648 173204 275654 173256
rect 1600 172944 583316 173040
rect 285158 172564 285164 172576
rect 285119 172536 285164 172564
rect 285158 172524 285164 172536
rect 285216 172524 285222 172576
rect 1600 172400 583316 172496
rect 1600 171856 583316 171952
rect 1600 171312 583316 171408
rect 278810 171136 278816 171148
rect 278771 171108 278816 171136
rect 278810 171096 278816 171108
rect 278868 171096 278874 171148
rect 1600 170768 583316 170864
rect 1600 170224 583316 170320
rect 1600 169680 583316 169776
rect 246889 169303 246947 169309
rect 246889 169269 246901 169303
rect 246935 169300 246947 169303
rect 246978 169300 246984 169312
rect 246935 169272 246984 169300
rect 246935 169269 246947 169272
rect 246889 169263 246947 169269
rect 246978 169260 246984 169272
rect 247036 169260 247042 169312
rect 1600 169136 583316 169232
rect 1600 168592 583316 168688
rect 273017 168351 273075 168357
rect 273017 168317 273029 168351
rect 273063 168348 273075 168351
rect 273106 168348 273112 168360
rect 273063 168320 273112 168348
rect 273063 168317 273075 168320
rect 273017 168311 273075 168317
rect 273106 168308 273112 168320
rect 273164 168308 273170 168360
rect 1600 168048 583316 168144
rect 1600 167504 583316 167600
rect 235481 167195 235539 167201
rect 235481 167161 235493 167195
rect 235527 167192 235539 167195
rect 235570 167192 235576 167204
rect 235527 167164 235576 167192
rect 235527 167161 235539 167164
rect 235481 167155 235539 167161
rect 235570 167152 235576 167164
rect 235628 167152 235634 167204
rect 239250 167084 239256 167136
rect 239308 167124 239314 167136
rect 239434 167124 239440 167136
rect 239308 167096 239440 167124
rect 239308 167084 239314 167096
rect 239434 167084 239440 167096
rect 239492 167084 239498 167136
rect 1600 166960 583316 167056
rect 235478 166920 235484 166932
rect 235439 166892 235484 166920
rect 235478 166880 235484 166892
rect 235536 166880 235542 166932
rect 239250 166880 239256 166932
rect 239308 166920 239314 166932
rect 239434 166920 239440 166932
rect 239308 166892 239440 166920
rect 239308 166880 239314 166892
rect 239434 166880 239440 166892
rect 239492 166880 239498 166932
rect 285710 166812 285716 166864
rect 285768 166812 285774 166864
rect 285728 166728 285756 166812
rect 285710 166676 285716 166728
rect 285768 166676 285774 166728
rect 1600 166416 583316 166512
rect 272922 166308 272928 166320
rect 272848 166280 272928 166308
rect 272848 166252 272876 166280
rect 272922 166268 272928 166280
rect 272980 166268 272986 166320
rect 272830 166200 272836 166252
rect 272888 166200 272894 166252
rect 1600 165872 583316 165968
rect 1600 165328 583316 165424
rect 1600 164784 583316 164880
rect 284790 164364 284796 164416
rect 284848 164404 284854 164416
rect 285618 164404 285624 164416
rect 284848 164376 285624 164404
rect 284848 164364 284854 164376
rect 285618 164364 285624 164376
rect 285676 164364 285682 164416
rect 382034 164364 382040 164416
rect 382092 164404 382098 164416
rect 385806 164404 385812 164416
rect 382092 164376 385812 164404
rect 382092 164364 382098 164376
rect 385806 164364 385812 164376
rect 385864 164364 385870 164416
rect 391694 164364 391700 164416
rect 391752 164404 391758 164416
rect 392706 164404 392712 164416
rect 391752 164376 392712 164404
rect 391752 164364 391758 164376
rect 392706 164364 392712 164376
rect 392764 164364 392770 164416
rect 526934 164364 526940 164416
rect 526992 164404 526998 164416
rect 529326 164404 529332 164416
rect 526992 164376 529332 164404
rect 526992 164364 526998 164376
rect 529326 164364 529332 164376
rect 529384 164364 529390 164416
rect 535674 164364 535680 164416
rect 535732 164404 535738 164416
rect 536594 164404 536600 164416
rect 535732 164376 536600 164404
rect 535732 164364 535738 164376
rect 536594 164364 536600 164376
rect 536652 164364 536658 164416
rect 552510 164364 552516 164416
rect 552568 164404 552574 164416
rect 552694 164404 552700 164416
rect 552568 164376 552700 164404
rect 552568 164364 552574 164376
rect 552694 164364 552700 164376
rect 552752 164364 552758 164416
rect 571554 164364 571560 164416
rect 571612 164404 571618 164416
rect 572106 164404 572112 164416
rect 571612 164376 572112 164404
rect 571612 164364 571618 164376
rect 572106 164364 572112 164376
rect 572164 164364 572170 164416
rect 1600 164240 583316 164336
rect 242102 164160 242108 164212
rect 242160 164160 242166 164212
rect 242654 164200 242660 164212
rect 242615 164172 242660 164200
rect 242654 164160 242660 164172
rect 242712 164160 242718 164212
rect 246518 164160 246524 164212
rect 246576 164160 246582 164212
rect 259306 164200 259312 164212
rect 259267 164172 259312 164200
rect 259306 164160 259312 164172
rect 259364 164160 259370 164212
rect 305122 164200 305128 164212
rect 305083 164172 305128 164200
rect 305122 164160 305128 164172
rect 305180 164160 305186 164212
rect 308986 164160 308992 164212
rect 309044 164200 309050 164212
rect 309078 164200 309084 164212
rect 309044 164172 309084 164200
rect 309044 164160 309050 164172
rect 309078 164160 309084 164172
rect 309136 164160 309142 164212
rect 331066 164160 331072 164212
rect 331124 164200 331130 164212
rect 331250 164200 331256 164212
rect 331124 164172 331256 164200
rect 331124 164160 331130 164172
rect 331250 164160 331256 164172
rect 331308 164160 331314 164212
rect 341002 164160 341008 164212
rect 341060 164200 341066 164212
rect 341094 164200 341100 164212
rect 341060 164172 341100 164200
rect 341060 164160 341066 164172
rect 341094 164160 341100 164172
rect 341152 164160 341158 164212
rect 553890 164200 553896 164212
rect 553851 164172 553896 164200
rect 553890 164160 553896 164172
rect 553948 164160 553954 164212
rect 242120 164132 242148 164160
rect 242194 164132 242200 164144
rect 242120 164104 242200 164132
rect 242194 164092 242200 164104
rect 242252 164092 242258 164144
rect 246536 164132 246564 164160
rect 246610 164132 246616 164144
rect 246536 164104 246616 164132
rect 246610 164092 246616 164104
rect 246668 164092 246674 164144
rect 320026 164092 320032 164144
rect 320084 164132 320090 164144
rect 320118 164132 320124 164144
rect 320084 164104 320124 164132
rect 320084 164092 320090 164104
rect 320118 164092 320124 164104
rect 320176 164092 320182 164144
rect 1600 163696 583316 163792
rect 273014 163520 273020 163532
rect 272975 163492 273020 163520
rect 273014 163480 273020 163492
rect 273072 163480 273078 163532
rect 275590 163520 275596 163532
rect 275551 163492 275596 163520
rect 275590 163480 275596 163492
rect 275648 163480 275654 163532
rect 1600 163152 583316 163248
rect 242562 162908 242568 162920
rect 242488 162880 242568 162908
rect 135658 162840 135664 162852
rect 135619 162812 135664 162840
rect 135658 162800 135664 162812
rect 135716 162800 135722 162852
rect 152218 162840 152224 162852
rect 152179 162812 152224 162840
rect 152218 162800 152224 162812
rect 152276 162800 152282 162852
rect 170158 162840 170164 162852
rect 170119 162812 170164 162840
rect 170158 162800 170164 162812
rect 170216 162800 170222 162852
rect 190858 162840 190864 162852
rect 190819 162812 190864 162840
rect 190858 162800 190864 162812
rect 190916 162800 190922 162852
rect 214318 162840 214324 162852
rect 214279 162812 214324 162840
rect 214318 162800 214324 162812
rect 214376 162800 214382 162852
rect 230050 162840 230056 162852
rect 230011 162812 230056 162840
rect 230050 162800 230056 162812
rect 230108 162800 230114 162852
rect 242010 162800 242016 162852
rect 242068 162840 242074 162852
rect 242194 162840 242200 162852
rect 242068 162812 242200 162840
rect 242068 162800 242074 162812
rect 242194 162800 242200 162812
rect 242252 162800 242258 162852
rect 242488 162849 242516 162880
rect 242562 162868 242568 162880
rect 242620 162868 242626 162920
rect 242473 162843 242531 162849
rect 242473 162809 242485 162843
rect 242519 162809 242531 162843
rect 246610 162840 246616 162852
rect 246571 162812 246616 162840
rect 242473 162803 242531 162809
rect 246610 162800 246616 162812
rect 246668 162800 246674 162852
rect 385530 162800 385536 162852
rect 385588 162840 385594 162852
rect 392430 162840 392436 162852
rect 385588 162812 385633 162840
rect 392391 162812 392436 162840
rect 385588 162800 385594 162812
rect 392430 162800 392436 162812
rect 392488 162800 392494 162852
rect 529050 162840 529056 162852
rect 529011 162812 529056 162840
rect 529050 162800 529056 162812
rect 529108 162800 529114 162852
rect 535950 162840 535956 162852
rect 535911 162812 535956 162840
rect 535950 162800 535956 162812
rect 536008 162800 536014 162852
rect 552510 162840 552516 162852
rect 552471 162812 552516 162840
rect 552510 162800 552516 162812
rect 552568 162800 552574 162852
rect 571830 162840 571836 162852
rect 571791 162812 571836 162840
rect 571830 162800 571836 162812
rect 571888 162800 571894 162852
rect 1600 162608 583316 162704
rect 1600 162064 583316 162160
rect 1600 161520 583316 161616
rect 246886 161480 246892 161492
rect 246847 161452 246892 161480
rect 246886 161440 246892 161452
rect 246944 161440 246950 161492
rect 285250 161440 285256 161492
rect 285308 161480 285314 161492
rect 285342 161480 285348 161492
rect 285308 161452 285348 161480
rect 285308 161440 285314 161452
rect 285342 161440 285348 161452
rect 285400 161440 285406 161492
rect 371917 161483 371975 161489
rect 371917 161449 371929 161483
rect 371963 161480 371975 161483
rect 372006 161480 372012 161492
rect 371963 161452 372012 161480
rect 371963 161449 371975 161452
rect 371917 161443 371975 161449
rect 372006 161440 372012 161452
rect 372064 161440 372070 161492
rect 268506 161276 268512 161288
rect 268467 161248 268512 161276
rect 268506 161236 268512 161248
rect 268564 161236 268570 161288
rect 1600 160976 583316 161072
rect 1600 160432 583316 160528
rect 1600 159888 583316 159984
rect 246797 159511 246855 159517
rect 246797 159477 246809 159511
rect 246843 159508 246855 159511
rect 246886 159508 246892 159520
rect 246843 159480 246892 159508
rect 246843 159477 246855 159480
rect 246797 159471 246855 159477
rect 246886 159468 246892 159480
rect 246944 159468 246950 159520
rect 1600 159344 583316 159440
rect 235478 159304 235484 159316
rect 235439 159276 235484 159304
rect 235478 159264 235484 159276
rect 235536 159264 235542 159316
rect 1600 158800 583316 158896
rect 273014 158652 273020 158704
rect 273072 158692 273078 158704
rect 273106 158692 273112 158704
rect 273072 158664 273112 158692
rect 273072 158652 273078 158664
rect 273106 158652 273112 158664
rect 273164 158652 273170 158704
rect 1600 158256 583316 158352
rect 319842 157972 319848 158024
rect 319900 158012 319906 158024
rect 320118 158012 320124 158024
rect 319900 157984 320124 158012
rect 319900 157972 319906 157984
rect 320118 157972 320124 157984
rect 320176 157972 320182 158024
rect 242470 157944 242476 157956
rect 242431 157916 242476 157944
rect 242470 157904 242476 157916
rect 242528 157904 242534 157956
rect 1600 157712 583316 157808
rect 285253 157403 285311 157409
rect 285253 157369 285265 157403
rect 285299 157400 285311 157403
rect 285342 157400 285348 157412
rect 285299 157372 285348 157400
rect 285299 157369 285311 157372
rect 285253 157363 285311 157369
rect 285342 157360 285348 157372
rect 285400 157360 285406 157412
rect 259306 157332 259312 157344
rect 259267 157304 259312 157332
rect 259306 157292 259312 157304
rect 259364 157292 259370 157344
rect 273017 157335 273075 157341
rect 273017 157301 273029 157335
rect 273063 157332 273075 157335
rect 273106 157332 273112 157344
rect 273063 157304 273112 157332
rect 273063 157301 273075 157304
rect 273017 157295 273075 157301
rect 273106 157292 273112 157304
rect 273164 157292 273170 157344
rect 275590 157332 275596 157344
rect 275551 157304 275596 157332
rect 275590 157292 275596 157304
rect 275648 157292 275654 157344
rect 305122 157332 305128 157344
rect 305083 157304 305128 157332
rect 305122 157292 305128 157304
rect 305180 157292 305186 157344
rect 1600 157168 583316 157264
rect 230050 157128 230056 157140
rect 230011 157100 230056 157128
rect 230050 157088 230056 157100
rect 230108 157088 230114 157140
rect 235481 157131 235539 157137
rect 235481 157097 235493 157131
rect 235527 157128 235539 157131
rect 235570 157128 235576 157140
rect 235527 157100 235576 157128
rect 235527 157097 235539 157100
rect 235481 157091 235539 157097
rect 235570 157088 235576 157100
rect 235628 157088 235634 157140
rect 242654 157128 242660 157140
rect 242615 157100 242660 157128
rect 242654 157088 242660 157100
rect 242712 157088 242718 157140
rect 246794 157128 246800 157140
rect 246755 157100 246800 157128
rect 246794 157088 246800 157100
rect 246852 157088 246858 157140
rect 268509 157131 268567 157137
rect 268509 157097 268521 157131
rect 268555 157128 268567 157131
rect 268690 157128 268696 157140
rect 268555 157100 268696 157128
rect 268555 157097 268567 157100
rect 268509 157091 268567 157097
rect 268690 157088 268696 157100
rect 268748 157088 268754 157140
rect 285069 156791 285127 156797
rect 285069 156757 285081 156791
rect 285115 156788 285127 156791
rect 285158 156788 285164 156800
rect 285115 156760 285164 156788
rect 285115 156757 285127 156760
rect 285069 156751 285127 156757
rect 285158 156748 285164 156760
rect 285216 156748 285222 156800
rect 1600 156624 583316 156720
rect 1600 156080 583316 156176
rect 1600 155536 583316 155632
rect 1600 154992 583316 155088
rect 553890 154680 553896 154692
rect 553851 154652 553896 154680
rect 553890 154640 553896 154652
rect 553948 154640 553954 154692
rect 1600 154448 583316 154544
rect 268690 154408 268696 154420
rect 268651 154380 268696 154408
rect 268690 154368 268696 154380
rect 268748 154368 268754 154420
rect 1600 153904 583316 154000
rect 1600 153360 583316 153456
rect 135658 153252 135664 153264
rect 135619 153224 135664 153252
rect 135658 153212 135664 153224
rect 135716 153212 135722 153264
rect 152218 153252 152224 153264
rect 152179 153224 152224 153252
rect 152218 153212 152224 153224
rect 152276 153212 152282 153264
rect 170158 153252 170164 153264
rect 170119 153224 170164 153252
rect 170158 153212 170164 153224
rect 170216 153212 170222 153264
rect 190858 153252 190864 153264
rect 190819 153224 190864 153252
rect 190858 153212 190864 153224
rect 190916 153212 190922 153264
rect 214318 153252 214324 153264
rect 214279 153224 214324 153252
rect 214318 153212 214324 153224
rect 214376 153212 214382 153264
rect 246610 153252 246616 153264
rect 246571 153224 246616 153252
rect 246610 153212 246616 153224
rect 246668 153212 246674 153264
rect 372006 153252 372012 153264
rect 371932 153224 372012 153252
rect 371932 153196 371960 153224
rect 372006 153212 372012 153224
rect 372064 153212 372070 153264
rect 385530 153212 385536 153264
rect 385588 153252 385594 153264
rect 392430 153252 392436 153264
rect 385588 153224 385633 153252
rect 392391 153224 392436 153252
rect 385588 153212 385594 153224
rect 392430 153212 392436 153224
rect 392488 153212 392494 153264
rect 529050 153252 529056 153264
rect 529011 153224 529056 153252
rect 529050 153212 529056 153224
rect 529108 153212 529114 153264
rect 535950 153252 535956 153264
rect 535911 153224 535956 153252
rect 535950 153212 535956 153224
rect 536008 153212 536014 153264
rect 552510 153252 552516 153264
rect 552471 153224 552516 153252
rect 552510 153212 552516 153224
rect 552568 153212 552574 153264
rect 571830 153252 571836 153264
rect 571791 153224 571836 153252
rect 571830 153212 571836 153224
rect 571888 153212 571894 153264
rect 371914 153144 371920 153196
rect 371972 153144 371978 153196
rect 373110 153184 373116 153196
rect 373071 153156 373116 153184
rect 373110 153144 373116 153156
rect 373168 153144 373174 153196
rect 1600 152816 583316 152912
rect 1600 152272 583316 152368
rect 1600 151728 583316 151824
rect 1600 151184 583316 151280
rect 1600 150640 583316 150736
rect 1600 150096 583316 150192
rect 278718 149852 278724 149864
rect 278679 149824 278724 149852
rect 278718 149812 278724 149824
rect 278776 149812 278782 149864
rect 1600 149552 583316 149648
rect 271450 149132 271456 149184
rect 271508 149172 271514 149184
rect 271542 149172 271548 149184
rect 271508 149144 271548 149172
rect 271508 149132 271514 149144
rect 271542 149132 271548 149144
rect 271600 149132 271606 149184
rect 1600 149008 583316 149104
rect 351674 148928 351680 148980
rect 351732 148968 351738 148980
rect 580386 148968 580392 148980
rect 351732 148940 580392 148968
rect 351732 148928 351738 148940
rect 580386 148928 580392 148940
rect 580444 148928 580450 148980
rect 1600 148464 583316 148560
rect 1600 147920 583316 148016
rect 246610 147744 246616 147756
rect 246536 147716 246616 147744
rect 246536 147620 246564 147716
rect 246610 147704 246616 147716
rect 246668 147704 246674 147756
rect 341186 147744 341192 147756
rect 341112 147716 341192 147744
rect 273014 147676 273020 147688
rect 272975 147648 273020 147676
rect 273014 147636 273020 147648
rect 273072 147636 273078 147688
rect 275593 147679 275651 147685
rect 275593 147645 275605 147679
rect 275639 147676 275651 147679
rect 275682 147676 275688 147688
rect 275639 147648 275688 147676
rect 275639 147645 275651 147648
rect 275593 147639 275651 147645
rect 275682 147636 275688 147648
rect 275740 147636 275746 147688
rect 285526 147636 285532 147688
rect 285584 147676 285590 147688
rect 285710 147676 285716 147688
rect 285584 147648 285716 147676
rect 285584 147636 285590 147648
rect 285710 147636 285716 147648
rect 285768 147636 285774 147688
rect 305030 147636 305036 147688
rect 305088 147676 305094 147688
rect 305214 147676 305220 147688
rect 305088 147648 305220 147676
rect 305088 147636 305094 147648
rect 305214 147636 305220 147648
rect 305272 147636 305278 147688
rect 341112 147620 341140 147716
rect 341186 147704 341192 147716
rect 341244 147704 341250 147756
rect 246518 147568 246524 147620
rect 246576 147568 246582 147620
rect 268690 147608 268696 147620
rect 268651 147580 268696 147608
rect 268690 147568 268696 147580
rect 268748 147568 268754 147620
rect 341094 147568 341100 147620
rect 341152 147568 341158 147620
rect 1600 147376 583316 147472
rect 1600 146832 583316 146928
rect 1600 146288 583316 146384
rect 1600 145744 583316 145840
rect 1600 145200 583316 145296
rect 373110 145160 373116 145172
rect 373071 145132 373116 145160
rect 373110 145120 373116 145132
rect 373168 145120 373174 145172
rect 320026 144984 320032 145036
rect 320084 145024 320090 145036
rect 320118 145024 320124 145036
rect 320084 144996 320124 145024
rect 320084 144984 320090 144996
rect 320118 144984 320124 144996
rect 320176 144984 320182 145036
rect 328306 144984 328312 145036
rect 328364 145024 328370 145036
rect 328398 145024 328404 145036
rect 328364 144996 328404 145024
rect 328364 144984 328370 144996
rect 328398 144984 328404 144996
rect 328456 144984 328462 145036
rect 225358 144888 225364 144900
rect 225319 144860 225364 144888
rect 225358 144848 225364 144860
rect 225416 144848 225422 144900
rect 242102 144848 242108 144900
rect 242160 144888 242166 144900
rect 242194 144888 242200 144900
rect 242160 144860 242200 144888
rect 242160 144848 242166 144860
rect 242194 144848 242200 144860
rect 242252 144848 242258 144900
rect 285618 144888 285624 144900
rect 285579 144860 285624 144888
rect 285618 144848 285624 144860
rect 285676 144848 285682 144900
rect 331066 144848 331072 144900
rect 331124 144888 331130 144900
rect 331250 144888 331256 144900
rect 331124 144860 331256 144888
rect 331124 144848 331130 144860
rect 331250 144848 331256 144860
rect 331308 144848 331314 144900
rect 341002 144848 341008 144900
rect 341060 144888 341066 144900
rect 341094 144888 341100 144900
rect 341060 144860 341100 144888
rect 341060 144848 341066 144860
rect 341094 144848 341100 144860
rect 341152 144848 341158 144900
rect 553890 144888 553896 144900
rect 553851 144860 553896 144888
rect 553890 144848 553896 144860
rect 553948 144848 553954 144900
rect 242654 144780 242660 144832
rect 242712 144820 242718 144832
rect 242746 144820 242752 144832
rect 242712 144792 242752 144820
rect 242712 144780 242718 144792
rect 242746 144780 242752 144792
rect 242804 144780 242810 144832
rect 1600 144656 583316 144752
rect 1600 144112 583316 144208
rect 273014 143732 273020 143744
rect 272975 143704 273020 143732
rect 273014 143692 273020 143704
rect 273072 143692 273078 143744
rect 1600 143568 583316 143664
rect 4006 143488 4012 143540
rect 4064 143528 4070 143540
rect 227474 143528 227480 143540
rect 4064 143500 227480 143528
rect 4064 143488 4070 143500
rect 227474 143488 227480 143500
rect 227532 143488 227538 143540
rect 242010 143488 242016 143540
rect 242068 143528 242074 143540
rect 242194 143528 242200 143540
rect 242068 143500 242200 143528
rect 242068 143488 242074 143500
rect 242194 143488 242200 143500
rect 242252 143488 242258 143540
rect 242470 143488 242476 143540
rect 242528 143528 242534 143540
rect 242562 143528 242568 143540
rect 242528 143500 242568 143528
rect 242528 143488 242534 143500
rect 242562 143488 242568 143500
rect 242620 143488 242626 143540
rect 276694 143488 276700 143540
rect 276752 143528 276758 143540
rect 276878 143528 276884 143540
rect 276752 143500 276884 143528
rect 276752 143488 276758 143500
rect 276878 143488 276884 143500
rect 276936 143488 276942 143540
rect 319937 143531 319995 143537
rect 319937 143497 319949 143531
rect 319983 143528 319995 143531
rect 320118 143528 320124 143540
rect 319983 143500 320124 143528
rect 319983 143497 319995 143500
rect 319937 143491 319995 143497
rect 320118 143488 320124 143500
rect 320176 143488 320182 143540
rect 328398 143528 328404 143540
rect 328359 143500 328404 143528
rect 328398 143488 328404 143500
rect 328456 143488 328462 143540
rect 373018 143488 373024 143540
rect 373076 143528 373082 143540
rect 373110 143528 373116 143540
rect 373076 143500 373116 143528
rect 373076 143488 373082 143500
rect 373110 143488 373116 143500
rect 373168 143488 373174 143540
rect 385530 143488 385536 143540
rect 385588 143528 385594 143540
rect 392430 143528 392436 143540
rect 385588 143500 385633 143528
rect 392391 143500 392436 143528
rect 385588 143488 385594 143500
rect 392430 143488 392436 143500
rect 392488 143488 392494 143540
rect 529050 143528 529056 143540
rect 529011 143500 529056 143528
rect 529050 143488 529056 143500
rect 529108 143488 529114 143540
rect 535950 143528 535956 143540
rect 535911 143500 535956 143528
rect 535950 143488 535956 143500
rect 536008 143488 536014 143540
rect 552237 143531 552295 143537
rect 552237 143497 552249 143531
rect 552283 143528 552295 143531
rect 552510 143528 552516 143540
rect 552283 143500 552516 143528
rect 552283 143497 552295 143500
rect 552237 143491 552295 143497
rect 552510 143488 552516 143500
rect 552568 143488 552574 143540
rect 571830 143528 571836 143540
rect 571791 143500 571836 143528
rect 571830 143488 571836 143500
rect 571888 143488 571894 143540
rect 135658 143460 135664 143472
rect 135619 143432 135664 143460
rect 135658 143420 135664 143432
rect 135716 143420 135722 143472
rect 152218 143460 152224 143472
rect 152179 143432 152224 143460
rect 152218 143420 152224 143432
rect 152276 143420 152282 143472
rect 170158 143460 170164 143472
rect 170119 143432 170164 143460
rect 170158 143420 170164 143432
rect 170216 143420 170222 143472
rect 190858 143460 190864 143472
rect 190819 143432 190864 143460
rect 190858 143420 190864 143432
rect 190916 143420 190922 143472
rect 214318 143460 214324 143472
rect 214279 143432 214324 143460
rect 214318 143420 214324 143432
rect 214376 143420 214382 143472
rect 1600 143024 583316 143120
rect 1600 142480 583316 142576
rect 278721 142171 278779 142177
rect 278721 142137 278733 142171
rect 278767 142168 278779 142171
rect 278810 142168 278816 142180
rect 278767 142140 278816 142168
rect 278767 142137 278779 142140
rect 278721 142131 278779 142137
rect 278810 142128 278816 142140
rect 278868 142128 278874 142180
rect 1600 141936 583316 142032
rect 1600 141392 583316 141488
rect 1600 140848 583316 140944
rect 309078 140740 309084 140752
rect 309039 140712 309084 140740
rect 309078 140700 309084 140712
rect 309136 140700 309142 140752
rect 1600 140304 583316 140400
rect 1600 139760 583316 139856
rect 275498 139544 275504 139596
rect 275556 139584 275562 139596
rect 275682 139584 275688 139596
rect 275556 139556 275688 139584
rect 275556 139544 275562 139556
rect 275682 139544 275688 139556
rect 275740 139544 275746 139596
rect 271450 139408 271456 139460
rect 271508 139448 271514 139460
rect 271542 139448 271548 139460
rect 271508 139420 271548 139448
rect 271508 139408 271514 139420
rect 271542 139408 271548 139420
rect 271600 139408 271606 139460
rect 273014 139448 273020 139460
rect 272975 139420 273020 139448
rect 273014 139408 273020 139420
rect 273072 139408 273078 139460
rect 279730 139380 279736 139392
rect 279691 139352 279736 139380
rect 279730 139340 279736 139352
rect 279788 139340 279794 139392
rect 1600 139216 583316 139312
rect 1600 138672 583316 138768
rect 1600 138128 583316 138224
rect 246886 138088 246892 138100
rect 246812 138060 246892 138088
rect 229866 137980 229872 138032
rect 229924 137980 229930 138032
rect 235478 137980 235484 138032
rect 235536 137980 235542 138032
rect 229774 137912 229780 137964
rect 229832 137952 229838 137964
rect 229884 137952 229912 137980
rect 229832 137924 229912 137952
rect 235496 137952 235524 137980
rect 246812 137964 246840 138060
rect 246886 138048 246892 138060
rect 246944 138048 246950 138100
rect 285253 138091 285311 138097
rect 285253 138057 285265 138091
rect 285299 138088 285311 138091
rect 285342 138088 285348 138100
rect 285299 138060 285348 138088
rect 285299 138057 285311 138060
rect 285253 138051 285311 138057
rect 285342 138048 285348 138060
rect 285400 138048 285406 138100
rect 259306 137980 259312 138032
rect 259364 138020 259370 138032
rect 268782 138020 268788 138032
rect 259364 137992 259444 138020
rect 259364 137980 259370 137992
rect 235570 137952 235576 137964
rect 235496 137924 235576 137952
rect 229832 137912 229838 137924
rect 235570 137912 235576 137924
rect 235628 137912 235634 137964
rect 246794 137912 246800 137964
rect 246852 137912 246858 137964
rect 259416 137828 259444 137992
rect 268708 137992 268788 138020
rect 268708 137964 268736 137992
rect 268782 137980 268788 137992
rect 268840 137980 268846 138032
rect 305030 137980 305036 138032
rect 305088 137980 305094 138032
rect 371822 137980 371828 138032
rect 371880 137980 371886 138032
rect 268690 137912 268696 137964
rect 268748 137912 268754 137964
rect 271450 137952 271456 137964
rect 271411 137924 271456 137952
rect 271450 137912 271456 137924
rect 271508 137912 271514 137964
rect 285618 137952 285624 137964
rect 285579 137924 285624 137952
rect 285618 137912 285624 137924
rect 285676 137912 285682 137964
rect 305048 137952 305076 137980
rect 305122 137952 305128 137964
rect 305048 137924 305128 137952
rect 305122 137912 305128 137924
rect 305180 137912 305186 137964
rect 371840 137952 371868 137980
rect 371914 137952 371920 137964
rect 371840 137924 371920 137952
rect 371914 137912 371920 137924
rect 371972 137912 371978 137964
rect 285069 137887 285127 137893
rect 285069 137853 285081 137887
rect 285115 137884 285127 137887
rect 285158 137884 285164 137896
rect 285115 137856 285164 137884
rect 285115 137853 285127 137856
rect 285069 137847 285127 137853
rect 285158 137844 285164 137856
rect 285216 137844 285222 137896
rect 259398 137776 259404 137828
rect 259456 137776 259462 137828
rect 1600 137584 583316 137680
rect 1600 137040 583316 137136
rect 1600 136496 583316 136592
rect 1600 135952 583316 136048
rect 285434 135572 285440 135584
rect 285395 135544 285440 135572
rect 285434 135532 285440 135544
rect 285492 135532 285498 135584
rect 1600 135408 583316 135504
rect 225358 135368 225364 135380
rect 225319 135340 225364 135368
rect 225358 135328 225364 135340
rect 225416 135328 225422 135380
rect 553890 135368 553896 135380
rect 553851 135340 553896 135368
rect 553890 135328 553896 135340
rect 553948 135328 553954 135380
rect 246518 135260 246524 135312
rect 246576 135260 246582 135312
rect 285437 135303 285495 135309
rect 285437 135269 285449 135303
rect 285483 135300 285495 135303
rect 285526 135300 285532 135312
rect 285483 135272 285532 135300
rect 285483 135269 285495 135272
rect 285437 135263 285495 135269
rect 285526 135260 285532 135272
rect 285584 135260 285590 135312
rect 91314 135192 91320 135244
rect 91372 135232 91378 135244
rect 91498 135232 91504 135244
rect 91372 135204 91504 135232
rect 91372 135192 91378 135204
rect 91498 135192 91504 135204
rect 91556 135192 91562 135244
rect 235570 135192 235576 135244
rect 235628 135232 235634 135244
rect 235754 135232 235760 135244
rect 235628 135204 235760 135232
rect 235628 135192 235634 135204
rect 235754 135192 235760 135204
rect 235812 135192 235818 135244
rect 246536 135176 246564 135260
rect 259398 135232 259404 135244
rect 259359 135204 259404 135232
rect 259398 135192 259404 135204
rect 259456 135192 259462 135244
rect 268690 135232 268696 135244
rect 268651 135204 268696 135232
rect 268690 135192 268696 135204
rect 268748 135192 268754 135244
rect 341186 135192 341192 135244
rect 341244 135232 341250 135244
rect 341370 135232 341376 135244
rect 341244 135204 341376 135232
rect 341244 135192 341250 135204
rect 341370 135192 341376 135204
rect 341428 135192 341434 135244
rect 371914 135232 371920 135244
rect 371875 135204 371920 135232
rect 371914 135192 371920 135204
rect 371972 135192 371978 135244
rect 553706 135192 553712 135244
rect 553764 135232 553770 135244
rect 553890 135232 553896 135244
rect 553764 135204 553896 135232
rect 553764 135192 553770 135204
rect 553890 135192 553896 135204
rect 553948 135192 553954 135244
rect 246518 135124 246524 135176
rect 246576 135124 246582 135176
rect 1600 134864 583316 134960
rect 309078 134688 309084 134700
rect 309039 134660 309084 134688
rect 309078 134648 309084 134660
rect 309136 134648 309142 134700
rect 1600 134320 583316 134416
rect 135658 133940 135664 133952
rect 135619 133912 135664 133940
rect 135658 133900 135664 133912
rect 135716 133900 135722 133952
rect 152218 133940 152224 133952
rect 152179 133912 152224 133940
rect 152218 133900 152224 133912
rect 152276 133900 152282 133952
rect 170158 133940 170164 133952
rect 170119 133912 170164 133940
rect 170158 133900 170164 133912
rect 170216 133900 170222 133952
rect 190858 133940 190864 133952
rect 190819 133912 190864 133940
rect 190858 133900 190864 133912
rect 190916 133900 190922 133952
rect 214318 133940 214324 133952
rect 214279 133912 214324 133940
rect 214318 133900 214324 133912
rect 214376 133900 214382 133952
rect 319934 133940 319940 133952
rect 319895 133912 319940 133940
rect 319934 133900 319940 133912
rect 319992 133900 319998 133952
rect 328398 133940 328404 133952
rect 328359 133912 328404 133940
rect 328398 133900 328404 133912
rect 328456 133900 328462 133952
rect 385530 133900 385536 133952
rect 385588 133940 385594 133952
rect 392430 133940 392436 133952
rect 385588 133912 385633 133940
rect 392391 133912 392436 133940
rect 385588 133900 385594 133912
rect 392430 133900 392436 133912
rect 392488 133900 392494 133952
rect 529050 133940 529056 133952
rect 529011 133912 529056 133940
rect 529050 133900 529056 133912
rect 529108 133900 529114 133952
rect 535950 133940 535956 133952
rect 535911 133912 535956 133940
rect 535950 133900 535956 133912
rect 536008 133900 536014 133952
rect 552234 133940 552240 133952
rect 552195 133912 552240 133940
rect 552234 133900 552240 133912
rect 552292 133900 552298 133952
rect 571830 133940 571836 133952
rect 571791 133912 571836 133940
rect 571830 133900 571836 133912
rect 571888 133900 571894 133952
rect 1600 133776 583316 133872
rect 552234 133736 552240 133748
rect 552195 133708 552240 133736
rect 552234 133696 552240 133708
rect 552292 133696 552298 133748
rect 1600 133232 583316 133328
rect 290310 132812 290316 132864
rect 290368 132852 290374 132864
rect 293254 132852 293260 132864
rect 290368 132824 293260 132852
rect 290368 132812 290374 132824
rect 293254 132812 293260 132824
rect 293312 132812 293318 132864
rect 399238 132812 399244 132864
rect 399296 132852 399302 132864
rect 406138 132852 406144 132864
rect 399296 132824 406144 132852
rect 399296 132812 399302 132824
rect 406138 132812 406144 132824
rect 406196 132812 406202 132864
rect 1600 132688 583316 132784
rect 375870 132540 375876 132592
rect 375928 132580 375934 132592
rect 385438 132580 385444 132592
rect 375928 132552 385444 132580
rect 375928 132540 375934 132552
rect 385438 132540 385444 132552
rect 385496 132540 385502 132592
rect 1600 132144 583316 132240
rect 1600 131600 583316 131696
rect 1600 131056 583316 131152
rect 1600 130512 583316 130608
rect 1600 129968 583316 130064
rect 275498 129820 275504 129872
rect 275556 129860 275562 129872
rect 275682 129860 275688 129872
rect 275556 129832 275688 129860
rect 275556 129820 275562 129832
rect 275682 129820 275688 129832
rect 275740 129820 275746 129872
rect 279733 129795 279791 129801
rect 279733 129761 279745 129795
rect 279779 129792 279791 129795
rect 279822 129792 279828 129804
rect 279779 129764 279828 129792
rect 279779 129761 279791 129764
rect 279733 129755 279791 129761
rect 279822 129752 279828 129764
rect 279880 129752 279886 129804
rect 275590 129684 275596 129736
rect 275648 129724 275654 129736
rect 275682 129724 275688 129736
rect 275648 129696 275688 129724
rect 275648 129684 275654 129696
rect 275682 129684 275688 129696
rect 275740 129684 275746 129736
rect 1600 129424 583316 129520
rect 1600 128880 583316 128976
rect 239250 128460 239256 128512
rect 239308 128500 239314 128512
rect 239434 128500 239440 128512
rect 239308 128472 239440 128500
rect 239308 128460 239314 128472
rect 239434 128460 239440 128472
rect 239492 128460 239498 128512
rect 271450 128500 271456 128512
rect 271411 128472 271456 128500
rect 271450 128460 271456 128472
rect 271508 128460 271514 128512
rect 1600 128336 583316 128432
rect 239250 128256 239256 128308
rect 239308 128296 239314 128308
rect 239434 128296 239440 128308
rect 239308 128268 239440 128296
rect 239308 128256 239314 128268
rect 239434 128256 239440 128268
rect 239492 128256 239498 128308
rect 259398 128296 259404 128308
rect 259359 128268 259404 128296
rect 259398 128256 259404 128268
rect 259456 128256 259462 128308
rect 268690 128296 268696 128308
rect 268651 128268 268696 128296
rect 268690 128256 268696 128268
rect 268748 128256 268754 128308
rect 371914 128296 371920 128308
rect 371875 128268 371920 128296
rect 371914 128256 371920 128268
rect 371972 128256 371978 128308
rect 1600 127792 583316 127888
rect 1600 127248 583316 127344
rect 1600 126704 583316 126800
rect 1600 126160 583316 126256
rect 1600 125616 583316 125712
rect 242838 125576 242844 125588
rect 242799 125548 242844 125576
rect 242838 125536 242844 125548
rect 242896 125536 242902 125588
rect 246518 125536 246524 125588
rect 246576 125536 246582 125588
rect 305122 125576 305128 125588
rect 305083 125548 305128 125576
rect 305122 125536 305128 125548
rect 305180 125536 305186 125588
rect 308986 125576 308992 125588
rect 308947 125548 308992 125576
rect 308986 125536 308992 125548
rect 309044 125536 309050 125588
rect 331066 125536 331072 125588
rect 331124 125576 331130 125588
rect 331250 125576 331256 125588
rect 331124 125548 331256 125576
rect 331124 125536 331130 125548
rect 331250 125536 331256 125548
rect 331308 125536 331314 125588
rect 341094 125576 341100 125588
rect 341055 125548 341100 125576
rect 341094 125536 341100 125548
rect 341152 125536 341158 125588
rect 246536 125508 246564 125536
rect 246610 125508 246616 125520
rect 246536 125480 246616 125508
rect 246610 125468 246616 125480
rect 246668 125468 246674 125520
rect 552237 125443 552295 125449
rect 552237 125409 552249 125443
rect 552283 125440 552295 125443
rect 552510 125440 552516 125452
rect 552283 125412 552516 125440
rect 552283 125409 552295 125412
rect 552237 125403 552295 125409
rect 552510 125400 552516 125412
rect 552568 125400 552574 125452
rect 1600 125072 583316 125168
rect 1600 124528 583316 124624
rect 135658 124148 135664 124160
rect 135619 124120 135664 124148
rect 135658 124108 135664 124120
rect 135716 124108 135722 124160
rect 152218 124148 152224 124160
rect 152179 124120 152224 124148
rect 152218 124108 152224 124120
rect 152276 124108 152282 124160
rect 170158 124148 170164 124160
rect 170119 124120 170164 124148
rect 170158 124108 170164 124120
rect 170216 124108 170222 124160
rect 190858 124148 190864 124160
rect 190819 124120 190864 124148
rect 190858 124108 190864 124120
rect 190916 124108 190922 124160
rect 214318 124148 214324 124160
rect 214279 124120 214324 124148
rect 214318 124108 214324 124120
rect 214376 124108 214382 124160
rect 373110 124148 373116 124160
rect 373071 124120 373116 124148
rect 373110 124108 373116 124120
rect 373168 124108 373174 124160
rect 385530 124108 385536 124160
rect 385588 124148 385594 124160
rect 392430 124148 392436 124160
rect 385588 124120 385633 124148
rect 392391 124120 392436 124148
rect 385588 124108 385594 124120
rect 392430 124108 392436 124120
rect 392488 124108 392494 124160
rect 529050 124148 529056 124160
rect 529011 124120 529056 124148
rect 529050 124108 529056 124120
rect 529108 124108 529114 124160
rect 535950 124148 535956 124160
rect 535911 124120 535956 124148
rect 535950 124108 535956 124120
rect 536008 124108 536014 124160
rect 571830 124148 571836 124160
rect 571791 124120 571836 124148
rect 571830 124108 571836 124120
rect 571888 124108 571894 124160
rect 1600 123984 583316 124080
rect 1600 123440 583316 123536
rect 1600 122896 583316 122992
rect 553430 122748 553436 122800
rect 553488 122788 553494 122800
rect 553890 122788 553896 122800
rect 553488 122760 553896 122788
rect 553488 122748 553494 122760
rect 553890 122748 553896 122760
rect 553948 122748 553954 122800
rect 1600 122352 583316 122448
rect 1600 121808 583316 121904
rect 272830 121428 272836 121440
rect 272791 121400 272836 121428
rect 272830 121388 272836 121400
rect 272888 121388 272894 121440
rect 273014 121388 273020 121440
rect 273072 121428 273078 121440
rect 273106 121428 273112 121440
rect 273072 121400 273112 121428
rect 273072 121388 273078 121400
rect 273106 121388 273112 121400
rect 273164 121388 273170 121440
rect 279730 121388 279736 121440
rect 279788 121428 279794 121440
rect 279822 121428 279828 121440
rect 279788 121400 279828 121428
rect 279788 121388 279794 121400
rect 279822 121388 279828 121400
rect 279880 121388 279886 121440
rect 1600 121264 583316 121360
rect 1600 120720 583316 120816
rect 1600 120176 583316 120272
rect 285618 120068 285624 120080
rect 285579 120040 285624 120068
rect 285618 120028 285624 120040
rect 285676 120028 285682 120080
rect 1600 119632 583316 119728
rect 242562 119348 242568 119400
rect 242620 119388 242626 119400
rect 242930 119388 242936 119400
rect 242620 119360 242936 119388
rect 242620 119348 242626 119360
rect 242930 119348 242936 119360
rect 242988 119348 242994 119400
rect 308989 119391 309047 119397
rect 308989 119357 309001 119391
rect 309035 119388 309047 119391
rect 309170 119388 309176 119400
rect 309035 119360 309176 119388
rect 309035 119357 309047 119360
rect 308989 119351 309047 119357
rect 309170 119348 309176 119360
rect 309228 119348 309234 119400
rect 1600 119088 583316 119184
rect 229777 118779 229835 118785
rect 229777 118745 229789 118779
rect 229823 118776 229835 118779
rect 229866 118776 229872 118788
rect 229823 118748 229872 118776
rect 229823 118745 229835 118748
rect 229777 118739 229835 118745
rect 229866 118736 229872 118748
rect 229924 118736 229930 118788
rect 1600 118544 583316 118640
rect 305122 118504 305128 118516
rect 305083 118476 305128 118504
rect 305122 118464 305128 118476
rect 305180 118464 305186 118516
rect 1600 118000 583316 118096
rect 1600 117456 583316 117552
rect 1600 116912 583316 117008
rect 242838 116736 242844 116748
rect 242799 116708 242844 116736
rect 242838 116696 242844 116708
rect 242896 116696 242902 116748
rect 1600 116368 583316 116464
rect 341097 116059 341155 116065
rect 341097 116025 341109 116059
rect 341143 116056 341155 116059
rect 341186 116056 341192 116068
rect 341143 116028 341192 116056
rect 341143 116025 341155 116028
rect 341097 116019 341155 116025
rect 341186 116016 341192 116028
rect 341244 116016 341250 116068
rect 259306 115948 259312 116000
rect 259364 115988 259370 116000
rect 259490 115988 259496 116000
rect 259364 115960 259496 115988
rect 259364 115948 259370 115960
rect 259490 115948 259496 115960
rect 259548 115948 259554 116000
rect 1600 115824 583316 115920
rect 91498 115784 91504 115796
rect 91459 115756 91504 115784
rect 91498 115744 91504 115756
rect 91556 115744 91562 115796
rect 235570 115784 235576 115796
rect 235531 115756 235576 115784
rect 235570 115744 235576 115756
rect 235628 115744 235634 115796
rect 357930 115744 357936 115796
rect 357988 115784 357994 115796
rect 357988 115756 358033 115784
rect 357988 115744 357994 115756
rect 1600 115280 583316 115376
rect 1600 114736 583316 114832
rect 229774 114696 229780 114708
rect 229735 114668 229780 114696
rect 229774 114656 229780 114668
rect 229832 114656 229838 114708
rect 135658 114560 135664 114572
rect 135619 114532 135664 114560
rect 135658 114520 135664 114532
rect 135716 114520 135722 114572
rect 152218 114560 152224 114572
rect 152179 114532 152224 114560
rect 152218 114520 152224 114532
rect 152276 114520 152282 114572
rect 170158 114560 170164 114572
rect 170119 114532 170164 114560
rect 170158 114520 170164 114532
rect 170216 114520 170222 114572
rect 190858 114560 190864 114572
rect 190819 114532 190864 114560
rect 190858 114520 190864 114532
rect 190916 114520 190922 114572
rect 214318 114560 214324 114572
rect 214279 114532 214324 114560
rect 214318 114520 214324 114532
rect 214376 114520 214382 114572
rect 319934 114520 319940 114572
rect 319992 114560 319998 114572
rect 320118 114560 320124 114572
rect 319992 114532 320124 114560
rect 319992 114520 319998 114532
rect 320118 114520 320124 114532
rect 320176 114520 320182 114572
rect 373110 114560 373116 114572
rect 373071 114532 373116 114560
rect 373110 114520 373116 114532
rect 373168 114520 373174 114572
rect 385530 114520 385536 114572
rect 385588 114560 385594 114572
rect 392430 114560 392436 114572
rect 385588 114532 385633 114560
rect 392391 114532 392436 114560
rect 385588 114520 385594 114532
rect 392430 114520 392436 114532
rect 392488 114520 392494 114572
rect 529050 114560 529056 114572
rect 529011 114532 529056 114560
rect 529050 114520 529056 114532
rect 529108 114520 529114 114572
rect 535950 114560 535956 114572
rect 535911 114532 535956 114560
rect 535950 114520 535956 114532
rect 536008 114520 536014 114572
rect 571830 114560 571836 114572
rect 571791 114532 571836 114560
rect 571830 114520 571836 114532
rect 571888 114520 571894 114572
rect 242838 114492 242844 114504
rect 242799 114464 242844 114492
rect 242838 114452 242844 114464
rect 242896 114452 242902 114504
rect 552510 114452 552516 114504
rect 552568 114492 552574 114504
rect 552602 114492 552608 114504
rect 552568 114464 552608 114492
rect 552568 114452 552574 114464
rect 552602 114452 552608 114464
rect 552660 114452 552666 114504
rect 1600 114192 583316 114288
rect 1600 113648 583316 113744
rect 1600 113104 583316 113200
rect 1600 112560 583316 112656
rect 1600 112016 583316 112112
rect 272830 111840 272836 111852
rect 272791 111812 272836 111840
rect 272830 111800 272836 111812
rect 272888 111800 272894 111852
rect 285250 111800 285256 111852
rect 285308 111840 285314 111852
rect 285342 111840 285348 111852
rect 285308 111812 285348 111840
rect 285308 111800 285314 111812
rect 285342 111800 285348 111812
rect 285400 111800 285406 111852
rect 1600 111472 583316 111568
rect 285618 111296 285624 111308
rect 285579 111268 285624 111296
rect 285618 111256 285624 111268
rect 285676 111256 285682 111308
rect 242657 111163 242715 111169
rect 242657 111129 242669 111163
rect 242703 111160 242715 111163
rect 242930 111160 242936 111172
rect 242703 111132 242936 111160
rect 242703 111129 242715 111132
rect 242657 111123 242715 111129
rect 242930 111120 242936 111132
rect 242988 111120 242994 111172
rect 1600 110928 583316 111024
rect 242841 110551 242899 110557
rect 242841 110517 242853 110551
rect 242887 110548 242899 110551
rect 242930 110548 242936 110560
rect 242887 110520 242936 110548
rect 242887 110517 242899 110520
rect 242841 110511 242899 110517
rect 242930 110508 242936 110520
rect 242988 110508 242994 110560
rect 1600 110384 583316 110480
rect 1600 109840 583316 109936
rect 553614 109692 553620 109744
rect 553672 109732 553678 109744
rect 553893 109735 553951 109741
rect 553893 109732 553905 109735
rect 553672 109704 553905 109732
rect 553672 109692 553678 109704
rect 553893 109701 553905 109704
rect 553939 109701 553951 109735
rect 553893 109695 553951 109701
rect 1600 109296 583316 109392
rect 229774 109012 229780 109064
rect 229832 109012 229838 109064
rect 275498 109012 275504 109064
rect 275556 109052 275562 109064
rect 275590 109052 275596 109064
rect 275556 109024 275596 109052
rect 275556 109012 275562 109024
rect 275590 109012 275596 109024
rect 275648 109012 275654 109064
rect 305030 109012 305036 109064
rect 305088 109052 305094 109064
rect 305214 109052 305220 109064
rect 305088 109024 305220 109052
rect 305088 109012 305094 109024
rect 305214 109012 305220 109024
rect 305272 109012 305278 109064
rect 320118 109052 320124 109064
rect 320079 109024 320124 109052
rect 320118 109012 320124 109024
rect 320176 109012 320182 109064
rect 328398 109052 328404 109064
rect 328359 109024 328404 109052
rect 328398 109012 328404 109024
rect 328456 109012 328462 109064
rect 229792 108984 229820 109012
rect 229866 108984 229872 108996
rect 229792 108956 229872 108984
rect 229866 108944 229872 108956
rect 229924 108944 229930 108996
rect 235570 108984 235576 108996
rect 235531 108956 235576 108984
rect 235570 108944 235576 108956
rect 235628 108944 235634 108996
rect 1600 108752 583316 108848
rect 1600 108208 583316 108304
rect 1600 107664 583316 107760
rect 1600 107120 583316 107216
rect 1600 106576 583316 106672
rect 91498 106332 91504 106344
rect 91459 106304 91504 106332
rect 91498 106292 91504 106304
rect 91556 106292 91562 106344
rect 275501 106335 275559 106341
rect 275501 106301 275513 106335
rect 275547 106332 275559 106335
rect 275590 106332 275596 106344
rect 275547 106304 275596 106332
rect 275547 106301 275559 106304
rect 275501 106295 275559 106301
rect 275590 106292 275596 106304
rect 275648 106292 275654 106344
rect 309170 106332 309176 106344
rect 309096 106304 309176 106332
rect 309096 106276 309124 106304
rect 309170 106292 309176 106304
rect 309228 106292 309234 106344
rect 357930 106292 357936 106344
rect 357988 106332 357994 106344
rect 357988 106304 358033 106332
rect 357988 106292 357994 106304
rect 235478 106264 235484 106276
rect 235439 106236 235484 106264
rect 235478 106224 235484 106236
rect 235536 106224 235542 106276
rect 239250 106224 239256 106276
rect 239308 106264 239314 106276
rect 239434 106264 239440 106276
rect 239308 106236 239440 106264
rect 239308 106224 239314 106236
rect 239434 106224 239440 106236
rect 239492 106224 239498 106276
rect 309078 106224 309084 106276
rect 309136 106224 309142 106276
rect 331066 106224 331072 106276
rect 331124 106264 331130 106276
rect 331250 106264 331256 106276
rect 331124 106236 331256 106264
rect 331124 106224 331130 106236
rect 331250 106224 331256 106236
rect 331308 106224 331314 106276
rect 341002 106224 341008 106276
rect 341060 106264 341066 106276
rect 341094 106264 341100 106276
rect 341060 106236 341100 106264
rect 341060 106224 341066 106236
rect 341094 106224 341100 106236
rect 341152 106224 341158 106276
rect 1600 106032 583316 106128
rect 1600 105488 583316 105584
rect 1600 104944 583316 105040
rect 242654 104904 242660 104916
rect 242615 104876 242660 104904
rect 242654 104864 242660 104876
rect 242712 104864 242718 104916
rect 320118 104904 320124 104916
rect 320079 104876 320124 104904
rect 320118 104864 320124 104876
rect 320176 104864 320182 104916
rect 328398 104904 328404 104916
rect 328359 104876 328404 104904
rect 328398 104864 328404 104876
rect 328456 104864 328462 104916
rect 371822 104864 371828 104916
rect 371880 104904 371886 104916
rect 371914 104904 371920 104916
rect 371880 104876 371920 104904
rect 371880 104864 371886 104876
rect 371914 104864 371920 104876
rect 371972 104864 371978 104916
rect 135658 104836 135664 104848
rect 135619 104808 135664 104836
rect 135658 104796 135664 104808
rect 135716 104796 135722 104848
rect 152218 104836 152224 104848
rect 152179 104808 152224 104836
rect 152218 104796 152224 104808
rect 152276 104796 152282 104848
rect 170158 104836 170164 104848
rect 170119 104808 170164 104836
rect 170158 104796 170164 104808
rect 170216 104796 170222 104848
rect 190858 104836 190864 104848
rect 190819 104808 190864 104836
rect 190858 104796 190864 104808
rect 190916 104796 190922 104848
rect 214318 104836 214324 104848
rect 214279 104808 214324 104836
rect 214318 104796 214324 104808
rect 214376 104796 214382 104848
rect 305030 104836 305036 104848
rect 304991 104808 305036 104836
rect 305030 104796 305036 104808
rect 305088 104796 305094 104848
rect 373110 104836 373116 104848
rect 373071 104808 373116 104836
rect 373110 104796 373116 104808
rect 373168 104796 373174 104848
rect 385530 104796 385536 104848
rect 385588 104836 385594 104848
rect 392430 104836 392436 104848
rect 385588 104808 385633 104836
rect 392391 104808 392436 104836
rect 385588 104796 385594 104808
rect 392430 104796 392436 104808
rect 392488 104796 392494 104848
rect 529050 104836 529056 104848
rect 529011 104808 529056 104836
rect 529050 104796 529056 104808
rect 529108 104796 529114 104848
rect 535950 104836 535956 104848
rect 535911 104808 535956 104836
rect 535950 104796 535956 104808
rect 536008 104796 536014 104848
rect 571830 104836 571836 104848
rect 571791 104808 571836 104836
rect 571830 104796 571836 104808
rect 571888 104796 571894 104848
rect 1600 104400 583316 104496
rect 1600 103856 583316 103952
rect 229777 103479 229835 103485
rect 229777 103445 229789 103479
rect 229823 103476 229835 103479
rect 229866 103476 229872 103488
rect 229823 103448 229872 103476
rect 229823 103445 229835 103448
rect 229777 103439 229835 103445
rect 229866 103436 229872 103448
rect 229924 103436 229930 103488
rect 308897 103479 308955 103485
rect 308897 103445 308909 103479
rect 308943 103476 308955 103479
rect 309078 103476 309084 103488
rect 308943 103448 309084 103476
rect 308943 103445 308955 103448
rect 308897 103439 308955 103445
rect 309078 103436 309084 103448
rect 309136 103436 309142 103488
rect 319937 103479 319995 103485
rect 319937 103445 319949 103479
rect 319983 103476 319995 103479
rect 320118 103476 320124 103488
rect 319983 103448 320124 103476
rect 319983 103445 319995 103448
rect 319937 103439 319995 103445
rect 320118 103436 320124 103448
rect 320176 103436 320182 103488
rect 552418 103436 552424 103488
rect 552476 103476 552482 103488
rect 552513 103479 552571 103485
rect 552513 103476 552525 103479
rect 552476 103448 552525 103476
rect 552476 103436 552482 103448
rect 552513 103445 552525 103448
rect 552559 103445 552571 103479
rect 552513 103439 552571 103445
rect 1600 103312 583316 103408
rect 1600 102768 583316 102864
rect 285253 102391 285311 102397
rect 285253 102357 285265 102391
rect 285299 102388 285311 102391
rect 285342 102388 285348 102400
rect 285299 102360 285348 102388
rect 285299 102357 285311 102360
rect 285253 102351 285311 102357
rect 285342 102348 285348 102360
rect 285400 102348 285406 102400
rect 1600 102224 583316 102320
rect 285250 102184 285256 102196
rect 285211 102156 285256 102184
rect 285250 102144 285256 102156
rect 285308 102144 285314 102196
rect 1600 101680 583316 101776
rect 242013 101439 242071 101445
rect 242013 101405 242025 101439
rect 242059 101436 242071 101439
rect 242102 101436 242108 101448
rect 242059 101408 242108 101436
rect 242059 101405 242071 101408
rect 242013 101399 242071 101405
rect 242102 101396 242108 101408
rect 242160 101396 242166 101448
rect 1600 101136 583316 101232
rect 360414 100920 360420 100972
rect 360472 100960 360478 100972
rect 366118 100960 366124 100972
rect 360472 100932 366124 100960
rect 360472 100920 360478 100932
rect 366118 100920 366124 100932
rect 366176 100920 366182 100972
rect 251670 100852 251676 100904
rect 251728 100892 251734 100904
rect 261146 100892 261152 100904
rect 251728 100864 261152 100892
rect 251728 100852 251734 100864
rect 261146 100852 261152 100864
rect 261204 100852 261210 100904
rect 275498 100756 275504 100768
rect 275459 100728 275504 100756
rect 275498 100716 275504 100728
rect 275556 100716 275562 100768
rect 279730 100716 279736 100768
rect 279788 100756 279794 100768
rect 280006 100756 280012 100768
rect 279788 100728 280012 100756
rect 279788 100716 279794 100728
rect 280006 100716 280012 100728
rect 280064 100716 280070 100768
rect 1600 100592 583316 100688
rect 1600 100048 583316 100144
rect 1600 99504 583316 99600
rect 246610 99424 246616 99476
rect 246668 99424 246674 99476
rect 246628 99340 246656 99424
rect 268690 99356 268696 99408
rect 268748 99356 268754 99408
rect 271450 99356 271456 99408
rect 271508 99396 271514 99408
rect 271634 99396 271640 99408
rect 271508 99368 271640 99396
rect 271508 99356 271514 99368
rect 271634 99356 271640 99368
rect 271692 99356 271698 99408
rect 246610 99288 246616 99340
rect 246668 99288 246674 99340
rect 268708 99272 268736 99356
rect 305033 99331 305091 99337
rect 305033 99297 305045 99331
rect 305079 99328 305091 99331
rect 305122 99328 305128 99340
rect 305079 99300 305128 99328
rect 305079 99297 305091 99300
rect 305033 99291 305091 99297
rect 305122 99288 305128 99300
rect 305180 99288 305186 99340
rect 268690 99220 268696 99272
rect 268748 99220 268754 99272
rect 1600 98960 583316 99056
rect 1600 98416 583316 98512
rect 1600 97872 583316 97968
rect 1600 97328 583316 97424
rect 1600 96784 583316 96880
rect 553890 96744 553896 96756
rect 553851 96716 553896 96744
rect 553890 96704 553896 96716
rect 553948 96704 553954 96756
rect 235478 96676 235484 96688
rect 235439 96648 235484 96676
rect 235478 96636 235484 96648
rect 235536 96636 235542 96688
rect 91314 96568 91320 96620
rect 91372 96608 91378 96620
rect 91498 96608 91504 96620
rect 91372 96580 91504 96608
rect 91372 96568 91378 96580
rect 91498 96568 91504 96580
rect 91556 96568 91562 96620
rect 235570 96608 235576 96620
rect 235531 96580 235576 96608
rect 235570 96568 235576 96580
rect 235628 96568 235634 96620
rect 268690 96608 268696 96620
rect 268651 96580 268696 96608
rect 268690 96568 268696 96580
rect 268748 96568 268754 96620
rect 307882 96568 307888 96620
rect 307940 96608 307946 96620
rect 308250 96608 308256 96620
rect 307940 96580 308256 96608
rect 307940 96568 307946 96580
rect 308250 96568 308256 96580
rect 308308 96568 308314 96620
rect 341186 96568 341192 96620
rect 341244 96608 341250 96620
rect 341370 96608 341376 96620
rect 341244 96580 341376 96608
rect 341244 96568 341250 96580
rect 341370 96568 341376 96580
rect 341428 96568 341434 96620
rect 357930 96568 357936 96620
rect 357988 96608 357994 96620
rect 358206 96608 358212 96620
rect 357988 96580 358212 96608
rect 357988 96568 357994 96580
rect 358206 96568 358212 96580
rect 358264 96568 358270 96620
rect 553706 96568 553712 96620
rect 553764 96608 553770 96620
rect 553890 96608 553896 96620
rect 553764 96580 553896 96608
rect 553764 96568 553770 96580
rect 553890 96568 553896 96580
rect 553948 96568 553954 96620
rect 1600 96240 583316 96336
rect 1600 95696 583316 95792
rect 135658 95316 135664 95328
rect 135619 95288 135664 95316
rect 135658 95276 135664 95288
rect 135716 95276 135722 95328
rect 152218 95316 152224 95328
rect 152179 95288 152224 95316
rect 152218 95276 152224 95288
rect 152276 95276 152282 95328
rect 170158 95316 170164 95328
rect 170119 95288 170164 95316
rect 170158 95276 170164 95288
rect 170216 95276 170222 95328
rect 190858 95316 190864 95328
rect 190819 95288 190864 95316
rect 190858 95276 190864 95288
rect 190916 95276 190922 95328
rect 214318 95316 214324 95328
rect 214279 95288 214324 95316
rect 214318 95276 214324 95288
rect 214376 95276 214382 95328
rect 371914 95276 371920 95328
rect 371972 95316 371978 95328
rect 372006 95316 372012 95328
rect 371972 95288 372012 95316
rect 371972 95276 371978 95288
rect 372006 95276 372012 95288
rect 372064 95276 372070 95328
rect 373110 95316 373116 95328
rect 373071 95288 373116 95316
rect 373110 95276 373116 95288
rect 373168 95276 373174 95328
rect 385530 95276 385536 95328
rect 385588 95316 385594 95328
rect 392430 95316 392436 95328
rect 385588 95288 385633 95316
rect 392391 95288 392436 95316
rect 385588 95276 385594 95288
rect 392430 95276 392436 95288
rect 392488 95276 392494 95328
rect 529050 95316 529056 95328
rect 529011 95288 529056 95316
rect 529050 95276 529056 95288
rect 529108 95276 529114 95328
rect 535950 95316 535956 95328
rect 535911 95288 535956 95316
rect 535950 95276 535956 95288
rect 536008 95276 536014 95328
rect 571830 95316 571836 95328
rect 571791 95288 571836 95316
rect 571830 95276 571836 95288
rect 571888 95276 571894 95328
rect 1600 95152 583316 95248
rect 328582 95072 328588 95124
rect 328640 95072 328646 95124
rect 371914 95112 371920 95124
rect 371875 95084 371920 95112
rect 371914 95072 371920 95084
rect 371972 95072 371978 95124
rect 328600 94988 328628 95072
rect 328582 94936 328588 94988
rect 328640 94936 328646 94988
rect 1600 94608 583316 94704
rect 1600 94064 583316 94160
rect 278810 93956 278816 93968
rect 278736 93928 278816 93956
rect 278736 93900 278764 93928
rect 278810 93916 278816 93928
rect 278868 93916 278874 93968
rect 242010 93888 242016 93900
rect 241971 93860 242016 93888
rect 242010 93848 242016 93860
rect 242068 93848 242074 93900
rect 276510 93848 276516 93900
rect 276568 93888 276574 93900
rect 276568 93860 276648 93888
rect 276568 93848 276574 93860
rect 276620 93832 276648 93860
rect 278718 93848 278724 93900
rect 278776 93848 278782 93900
rect 285250 93848 285256 93900
rect 285308 93888 285314 93900
rect 285342 93888 285348 93900
rect 285308 93860 285348 93888
rect 285308 93848 285314 93860
rect 285342 93848 285348 93860
rect 285400 93848 285406 93900
rect 308894 93888 308900 93900
rect 308855 93860 308900 93888
rect 308894 93848 308900 93860
rect 308952 93848 308958 93900
rect 319934 93888 319940 93900
rect 319895 93860 319940 93888
rect 319934 93848 319940 93860
rect 319992 93848 319998 93900
rect 552418 93848 552424 93900
rect 552476 93888 552482 93900
rect 552513 93891 552571 93897
rect 552513 93888 552525 93891
rect 552476 93860 552525 93888
rect 552476 93848 552482 93860
rect 552513 93857 552525 93860
rect 552559 93857 552571 93891
rect 552513 93851 552571 93857
rect 276602 93780 276608 93832
rect 276660 93780 276666 93832
rect 1600 93520 583316 93616
rect 1600 92976 583316 93072
rect 1600 92432 583316 92528
rect 1600 91888 583316 91984
rect 1600 91344 583316 91440
rect 275498 91060 275504 91112
rect 275556 91100 275562 91112
rect 275682 91100 275688 91112
rect 275556 91072 275688 91100
rect 275556 91060 275562 91072
rect 275682 91060 275688 91072
rect 275740 91060 275746 91112
rect 279822 91060 279828 91112
rect 279880 91100 279886 91112
rect 280006 91100 280012 91112
rect 279880 91072 280012 91100
rect 279880 91060 279886 91072
rect 280006 91060 280012 91072
rect 280064 91060 280070 91112
rect 1600 90800 583316 90896
rect 1600 90256 583316 90352
rect 246521 90083 246579 90089
rect 246521 90049 246533 90083
rect 246567 90080 246579 90083
rect 246610 90080 246616 90092
rect 246567 90052 246616 90080
rect 246567 90049 246579 90052
rect 246521 90043 246579 90049
rect 246610 90040 246616 90052
rect 246668 90040 246674 90092
rect 1600 89712 583316 89808
rect 235570 89672 235576 89684
rect 235531 89644 235576 89672
rect 235570 89632 235576 89644
rect 235628 89632 235634 89684
rect 268690 89672 268696 89684
rect 268651 89644 268696 89672
rect 268690 89632 268696 89644
rect 268748 89632 268754 89684
rect 1600 89168 583316 89264
rect 97018 88952 97024 89004
rect 97076 88992 97082 89004
rect 249002 88992 249008 89004
rect 97076 88964 249008 88992
rect 97076 88952 97082 88964
rect 249002 88952 249008 88964
rect 249060 88952 249066 89004
rect 1600 88624 583316 88720
rect 246518 88448 246524 88460
rect 246479 88420 246524 88448
rect 246518 88408 246524 88420
rect 246576 88408 246582 88460
rect 1600 88080 583316 88176
rect 1600 87536 583316 87632
rect 242470 87224 242476 87236
rect 242431 87196 242476 87224
rect 242470 87184 242476 87196
rect 242528 87184 242534 87236
rect 552418 87156 552424 87168
rect 552379 87128 552424 87156
rect 552418 87116 552424 87128
rect 552476 87116 552482 87168
rect 1600 86992 583316 87088
rect 242838 86912 242844 86964
rect 242896 86952 242902 86964
rect 242930 86952 242936 86964
rect 242896 86924 242936 86952
rect 242896 86912 242902 86924
rect 242930 86912 242936 86924
rect 242988 86912 242994 86964
rect 305122 86952 305128 86964
rect 305083 86924 305128 86952
rect 305122 86912 305128 86924
rect 305180 86912 305186 86964
rect 331066 86912 331072 86964
rect 331124 86952 331130 86964
rect 331250 86952 331256 86964
rect 331124 86924 331256 86952
rect 331124 86912 331130 86924
rect 331250 86912 331256 86924
rect 331308 86912 331314 86964
rect 341094 86952 341100 86964
rect 341055 86924 341100 86952
rect 341094 86912 341100 86924
rect 341152 86912 341158 86964
rect 361334 86912 361340 86964
rect 361392 86952 361398 86964
rect 580662 86952 580668 86964
rect 361392 86924 580668 86952
rect 361392 86912 361398 86924
rect 580662 86912 580668 86924
rect 580720 86912 580726 86964
rect 242470 86884 242476 86896
rect 242431 86856 242476 86884
rect 242470 86844 242476 86856
rect 242528 86844 242534 86896
rect 552418 86884 552424 86896
rect 552379 86856 552424 86884
rect 552418 86844 552424 86856
rect 552476 86844 552482 86896
rect 279822 86776 279828 86828
rect 279880 86816 279886 86828
rect 280006 86816 280012 86828
rect 279880 86788 280012 86816
rect 279880 86776 279886 86788
rect 280006 86776 280012 86788
rect 280064 86776 280070 86828
rect 1600 86448 583316 86544
rect 1600 85904 583316 86000
rect 229869 85595 229927 85601
rect 229869 85561 229881 85595
rect 229915 85592 229927 85595
rect 230050 85592 230056 85604
rect 229915 85564 230056 85592
rect 229915 85561 229927 85564
rect 229869 85555 229927 85561
rect 230050 85552 230056 85564
rect 230108 85552 230114 85604
rect 371917 85595 371975 85601
rect 371917 85561 371929 85595
rect 371963 85592 371975 85595
rect 372006 85592 372012 85604
rect 371963 85564 372012 85592
rect 371963 85561 371975 85564
rect 371917 85555 371975 85561
rect 372006 85552 372012 85564
rect 372064 85552 372070 85604
rect 135658 85524 135664 85536
rect 135619 85496 135664 85524
rect 135658 85484 135664 85496
rect 135716 85484 135722 85536
rect 152218 85524 152224 85536
rect 152179 85496 152224 85524
rect 152218 85484 152224 85496
rect 152276 85484 152282 85536
rect 170158 85524 170164 85536
rect 170119 85496 170164 85524
rect 170158 85484 170164 85496
rect 170216 85484 170222 85536
rect 190858 85524 190864 85536
rect 190819 85496 190864 85524
rect 190858 85484 190864 85496
rect 190916 85484 190922 85536
rect 214318 85524 214324 85536
rect 214279 85496 214324 85524
rect 214318 85484 214324 85496
rect 214376 85484 214382 85536
rect 242470 85524 242476 85536
rect 242431 85496 242476 85524
rect 242470 85484 242476 85496
rect 242528 85484 242534 85536
rect 319934 85524 319940 85536
rect 319895 85496 319940 85524
rect 319934 85484 319940 85496
rect 319992 85484 319998 85536
rect 373110 85524 373116 85536
rect 373071 85496 373116 85524
rect 373110 85484 373116 85496
rect 373168 85484 373174 85536
rect 385530 85484 385536 85536
rect 385588 85524 385594 85536
rect 392430 85524 392436 85536
rect 385588 85496 385633 85524
rect 392391 85496 392436 85524
rect 385588 85484 385594 85496
rect 392430 85484 392436 85496
rect 392488 85484 392494 85536
rect 529050 85524 529056 85536
rect 529011 85496 529056 85524
rect 529050 85484 529056 85496
rect 529108 85484 529114 85536
rect 535950 85524 535956 85536
rect 535911 85496 535956 85524
rect 535950 85484 535956 85496
rect 536008 85484 536014 85536
rect 552329 85527 552387 85533
rect 552329 85493 552341 85527
rect 552375 85524 552387 85527
rect 552418 85524 552424 85536
rect 552375 85496 552424 85524
rect 552375 85493 552387 85496
rect 552329 85487 552387 85493
rect 552418 85484 552424 85496
rect 552476 85484 552482 85536
rect 571830 85524 571836 85536
rect 571791 85496 571836 85524
rect 571830 85484 571836 85496
rect 571888 85484 571894 85536
rect 1600 85360 583316 85456
rect 242473 85323 242531 85329
rect 242473 85289 242485 85323
rect 242519 85320 242531 85323
rect 242562 85320 242568 85332
rect 242519 85292 242568 85320
rect 242519 85289 242531 85292
rect 242473 85283 242531 85289
rect 242562 85280 242568 85292
rect 242620 85280 242626 85332
rect 1600 84816 583316 84912
rect 1600 84272 583316 84368
rect 280006 84232 280012 84244
rect 279932 84204 280012 84232
rect 279932 84176 279960 84204
rect 280006 84192 280012 84204
rect 280064 84192 280070 84244
rect 279914 84124 279920 84176
rect 279972 84124 279978 84176
rect 1600 83728 583316 83824
rect 1600 83184 583316 83280
rect 276970 82900 276976 82952
rect 277028 82940 277034 82952
rect 277028 82912 277108 82940
rect 277028 82900 277034 82912
rect 277080 82884 277108 82912
rect 277062 82832 277068 82884
rect 277120 82832 277126 82884
rect 276602 82804 276608 82816
rect 276563 82776 276608 82804
rect 276602 82764 276608 82776
rect 276660 82764 276666 82816
rect 279822 82764 279828 82816
rect 279880 82804 279886 82816
rect 280098 82804 280104 82816
rect 279880 82776 280104 82804
rect 279880 82764 279886 82776
rect 280098 82764 280104 82776
rect 280156 82764 280162 82816
rect 285250 82804 285256 82816
rect 285211 82776 285256 82804
rect 285250 82764 285256 82776
rect 285308 82764 285314 82816
rect 1600 82640 583316 82736
rect 1600 82096 583316 82192
rect 1600 81552 583316 81648
rect 271361 81515 271419 81521
rect 271361 81481 271373 81515
rect 271407 81512 271419 81515
rect 271450 81512 271456 81524
rect 271407 81484 271456 81512
rect 271407 81481 271419 81484
rect 271361 81475 271419 81481
rect 271450 81472 271456 81484
rect 271508 81472 271514 81524
rect 1600 81008 583316 81104
rect 1600 80464 583316 80560
rect 229961 80155 230019 80161
rect 229961 80121 229973 80155
rect 230007 80152 230019 80155
rect 230050 80152 230056 80164
rect 230007 80124 230056 80152
rect 230007 80121 230019 80124
rect 229961 80115 230019 80121
rect 230050 80112 230056 80124
rect 230108 80112 230114 80164
rect 271358 80084 271364 80096
rect 271319 80056 271364 80084
rect 271358 80044 271364 80056
rect 271416 80044 271422 80096
rect 1600 79920 583316 80016
rect 229958 79880 229964 79892
rect 229919 79852 229964 79880
rect 229958 79840 229964 79852
rect 230016 79840 230022 79892
rect 305122 79880 305128 79892
rect 305083 79852 305128 79880
rect 305122 79840 305128 79852
rect 305180 79840 305186 79892
rect 1600 79376 583316 79472
rect 1600 78832 583316 78928
rect 1600 78288 583316 78384
rect 285250 77976 285256 77988
rect 285211 77948 285256 77976
rect 285250 77936 285256 77948
rect 285308 77936 285314 77988
rect 1600 77744 583316 77840
rect 341097 77435 341155 77441
rect 341097 77401 341109 77435
rect 341143 77432 341155 77435
rect 341186 77432 341192 77444
rect 341143 77404 341192 77432
rect 341143 77401 341155 77404
rect 341097 77395 341155 77401
rect 341186 77392 341192 77404
rect 341244 77392 341250 77444
rect 1600 77200 583316 77296
rect 91498 77160 91504 77172
rect 91459 77132 91504 77160
rect 91498 77120 91504 77132
rect 91556 77120 91562 77172
rect 235481 77163 235539 77169
rect 235481 77129 235493 77163
rect 235527 77160 235539 77163
rect 235570 77160 235576 77172
rect 235527 77132 235576 77160
rect 235527 77129 235539 77132
rect 235481 77123 235539 77129
rect 235570 77120 235576 77132
rect 235628 77120 235634 77172
rect 341097 77163 341155 77169
rect 341097 77129 341109 77163
rect 341143 77160 341155 77163
rect 341186 77160 341192 77172
rect 341143 77132 341192 77160
rect 341143 77129 341155 77132
rect 341097 77123 341155 77129
rect 341186 77120 341192 77132
rect 341244 77120 341250 77172
rect 357930 77120 357936 77172
rect 357988 77160 357994 77172
rect 552326 77160 552332 77172
rect 357988 77132 358033 77160
rect 552287 77132 552332 77160
rect 357988 77120 357994 77132
rect 552326 77120 552332 77132
rect 552384 77120 552390 77172
rect 1600 76656 583316 76752
rect 271358 76576 271364 76628
rect 271416 76616 271422 76628
rect 271453 76619 271511 76625
rect 271453 76616 271465 76619
rect 271416 76588 271465 76616
rect 271416 76576 271422 76588
rect 271453 76585 271465 76588
rect 271499 76585 271511 76619
rect 271453 76579 271511 76585
rect 1600 76112 583316 76208
rect 135658 75936 135664 75948
rect 135619 75908 135664 75936
rect 135658 75896 135664 75908
rect 135716 75896 135722 75948
rect 152218 75936 152224 75948
rect 152179 75908 152224 75936
rect 152218 75896 152224 75908
rect 152276 75896 152282 75948
rect 170158 75936 170164 75948
rect 170119 75908 170164 75936
rect 170158 75896 170164 75908
rect 170216 75896 170222 75948
rect 190858 75936 190864 75948
rect 190819 75908 190864 75936
rect 190858 75896 190864 75908
rect 190916 75896 190922 75948
rect 214318 75936 214324 75948
rect 214279 75908 214324 75936
rect 214318 75896 214324 75908
rect 214376 75896 214382 75948
rect 319937 75939 319995 75945
rect 319937 75905 319949 75939
rect 319983 75936 319995 75939
rect 320118 75936 320124 75948
rect 319983 75908 320124 75936
rect 319983 75905 319995 75908
rect 319937 75899 319995 75905
rect 320118 75896 320124 75908
rect 320176 75896 320182 75948
rect 373110 75936 373116 75948
rect 373071 75908 373116 75936
rect 373110 75896 373116 75908
rect 373168 75896 373174 75948
rect 385530 75896 385536 75948
rect 385588 75936 385594 75948
rect 392430 75936 392436 75948
rect 385588 75908 385633 75936
rect 392391 75908 392436 75936
rect 385588 75896 385594 75908
rect 392430 75896 392436 75908
rect 392488 75896 392494 75948
rect 529050 75936 529056 75948
rect 529011 75908 529056 75936
rect 529050 75896 529056 75908
rect 529108 75896 529114 75948
rect 535950 75936 535956 75948
rect 535911 75908 535956 75936
rect 535950 75896 535956 75908
rect 536008 75896 536014 75948
rect 571830 75936 571836 75948
rect 571791 75908 571836 75936
rect 571830 75896 571836 75908
rect 571888 75896 571894 75948
rect 1600 75568 583316 75664
rect 1600 75024 583316 75120
rect 279914 74644 279920 74656
rect 279875 74616 279920 74644
rect 279914 74604 279920 74616
rect 279972 74604 279978 74656
rect 1600 74480 583316 74576
rect 279914 74440 279920 74452
rect 279875 74412 279920 74440
rect 279914 74400 279920 74412
rect 279972 74400 279978 74452
rect 1600 73936 583316 74032
rect 1600 73392 583316 73488
rect 276602 73216 276608 73228
rect 276563 73188 276608 73216
rect 276602 73176 276608 73188
rect 276660 73176 276666 73228
rect 275593 73151 275651 73157
rect 275593 73117 275605 73151
rect 275639 73148 275651 73151
rect 275682 73148 275688 73160
rect 275639 73120 275688 73148
rect 275639 73117 275651 73120
rect 275593 73111 275651 73117
rect 275682 73108 275688 73120
rect 275740 73108 275746 73160
rect 1600 72848 583316 72944
rect 1600 72304 583316 72400
rect 371914 72156 371920 72208
rect 371972 72196 371978 72208
rect 372098 72196 372104 72208
rect 371972 72168 372104 72196
rect 371972 72156 371978 72168
rect 372098 72156 372104 72168
rect 372156 72156 372162 72208
rect 1600 71760 583316 71856
rect 1600 71216 583316 71312
rect 1600 70672 583316 70768
rect 246702 70496 246708 70508
rect 246663 70468 246708 70496
rect 246702 70456 246708 70468
rect 246760 70456 246766 70508
rect 1600 70128 583316 70224
rect 1600 69584 583316 69680
rect 1600 69040 583316 69136
rect 1600 68496 583316 68592
rect 1600 67952 583316 68048
rect 278718 67708 278724 67720
rect 278644 67680 278724 67708
rect 91498 67640 91504 67652
rect 91459 67612 91504 67640
rect 91498 67600 91504 67612
rect 91556 67600 91562 67652
rect 235478 67640 235484 67652
rect 235439 67612 235484 67640
rect 235478 67600 235484 67612
rect 235536 67600 235542 67652
rect 242010 67600 242016 67652
rect 242068 67640 242074 67652
rect 242102 67640 242108 67652
rect 242068 67612 242108 67640
rect 242068 67600 242074 67612
rect 242102 67600 242108 67612
rect 242160 67600 242166 67652
rect 276970 67600 276976 67652
rect 277028 67640 277034 67652
rect 277065 67643 277123 67649
rect 277065 67640 277077 67643
rect 277028 67612 277077 67640
rect 277028 67600 277034 67612
rect 277065 67609 277077 67612
rect 277111 67609 277123 67643
rect 277065 67603 277123 67609
rect 278644 67584 278672 67680
rect 278718 67668 278724 67680
rect 278776 67668 278782 67720
rect 341094 67640 341100 67652
rect 341055 67612 341100 67640
rect 341094 67600 341100 67612
rect 341152 67600 341158 67652
rect 357930 67600 357936 67652
rect 357988 67640 357994 67652
rect 357988 67612 358033 67640
rect 357988 67600 357994 67612
rect 553890 67600 553896 67652
rect 553948 67640 553954 67652
rect 553982 67640 553988 67652
rect 553948 67612 553988 67640
rect 553948 67600 553954 67612
rect 553982 67600 553988 67612
rect 554040 67600 554046 67652
rect 278626 67532 278632 67584
rect 278684 67532 278690 67584
rect 331250 67572 331256 67584
rect 331211 67544 331256 67572
rect 331250 67532 331256 67544
rect 331308 67532 331314 67584
rect 1600 67408 583316 67504
rect 1600 66864 583316 66960
rect 1600 66320 583316 66416
rect 229866 66240 229872 66292
rect 229924 66280 229930 66292
rect 229958 66280 229964 66292
rect 229924 66252 229964 66280
rect 229924 66240 229930 66252
rect 229958 66240 229964 66252
rect 230016 66240 230022 66292
rect 246702 66280 246708 66292
rect 246663 66252 246708 66280
rect 246702 66240 246708 66252
rect 246760 66240 246766 66292
rect 285618 66240 285624 66292
rect 285676 66280 285682 66292
rect 285802 66280 285808 66292
rect 285676 66252 285808 66280
rect 285676 66240 285682 66252
rect 285802 66240 285808 66252
rect 285860 66240 285866 66292
rect 373202 66240 373208 66292
rect 373260 66280 373266 66292
rect 373294 66280 373300 66292
rect 373260 66252 373300 66280
rect 373260 66240 373266 66252
rect 373294 66240 373300 66252
rect 373352 66240 373358 66292
rect 135658 66212 135664 66224
rect 135619 66184 135664 66212
rect 135658 66172 135664 66184
rect 135716 66172 135722 66224
rect 152218 66212 152224 66224
rect 152179 66184 152224 66212
rect 152218 66172 152224 66184
rect 152276 66172 152282 66224
rect 170158 66212 170164 66224
rect 170119 66184 170164 66212
rect 170158 66172 170164 66184
rect 170216 66172 170222 66224
rect 190858 66212 190864 66224
rect 190819 66184 190864 66212
rect 190858 66172 190864 66184
rect 190916 66172 190922 66224
rect 214318 66212 214324 66224
rect 214279 66184 214324 66212
rect 214318 66172 214324 66184
rect 214376 66172 214382 66224
rect 308897 66215 308955 66221
rect 308897 66181 308909 66215
rect 308943 66212 308955 66215
rect 309078 66212 309084 66224
rect 308943 66184 309084 66212
rect 308943 66181 308955 66184
rect 308897 66175 308955 66181
rect 309078 66172 309084 66184
rect 309136 66172 309142 66224
rect 320118 66212 320124 66224
rect 320079 66184 320124 66212
rect 320118 66172 320124 66184
rect 320176 66172 320182 66224
rect 385530 66172 385536 66224
rect 385588 66212 385594 66224
rect 392430 66212 392436 66224
rect 385588 66184 385633 66212
rect 392391 66184 392436 66212
rect 385588 66172 385594 66184
rect 392430 66172 392436 66184
rect 392488 66172 392494 66224
rect 529050 66212 529056 66224
rect 529011 66184 529056 66212
rect 529050 66172 529056 66184
rect 529108 66172 529114 66224
rect 535950 66212 535956 66224
rect 535911 66184 535956 66212
rect 535950 66172 535956 66184
rect 536008 66172 536014 66224
rect 552510 66212 552516 66224
rect 552471 66184 552516 66212
rect 552510 66172 552516 66184
rect 552568 66172 552574 66224
rect 571830 66212 571836 66224
rect 571791 66184 571836 66212
rect 571830 66172 571836 66184
rect 571888 66172 571894 66224
rect 1600 65776 583316 65872
rect 1600 65232 583316 65328
rect 242562 64988 242568 65000
rect 242488 64960 242568 64988
rect 242488 64932 242516 64960
rect 242562 64948 242568 64960
rect 242620 64948 242626 65000
rect 242470 64880 242476 64932
rect 242528 64880 242534 64932
rect 278626 64852 278632 64864
rect 278587 64824 278632 64852
rect 278626 64812 278632 64824
rect 278684 64812 278690 64864
rect 279730 64852 279736 64864
rect 279691 64824 279736 64852
rect 279730 64812 279736 64824
rect 279788 64812 279794 64864
rect 285250 64852 285256 64864
rect 285211 64824 285256 64852
rect 285250 64812 285256 64824
rect 285308 64812 285314 64864
rect 371917 64855 371975 64861
rect 371917 64821 371929 64855
rect 371963 64852 371975 64855
rect 372006 64852 372012 64864
rect 371963 64824 372012 64852
rect 371963 64821 371975 64824
rect 371917 64815 371975 64821
rect 372006 64812 372012 64824
rect 372064 64812 372070 64864
rect 1600 64688 583316 64784
rect 1600 64144 583316 64240
rect 1600 63600 583316 63696
rect 271450 63560 271456 63572
rect 271411 63532 271456 63560
rect 271450 63520 271456 63532
rect 271508 63520 271514 63572
rect 275590 63560 275596 63572
rect 275551 63532 275596 63560
rect 275590 63520 275596 63532
rect 275648 63520 275654 63572
rect 242470 63492 242476 63504
rect 242431 63464 242476 63492
rect 242470 63452 242476 63464
rect 242528 63452 242534 63504
rect 1600 63056 583316 63152
rect 331250 62812 331256 62824
rect 331211 62784 331256 62812
rect 331250 62772 331256 62784
rect 331308 62772 331314 62824
rect 277062 62744 277068 62756
rect 277023 62716 277068 62744
rect 277062 62704 277068 62716
rect 277120 62704 277126 62756
rect 1600 62512 583316 62608
rect 273014 62092 273020 62144
rect 273072 62132 273078 62144
rect 273106 62132 273112 62144
rect 273072 62104 273112 62132
rect 273072 62092 273078 62104
rect 273106 62092 273112 62104
rect 273164 62092 273170 62144
rect 1600 61968 583316 62064
rect 1600 61424 583316 61520
rect 1600 60880 583316 60976
rect 229866 60840 229872 60852
rect 229792 60812 229872 60840
rect 229792 60716 229820 60812
rect 229866 60800 229872 60812
rect 229924 60800 229930 60852
rect 235478 60732 235484 60784
rect 235536 60732 235542 60784
rect 341186 60772 341192 60784
rect 341112 60744 341192 60772
rect 229774 60664 229780 60716
rect 229832 60664 229838 60716
rect 235496 60636 235524 60732
rect 341112 60716 341140 60744
rect 341186 60732 341192 60744
rect 341244 60732 341250 60784
rect 341094 60664 341100 60716
rect 341152 60664 341158 60716
rect 235570 60636 235576 60648
rect 235496 60608 235576 60636
rect 235570 60596 235576 60608
rect 235628 60596 235634 60648
rect 1600 60336 583316 60432
rect 1600 59792 583316 59888
rect 1600 59248 583316 59344
rect 3638 59168 3644 59220
rect 3696 59208 3702 59220
rect 219194 59208 219200 59220
rect 3696 59180 219200 59208
rect 3696 59168 3702 59180
rect 219194 59168 219200 59180
rect 219252 59168 219258 59220
rect 1600 58704 583316 58800
rect 1600 58160 583316 58256
rect 553890 58012 553896 58064
rect 553948 58012 553954 58064
rect 275590 57984 275596 57996
rect 275551 57956 275596 57984
rect 275590 57944 275596 57956
rect 275648 57944 275654 57996
rect 91498 57916 91504 57928
rect 91459 57888 91504 57916
rect 91498 57876 91504 57888
rect 91556 57876 91562 57928
rect 225174 57876 225180 57928
rect 225232 57916 225238 57928
rect 225358 57916 225364 57928
rect 225232 57888 225364 57916
rect 225232 57876 225238 57888
rect 225358 57876 225364 57888
rect 225416 57876 225422 57928
rect 235389 57919 235447 57925
rect 235389 57885 235401 57919
rect 235435 57916 235447 57919
rect 235570 57916 235576 57928
rect 235435 57888 235576 57916
rect 235435 57885 235447 57888
rect 235389 57879 235447 57885
rect 235570 57876 235576 57888
rect 235628 57876 235634 57928
rect 272830 57916 272836 57928
rect 272791 57888 272836 57916
rect 272830 57876 272836 57888
rect 272888 57876 272894 57928
rect 340910 57876 340916 57928
rect 340968 57916 340974 57928
rect 341186 57916 341192 57928
rect 340968 57888 341192 57916
rect 340968 57876 340974 57888
rect 341186 57876 341192 57888
rect 341244 57876 341250 57928
rect 357930 57876 357936 57928
rect 357988 57916 357994 57928
rect 553908 57916 553936 58012
rect 553982 57916 553988 57928
rect 357988 57888 358033 57916
rect 553908 57888 553988 57916
rect 357988 57876 357994 57888
rect 553982 57876 553988 57888
rect 554040 57876 554046 57928
rect 1600 57616 583316 57712
rect 276418 57264 276424 57316
rect 276476 57304 276482 57316
rect 276513 57307 276571 57313
rect 276513 57304 276525 57307
rect 276476 57276 276525 57304
rect 276476 57264 276482 57276
rect 276513 57273 276525 57276
rect 276559 57273 276571 57307
rect 276513 57267 276571 57273
rect 1600 57072 583316 57168
rect 135658 56692 135664 56704
rect 135619 56664 135664 56692
rect 135658 56652 135664 56664
rect 135716 56652 135722 56704
rect 152218 56692 152224 56704
rect 152179 56664 152224 56692
rect 152218 56652 152224 56664
rect 152276 56652 152282 56704
rect 170158 56692 170164 56704
rect 170119 56664 170164 56692
rect 170158 56652 170164 56664
rect 170216 56652 170222 56704
rect 190858 56692 190864 56704
rect 190819 56664 190864 56692
rect 190858 56652 190864 56664
rect 190916 56652 190922 56704
rect 214318 56692 214324 56704
rect 214279 56664 214324 56692
rect 214318 56652 214324 56664
rect 214376 56652 214382 56704
rect 308894 56692 308900 56704
rect 308855 56664 308900 56692
rect 308894 56652 308900 56664
rect 308952 56652 308958 56704
rect 320118 56692 320124 56704
rect 320079 56664 320124 56692
rect 320118 56652 320124 56664
rect 320176 56652 320182 56704
rect 373110 56652 373116 56704
rect 373168 56692 373174 56704
rect 373294 56692 373300 56704
rect 373168 56664 373300 56692
rect 373168 56652 373174 56664
rect 373294 56652 373300 56664
rect 373352 56652 373358 56704
rect 385530 56652 385536 56704
rect 385588 56692 385594 56704
rect 392430 56692 392436 56704
rect 385588 56664 385633 56692
rect 392391 56664 392436 56692
rect 385588 56652 385594 56664
rect 392430 56652 392436 56664
rect 392488 56652 392494 56704
rect 529050 56692 529056 56704
rect 529011 56664 529056 56692
rect 529050 56652 529056 56664
rect 529108 56652 529114 56704
rect 535950 56692 535956 56704
rect 535911 56664 535956 56692
rect 535950 56652 535956 56664
rect 536008 56652 536014 56704
rect 552510 56692 552516 56704
rect 552471 56664 552516 56692
rect 552510 56652 552516 56664
rect 552568 56652 552574 56704
rect 571830 56692 571836 56704
rect 571791 56664 571836 56692
rect 571830 56652 571836 56664
rect 571888 56652 571894 56704
rect 1600 56528 583316 56624
rect 285250 56488 285256 56500
rect 285211 56460 285256 56488
rect 285250 56448 285256 56460
rect 285308 56448 285314 56500
rect 1600 55984 583316 56080
rect 1600 55440 583316 55536
rect 278629 55267 278687 55273
rect 278629 55233 278641 55267
rect 278675 55264 278687 55267
rect 278718 55264 278724 55276
rect 278675 55236 278724 55264
rect 278675 55233 278687 55236
rect 278629 55227 278687 55233
rect 278718 55224 278724 55236
rect 278776 55224 278782 55276
rect 279730 55264 279736 55276
rect 279691 55236 279736 55264
rect 279730 55224 279736 55236
rect 279788 55224 279794 55276
rect 371914 55264 371920 55276
rect 371875 55236 371920 55264
rect 371914 55224 371920 55236
rect 371972 55224 371978 55276
rect 246886 55196 246892 55208
rect 246847 55168 246892 55196
rect 246886 55156 246892 55168
rect 246944 55156 246950 55208
rect 1600 54896 583316 54992
rect 1600 54352 583316 54448
rect 1600 53808 583316 53904
rect 1600 53264 583316 53360
rect 1600 52720 583316 52816
rect 268598 52504 268604 52556
rect 268656 52544 268662 52556
rect 268690 52544 268696 52556
rect 268656 52516 268696 52544
rect 268656 52504 268662 52516
rect 268690 52504 268696 52516
rect 268748 52504 268754 52556
rect 275590 52476 275596 52488
rect 275551 52448 275596 52476
rect 275590 52436 275596 52448
rect 275648 52436 275654 52488
rect 1600 52176 583316 52272
rect 279730 51756 279736 51808
rect 279788 51796 279794 51808
rect 280006 51796 280012 51808
rect 279788 51768 280012 51796
rect 279788 51756 279794 51768
rect 280006 51756 280012 51768
rect 280064 51756 280070 51808
rect 1600 51632 583316 51728
rect 1600 51088 583316 51184
rect 239250 51008 239256 51060
rect 239308 51048 239314 51060
rect 239434 51048 239440 51060
rect 239308 51020 239440 51048
rect 239308 51008 239314 51020
rect 239434 51008 239440 51020
rect 239492 51008 239498 51060
rect 259214 51008 259220 51060
rect 259272 51048 259278 51060
rect 259398 51048 259404 51060
rect 259272 51020 259404 51048
rect 259272 51008 259278 51020
rect 259398 51008 259404 51020
rect 259456 51008 259462 51060
rect 271358 51008 271364 51060
rect 271416 51048 271422 51060
rect 271542 51048 271548 51060
rect 271416 51020 271548 51048
rect 271416 51008 271422 51020
rect 271542 51008 271548 51020
rect 271600 51008 271606 51060
rect 1600 50544 583316 50640
rect 1600 50000 583316 50096
rect 1600 49456 583316 49552
rect 1600 48912 583316 49008
rect 1600 48368 583316 48464
rect 91498 48328 91504 48340
rect 91459 48300 91504 48328
rect 91498 48288 91504 48300
rect 91556 48288 91562 48340
rect 235386 48328 235392 48340
rect 235347 48300 235392 48328
rect 235386 48288 235392 48300
rect 235444 48288 235450 48340
rect 242746 48288 242752 48340
rect 242804 48328 242810 48340
rect 242838 48328 242844 48340
rect 242804 48300 242844 48328
rect 242804 48288 242810 48300
rect 242838 48288 242844 48300
rect 242896 48288 242902 48340
rect 272830 48328 272836 48340
rect 272791 48300 272836 48328
rect 272830 48288 272836 48300
rect 272888 48288 272894 48340
rect 278721 48331 278779 48337
rect 278721 48297 278733 48331
rect 278767 48328 278779 48331
rect 278810 48328 278816 48340
rect 278767 48300 278816 48328
rect 278767 48297 278779 48300
rect 278721 48291 278779 48297
rect 278810 48288 278816 48300
rect 278868 48288 278874 48340
rect 357930 48288 357936 48340
rect 357988 48328 357994 48340
rect 357988 48300 358033 48328
rect 357988 48288 357994 48300
rect 259309 48263 259367 48269
rect 259309 48229 259321 48263
rect 259355 48260 259367 48263
rect 259398 48260 259404 48272
rect 259355 48232 259404 48260
rect 259355 48229 259367 48232
rect 259309 48223 259367 48229
rect 259398 48220 259404 48232
rect 259456 48220 259462 48272
rect 341002 48220 341008 48272
rect 341060 48260 341066 48272
rect 341094 48260 341100 48272
rect 341060 48232 341100 48260
rect 341060 48220 341066 48232
rect 341094 48220 341100 48232
rect 341152 48220 341158 48272
rect 553798 48220 553804 48272
rect 553856 48260 553862 48272
rect 553890 48260 553896 48272
rect 553856 48232 553896 48260
rect 553856 48220 553862 48232
rect 553890 48220 553896 48232
rect 553948 48220 553954 48272
rect 1600 47824 583316 47920
rect 1600 47280 583316 47376
rect 319842 46996 319848 47048
rect 319900 47036 319906 47048
rect 320026 47036 320032 47048
rect 319900 47008 320032 47036
rect 319900 46996 319906 47008
rect 320026 46996 320032 47008
rect 320084 46996 320090 47048
rect 275590 46968 275596 46980
rect 275551 46940 275596 46968
rect 275590 46928 275596 46940
rect 275648 46928 275654 46980
rect 135658 46900 135664 46912
rect 135619 46872 135664 46900
rect 135658 46860 135664 46872
rect 135716 46860 135722 46912
rect 152218 46900 152224 46912
rect 152179 46872 152224 46900
rect 152218 46860 152224 46872
rect 152276 46860 152282 46912
rect 170158 46900 170164 46912
rect 170119 46872 170164 46900
rect 170158 46860 170164 46872
rect 170216 46860 170222 46912
rect 190858 46900 190864 46912
rect 190819 46872 190864 46900
rect 190858 46860 190864 46872
rect 190916 46860 190922 46912
rect 214318 46900 214324 46912
rect 214279 46872 214324 46900
rect 214318 46860 214324 46872
rect 214376 46860 214382 46912
rect 225358 46900 225364 46912
rect 225319 46872 225364 46900
rect 225358 46860 225364 46872
rect 225416 46860 225422 46912
rect 242010 46860 242016 46912
rect 242068 46900 242074 46912
rect 242102 46900 242108 46912
rect 242068 46872 242108 46900
rect 242068 46860 242074 46872
rect 242102 46860 242108 46872
rect 242160 46860 242166 46912
rect 272830 46900 272836 46912
rect 272791 46872 272836 46900
rect 272830 46860 272836 46872
rect 272888 46860 272894 46912
rect 285066 46860 285072 46912
rect 285124 46900 285130 46912
rect 285250 46900 285256 46912
rect 285124 46872 285256 46900
rect 285124 46860 285130 46872
rect 285250 46860 285256 46872
rect 285308 46860 285314 46912
rect 308986 46860 308992 46912
rect 309044 46900 309050 46912
rect 309170 46900 309176 46912
rect 309044 46872 309176 46900
rect 309044 46860 309050 46872
rect 309170 46860 309176 46872
rect 309228 46860 309234 46912
rect 319937 46903 319995 46909
rect 319937 46869 319949 46903
rect 319983 46900 319995 46903
rect 320026 46900 320032 46912
rect 319983 46872 320032 46900
rect 319983 46869 319995 46872
rect 319937 46863 319995 46869
rect 320026 46860 320032 46872
rect 320084 46860 320090 46912
rect 328217 46903 328275 46909
rect 328217 46869 328229 46903
rect 328263 46900 328275 46903
rect 328398 46900 328404 46912
rect 328263 46872 328404 46900
rect 328263 46869 328275 46872
rect 328217 46863 328275 46869
rect 328398 46860 328404 46872
rect 328456 46860 328462 46912
rect 385530 46860 385536 46912
rect 385588 46900 385594 46912
rect 392430 46900 392436 46912
rect 385588 46872 385633 46900
rect 392391 46872 392436 46900
rect 385588 46860 385594 46872
rect 392430 46860 392436 46872
rect 392488 46860 392494 46912
rect 529050 46900 529056 46912
rect 529011 46872 529056 46900
rect 529050 46860 529056 46872
rect 529108 46860 529114 46912
rect 535950 46900 535956 46912
rect 535911 46872 535956 46900
rect 535950 46860 535956 46872
rect 536008 46860 536014 46912
rect 552510 46900 552516 46912
rect 552471 46872 552516 46900
rect 552510 46860 552516 46872
rect 552568 46860 552574 46912
rect 553798 46900 553804 46912
rect 553759 46872 553804 46900
rect 553798 46860 553804 46872
rect 553856 46860 553862 46912
rect 571830 46900 571836 46912
rect 571791 46872 571836 46900
rect 571830 46860 571836 46872
rect 571888 46860 571894 46912
rect 1600 46736 583316 46832
rect 392433 46699 392491 46705
rect 392433 46665 392445 46699
rect 392479 46696 392491 46699
rect 392522 46696 392528 46708
rect 392479 46668 392528 46696
rect 392479 46665 392491 46668
rect 392433 46659 392491 46665
rect 392522 46656 392528 46668
rect 392580 46656 392586 46708
rect 1600 46192 583316 46288
rect 1600 45648 583316 45744
rect 242473 45611 242531 45617
rect 242473 45577 242485 45611
rect 242519 45608 242531 45611
rect 242562 45608 242568 45620
rect 242519 45580 242568 45608
rect 242519 45577 242531 45580
rect 242473 45571 242531 45577
rect 242562 45568 242568 45580
rect 242620 45568 242626 45620
rect 246886 45608 246892 45620
rect 246847 45580 246892 45608
rect 246886 45568 246892 45580
rect 246944 45568 246950 45620
rect 278718 45608 278724 45620
rect 278679 45580 278724 45608
rect 278718 45568 278724 45580
rect 278776 45568 278782 45620
rect 1600 45104 583316 45200
rect 1600 44560 583316 44656
rect 276513 44183 276571 44189
rect 276513 44149 276525 44183
rect 276559 44180 276571 44183
rect 276602 44180 276608 44192
rect 276559 44152 276608 44180
rect 276559 44149 276571 44152
rect 276513 44143 276571 44149
rect 276602 44140 276608 44152
rect 276660 44140 276666 44192
rect 1600 44016 583316 44112
rect 1600 43472 583316 43568
rect 1600 42928 583316 43024
rect 273106 42780 273112 42832
rect 273164 42820 273170 42832
rect 273290 42820 273296 42832
rect 273164 42792 273296 42820
rect 273164 42780 273170 42792
rect 273290 42780 273296 42792
rect 273348 42780 273354 42832
rect 275590 42820 275596 42832
rect 275551 42792 275596 42820
rect 275590 42780 275596 42792
rect 275648 42780 275654 42832
rect 273106 42644 273112 42696
rect 273164 42644 273170 42696
rect 273014 42576 273020 42628
rect 273072 42616 273078 42628
rect 273124 42616 273152 42644
rect 273072 42588 273152 42616
rect 273072 42576 273078 42588
rect 1600 42384 583316 42480
rect 285618 42032 285624 42084
rect 285676 42072 285682 42084
rect 285713 42075 285771 42081
rect 285713 42072 285725 42075
rect 285676 42044 285725 42072
rect 285676 42032 285682 42044
rect 285713 42041 285725 42044
rect 285759 42041 285771 42075
rect 285713 42035 285771 42041
rect 1600 41840 583316 41936
rect 1600 41296 583316 41392
rect 1600 40752 583316 40848
rect 1600 40208 583316 40304
rect 1600 39664 583316 39760
rect 1600 39120 583316 39216
rect 399238 38836 399244 38888
rect 399296 38876 399302 38888
rect 406138 38876 406144 38888
rect 399296 38848 406144 38876
rect 399296 38836 399302 38848
rect 406138 38836 406144 38848
rect 406196 38836 406202 38888
rect 298590 38768 298596 38820
rect 298648 38808 298654 38820
rect 308158 38808 308164 38820
rect 298648 38780 308164 38808
rect 298648 38768 298654 38780
rect 308158 38768 308164 38780
rect 308216 38768 308222 38820
rect 259306 38740 259312 38752
rect 259267 38712 259312 38740
rect 259306 38700 259312 38712
rect 259364 38700 259370 38752
rect 261054 38700 261060 38752
rect 261112 38740 261118 38752
rect 268138 38740 268144 38752
rect 261112 38712 268144 38740
rect 261112 38700 261118 38712
rect 268138 38700 268144 38712
rect 268196 38700 268202 38752
rect 377342 38700 377348 38752
rect 377400 38740 377406 38752
rect 382034 38740 382040 38752
rect 377400 38712 382040 38740
rect 377400 38700 377406 38712
rect 382034 38700 382040 38712
rect 382092 38700 382098 38752
rect 1600 38576 583316 38672
rect 91498 38536 91504 38548
rect 91459 38508 91504 38536
rect 91498 38496 91504 38508
rect 91556 38496 91562 38548
rect 320302 38536 320308 38548
rect 320263 38508 320308 38536
rect 320302 38496 320308 38508
rect 320360 38496 320366 38548
rect 357930 38496 357936 38548
rect 357988 38536 357994 38548
rect 357988 38508 358033 38536
rect 357988 38496 357994 38508
rect 553798 38400 553804 38412
rect 553759 38372 553804 38400
rect 553798 38360 553804 38372
rect 553856 38360 553862 38412
rect 1600 38032 583316 38128
rect 275498 37952 275504 38004
rect 275556 37992 275562 38004
rect 275593 37995 275651 38001
rect 275593 37992 275605 37995
rect 275556 37964 275605 37992
rect 275556 37952 275562 37964
rect 275593 37961 275605 37964
rect 275639 37961 275651 37995
rect 275593 37955 275651 37961
rect 276234 37952 276240 38004
rect 276292 37992 276298 38004
rect 276602 37992 276608 38004
rect 276292 37964 276608 37992
rect 276292 37952 276298 37964
rect 276602 37952 276608 37964
rect 276660 37952 276666 38004
rect 1600 37488 583316 37584
rect 135658 37312 135664 37324
rect 135619 37284 135664 37312
rect 135658 37272 135664 37284
rect 135716 37272 135722 37324
rect 152218 37312 152224 37324
rect 152179 37284 152224 37312
rect 152218 37272 152224 37284
rect 152276 37272 152282 37324
rect 170158 37312 170164 37324
rect 170119 37284 170164 37312
rect 170158 37272 170164 37284
rect 170216 37272 170222 37324
rect 190858 37312 190864 37324
rect 190819 37284 190864 37312
rect 190858 37272 190864 37284
rect 190916 37272 190922 37324
rect 214318 37312 214324 37324
rect 214279 37284 214324 37312
rect 214318 37272 214324 37284
rect 214376 37272 214382 37324
rect 225361 37315 225419 37321
rect 225361 37281 225373 37315
rect 225407 37312 225419 37315
rect 225450 37312 225456 37324
rect 225407 37284 225456 37312
rect 225407 37281 225419 37284
rect 225361 37275 225419 37281
rect 225450 37272 225456 37284
rect 225508 37272 225514 37324
rect 271450 37272 271456 37324
rect 271508 37312 271514 37324
rect 271542 37312 271548 37324
rect 271508 37284 271548 37312
rect 271508 37272 271514 37284
rect 271542 37272 271548 37284
rect 271600 37272 271606 37324
rect 272830 37312 272836 37324
rect 272791 37284 272836 37312
rect 272830 37272 272836 37284
rect 272888 37272 272894 37324
rect 276970 37272 276976 37324
rect 277028 37312 277034 37324
rect 277062 37312 277068 37324
rect 277028 37284 277068 37312
rect 277028 37272 277034 37284
rect 277062 37272 277068 37284
rect 277120 37272 277126 37324
rect 280006 37312 280012 37324
rect 279840 37284 280012 37312
rect 279840 37256 279868 37284
rect 280006 37272 280012 37284
rect 280064 37272 280070 37324
rect 319934 37312 319940 37324
rect 319895 37284 319940 37312
rect 319934 37272 319940 37284
rect 319992 37272 319998 37324
rect 328214 37312 328220 37324
rect 328175 37284 328220 37312
rect 328214 37272 328220 37284
rect 328272 37272 328278 37324
rect 371914 37272 371920 37324
rect 371972 37312 371978 37324
rect 372006 37312 372012 37324
rect 371972 37284 372012 37312
rect 371972 37272 371978 37284
rect 372006 37272 372012 37284
rect 372064 37272 372070 37324
rect 373018 37272 373024 37324
rect 373076 37312 373082 37324
rect 373110 37312 373116 37324
rect 373076 37284 373116 37312
rect 373076 37272 373082 37284
rect 373110 37272 373116 37284
rect 373168 37272 373174 37324
rect 385530 37272 385536 37324
rect 385588 37312 385594 37324
rect 529050 37312 529056 37324
rect 385588 37284 385633 37312
rect 529011 37284 529056 37312
rect 385588 37272 385594 37284
rect 529050 37272 529056 37284
rect 529108 37272 529114 37324
rect 535950 37312 535956 37324
rect 535911 37284 535956 37312
rect 535950 37272 535956 37284
rect 536008 37272 536014 37324
rect 552513 37315 552571 37321
rect 552513 37281 552525 37315
rect 552559 37312 552571 37315
rect 552602 37312 552608 37324
rect 552559 37284 552608 37312
rect 552559 37281 552571 37284
rect 552513 37275 552571 37281
rect 552602 37272 552608 37284
rect 552660 37272 552666 37324
rect 571830 37312 571836 37324
rect 571791 37284 571836 37312
rect 571830 37272 571836 37284
rect 571888 37272 571894 37324
rect 242010 37204 242016 37256
rect 242068 37244 242074 37256
rect 242102 37244 242108 37256
rect 242068 37216 242108 37244
rect 242068 37204 242074 37216
rect 242102 37204 242108 37216
rect 242160 37204 242166 37256
rect 278718 37204 278724 37256
rect 278776 37244 278782 37256
rect 278902 37244 278908 37256
rect 278776 37216 278908 37244
rect 278776 37204 278782 37216
rect 278902 37204 278908 37216
rect 278960 37204 278966 37256
rect 279822 37204 279828 37256
rect 279880 37204 279886 37256
rect 1600 36944 583316 37040
rect 1600 36400 583316 36496
rect 1600 35856 583316 35952
rect 1600 35312 583316 35408
rect 1600 34768 583316 34864
rect 1600 34224 583316 34320
rect 1600 33680 583316 33776
rect 1600 33136 583316 33232
rect 1600 32592 583316 32688
rect 1600 32048 583316 32144
rect 320302 31872 320308 31884
rect 320263 31844 320308 31872
rect 320302 31832 320308 31844
rect 320360 31832 320366 31884
rect 341005 31875 341063 31881
rect 341005 31841 341017 31875
rect 341051 31872 341063 31875
rect 341094 31872 341100 31884
rect 341051 31844 341100 31872
rect 341051 31841 341063 31844
rect 341005 31835 341063 31841
rect 341094 31832 341100 31844
rect 341152 31832 341158 31884
rect 229958 31764 229964 31816
rect 230016 31764 230022 31816
rect 235478 31804 235484 31816
rect 235439 31776 235484 31804
rect 235478 31764 235484 31776
rect 235536 31764 235542 31816
rect 229976 31680 230004 31764
rect 229958 31628 229964 31680
rect 230016 31628 230022 31680
rect 1600 31504 583316 31600
rect 1600 30960 583316 31056
rect 1600 30416 583316 30512
rect 1600 29872 583316 29968
rect 1600 29328 583316 29424
rect 242654 29084 242660 29096
rect 242580 29056 242660 29084
rect 91498 29016 91504 29028
rect 91459 28988 91504 29016
rect 91498 28976 91504 28988
rect 91556 28976 91562 29028
rect 235478 29016 235484 29028
rect 235439 28988 235484 29016
rect 235478 28976 235484 28988
rect 235536 28976 235542 29028
rect 242580 28960 242608 29056
rect 242654 29044 242660 29056
rect 242712 29044 242718 29096
rect 246886 29084 246892 29096
rect 246720 29056 246892 29084
rect 246720 29028 246748 29056
rect 246886 29044 246892 29056
rect 246944 29044 246950 29096
rect 242746 28976 242752 29028
rect 242804 29016 242810 29028
rect 242838 29016 242844 29028
rect 242804 28988 242844 29016
rect 242804 28976 242810 28988
rect 242838 28976 242844 28988
rect 242896 28976 242902 29028
rect 246518 28976 246524 29028
rect 246576 29016 246582 29028
rect 246610 29016 246616 29028
rect 246576 28988 246616 29016
rect 246576 28976 246582 28988
rect 246610 28976 246616 28988
rect 246668 28976 246674 29028
rect 246702 28976 246708 29028
rect 246760 28976 246766 29028
rect 285066 28976 285072 29028
rect 285124 29016 285130 29028
rect 285250 29016 285256 29028
rect 285124 28988 285256 29016
rect 285124 28976 285130 28988
rect 285250 28976 285256 28988
rect 285308 28976 285314 29028
rect 285713 29019 285771 29025
rect 285713 28985 285725 29019
rect 285759 29016 285771 29019
rect 285802 29016 285808 29028
rect 285759 28988 285808 29016
rect 285759 28985 285771 28988
rect 285713 28979 285771 28985
rect 285802 28976 285808 28988
rect 285860 28976 285866 29028
rect 308986 28976 308992 29028
rect 309044 29016 309050 29028
rect 309170 29016 309176 29028
rect 309044 28988 309176 29016
rect 309044 28976 309050 28988
rect 309170 28976 309176 28988
rect 309228 28976 309234 29028
rect 341002 29016 341008 29028
rect 340963 28988 341008 29016
rect 341002 28976 341008 28988
rect 341060 28976 341066 29028
rect 357930 28976 357936 29028
rect 357988 29016 357994 29028
rect 357988 28988 358033 29016
rect 357988 28976 357994 28988
rect 553798 28976 553804 29028
rect 553856 29016 553862 29028
rect 553890 29016 553896 29028
rect 553856 28988 553896 29016
rect 553856 28976 553862 28988
rect 553890 28976 553896 28988
rect 553948 28976 553954 29028
rect 242562 28908 242568 28960
rect 242620 28908 242626 28960
rect 254801 28951 254859 28957
rect 254801 28917 254813 28951
rect 254847 28948 254859 28951
rect 254890 28948 254896 28960
rect 254847 28920 254896 28948
rect 254847 28917 254859 28920
rect 254801 28911 254859 28917
rect 254890 28908 254896 28920
rect 254948 28908 254954 28960
rect 285158 28948 285164 28960
rect 285119 28920 285164 28948
rect 285158 28908 285164 28920
rect 285216 28908 285222 28960
rect 1600 28784 583316 28880
rect 1600 28240 583316 28336
rect 1600 27696 583316 27792
rect 276234 27616 276240 27668
rect 276292 27656 276298 27668
rect 276510 27656 276516 27668
rect 276292 27628 276516 27656
rect 276292 27616 276298 27628
rect 276510 27616 276516 27628
rect 276568 27616 276574 27668
rect 278810 27656 278816 27668
rect 278771 27628 278816 27656
rect 278810 27616 278816 27628
rect 278868 27616 278874 27668
rect 135293 27591 135351 27597
rect 135293 27557 135305 27591
rect 135339 27588 135351 27591
rect 135658 27588 135664 27600
rect 135339 27560 135664 27588
rect 135339 27557 135351 27560
rect 135293 27551 135351 27557
rect 135658 27548 135664 27560
rect 135716 27548 135722 27600
rect 151853 27591 151911 27597
rect 151853 27557 151865 27591
rect 151899 27588 151911 27591
rect 152218 27588 152224 27600
rect 151899 27560 152224 27588
rect 151899 27557 151911 27560
rect 151853 27551 151911 27557
rect 152218 27548 152224 27560
rect 152276 27548 152282 27600
rect 169701 27591 169759 27597
rect 169701 27557 169713 27591
rect 169747 27588 169759 27591
rect 170158 27588 170164 27600
rect 169747 27560 170164 27588
rect 169747 27557 169759 27560
rect 169701 27551 169759 27557
rect 170158 27548 170164 27560
rect 170216 27548 170222 27600
rect 190214 27548 190220 27600
rect 190272 27588 190278 27600
rect 190858 27588 190864 27600
rect 190272 27560 190864 27588
rect 190272 27548 190278 27560
rect 190858 27548 190864 27560
rect 190916 27548 190922 27600
rect 214318 27548 214324 27600
rect 214376 27588 214382 27600
rect 214502 27588 214508 27600
rect 214376 27560 214508 27588
rect 214376 27548 214382 27560
rect 214502 27548 214508 27560
rect 214560 27548 214566 27600
rect 225085 27591 225143 27597
rect 225085 27557 225097 27591
rect 225131 27588 225143 27591
rect 225358 27588 225364 27600
rect 225131 27560 225364 27588
rect 225131 27557 225143 27560
rect 225085 27551 225143 27557
rect 225358 27548 225364 27560
rect 225416 27548 225422 27600
rect 242562 27588 242568 27600
rect 242523 27560 242568 27588
rect 242562 27548 242568 27560
rect 242620 27548 242626 27600
rect 246518 27548 246524 27600
rect 246576 27588 246582 27600
rect 246610 27588 246616 27600
rect 246576 27560 246616 27588
rect 246576 27548 246582 27560
rect 246610 27548 246616 27560
rect 246668 27548 246674 27600
rect 272830 27588 272836 27600
rect 272791 27560 272836 27588
rect 272830 27548 272836 27560
rect 272888 27548 272894 27600
rect 305122 27588 305128 27600
rect 305083 27560 305128 27588
rect 305122 27548 305128 27560
rect 305180 27548 305186 27600
rect 385530 27548 385536 27600
rect 385588 27588 385594 27600
rect 385990 27588 385996 27600
rect 385588 27560 385996 27588
rect 385588 27548 385594 27560
rect 385990 27548 385996 27560
rect 386048 27548 386054 27600
rect 392430 27548 392436 27600
rect 392488 27588 392494 27600
rect 392614 27588 392620 27600
rect 392488 27560 392620 27588
rect 392488 27548 392494 27560
rect 392614 27548 392620 27560
rect 392672 27548 392678 27600
rect 529050 27588 529056 27600
rect 529011 27560 529056 27588
rect 529050 27548 529056 27560
rect 529108 27548 529114 27600
rect 535950 27588 535956 27600
rect 535911 27560 535956 27588
rect 535950 27548 535956 27560
rect 536008 27548 536014 27600
rect 552510 27588 552516 27600
rect 552471 27560 552516 27588
rect 552510 27548 552516 27560
rect 552568 27548 552574 27600
rect 571830 27588 571836 27600
rect 571791 27560 571836 27588
rect 571830 27548 571836 27560
rect 571888 27548 571894 27600
rect 1600 27152 583316 27248
rect 1600 26608 583316 26704
rect 278810 26296 278816 26308
rect 278771 26268 278816 26296
rect 278810 26256 278816 26268
rect 278868 26256 278874 26308
rect 3914 26188 3920 26240
rect 3972 26228 3978 26240
rect 268417 26231 268475 26237
rect 268417 26228 268429 26231
rect 3972 26200 268429 26228
rect 3972 26188 3978 26200
rect 268417 26197 268429 26200
rect 268463 26197 268475 26231
rect 268417 26191 268475 26197
rect 273017 26231 273075 26237
rect 273017 26197 273029 26231
rect 273063 26228 273075 26231
rect 350018 26228 350024 26240
rect 273063 26200 350024 26228
rect 273063 26197 273075 26200
rect 273017 26191 273075 26197
rect 350018 26188 350024 26200
rect 350076 26188 350082 26240
rect 1600 26064 583316 26160
rect 268417 26027 268475 26033
rect 268417 25993 268429 26027
rect 268463 26024 268475 26027
rect 273017 26027 273075 26033
rect 273017 26024 273029 26027
rect 268463 25996 273029 26024
rect 268463 25993 268475 25996
rect 268417 25987 268475 25993
rect 273017 25993 273029 25996
rect 273063 25993 273075 26027
rect 273017 25987 273075 25993
rect 1600 25520 583316 25616
rect 1600 24976 583316 25072
rect 275593 24871 275651 24877
rect 275593 24837 275605 24871
rect 275639 24868 275651 24871
rect 275682 24868 275688 24880
rect 275639 24840 275688 24868
rect 275639 24837 275651 24840
rect 275593 24831 275651 24837
rect 275682 24828 275688 24840
rect 275740 24828 275746 24880
rect 1600 24432 583316 24528
rect 229958 24148 229964 24200
rect 230016 24188 230022 24200
rect 230142 24188 230148 24200
rect 230016 24160 230148 24188
rect 230016 24148 230022 24160
rect 230142 24148 230148 24160
rect 230200 24148 230206 24200
rect 285713 24191 285771 24197
rect 285713 24157 285725 24191
rect 285759 24188 285771 24191
rect 285802 24188 285808 24200
rect 285759 24160 285808 24188
rect 285759 24157 285771 24160
rect 285713 24151 285771 24157
rect 285802 24148 285808 24160
rect 285860 24148 285866 24200
rect 319934 24148 319940 24200
rect 319992 24188 319998 24200
rect 320118 24188 320124 24200
rect 319992 24160 320124 24188
rect 319992 24148 319998 24160
rect 320118 24148 320124 24160
rect 320176 24148 320182 24200
rect 1600 23888 583316 23984
rect 1600 23344 583316 23440
rect 1600 22800 583316 22896
rect 242562 22692 242568 22704
rect 242523 22664 242568 22692
rect 242562 22652 242568 22664
rect 242620 22652 242626 22704
rect 1600 22256 583316 22352
rect 235478 22108 235484 22160
rect 235536 22108 235542 22160
rect 277062 22148 277068 22160
rect 276988 22120 277068 22148
rect 235496 22012 235524 22108
rect 276988 22092 277016 22120
rect 277062 22108 277068 22120
rect 277120 22108 277126 22160
rect 276970 22040 276976 22092
rect 277028 22040 277034 22092
rect 367590 22040 367596 22092
rect 367648 22080 367654 22092
rect 368326 22080 368332 22092
rect 367648 22052 368332 22080
rect 367648 22040 367654 22052
rect 368326 22040 368332 22052
rect 368384 22040 368390 22092
rect 368970 22040 368976 22092
rect 369028 22080 369034 22092
rect 369522 22080 369528 22092
rect 369028 22052 369528 22080
rect 369028 22040 369034 22052
rect 369522 22040 369528 22052
rect 369580 22040 369586 22092
rect 235570 22012 235576 22024
rect 235496 21984 235576 22012
rect 235570 21972 235576 21984
rect 235628 21972 235634 22024
rect 1600 21712 583316 21808
rect 254798 21400 254804 21412
rect 254759 21372 254804 21400
rect 254798 21360 254804 21372
rect 254856 21360 254862 21412
rect 313034 21360 313040 21412
rect 313092 21400 313098 21412
rect 346890 21400 346896 21412
rect 313092 21372 346896 21400
rect 313092 21360 313098 21372
rect 346890 21360 346896 21372
rect 346948 21360 346954 21412
rect 1600 21168 583316 21264
rect 1600 20624 583316 20720
rect 1600 20080 583316 20176
rect 1600 19536 583316 19632
rect 285066 19388 285072 19440
rect 285124 19428 285130 19440
rect 285124 19400 285296 19428
rect 285124 19388 285130 19400
rect 285158 19360 285164 19372
rect 285119 19332 285164 19360
rect 285158 19320 285164 19332
rect 285216 19320 285222 19372
rect 285268 19360 285296 19400
rect 285342 19360 285348 19372
rect 285268 19332 285348 19360
rect 285342 19320 285348 19332
rect 285400 19320 285406 19372
rect 285710 19360 285716 19372
rect 285671 19332 285716 19360
rect 285710 19320 285716 19332
rect 285768 19320 285774 19372
rect 91498 19292 91504 19304
rect 91459 19264 91504 19292
rect 91498 19252 91504 19264
rect 91556 19252 91562 19304
rect 145318 19252 145324 19304
rect 145376 19252 145382 19304
rect 308250 19292 308256 19304
rect 308211 19264 308256 19292
rect 308250 19252 308256 19264
rect 308308 19252 308314 19304
rect 340726 19252 340732 19304
rect 340784 19292 340790 19304
rect 341002 19292 341008 19304
rect 340784 19264 341008 19292
rect 340784 19252 340790 19264
rect 341002 19252 341008 19264
rect 341060 19252 341066 19304
rect 346890 19252 346896 19304
rect 346948 19292 346954 19304
rect 347074 19292 347080 19304
rect 346948 19264 347080 19292
rect 346948 19252 346954 19264
rect 347074 19252 347080 19264
rect 347132 19252 347138 19304
rect 351030 19252 351036 19304
rect 351088 19292 351094 19304
rect 351306 19292 351312 19304
rect 351088 19264 351312 19292
rect 351088 19252 351094 19264
rect 351306 19252 351312 19264
rect 351364 19252 351370 19304
rect 414510 19252 414516 19304
rect 414568 19292 414574 19304
rect 414878 19292 414884 19304
rect 414568 19264 414884 19292
rect 414568 19252 414574 19264
rect 414878 19252 414884 19264
rect 414936 19252 414942 19304
rect 541470 19252 541476 19304
rect 541528 19292 541534 19304
rect 541528 19264 541573 19292
rect 541528 19252 541534 19264
rect 560790 19252 560796 19304
rect 560848 19292 560854 19304
rect 560848 19264 560893 19292
rect 560848 19252 560854 19264
rect 145226 19184 145232 19236
rect 145284 19224 145290 19236
rect 145336 19224 145364 19252
rect 145284 19196 145364 19224
rect 145284 19184 145290 19196
rect 1600 18992 583316 19088
rect 273014 18776 273020 18828
rect 273072 18816 273078 18828
rect 273198 18816 273204 18828
rect 273072 18788 273204 18816
rect 273072 18776 273078 18788
rect 273198 18776 273204 18788
rect 273256 18776 273262 18828
rect 236398 18572 236404 18624
rect 236456 18612 236462 18624
rect 275774 18612 275780 18624
rect 236456 18584 275780 18612
rect 236456 18572 236462 18584
rect 275774 18572 275780 18584
rect 275832 18572 275838 18624
rect 299602 18572 299608 18624
rect 299660 18612 299666 18624
rect 336126 18612 336132 18624
rect 299660 18584 336132 18612
rect 299660 18572 299666 18584
rect 336126 18572 336132 18584
rect 336184 18572 336190 18624
rect 1600 18448 583316 18544
rect 242746 18136 242752 18148
rect 242672 18108 242752 18136
rect 242672 18080 242700 18108
rect 242746 18096 242752 18108
rect 242804 18096 242810 18148
rect 135290 18068 135296 18080
rect 135251 18040 135296 18068
rect 135290 18028 135296 18040
rect 135348 18028 135354 18080
rect 151850 18068 151856 18080
rect 151811 18040 151856 18068
rect 151850 18028 151856 18040
rect 151908 18028 151914 18080
rect 169698 18068 169704 18080
rect 169659 18040 169704 18068
rect 169698 18028 169704 18040
rect 169756 18028 169762 18080
rect 225082 18068 225088 18080
rect 225043 18040 225088 18068
rect 225082 18028 225088 18040
rect 225140 18028 225146 18080
rect 242654 18028 242660 18080
rect 242712 18028 242718 18080
rect 272830 18068 272836 18080
rect 272791 18040 272836 18068
rect 272830 18028 272836 18040
rect 272888 18028 272894 18080
rect 305122 18068 305128 18080
rect 305083 18040 305128 18068
rect 305122 18028 305128 18040
rect 305180 18028 305186 18080
rect 1600 17904 583316 18000
rect 373110 17864 373116 17876
rect 373071 17836 373116 17864
rect 373110 17824 373116 17836
rect 373168 17824 373174 17876
rect 1600 17360 583316 17456
rect 239250 17280 239256 17332
rect 239308 17320 239314 17332
rect 239526 17320 239532 17332
rect 239308 17292 239532 17320
rect 239308 17280 239314 17292
rect 239526 17280 239532 17292
rect 239584 17280 239590 17332
rect 242470 17280 242476 17332
rect 242528 17320 242534 17332
rect 242654 17320 242660 17332
rect 242528 17292 242660 17320
rect 242528 17280 242534 17292
rect 242654 17280 242660 17292
rect 242712 17280 242718 17332
rect 232166 17212 232172 17264
rect 232224 17252 232230 17264
rect 277154 17252 277160 17264
rect 232224 17224 277160 17252
rect 232224 17212 232230 17224
rect 277154 17212 277160 17224
rect 277212 17212 277218 17264
rect 306134 17212 306140 17264
rect 306192 17252 306198 17264
rect 328950 17252 328956 17264
rect 306192 17224 328956 17252
rect 306192 17212 306198 17224
rect 328950 17212 328956 17224
rect 329008 17212 329014 17264
rect 1600 16816 583316 16912
rect 278626 16600 278632 16652
rect 278684 16640 278690 16652
rect 278810 16640 278816 16652
rect 278684 16612 278816 16640
rect 278684 16600 278690 16612
rect 278810 16600 278816 16612
rect 278868 16600 278874 16652
rect 347902 16532 347908 16584
rect 347960 16572 347966 16584
rect 348178 16572 348184 16584
rect 347960 16544 348184 16572
rect 347960 16532 347966 16544
rect 348178 16532 348184 16544
rect 348236 16532 348242 16584
rect 1600 16272 583316 16368
rect 1600 15728 583316 15824
rect 392338 15444 392344 15496
rect 392396 15484 392402 15496
rect 393534 15484 393540 15496
rect 392396 15456 393540 15484
rect 392396 15444 392402 15456
rect 393534 15444 393540 15456
rect 393592 15444 393598 15496
rect 1600 15184 583316 15280
rect 1600 14640 583316 14736
rect 483510 14560 483516 14612
rect 483568 14600 483574 14612
rect 483970 14600 483976 14612
rect 483568 14572 483976 14600
rect 483568 14560 483574 14572
rect 483970 14560 483976 14572
rect 484028 14560 484034 14612
rect 246058 14492 246064 14544
rect 246116 14532 246122 14544
rect 264734 14532 264740 14544
rect 246116 14504 264740 14532
rect 246116 14492 246122 14504
rect 264734 14492 264740 14504
rect 264792 14492 264798 14544
rect 252958 14424 252964 14476
rect 253016 14464 253022 14476
rect 282214 14464 282220 14476
rect 253016 14436 282220 14464
rect 253016 14424 253022 14436
rect 282214 14424 282220 14436
rect 282272 14424 282278 14476
rect 303374 14424 303380 14476
rect 303432 14464 303438 14476
rect 322050 14464 322056 14476
rect 303432 14436 322056 14464
rect 303432 14424 303438 14436
rect 322050 14424 322056 14436
rect 322108 14424 322114 14476
rect 1600 14096 583316 14192
rect 1600 13552 583316 13648
rect 1600 13008 583316 13104
rect 1600 12464 583316 12560
rect 114958 12384 114964 12436
rect 115016 12424 115022 12436
rect 253326 12424 253332 12436
rect 115016 12396 253332 12424
rect 115016 12384 115022 12396
rect 253326 12384 253332 12396
rect 253384 12384 253390 12436
rect 332906 12384 332912 12436
rect 332964 12424 332970 12436
rect 493170 12424 493176 12436
rect 332964 12396 493176 12424
rect 332964 12384 332970 12396
rect 493170 12384 493176 12396
rect 493228 12384 493234 12436
rect 513870 12384 513876 12436
rect 513928 12424 513934 12436
rect 514882 12424 514888 12436
rect 513928 12396 514888 12424
rect 513928 12384 513934 12396
rect 514882 12384 514888 12396
rect 514940 12384 514946 12436
rect 530430 12384 530436 12436
rect 530488 12424 530494 12436
rect 531534 12424 531540 12436
rect 530488 12396 531540 12424
rect 530488 12384 530494 12396
rect 531534 12384 531540 12396
rect 531592 12384 531598 12436
rect 534570 12384 534576 12436
rect 534628 12424 534634 12436
rect 535030 12424 535036 12436
rect 534628 12396 535036 12424
rect 534628 12384 534634 12396
rect 535030 12384 535036 12396
rect 535088 12384 535094 12436
rect 542850 12384 542856 12436
rect 542908 12424 542914 12436
rect 543402 12424 543408 12436
rect 542908 12396 543408 12424
rect 542908 12384 542914 12396
rect 543402 12384 543408 12396
rect 543460 12384 543466 12436
rect 548370 12384 548376 12436
rect 548428 12424 548434 12436
rect 549382 12424 549388 12436
rect 548428 12396 549388 12424
rect 548428 12384 548434 12396
rect 549382 12384 549388 12396
rect 549440 12384 549446 12436
rect 549750 12384 549756 12436
rect 549808 12424 549814 12436
rect 550578 12424 550584 12436
rect 549808 12396 550584 12424
rect 549808 12384 549814 12396
rect 550578 12384 550584 12396
rect 550636 12384 550642 12436
rect 556650 12384 556656 12436
rect 556708 12424 556714 12436
rect 557662 12424 557668 12436
rect 556708 12396 557668 12424
rect 556708 12384 556714 12396
rect 557662 12384 557668 12396
rect 557720 12384 557726 12436
rect 567690 12384 567696 12436
rect 567748 12424 567754 12436
rect 568334 12424 568340 12436
rect 567748 12396 568340 12424
rect 567748 12384 567754 12396
rect 568334 12384 568340 12396
rect 568392 12384 568398 12436
rect 574590 12384 574596 12436
rect 574648 12424 574654 12436
rect 575510 12424 575516 12436
rect 574648 12396 575516 12424
rect 574648 12384 574654 12396
rect 575510 12384 575516 12396
rect 575568 12384 575574 12436
rect 575970 12384 575976 12436
rect 576028 12424 576034 12436
rect 576706 12424 576712 12436
rect 576028 12396 576712 12424
rect 576028 12384 576034 12396
rect 576706 12384 576712 12396
rect 576764 12384 576770 12436
rect 107966 12316 107972 12368
rect 108024 12356 108030 12368
rect 251946 12356 251952 12368
rect 108024 12328 251952 12356
rect 108024 12316 108030 12328
rect 251946 12316 251952 12328
rect 252004 12316 252010 12368
rect 332814 12316 332820 12368
rect 332872 12356 332878 12368
rect 495930 12356 495936 12368
rect 332872 12328 495936 12356
rect 332872 12316 332878 12328
rect 495930 12316 495936 12328
rect 495988 12316 495994 12368
rect 99502 12248 99508 12300
rect 99560 12288 99566 12300
rect 250474 12288 250480 12300
rect 99560 12260 250480 12288
rect 99560 12248 99566 12260
rect 250474 12248 250480 12260
rect 250532 12248 250538 12300
rect 334194 12248 334200 12300
rect 334252 12288 334258 12300
rect 500070 12288 500076 12300
rect 334252 12260 500076 12288
rect 334252 12248 334258 12260
rect 500070 12248 500076 12260
rect 500128 12248 500134 12300
rect 92602 12180 92608 12232
rect 92660 12220 92666 12232
rect 249278 12220 249284 12232
rect 92660 12192 249284 12220
rect 92660 12180 92666 12192
rect 249278 12180 249284 12192
rect 249336 12180 249342 12232
rect 334102 12180 334108 12232
rect 334160 12220 334166 12232
rect 504118 12220 504124 12232
rect 334160 12192 504124 12220
rect 334160 12180 334166 12192
rect 504118 12180 504124 12192
rect 504176 12180 504182 12232
rect 85978 12112 85984 12164
rect 86036 12152 86042 12164
rect 248174 12152 248180 12164
rect 86036 12124 248180 12152
rect 86036 12112 86042 12124
rect 248174 12112 248180 12124
rect 248232 12112 248238 12164
rect 335482 12112 335488 12164
rect 335540 12152 335546 12164
rect 511294 12152 511300 12164
rect 335540 12124 511300 12152
rect 335540 12112 335546 12124
rect 511294 12112 511300 12124
rect 511352 12112 511358 12164
rect 83126 12044 83132 12096
rect 83184 12084 83190 12096
rect 246702 12084 246708 12096
rect 83184 12056 246708 12084
rect 83184 12044 83190 12056
rect 246702 12044 246708 12056
rect 246760 12044 246766 12096
rect 336862 12044 336868 12096
rect 336920 12084 336926 12096
rect 518378 12084 518384 12096
rect 336920 12056 518384 12084
rect 336920 12044 336926 12056
rect 518378 12044 518384 12056
rect 518436 12044 518442 12096
rect 1600 11920 583316 12016
rect 79078 11840 79084 11892
rect 79136 11880 79142 11892
rect 246242 11880 246248 11892
rect 79136 11852 246248 11880
rect 79136 11840 79142 11852
rect 246242 11840 246248 11852
rect 246300 11840 246306 11892
rect 338150 11840 338156 11892
rect 338208 11880 338214 11892
rect 525554 11880 525560 11892
rect 338208 11852 525560 11880
rect 338208 11840 338214 11852
rect 525554 11840 525560 11852
rect 525612 11840 525618 11892
rect 74938 11772 74944 11824
rect 74996 11812 75002 11824
rect 244862 11812 244868 11824
rect 74996 11784 244868 11812
rect 74996 11772 75002 11784
rect 244862 11772 244868 11784
rect 244920 11772 244926 11824
rect 295554 11772 295560 11824
rect 295612 11812 295618 11824
rect 316162 11812 316168 11824
rect 295612 11784 316168 11812
rect 295612 11772 295618 11784
rect 316162 11772 316168 11784
rect 316220 11772 316226 11824
rect 339622 11772 339628 11824
rect 339680 11812 339686 11824
rect 532730 11812 532736 11824
rect 339680 11784 532736 11812
rect 339680 11772 339686 11784
rect 532730 11772 532736 11784
rect 532788 11772 532794 11824
rect 72178 11704 72184 11756
rect 72236 11744 72242 11756
rect 244954 11744 244960 11756
rect 72236 11716 244960 11744
rect 72236 11704 72242 11716
rect 244954 11704 244960 11716
rect 245012 11704 245018 11756
rect 248818 11704 248824 11756
rect 248876 11744 248882 11756
rect 281294 11744 281300 11756
rect 248876 11716 281300 11744
rect 248876 11704 248882 11716
rect 281294 11704 281300 11716
rect 281352 11704 281358 11756
rect 304754 11704 304760 11756
rect 304812 11744 304818 11756
rect 324810 11744 324816 11756
rect 304812 11716 324816 11744
rect 304812 11704 304818 11716
rect 324810 11704 324816 11716
rect 324868 11704 324874 11756
rect 342474 11704 342480 11756
rect 342532 11744 342538 11756
rect 539814 11744 539820 11756
rect 342532 11716 539820 11744
rect 342532 11704 342538 11716
rect 539814 11704 539820 11716
rect 539872 11704 539878 11756
rect 331342 11636 331348 11688
rect 331400 11676 331406 11688
rect 489858 11676 489864 11688
rect 331400 11648 489864 11676
rect 331400 11636 331406 11648
rect 489858 11636 489864 11648
rect 489916 11636 489922 11688
rect 1600 11376 583316 11472
rect 176693 11339 176751 11345
rect 176693 11305 176705 11339
rect 176739 11336 176751 11339
rect 179177 11339 179235 11345
rect 179177 11336 179189 11339
rect 176739 11308 179189 11336
rect 176739 11305 176751 11308
rect 176693 11299 176751 11305
rect 179177 11305 179189 11308
rect 179223 11305 179235 11339
rect 179177 11299 179235 11305
rect 331437 11339 331495 11345
rect 331437 11305 331449 11339
rect 331483 11336 331495 11339
rect 333737 11339 333795 11345
rect 333737 11336 333749 11339
rect 331483 11308 333749 11336
rect 331483 11305 331495 11308
rect 331437 11299 331495 11305
rect 333737 11305 333749 11308
rect 333783 11305 333795 11339
rect 333737 11299 333795 11305
rect 340913 11339 340971 11345
rect 340913 11305 340925 11339
rect 340959 11336 340971 11339
rect 340959 11308 343164 11336
rect 340959 11305 340971 11308
rect 340913 11299 340971 11305
rect 234745 11271 234803 11277
rect 234745 11237 234757 11271
rect 234791 11268 234803 11271
rect 235294 11268 235300 11280
rect 234791 11240 235300 11268
rect 234791 11237 234803 11240
rect 234745 11231 234803 11237
rect 235294 11228 235300 11240
rect 235352 11228 235358 11280
rect 331529 11271 331587 11277
rect 331529 11237 331541 11271
rect 331575 11268 331587 11271
rect 341281 11271 341339 11277
rect 341281 11268 341293 11271
rect 331575 11240 341293 11268
rect 331575 11237 331587 11240
rect 331529 11231 331587 11237
rect 341281 11237 341293 11240
rect 341327 11237 341339 11271
rect 341281 11231 341339 11237
rect 129037 11203 129095 11209
rect 129037 11200 129049 11203
rect 123532 11172 129049 11200
rect 117626 11092 117632 11144
rect 117684 11132 117690 11144
rect 123532 11132 123560 11172
rect 129037 11169 129049 11172
rect 129083 11169 129095 11203
rect 129037 11163 129095 11169
rect 148265 11203 148323 11209
rect 148265 11169 148277 11203
rect 148311 11200 148323 11203
rect 157741 11203 157799 11209
rect 157741 11200 157753 11203
rect 148311 11172 157753 11200
rect 148311 11169 148323 11172
rect 148265 11163 148323 11169
rect 157741 11169 157753 11172
rect 157787 11169 157799 11203
rect 157741 11163 157799 11169
rect 167582 11160 167588 11212
rect 167640 11200 167646 11212
rect 177061 11203 177119 11209
rect 177061 11200 177073 11203
rect 167640 11172 177073 11200
rect 167640 11160 167646 11172
rect 177061 11169 177073 11172
rect 177107 11169 177119 11203
rect 177061 11163 177119 11169
rect 215974 11160 215980 11212
rect 216032 11200 216038 11212
rect 238333 11203 238391 11209
rect 238333 11200 238345 11203
rect 216032 11172 238345 11200
rect 216032 11160 216038 11172
rect 238333 11169 238345 11172
rect 238379 11169 238391 11203
rect 238333 11163 238391 11169
rect 331253 11203 331311 11209
rect 331253 11169 331265 11203
rect 331299 11200 331311 11203
rect 341005 11203 341063 11209
rect 341005 11200 341017 11203
rect 331299 11172 341017 11200
rect 331299 11169 331311 11172
rect 331253 11163 331311 11169
rect 341005 11169 341017 11172
rect 341051 11169 341063 11203
rect 341462 11200 341468 11212
rect 341005 11163 341063 11169
rect 341112 11172 341468 11200
rect 128945 11135 129003 11141
rect 128945 11132 128957 11135
rect 117684 11104 123560 11132
rect 125188 11104 128957 11132
rect 117684 11092 117690 11104
rect 123333 11067 123391 11073
rect 123333 11033 123345 11067
rect 123379 11064 123391 11067
rect 125188 11064 125216 11104
rect 128945 11101 128957 11104
rect 128991 11101 129003 11135
rect 138237 11135 138295 11141
rect 138237 11132 138249 11135
rect 128945 11095 129003 11101
rect 129144 11104 138249 11132
rect 129144 11064 129172 11104
rect 138237 11101 138249 11104
rect 138283 11101 138295 11135
rect 138237 11095 138295 11101
rect 147897 11135 147955 11141
rect 147897 11101 147909 11135
rect 147943 11132 147955 11135
rect 148357 11135 148415 11141
rect 148357 11132 148369 11135
rect 147943 11104 148369 11132
rect 147943 11101 147955 11104
rect 147897 11095 147955 11101
rect 148357 11101 148369 11104
rect 148403 11101 148415 11135
rect 148357 11095 148415 11101
rect 176877 11135 176935 11141
rect 176877 11101 176889 11135
rect 176923 11132 176935 11135
rect 177242 11132 177248 11144
rect 176923 11104 177248 11132
rect 176923 11101 176935 11104
rect 176877 11095 176935 11101
rect 177242 11092 177248 11104
rect 177300 11092 177306 11144
rect 179177 11135 179235 11141
rect 179177 11101 179189 11135
rect 179223 11132 179235 11135
rect 186997 11135 187055 11141
rect 186997 11132 187009 11135
rect 179223 11104 187009 11132
rect 179223 11101 179235 11104
rect 179177 11095 179235 11101
rect 186997 11101 187009 11104
rect 187043 11101 187055 11135
rect 186997 11095 187055 11101
rect 225545 11135 225603 11141
rect 225545 11101 225557 11135
rect 225591 11132 225603 11135
rect 331897 11135 331955 11141
rect 331897 11132 331909 11135
rect 225591 11104 236904 11132
rect 225591 11101 225603 11104
rect 225545 11095 225603 11101
rect 133821 11067 133879 11073
rect 133821 11064 133833 11067
rect 123379 11036 125216 11064
rect 128960 11036 129172 11064
rect 133560 11036 133833 11064
rect 123379 11033 123391 11036
rect 123333 11027 123391 11033
rect 56906 10956 56912 11008
rect 56964 10996 56970 11008
rect 128960 10996 128988 11036
rect 56964 10968 128988 10996
rect 129037 10999 129095 11005
rect 56964 10956 56970 10968
rect 129037 10965 129049 10999
rect 129083 10996 129095 10999
rect 133560 10996 133588 11036
rect 133821 11033 133833 11036
rect 133867 11033 133879 11067
rect 133821 11027 133879 11033
rect 138513 11067 138571 11073
rect 138513 11033 138525 11067
rect 138559 11064 138571 11067
rect 148081 11067 148139 11073
rect 148081 11064 148093 11067
rect 138559 11036 148093 11064
rect 138559 11033 138571 11036
rect 138513 11027 138571 11033
rect 148081 11033 148093 11036
rect 148127 11033 148139 11067
rect 148081 11027 148139 11033
rect 148173 11067 148231 11073
rect 148173 11033 148185 11067
rect 148219 11064 148231 11067
rect 157649 11067 157707 11073
rect 157649 11064 157661 11067
rect 148219 11036 157661 11064
rect 148219 11033 148231 11036
rect 148173 11027 148231 11033
rect 157649 11033 157661 11036
rect 157695 11033 157707 11067
rect 157649 11027 157707 11033
rect 157833 11067 157891 11073
rect 157833 11033 157845 11067
rect 157879 11064 157891 11067
rect 167490 11064 167496 11076
rect 157879 11036 167496 11064
rect 157879 11033 157891 11036
rect 157833 11027 157891 11033
rect 167490 11024 167496 11036
rect 167548 11024 167554 11076
rect 167585 11067 167643 11073
rect 167585 11033 167597 11067
rect 167631 11064 167643 11067
rect 176785 11067 176843 11073
rect 176785 11064 176797 11067
rect 167631 11036 176797 11064
rect 167631 11033 167643 11036
rect 167585 11027 167643 11033
rect 176785 11033 176797 11036
rect 176831 11033 176843 11067
rect 176785 11027 176843 11033
rect 186905 11067 186963 11073
rect 186905 11033 186917 11067
rect 186951 11064 186963 11067
rect 196197 11067 196255 11073
rect 196197 11064 196209 11067
rect 186951 11036 196209 11064
rect 186951 11033 186963 11036
rect 186905 11027 186963 11033
rect 196197 11033 196209 11036
rect 196243 11033 196255 11067
rect 196197 11027 196255 11033
rect 196565 11067 196623 11073
rect 196565 11033 196577 11067
rect 196611 11064 196623 11067
rect 215790 11064 215796 11076
rect 196611 11036 215796 11064
rect 196611 11033 196623 11036
rect 196565 11027 196623 11033
rect 215790 11024 215796 11036
rect 215848 11024 215854 11076
rect 234926 11024 234932 11076
rect 234984 11064 234990 11076
rect 235481 11067 235539 11073
rect 235481 11064 235493 11067
rect 234984 11036 235493 11064
rect 234984 11024 234990 11036
rect 235481 11033 235493 11036
rect 235527 11033 235539 11067
rect 235481 11027 235539 11033
rect 129083 10968 133588 10996
rect 133637 10999 133695 11005
rect 129083 10965 129095 10968
rect 129037 10959 129095 10965
rect 133637 10965 133649 10999
rect 133683 10996 133695 10999
rect 236766 10996 236772 11008
rect 133683 10968 236772 10996
rect 133683 10965 133695 10968
rect 133637 10959 133695 10965
rect 236766 10956 236772 10968
rect 236824 10956 236830 11008
rect 236876 10996 236904 11104
rect 331544 11104 331909 11132
rect 331342 11064 331348 11076
rect 328140 11036 331348 11064
rect 242286 10996 242292 11008
rect 236876 10968 242292 10996
rect 242286 10956 242292 10968
rect 242344 10956 242350 11008
rect 323154 10956 323160 11008
rect 323212 10996 323218 11008
rect 328140 10996 328168 11036
rect 331342 11024 331348 11036
rect 331400 11024 331406 11076
rect 323212 10968 328168 10996
rect 323212 10956 323218 10968
rect 328398 10956 328404 11008
rect 328456 10996 328462 11008
rect 331544 10996 331572 11104
rect 331897 11101 331909 11104
rect 331943 11101 331955 11135
rect 341112 11132 341140 11172
rect 341462 11160 341468 11172
rect 341520 11160 341526 11212
rect 331897 11095 331955 11101
rect 332004 11104 341140 11132
rect 343136 11132 343164 11308
rect 348086 11228 348092 11280
rect 348144 11268 348150 11280
rect 350941 11271 350999 11277
rect 350941 11268 350953 11271
rect 348144 11240 350953 11268
rect 348144 11228 348150 11240
rect 350941 11237 350953 11240
rect 350987 11237 350999 11271
rect 350941 11231 350999 11237
rect 346522 11160 346528 11212
rect 346580 11200 346586 11212
rect 351309 11203 351367 11209
rect 351309 11200 351321 11203
rect 346580 11172 351321 11200
rect 346580 11160 346586 11172
rect 351309 11169 351321 11172
rect 351355 11169 351367 11203
rect 351309 11163 351367 11169
rect 408990 11160 408996 11212
rect 409048 11200 409054 11212
rect 410186 11200 410192 11212
rect 409048 11172 410192 11200
rect 409048 11160 409054 11172
rect 410186 11160 410192 11172
rect 410244 11160 410250 11212
rect 409085 11135 409143 11141
rect 409085 11132 409097 11135
rect 343136 11104 409097 11132
rect 331713 11067 331771 11073
rect 331713 11033 331725 11067
rect 331759 11064 331771 11067
rect 332004 11064 332032 11104
rect 409085 11101 409097 11104
rect 409131 11101 409143 11135
rect 409085 11095 409143 11101
rect 418469 11135 418527 11141
rect 418469 11101 418481 11135
rect 418515 11132 418527 11135
rect 418745 11135 418803 11141
rect 418745 11132 418757 11135
rect 418515 11104 418757 11132
rect 418515 11101 418527 11104
rect 418469 11095 418527 11101
rect 418745 11101 418757 11104
rect 418791 11101 418803 11135
rect 418745 11095 418803 11101
rect 331759 11036 332032 11064
rect 341097 11067 341155 11073
rect 331759 11033 331771 11036
rect 331713 11027 331771 11033
rect 341097 11033 341109 11067
rect 341143 11064 341155 11067
rect 418561 11067 418619 11073
rect 418561 11064 418573 11067
rect 341143 11036 418573 11064
rect 341143 11033 341155 11036
rect 341097 11027 341155 11033
rect 418561 11033 418573 11036
rect 418607 11033 418619 11067
rect 418561 11027 418619 11033
rect 328456 10968 331572 10996
rect 333737 10999 333795 11005
rect 328456 10956 328462 10968
rect 333737 10965 333749 10999
rect 333783 10996 333795 10999
rect 460142 10996 460148 11008
rect 333783 10968 460148 10996
rect 333783 10965 333795 10968
rect 333737 10959 333795 10965
rect 460142 10956 460148 10968
rect 460200 10956 460206 11008
rect 1600 10832 583316 10928
rect 53318 10752 53324 10804
rect 53376 10792 53382 10804
rect 128853 10795 128911 10801
rect 128853 10792 128865 10795
rect 53376 10764 128865 10792
rect 53376 10752 53382 10764
rect 128853 10761 128865 10764
rect 128899 10761 128911 10795
rect 128853 10755 128911 10761
rect 128945 10795 129003 10801
rect 128945 10761 128957 10795
rect 128991 10792 129003 10795
rect 147802 10792 147808 10804
rect 128991 10764 147808 10792
rect 128991 10761 129003 10764
rect 128945 10755 129003 10761
rect 147802 10752 147808 10764
rect 147860 10752 147866 10804
rect 148081 10795 148139 10801
rect 148081 10761 148093 10795
rect 148127 10792 148139 10795
rect 148265 10795 148323 10801
rect 148265 10792 148277 10795
rect 148127 10764 148277 10792
rect 148127 10761 148139 10764
rect 148081 10755 148139 10761
rect 148265 10761 148277 10764
rect 148311 10761 148323 10795
rect 148265 10755 148323 10761
rect 148446 10752 148452 10804
rect 148504 10792 148510 10804
rect 153046 10792 153052 10804
rect 148504 10764 153052 10792
rect 148504 10752 148510 10764
rect 153046 10752 153052 10764
rect 153104 10752 153110 10804
rect 153141 10795 153199 10801
rect 153141 10761 153153 10795
rect 153187 10792 153199 10795
rect 176693 10795 176751 10801
rect 176693 10792 176705 10795
rect 153187 10764 176705 10792
rect 153187 10761 153199 10764
rect 153141 10755 153199 10761
rect 176693 10761 176705 10764
rect 176739 10761 176751 10795
rect 176693 10755 176751 10761
rect 177061 10795 177119 10801
rect 177061 10761 177073 10795
rect 177107 10792 177119 10795
rect 186905 10795 186963 10801
rect 186905 10792 186917 10795
rect 177107 10764 186917 10792
rect 177107 10761 177119 10764
rect 177061 10755 177119 10761
rect 186905 10761 186917 10764
rect 186951 10761 186963 10795
rect 186905 10755 186963 10761
rect 187086 10752 187092 10804
rect 187144 10792 187150 10804
rect 191686 10792 191692 10804
rect 187144 10764 191692 10792
rect 187144 10752 187150 10764
rect 191686 10752 191692 10764
rect 191744 10752 191750 10804
rect 191781 10795 191839 10801
rect 191781 10761 191793 10795
rect 191827 10792 191839 10795
rect 230053 10795 230111 10801
rect 230053 10792 230065 10795
rect 191827 10764 230065 10792
rect 191827 10761 191839 10764
rect 191781 10755 191839 10761
rect 230053 10761 230065 10764
rect 230099 10761 230111 10795
rect 230053 10755 230111 10761
rect 230145 10795 230203 10801
rect 230145 10761 230157 10795
rect 230191 10792 230203 10795
rect 234650 10792 234656 10804
rect 230191 10764 234656 10792
rect 230191 10761 230203 10764
rect 230145 10755 230203 10761
rect 234650 10752 234656 10764
rect 234708 10752 234714 10804
rect 235018 10752 235024 10804
rect 235076 10792 235082 10804
rect 235389 10795 235447 10801
rect 235389 10792 235401 10795
rect 235076 10764 235401 10792
rect 235076 10752 235082 10764
rect 235389 10761 235401 10764
rect 235435 10761 235447 10795
rect 235389 10755 235447 10761
rect 235481 10795 235539 10801
rect 235481 10761 235493 10795
rect 235527 10792 235539 10795
rect 238146 10792 238152 10804
rect 235527 10764 238152 10792
rect 235527 10761 235539 10764
rect 235481 10755 235539 10761
rect 238146 10752 238152 10764
rect 238204 10752 238210 10804
rect 238514 10752 238520 10804
rect 238572 10792 238578 10804
rect 244126 10792 244132 10804
rect 238572 10764 244132 10792
rect 238572 10752 238578 10764
rect 244126 10752 244132 10764
rect 244184 10752 244190 10804
rect 327202 10752 327208 10804
rect 327260 10792 327266 10804
rect 331529 10795 331587 10801
rect 331529 10792 331541 10795
rect 327260 10764 331541 10792
rect 327260 10752 327266 10764
rect 331529 10761 331541 10764
rect 331575 10761 331587 10795
rect 331529 10755 331587 10761
rect 331621 10795 331679 10801
rect 331621 10761 331633 10795
rect 331667 10792 331679 10795
rect 462810 10792 462816 10804
rect 331667 10764 462816 10792
rect 331667 10761 331679 10764
rect 331621 10755 331679 10761
rect 462810 10752 462816 10764
rect 462868 10752 462874 10804
rect 50098 10684 50104 10736
rect 50156 10724 50162 10736
rect 133545 10727 133603 10733
rect 133545 10724 133557 10727
rect 50156 10696 133557 10724
rect 50156 10684 50162 10696
rect 133545 10693 133557 10696
rect 133591 10693 133603 10727
rect 143297 10727 143355 10733
rect 143297 10724 143309 10727
rect 133545 10687 133603 10693
rect 133652 10696 143309 10724
rect 45958 10616 45964 10668
rect 46016 10656 46022 10668
rect 133652 10656 133680 10696
rect 143297 10693 143309 10696
rect 143343 10693 143355 10727
rect 147897 10727 147955 10733
rect 147897 10724 147909 10727
rect 143297 10687 143355 10693
rect 143404 10696 147909 10724
rect 46016 10628 133680 10656
rect 133729 10659 133787 10665
rect 46016 10616 46022 10628
rect 133729 10625 133741 10659
rect 133775 10656 133787 10659
rect 143404 10656 143432 10696
rect 147897 10693 147909 10696
rect 147943 10693 147955 10727
rect 147897 10687 147955 10693
rect 147989 10727 148047 10733
rect 147989 10693 148001 10727
rect 148035 10724 148047 10727
rect 148173 10727 148231 10733
rect 148173 10724 148185 10727
rect 148035 10696 148185 10724
rect 148035 10693 148047 10696
rect 147989 10687 148047 10693
rect 148173 10693 148185 10696
rect 148219 10693 148231 10727
rect 148173 10687 148231 10693
rect 148357 10727 148415 10733
rect 148357 10693 148369 10727
rect 148403 10724 148415 10727
rect 152865 10727 152923 10733
rect 152865 10724 152877 10727
rect 148403 10696 152877 10724
rect 148403 10693 148415 10696
rect 148357 10687 148415 10693
rect 152865 10693 152877 10696
rect 152911 10693 152923 10727
rect 172369 10727 172427 10733
rect 152865 10687 152923 10693
rect 152972 10696 172320 10724
rect 133775 10628 143432 10656
rect 143481 10659 143539 10665
rect 133775 10625 133787 10628
rect 133729 10619 133787 10625
rect 143481 10625 143493 10659
rect 143527 10656 143539 10659
rect 152972 10656 153000 10696
rect 143527 10628 153000 10656
rect 143527 10625 143539 10628
rect 143481 10619 143539 10625
rect 153046 10616 153052 10668
rect 153104 10656 153110 10668
rect 172185 10659 172243 10665
rect 172185 10656 172197 10659
rect 153104 10628 172197 10656
rect 153104 10616 153110 10628
rect 172185 10625 172197 10628
rect 172231 10625 172243 10659
rect 172292 10656 172320 10696
rect 172369 10693 172381 10727
rect 172415 10724 172427 10727
rect 176877 10727 176935 10733
rect 176877 10724 176889 10727
rect 172415 10696 176889 10724
rect 172415 10693 172427 10696
rect 172369 10687 172427 10693
rect 176877 10693 176889 10696
rect 176923 10693 176935 10727
rect 176877 10687 176935 10693
rect 176969 10727 177027 10733
rect 176969 10693 176981 10727
rect 177015 10724 177027 10727
rect 186810 10724 186816 10736
rect 177015 10696 186816 10724
rect 177015 10693 177027 10696
rect 176969 10687 177027 10693
rect 186810 10684 186816 10696
rect 186868 10684 186874 10736
rect 186997 10727 187055 10733
rect 186997 10693 187009 10727
rect 187043 10724 187055 10727
rect 191505 10727 191563 10733
rect 191505 10724 191517 10727
rect 187043 10696 191517 10724
rect 187043 10693 187055 10696
rect 186997 10687 187055 10693
rect 191505 10693 191517 10696
rect 191551 10693 191563 10727
rect 230329 10727 230387 10733
rect 191505 10687 191563 10693
rect 191612 10696 230280 10724
rect 191612 10656 191640 10696
rect 172292 10628 191640 10656
rect 172185 10619 172243 10625
rect 191686 10616 191692 10668
rect 191744 10656 191750 10668
rect 230145 10659 230203 10665
rect 230145 10656 230157 10659
rect 191744 10628 230157 10656
rect 191744 10616 191750 10628
rect 230145 10625 230157 10628
rect 230191 10625 230203 10659
rect 230252 10656 230280 10696
rect 230329 10693 230341 10727
rect 230375 10724 230387 10727
rect 234834 10724 234840 10736
rect 230375 10696 234840 10724
rect 230375 10693 230387 10696
rect 230329 10687 230387 10693
rect 234834 10684 234840 10696
rect 234892 10684 234898 10736
rect 234929 10727 234987 10733
rect 234929 10693 234941 10727
rect 234975 10724 234987 10727
rect 235113 10727 235171 10733
rect 235113 10724 235125 10727
rect 234975 10696 235125 10724
rect 234975 10693 234987 10696
rect 234929 10687 234987 10693
rect 235113 10693 235125 10696
rect 235159 10693 235171 10727
rect 239250 10724 239256 10736
rect 235113 10687 235171 10693
rect 235220 10696 239256 10724
rect 235220 10656 235248 10696
rect 239250 10684 239256 10696
rect 239308 10684 239314 10736
rect 323062 10684 323068 10736
rect 323120 10724 323126 10736
rect 328398 10724 328404 10736
rect 323120 10696 328404 10724
rect 323120 10684 323126 10696
rect 328398 10684 328404 10696
rect 328456 10684 328462 10736
rect 328490 10684 328496 10736
rect 328548 10724 328554 10736
rect 331897 10727 331955 10733
rect 328548 10696 331848 10724
rect 328548 10684 328554 10696
rect 230252 10628 235248 10656
rect 230145 10619 230203 10625
rect 235386 10616 235392 10668
rect 235444 10656 235450 10668
rect 238238 10656 238244 10668
rect 235444 10628 238244 10656
rect 235444 10616 235450 10628
rect 238238 10616 238244 10628
rect 238296 10616 238302 10668
rect 238333 10659 238391 10665
rect 238333 10625 238345 10659
rect 238379 10656 238391 10659
rect 243758 10656 243764 10668
rect 238379 10628 243764 10656
rect 238379 10625 238391 10628
rect 238333 10619 238391 10625
rect 243758 10616 243764 10628
rect 243816 10616 243822 10668
rect 324442 10616 324448 10668
rect 324500 10656 324506 10668
rect 329870 10656 329876 10668
rect 324500 10628 329876 10656
rect 324500 10616 324506 10628
rect 329870 10616 329876 10628
rect 329928 10616 329934 10668
rect 329962 10616 329968 10668
rect 330020 10656 330026 10668
rect 331713 10659 331771 10665
rect 331713 10656 331725 10659
rect 330020 10628 331725 10656
rect 330020 10616 330026 10628
rect 331713 10625 331725 10628
rect 331759 10625 331771 10659
rect 331820 10656 331848 10696
rect 331897 10693 331909 10727
rect 331943 10724 331955 10727
rect 340913 10727 340971 10733
rect 340913 10724 340925 10727
rect 331943 10696 340925 10724
rect 331943 10693 331955 10696
rect 331897 10687 331955 10693
rect 340913 10693 340925 10696
rect 340959 10693 340971 10727
rect 340913 10687 340971 10693
rect 341281 10727 341339 10733
rect 341281 10693 341293 10727
rect 341327 10724 341339 10727
rect 466950 10724 466956 10736
rect 341327 10696 466956 10724
rect 341327 10693 341339 10696
rect 341281 10687 341339 10693
rect 466950 10684 466956 10696
rect 467008 10684 467014 10736
rect 341097 10659 341155 10665
rect 341097 10656 341109 10659
rect 331820 10628 341109 10656
rect 331713 10619 331771 10625
rect 341097 10625 341109 10628
rect 341143 10625 341155 10659
rect 341097 10619 341155 10625
rect 341189 10659 341247 10665
rect 341189 10625 341201 10659
rect 341235 10656 341247 10659
rect 469710 10656 469716 10668
rect 341235 10628 469716 10656
rect 341235 10625 341247 10628
rect 341189 10619 341247 10625
rect 469710 10616 469716 10628
rect 469768 10616 469774 10668
rect 41818 10548 41824 10600
rect 41876 10588 41882 10600
rect 41876 10560 123468 10588
rect 41876 10548 41882 10560
rect 39058 10480 39064 10532
rect 39116 10520 39122 10532
rect 123333 10523 123391 10529
rect 123333 10520 123345 10523
rect 39116 10492 123345 10520
rect 39116 10480 39122 10492
rect 123333 10489 123345 10492
rect 123379 10489 123391 10523
rect 123440 10520 123468 10560
rect 123514 10548 123520 10600
rect 123572 10588 123578 10600
rect 254982 10588 254988 10600
rect 123572 10560 254988 10588
rect 123572 10548 123578 10560
rect 254982 10548 254988 10560
rect 255040 10548 255046 10600
rect 318830 10548 318836 10600
rect 318888 10588 318894 10600
rect 418653 10591 418711 10597
rect 418653 10588 418665 10591
rect 318888 10560 418665 10588
rect 318888 10548 318894 10560
rect 418653 10557 418665 10560
rect 418699 10557 418711 10591
rect 418653 10551 418711 10557
rect 418745 10591 418803 10597
rect 418745 10557 418757 10591
rect 418791 10588 418803 10591
rect 423345 10591 423403 10597
rect 423345 10588 423357 10591
rect 418791 10560 423357 10588
rect 418791 10557 418803 10560
rect 418745 10551 418803 10557
rect 423345 10557 423357 10560
rect 423391 10557 423403 10591
rect 474402 10588 474408 10600
rect 423345 10551 423403 10557
rect 423452 10560 474408 10588
rect 133729 10523 133787 10529
rect 133729 10520 133741 10523
rect 123440 10492 133741 10520
rect 123333 10483 123391 10489
rect 133729 10489 133741 10492
rect 133775 10489 133787 10523
rect 133729 10483 133787 10489
rect 133913 10523 133971 10529
rect 133913 10489 133925 10523
rect 133959 10520 133971 10523
rect 138329 10523 138387 10529
rect 138329 10520 138341 10523
rect 133959 10492 138341 10520
rect 133959 10489 133971 10492
rect 133913 10483 133971 10489
rect 138329 10489 138341 10492
rect 138375 10489 138387 10523
rect 138329 10483 138387 10489
rect 138418 10480 138424 10532
rect 138476 10520 138482 10532
rect 254614 10520 254620 10532
rect 138476 10492 254620 10520
rect 138476 10480 138482 10492
rect 254614 10480 254620 10492
rect 254672 10480 254678 10532
rect 317542 10480 317548 10532
rect 317600 10520 317606 10532
rect 408990 10520 408996 10532
rect 317600 10492 408996 10520
rect 317600 10480 317606 10492
rect 408990 10480 408996 10492
rect 409048 10480 409054 10532
rect 409085 10523 409143 10529
rect 409085 10489 409097 10523
rect 409131 10520 409143 10523
rect 418469 10523 418527 10529
rect 418469 10520 418481 10523
rect 409131 10492 418481 10520
rect 409131 10489 409143 10492
rect 409085 10483 409143 10489
rect 418469 10489 418481 10492
rect 418515 10489 418527 10523
rect 418469 10483 418527 10489
rect 418561 10523 418619 10529
rect 418561 10489 418573 10523
rect 418607 10520 418619 10523
rect 423452 10520 423480 10560
rect 474402 10548 474408 10560
rect 474460 10548 474466 10600
rect 418607 10492 423480 10520
rect 423529 10523 423587 10529
rect 418607 10489 418619 10492
rect 418561 10483 418619 10489
rect 423529 10489 423541 10523
rect 423575 10520 423587 10523
rect 477990 10520 477996 10532
rect 423575 10492 477996 10520
rect 423575 10489 423587 10492
rect 423529 10483 423587 10489
rect 477990 10480 477996 10492
rect 478048 10480 478054 10532
rect 34918 10412 34924 10464
rect 34976 10452 34982 10464
rect 133637 10455 133695 10461
rect 133637 10452 133649 10455
rect 34976 10424 133649 10452
rect 34976 10412 34982 10424
rect 133637 10421 133649 10424
rect 133683 10421 133695 10455
rect 133637 10415 133695 10421
rect 133821 10455 133879 10461
rect 133821 10421 133833 10455
rect 133867 10452 133879 10455
rect 253142 10452 253148 10464
rect 133867 10424 253148 10452
rect 133867 10421 133879 10424
rect 133821 10415 133879 10421
rect 253142 10412 253148 10424
rect 253200 10412 253206 10464
rect 255718 10412 255724 10464
rect 255776 10452 255782 10464
rect 282490 10452 282496 10464
rect 255776 10424 282496 10452
rect 255776 10412 255782 10424
rect 282490 10412 282496 10424
rect 282548 10412 282554 10464
rect 318646 10412 318652 10464
rect 318704 10452 318710 10464
rect 418653 10455 418711 10461
rect 418653 10452 418665 10455
rect 318704 10424 418665 10452
rect 318704 10412 318710 10424
rect 418653 10421 418665 10424
rect 418699 10421 418711 10455
rect 418653 10415 418711 10421
rect 418742 10412 418748 10464
rect 418800 10452 418806 10464
rect 481578 10452 481584 10464
rect 418800 10424 481584 10452
rect 418800 10412 418806 10424
rect 481578 10412 481584 10424
rect 481636 10412 481642 10464
rect 1600 10288 583316 10384
rect 60494 10208 60500 10260
rect 60552 10248 60558 10260
rect 133545 10251 133603 10257
rect 60552 10220 133496 10248
rect 60552 10208 60558 10220
rect 65278 10140 65284 10192
rect 65336 10180 65342 10192
rect 128850 10180 128856 10192
rect 65336 10152 128856 10180
rect 65336 10140 65342 10152
rect 128850 10140 128856 10152
rect 128908 10140 128914 10192
rect 128945 10183 129003 10189
rect 128945 10149 128957 10183
rect 128991 10180 129003 10183
rect 133361 10183 133419 10189
rect 133361 10180 133373 10183
rect 128991 10152 133373 10180
rect 128991 10149 129003 10152
rect 128945 10143 129003 10149
rect 133361 10149 133373 10152
rect 133407 10149 133419 10183
rect 133468 10180 133496 10220
rect 133545 10217 133557 10251
rect 133591 10248 133603 10251
rect 143205 10251 143263 10257
rect 143205 10248 143217 10251
rect 133591 10220 143217 10248
rect 133591 10217 133603 10220
rect 133545 10211 133603 10217
rect 143205 10217 143217 10220
rect 143251 10217 143263 10251
rect 143205 10211 143263 10217
rect 143294 10208 143300 10260
rect 143352 10248 143358 10260
rect 157649 10251 157707 10257
rect 143352 10220 157600 10248
rect 143352 10208 143358 10220
rect 138145 10183 138203 10189
rect 138145 10180 138157 10183
rect 133468 10152 138157 10180
rect 133361 10143 133419 10149
rect 138145 10149 138157 10152
rect 138191 10149 138203 10183
rect 138145 10143 138203 10149
rect 138421 10183 138479 10189
rect 138421 10149 138433 10183
rect 138467 10180 138479 10183
rect 138513 10183 138571 10189
rect 138513 10180 138525 10183
rect 138467 10152 138525 10180
rect 138467 10149 138479 10152
rect 138421 10143 138479 10149
rect 138513 10149 138525 10152
rect 138559 10149 138571 10183
rect 138513 10143 138571 10149
rect 138602 10140 138608 10192
rect 138660 10180 138666 10192
rect 147989 10183 148047 10189
rect 147989 10180 148001 10183
rect 138660 10152 148001 10180
rect 138660 10140 138666 10152
rect 147989 10149 148001 10152
rect 148035 10149 148047 10183
rect 147989 10143 148047 10149
rect 148081 10183 148139 10189
rect 148081 10149 148093 10183
rect 148127 10180 148139 10183
rect 157462 10180 157468 10192
rect 148127 10152 157468 10180
rect 148127 10149 148139 10152
rect 148081 10143 148139 10149
rect 157462 10140 157468 10152
rect 157520 10140 157526 10192
rect 157572 10180 157600 10220
rect 157649 10217 157661 10251
rect 157695 10248 157707 10251
rect 167493 10251 167551 10257
rect 167493 10248 167505 10251
rect 157695 10220 167505 10248
rect 157695 10217 157707 10220
rect 157649 10211 157707 10217
rect 167493 10217 167505 10220
rect 167539 10217 167551 10251
rect 167493 10211 167551 10217
rect 167692 10220 196148 10248
rect 157741 10183 157799 10189
rect 157572 10152 157692 10180
rect 68038 10072 68044 10124
rect 68096 10112 68102 10124
rect 138234 10112 138240 10124
rect 68096 10084 138240 10112
rect 68096 10072 68102 10084
rect 138234 10072 138240 10084
rect 138292 10072 138298 10124
rect 138329 10115 138387 10121
rect 138329 10081 138341 10115
rect 138375 10112 138387 10115
rect 143294 10112 143300 10124
rect 138375 10084 143300 10112
rect 138375 10081 138387 10084
rect 138329 10075 138387 10081
rect 143294 10072 143300 10084
rect 143352 10072 143358 10124
rect 143389 10115 143447 10121
rect 143389 10081 143401 10115
rect 143435 10112 143447 10115
rect 147805 10115 147863 10121
rect 147805 10112 147817 10115
rect 143435 10084 147817 10112
rect 143435 10081 143447 10084
rect 143389 10075 143447 10081
rect 147805 10081 147817 10084
rect 147851 10081 147863 10115
rect 147805 10075 147863 10081
rect 147897 10115 147955 10121
rect 147897 10081 147909 10115
rect 147943 10112 147955 10115
rect 157554 10112 157560 10124
rect 147943 10084 157560 10112
rect 147943 10081 147955 10084
rect 147897 10075 147955 10081
rect 157554 10072 157560 10084
rect 157612 10072 157618 10124
rect 157664 10112 157692 10152
rect 157741 10149 157753 10183
rect 157787 10180 157799 10183
rect 167582 10180 167588 10192
rect 157787 10152 167588 10180
rect 157787 10149 157799 10152
rect 157741 10143 157799 10149
rect 167582 10140 167588 10152
rect 167640 10140 167646 10192
rect 167692 10112 167720 10220
rect 167858 10140 167864 10192
rect 167916 10180 167922 10192
rect 195918 10180 195924 10192
rect 167916 10152 195924 10180
rect 167916 10140 167922 10152
rect 195918 10140 195924 10152
rect 195976 10140 195982 10192
rect 157664 10084 167720 10112
rect 167766 10072 167772 10124
rect 167824 10112 167830 10124
rect 196010 10112 196016 10124
rect 167824 10084 196016 10112
rect 167824 10072 167830 10084
rect 196010 10072 196016 10084
rect 196068 10072 196074 10124
rect 196120 10112 196148 10220
rect 196378 10208 196384 10260
rect 196436 10248 196442 10260
rect 196436 10220 225588 10248
rect 196436 10208 196442 10220
rect 196197 10183 196255 10189
rect 196197 10149 196209 10183
rect 196243 10180 196255 10183
rect 225450 10180 225456 10192
rect 196243 10152 225456 10180
rect 196243 10149 196255 10152
rect 196197 10143 196255 10149
rect 225450 10140 225456 10152
rect 225508 10140 225514 10192
rect 225560 10180 225588 10220
rect 225634 10208 225640 10260
rect 225692 10248 225698 10260
rect 232353 10251 232411 10257
rect 232353 10248 232365 10251
rect 225692 10220 232365 10248
rect 225692 10208 225698 10220
rect 232353 10217 232365 10220
rect 232399 10217 232411 10251
rect 232353 10211 232411 10217
rect 232442 10208 232448 10260
rect 232500 10248 232506 10260
rect 235297 10251 235355 10257
rect 232500 10220 232545 10248
rect 232500 10208 232506 10220
rect 235297 10217 235309 10251
rect 235343 10248 235355 10251
rect 239618 10248 239624 10260
rect 235343 10220 239624 10248
rect 235343 10217 235355 10220
rect 235297 10211 235355 10217
rect 239618 10208 239624 10220
rect 239676 10208 239682 10260
rect 327110 10208 327116 10260
rect 327168 10248 327174 10260
rect 331253 10251 331311 10257
rect 331253 10248 331265 10251
rect 327168 10220 331265 10248
rect 327168 10208 327174 10220
rect 331253 10217 331265 10220
rect 331299 10217 331311 10251
rect 455910 10248 455916 10260
rect 331253 10211 331311 10217
rect 331544 10220 455916 10248
rect 234929 10183 234987 10189
rect 234929 10180 234941 10183
rect 225560 10152 234941 10180
rect 234929 10149 234941 10152
rect 234975 10149 234987 10183
rect 234929 10143 234987 10149
rect 235389 10183 235447 10189
rect 235389 10149 235401 10183
rect 235435 10180 235447 10183
rect 240906 10180 240912 10192
rect 235435 10152 240912 10180
rect 235435 10149 235447 10152
rect 235389 10143 235447 10149
rect 240906 10140 240912 10152
rect 240964 10140 240970 10192
rect 244865 10183 244923 10189
rect 244865 10149 244877 10183
rect 244911 10180 244923 10183
rect 253510 10180 253516 10192
rect 244911 10152 253516 10180
rect 244911 10149 244923 10152
rect 244865 10143 244923 10149
rect 253510 10140 253516 10152
rect 253568 10140 253574 10192
rect 325822 10140 325828 10192
rect 325880 10180 325886 10192
rect 331544 10189 331572 10220
rect 455910 10208 455916 10220
rect 455968 10208 455974 10260
rect 331437 10183 331495 10189
rect 331437 10180 331449 10183
rect 325880 10152 331449 10180
rect 325880 10140 325886 10152
rect 331437 10149 331449 10152
rect 331483 10149 331495 10183
rect 331437 10143 331495 10149
rect 331529 10183 331587 10189
rect 331529 10149 331541 10183
rect 331575 10149 331587 10183
rect 331529 10143 331587 10149
rect 331618 10140 331624 10192
rect 331676 10180 331682 10192
rect 451862 10180 451868 10192
rect 331676 10152 451868 10180
rect 331676 10140 331682 10152
rect 451862 10140 451868 10152
rect 451920 10140 451926 10192
rect 225545 10115 225603 10121
rect 225545 10112 225557 10115
rect 196120 10084 225557 10112
rect 225545 10081 225557 10084
rect 225591 10081 225603 10115
rect 225545 10075 225603 10081
rect 225634 10072 225640 10124
rect 225692 10112 225698 10124
rect 235018 10112 235024 10124
rect 225692 10084 235024 10112
rect 225692 10072 225698 10084
rect 235018 10072 235024 10084
rect 235076 10072 235082 10124
rect 241918 10072 241924 10124
rect 241976 10112 241982 10124
rect 242378 10112 242384 10124
rect 241976 10084 242384 10112
rect 241976 10072 241982 10084
rect 242378 10072 242384 10084
rect 242436 10072 242442 10124
rect 244770 10072 244776 10124
rect 244828 10112 244834 10124
rect 254525 10115 254583 10121
rect 254525 10112 254537 10115
rect 244828 10084 254537 10112
rect 244828 10072 244834 10084
rect 254525 10081 254537 10084
rect 254571 10081 254583 10115
rect 254525 10075 254583 10081
rect 325914 10072 325920 10124
rect 325972 10112 325978 10124
rect 325972 10084 331296 10112
rect 325972 10072 325978 10084
rect 102538 10004 102544 10056
rect 102596 10044 102602 10056
rect 250382 10044 250388 10056
rect 102596 10016 250388 10044
rect 102596 10004 102602 10016
rect 250382 10004 250388 10016
rect 250440 10004 250446 10056
rect 324534 10004 324540 10056
rect 324592 10044 324598 10056
rect 331161 10047 331219 10053
rect 331161 10044 331173 10047
rect 324592 10016 331173 10044
rect 324592 10004 324598 10016
rect 331161 10013 331173 10016
rect 331207 10013 331219 10047
rect 331268 10044 331296 10084
rect 331342 10072 331348 10124
rect 331400 10112 331406 10124
rect 449010 10112 449016 10124
rect 331400 10084 449016 10112
rect 331400 10072 331406 10084
rect 449010 10072 449016 10084
rect 449068 10072 449074 10124
rect 331529 10047 331587 10053
rect 331529 10044 331541 10047
rect 331268 10016 331541 10044
rect 331161 10007 331219 10013
rect 331529 10013 331541 10016
rect 331575 10013 331587 10047
rect 331529 10007 331587 10013
rect 331618 10004 331624 10056
rect 331676 10044 331682 10056
rect 444870 10044 444876 10056
rect 331676 10016 444876 10044
rect 331676 10004 331682 10016
rect 444870 10004 444876 10016
rect 444928 10004 444934 10056
rect 106678 9936 106684 9988
rect 106736 9976 106742 9988
rect 252314 9976 252320 9988
rect 106736 9948 252320 9976
rect 106736 9936 106742 9948
rect 252314 9936 252320 9948
rect 252372 9936 252378 9988
rect 321774 9936 321780 9988
rect 321832 9976 321838 9988
rect 442110 9976 442116 9988
rect 321832 9948 442116 9976
rect 321832 9936 321838 9948
rect 442110 9936 442116 9948
rect 442168 9936 442174 9988
rect 109438 9868 109444 9920
rect 109496 9908 109502 9920
rect 251854 9908 251860 9920
rect 109496 9880 251860 9908
rect 109496 9868 109502 9880
rect 251854 9868 251860 9880
rect 251912 9868 251918 9920
rect 254617 9911 254675 9917
rect 254617 9877 254629 9911
rect 254663 9908 254675 9911
rect 259125 9911 259183 9917
rect 259125 9908 259137 9911
rect 254663 9880 259137 9908
rect 254663 9877 254675 9880
rect 254617 9871 254675 9877
rect 259125 9877 259137 9880
rect 259171 9877 259183 9911
rect 259125 9871 259183 9877
rect 320210 9868 320216 9920
rect 320268 9908 320274 9920
rect 437970 9908 437976 9920
rect 320268 9880 437976 9908
rect 320268 9868 320274 9880
rect 437970 9868 437976 9880
rect 438028 9868 438034 9920
rect 1600 9744 583316 9840
rect 91498 9704 91504 9716
rect 91459 9676 91504 9704
rect 91498 9664 91504 9676
rect 91556 9664 91562 9716
rect 113578 9664 113584 9716
rect 113636 9704 113642 9716
rect 244865 9707 244923 9713
rect 244865 9704 244877 9707
rect 113636 9676 244877 9704
rect 113636 9664 113642 9676
rect 244865 9673 244877 9676
rect 244911 9673 244923 9707
rect 244865 9667 244923 9673
rect 244957 9707 245015 9713
rect 244957 9673 244969 9707
rect 245003 9704 245015 9707
rect 254341 9707 254399 9713
rect 254341 9704 254353 9707
rect 245003 9676 254353 9704
rect 245003 9673 245015 9676
rect 244957 9667 245015 9673
rect 254341 9673 254353 9676
rect 254387 9673 254399 9707
rect 254709 9707 254767 9713
rect 254709 9704 254721 9707
rect 254341 9667 254399 9673
rect 254448 9676 254721 9704
rect 124618 9596 124624 9648
rect 124676 9636 124682 9648
rect 138234 9636 138240 9648
rect 124676 9608 138240 9636
rect 124676 9596 124682 9608
rect 138234 9596 138240 9608
rect 138292 9596 138298 9648
rect 138329 9639 138387 9645
rect 138329 9605 138341 9639
rect 138375 9636 138387 9639
rect 138697 9639 138755 9645
rect 138375 9608 138648 9636
rect 138375 9605 138387 9608
rect 138329 9599 138387 9605
rect 128850 9528 128856 9580
rect 128908 9568 128914 9580
rect 138513 9571 138571 9577
rect 138513 9568 138525 9571
rect 128908 9540 138525 9568
rect 128908 9528 128914 9540
rect 138513 9537 138525 9540
rect 138559 9537 138571 9571
rect 138620 9568 138648 9608
rect 138697 9605 138709 9639
rect 138743 9636 138755 9639
rect 147897 9639 147955 9645
rect 147897 9636 147909 9639
rect 138743 9608 147909 9636
rect 138743 9605 138755 9608
rect 138697 9599 138755 9605
rect 147897 9605 147909 9608
rect 147943 9605 147955 9639
rect 147897 9599 147955 9605
rect 147989 9639 148047 9645
rect 147989 9605 148001 9639
rect 148035 9636 148047 9639
rect 148265 9639 148323 9645
rect 148265 9636 148277 9639
rect 148035 9608 148277 9636
rect 148035 9605 148047 9608
rect 147989 9599 148047 9605
rect 148265 9605 148277 9608
rect 148311 9605 148323 9639
rect 148265 9599 148323 9605
rect 162525 9639 162583 9645
rect 162525 9605 162537 9639
rect 162571 9636 162583 9639
rect 169514 9636 169520 9648
rect 162571 9608 169520 9636
rect 162571 9605 162583 9608
rect 162525 9599 162583 9605
rect 169514 9596 169520 9608
rect 169572 9596 169578 9648
rect 170158 9596 170164 9648
rect 170216 9636 170222 9648
rect 254448 9636 254476 9676
rect 254709 9673 254721 9676
rect 254755 9673 254767 9707
rect 254709 9667 254767 9673
rect 254801 9707 254859 9713
rect 254801 9673 254813 9707
rect 254847 9704 254859 9707
rect 254847 9676 257604 9704
rect 254847 9673 254859 9676
rect 254801 9667 254859 9673
rect 170216 9608 254476 9636
rect 254525 9639 254583 9645
rect 170216 9596 170222 9608
rect 254525 9605 254537 9639
rect 254571 9636 254583 9639
rect 257466 9636 257472 9648
rect 254571 9608 257472 9636
rect 254571 9605 254583 9608
rect 254525 9599 254583 9605
rect 257466 9596 257472 9608
rect 257524 9596 257530 9648
rect 257576 9636 257604 9676
rect 285066 9664 285072 9716
rect 285124 9704 285130 9716
rect 285250 9704 285256 9716
rect 285124 9676 285256 9704
rect 285124 9664 285130 9676
rect 285250 9664 285256 9676
rect 285308 9664 285314 9716
rect 305030 9664 305036 9716
rect 305088 9704 305094 9716
rect 305122 9704 305128 9716
rect 305088 9676 305128 9704
rect 305088 9664 305094 9676
rect 305122 9664 305128 9676
rect 305180 9664 305186 9716
rect 308250 9704 308256 9716
rect 308211 9676 308256 9704
rect 308250 9664 308256 9676
rect 308308 9664 308314 9716
rect 320118 9664 320124 9716
rect 320176 9704 320182 9716
rect 428313 9707 428371 9713
rect 428313 9704 428325 9707
rect 320176 9676 428325 9704
rect 320176 9664 320182 9676
rect 428313 9673 428325 9676
rect 428359 9673 428371 9707
rect 435118 9704 435124 9716
rect 428313 9667 428371 9673
rect 431272 9676 435124 9704
rect 262802 9636 262808 9648
rect 257576 9608 262808 9636
rect 262802 9596 262808 9608
rect 262860 9596 262866 9648
rect 309170 9596 309176 9648
rect 309228 9636 309234 9648
rect 385162 9636 385168 9648
rect 309228 9608 385168 9636
rect 309228 9596 309234 9608
rect 385162 9596 385168 9608
rect 385220 9596 385226 9648
rect 418653 9639 418711 9645
rect 418653 9605 418665 9639
rect 418699 9636 418711 9639
rect 431070 9636 431076 9648
rect 418699 9608 431076 9636
rect 418699 9605 418711 9608
rect 418653 9599 418711 9605
rect 431070 9596 431076 9608
rect 431128 9596 431134 9648
rect 148081 9571 148139 9577
rect 148081 9568 148093 9571
rect 138620 9540 148093 9568
rect 138513 9531 138571 9537
rect 148081 9537 148093 9540
rect 148127 9537 148139 9571
rect 148081 9531 148139 9537
rect 150930 9528 150936 9580
rect 150988 9568 150994 9580
rect 261606 9568 261612 9580
rect 150988 9540 261612 9568
rect 150988 9528 150994 9540
rect 261606 9528 261612 9540
rect 261664 9528 261670 9580
rect 310642 9528 310648 9580
rect 310700 9568 310706 9580
rect 388750 9568 388756 9580
rect 310700 9540 388756 9568
rect 310700 9528 310706 9540
rect 388750 9528 388756 9540
rect 388808 9528 388814 9580
rect 418745 9571 418803 9577
rect 418745 9537 418757 9571
rect 418791 9568 418803 9571
rect 426930 9568 426936 9580
rect 418791 9540 426936 9568
rect 418791 9537 418803 9540
rect 418745 9531 418803 9537
rect 426930 9528 426936 9540
rect 426988 9528 426994 9580
rect 147342 9460 147348 9512
rect 147400 9500 147406 9512
rect 244773 9503 244831 9509
rect 244773 9500 244785 9503
rect 147400 9472 244785 9500
rect 147400 9460 147406 9472
rect 244773 9469 244785 9472
rect 244819 9469 244831 9503
rect 244773 9463 244831 9469
rect 244865 9503 244923 9509
rect 244865 9469 244877 9503
rect 244911 9500 244923 9503
rect 259030 9500 259036 9512
rect 244911 9472 259036 9500
rect 244911 9469 244923 9472
rect 244865 9463 244923 9469
rect 259030 9460 259036 9472
rect 259088 9460 259094 9512
rect 259125 9503 259183 9509
rect 259125 9469 259137 9503
rect 259171 9500 259183 9503
rect 262894 9500 262900 9512
rect 259171 9472 262900 9500
rect 259171 9469 259183 9472
rect 259125 9463 259183 9469
rect 262894 9460 262900 9472
rect 262952 9460 262958 9512
rect 312022 9460 312028 9512
rect 312080 9500 312086 9512
rect 392338 9500 392344 9512
rect 312080 9472 392344 9500
rect 312080 9460 312086 9472
rect 392338 9460 392344 9472
rect 392396 9460 392402 9512
rect 428313 9503 428371 9509
rect 428313 9469 428325 9503
rect 428359 9500 428371 9503
rect 431272 9500 431300 9676
rect 435118 9664 435124 9676
rect 435176 9664 435182 9716
rect 529053 9707 529111 9713
rect 529053 9673 529065 9707
rect 529099 9704 529111 9707
rect 529142 9704 529148 9716
rect 529099 9676 529148 9704
rect 529099 9673 529111 9676
rect 529053 9667 529111 9673
rect 529142 9664 529148 9676
rect 529200 9664 529206 9716
rect 535953 9707 536011 9713
rect 535953 9673 535965 9707
rect 535999 9704 536011 9707
rect 536226 9704 536232 9716
rect 535999 9676 536232 9704
rect 535999 9673 536011 9676
rect 535953 9667 536011 9673
rect 536226 9664 536232 9676
rect 536284 9664 536290 9716
rect 541473 9707 541531 9713
rect 541473 9673 541485 9707
rect 541519 9704 541531 9707
rect 542206 9704 542212 9716
rect 541519 9676 542212 9704
rect 541519 9673 541531 9676
rect 541473 9667 541531 9673
rect 542206 9664 542212 9676
rect 542264 9664 542270 9716
rect 545518 9664 545524 9716
rect 545576 9704 545582 9716
rect 545794 9704 545800 9716
rect 545576 9676 545800 9704
rect 545576 9664 545582 9676
rect 545794 9664 545800 9676
rect 545852 9664 545858 9716
rect 552513 9707 552571 9713
rect 552513 9673 552525 9707
rect 552559 9704 552571 9707
rect 552878 9704 552884 9716
rect 552559 9676 552884 9704
rect 552559 9673 552571 9676
rect 552513 9667 552571 9673
rect 552878 9664 552884 9676
rect 552936 9664 552942 9716
rect 560793 9707 560851 9713
rect 560793 9673 560805 9707
rect 560839 9704 560851 9707
rect 561250 9704 561256 9716
rect 560839 9676 561256 9704
rect 560839 9673 560851 9676
rect 560793 9667 560851 9673
rect 561250 9664 561256 9676
rect 561308 9664 561314 9716
rect 571833 9707 571891 9713
rect 571833 9673 571845 9707
rect 571879 9704 571891 9707
rect 571922 9704 571928 9716
rect 571879 9676 571928 9704
rect 571879 9673 571891 9676
rect 571833 9667 571891 9673
rect 571922 9664 571928 9676
rect 571980 9664 571986 9716
rect 428359 9472 431300 9500
rect 428359 9469 428371 9472
rect 428313 9463 428371 9469
rect 259214 9432 259220 9444
rect 148004 9404 259220 9432
rect 143754 9324 143760 9376
rect 143812 9364 143818 9376
rect 148004 9364 148032 9404
rect 259214 9392 259220 9404
rect 259272 9392 259278 9444
rect 349374 9392 349380 9444
rect 349432 9432 349438 9444
rect 350757 9435 350815 9441
rect 350757 9432 350769 9435
rect 349432 9404 350769 9432
rect 349432 9392 349438 9404
rect 350757 9401 350769 9404
rect 350803 9401 350815 9435
rect 350757 9395 350815 9401
rect 350846 9392 350852 9444
rect 350904 9432 350910 9444
rect 351033 9435 351091 9441
rect 351033 9432 351045 9435
rect 350904 9404 351045 9432
rect 350904 9392 350910 9404
rect 351033 9401 351045 9404
rect 351079 9401 351091 9435
rect 351033 9395 351091 9401
rect 351122 9392 351128 9444
rect 351180 9432 351186 9444
rect 560054 9432 560060 9444
rect 351180 9404 560060 9432
rect 351180 9392 351186 9404
rect 560054 9392 560060 9404
rect 560112 9392 560118 9444
rect 143812 9336 148032 9364
rect 148081 9367 148139 9373
rect 143812 9324 143818 9336
rect 148081 9333 148093 9367
rect 148127 9364 148139 9367
rect 244773 9367 244831 9373
rect 244773 9364 244785 9367
rect 148127 9336 244785 9364
rect 148127 9333 148139 9336
rect 148081 9327 148139 9333
rect 244773 9333 244785 9336
rect 244819 9333 244831 9367
rect 244773 9327 244831 9333
rect 244862 9324 244868 9376
rect 244920 9364 244926 9376
rect 279638 9364 279644 9376
rect 244920 9336 279644 9364
rect 244920 9324 244926 9336
rect 279638 9324 279644 9336
rect 279696 9324 279702 9376
rect 341278 9324 341284 9376
rect 341336 9364 341342 9376
rect 346525 9367 346583 9373
rect 346525 9364 346537 9367
rect 341336 9336 346537 9364
rect 341336 9324 341342 9336
rect 346525 9333 346537 9336
rect 346571 9333 346583 9367
rect 346525 9327 346583 9333
rect 346614 9324 346620 9376
rect 346672 9364 346678 9376
rect 349282 9364 349288 9376
rect 346672 9336 349288 9364
rect 346672 9324 346678 9336
rect 349282 9324 349288 9336
rect 349340 9324 349346 9376
rect 349466 9324 349472 9376
rect 349524 9364 349530 9376
rect 350665 9367 350723 9373
rect 350665 9364 350677 9367
rect 349524 9336 350677 9364
rect 349524 9324 349530 9336
rect 350665 9333 350677 9336
rect 350711 9333 350723 9367
rect 350665 9327 350723 9333
rect 350941 9367 350999 9373
rect 350941 9333 350953 9367
rect 350987 9364 350999 9367
rect 355909 9367 355967 9373
rect 355909 9364 355921 9367
rect 350987 9336 355921 9364
rect 350987 9333 350999 9336
rect 350941 9327 350999 9333
rect 355909 9333 355921 9336
rect 355955 9333 355967 9367
rect 355909 9327 355967 9333
rect 356001 9367 356059 9373
rect 356001 9333 356013 9367
rect 356047 9364 356059 9367
rect 563642 9364 563648 9376
rect 356047 9336 563648 9364
rect 356047 9333 356059 9336
rect 356001 9327 356059 9333
rect 563642 9324 563648 9336
rect 563700 9324 563706 9376
rect 1600 9200 583316 9296
rect 18453 9163 18511 9169
rect 18453 9129 18465 9163
rect 18499 9160 18511 9163
rect 28021 9163 28079 9169
rect 28021 9160 28033 9163
rect 18499 9132 28033 9160
rect 18499 9129 18511 9132
rect 18453 9123 18511 9129
rect 28021 9129 28033 9132
rect 28067 9129 28079 9163
rect 28021 9123 28079 9129
rect 36393 9163 36451 9169
rect 36393 9129 36405 9163
rect 36439 9160 36451 9163
rect 42649 9163 42707 9169
rect 42649 9160 42661 9163
rect 36439 9132 42661 9160
rect 36439 9129 36451 9132
rect 36393 9123 36451 9129
rect 42649 9129 42661 9132
rect 42695 9129 42707 9163
rect 42649 9123 42707 9129
rect 54241 9163 54299 9169
rect 54241 9129 54253 9163
rect 54287 9160 54299 9163
rect 65373 9163 65431 9169
rect 65373 9160 65385 9163
rect 54287 9132 65385 9160
rect 54287 9129 54299 9132
rect 54241 9123 54299 9129
rect 65373 9129 65385 9132
rect 65419 9129 65431 9163
rect 65373 9123 65431 9129
rect 75033 9163 75091 9169
rect 75033 9129 75045 9163
rect 75079 9160 75091 9163
rect 81197 9163 81255 9169
rect 81197 9160 81209 9163
rect 75079 9132 81209 9160
rect 75079 9129 75091 9132
rect 75033 9123 75091 9129
rect 81197 9129 81209 9132
rect 81243 9129 81255 9163
rect 81197 9123 81255 9129
rect 92881 9163 92939 9169
rect 92881 9129 92893 9163
rect 92927 9160 92939 9163
rect 104013 9163 104071 9169
rect 104013 9160 104025 9163
rect 92927 9132 104025 9160
rect 92927 9129 92939 9132
rect 92881 9123 92939 9129
rect 104013 9129 104025 9132
rect 104059 9129 104071 9163
rect 104013 9123 104071 9129
rect 113673 9163 113731 9169
rect 113673 9129 113685 9163
rect 113719 9160 113731 9163
rect 116249 9163 116307 9169
rect 116249 9160 116261 9163
rect 113719 9132 116261 9160
rect 113719 9129 113731 9132
rect 113673 9123 113731 9129
rect 116249 9129 116261 9132
rect 116295 9129 116307 9163
rect 116249 9123 116307 9129
rect 136578 9120 136584 9172
rect 136636 9160 136642 9172
rect 244770 9160 244776 9172
rect 136636 9132 244776 9160
rect 136636 9120 136642 9132
rect 244770 9120 244776 9132
rect 244828 9120 244834 9172
rect 244862 9120 244868 9172
rect 244920 9160 244926 9172
rect 254246 9160 254252 9172
rect 244920 9132 254252 9160
rect 244920 9120 244926 9132
rect 254246 9120 254252 9132
rect 254304 9120 254310 9172
rect 254341 9163 254399 9169
rect 254341 9129 254353 9163
rect 254387 9160 254399 9163
rect 254430 9160 254436 9172
rect 254387 9132 254436 9160
rect 254387 9129 254399 9132
rect 254341 9123 254399 9129
rect 254430 9120 254436 9132
rect 254488 9120 254494 9172
rect 254522 9120 254528 9172
rect 254580 9160 254586 9172
rect 278074 9160 278080 9172
rect 254580 9132 278080 9160
rect 254580 9120 254586 9132
rect 278074 9120 278080 9132
rect 278132 9120 278138 9172
rect 341281 9163 341339 9169
rect 341281 9129 341293 9163
rect 341327 9160 341339 9163
rect 350665 9163 350723 9169
rect 350665 9160 350677 9163
rect 341327 9132 350677 9160
rect 341327 9129 341339 9132
rect 341281 9123 341339 9129
rect 350665 9129 350677 9132
rect 350711 9129 350723 9163
rect 350665 9123 350723 9129
rect 350849 9163 350907 9169
rect 350849 9129 350861 9163
rect 350895 9160 350907 9163
rect 351033 9163 351091 9169
rect 351033 9160 351045 9163
rect 350895 9132 351045 9160
rect 350895 9129 350907 9132
rect 350849 9123 350907 9129
rect 351033 9129 351045 9132
rect 351079 9129 351091 9163
rect 351033 9123 351091 9129
rect 351125 9163 351183 9169
rect 351125 9129 351137 9163
rect 351171 9160 351183 9163
rect 567230 9160 567236 9172
rect 351171 9132 567236 9160
rect 351171 9129 351183 9132
rect 351125 9123 351183 9129
rect 567230 9120 567236 9132
rect 567288 9120 567294 9172
rect 27190 9052 27196 9104
rect 27248 9092 27254 9104
rect 234745 9095 234803 9101
rect 234745 9092 234757 9095
rect 27248 9064 234757 9092
rect 27248 9052 27254 9064
rect 234745 9061 234757 9064
rect 234791 9061 234803 9095
rect 278166 9092 278172 9104
rect 234745 9055 234803 9061
rect 234852 9064 278172 9092
rect 31517 9027 31575 9033
rect 31517 8993 31529 9027
rect 31563 9024 31575 9027
rect 36393 9027 36451 9033
rect 36393 9024 36405 9027
rect 31563 8996 36405 9024
rect 31563 8993 31575 8996
rect 31517 8987 31575 8993
rect 36393 8993 36405 8996
rect 36439 8993 36451 9027
rect 36393 8987 36451 8993
rect 65373 9027 65431 9033
rect 65373 8993 65385 9027
rect 65419 9024 65431 9027
rect 75033 9027 75091 9033
rect 75033 9024 75045 9027
rect 65419 8996 75045 9024
rect 65419 8993 65431 8996
rect 65373 8987 65431 8993
rect 75033 8993 75045 8996
rect 75079 8993 75091 9027
rect 75033 8987 75091 8993
rect 85981 9027 86039 9033
rect 85981 8993 85993 9027
rect 86027 8993 86039 9027
rect 85981 8987 86039 8993
rect 104013 9027 104071 9033
rect 104013 8993 104025 9027
rect 104059 9024 104071 9027
rect 113673 9027 113731 9033
rect 113673 9024 113685 9027
rect 104059 8996 113685 9024
rect 104059 8993 104071 8996
rect 104013 8987 104071 8993
rect 113673 8993 113685 8996
rect 113719 8993 113731 9027
rect 113673 8987 113731 8993
rect 116249 9027 116307 9033
rect 116249 8993 116261 9027
rect 116295 9024 116307 9027
rect 140077 9027 140135 9033
rect 140077 9024 140089 9027
rect 116295 8996 140089 9024
rect 116295 8993 116307 8996
rect 116249 8987 116307 8993
rect 140077 8993 140089 8996
rect 140123 8993 140135 9027
rect 140077 8987 140135 8993
rect 9342 8916 9348 8968
rect 9400 8956 9406 8968
rect 18453 8959 18511 8965
rect 18453 8956 18465 8959
rect 9400 8928 18465 8956
rect 9400 8916 9406 8928
rect 18453 8925 18465 8928
rect 18499 8925 18511 8959
rect 18453 8919 18511 8925
rect 28021 8959 28079 8965
rect 28021 8925 28033 8959
rect 28067 8956 28079 8959
rect 37773 8959 37831 8965
rect 37773 8956 37785 8959
rect 28067 8928 37785 8956
rect 28067 8925 28079 8928
rect 28021 8919 28079 8925
rect 37773 8925 37785 8928
rect 37819 8925 37831 8959
rect 37773 8919 37831 8925
rect 47341 8959 47399 8965
rect 47341 8925 47353 8959
rect 47387 8956 47399 8959
rect 57093 8959 57151 8965
rect 57093 8956 57105 8959
rect 47387 8928 57105 8956
rect 47387 8925 47399 8928
rect 47341 8919 47399 8925
rect 57093 8925 57105 8928
rect 57139 8925 57151 8959
rect 57093 8919 57151 8925
rect 66661 8959 66719 8965
rect 66661 8925 66673 8959
rect 66707 8956 66719 8959
rect 68133 8959 68191 8965
rect 68133 8956 68145 8959
rect 66707 8928 68145 8956
rect 66707 8925 66719 8928
rect 66661 8919 66719 8925
rect 68133 8925 68145 8928
rect 68179 8925 68191 8959
rect 85996 8956 86024 8987
rect 140166 8984 140172 9036
rect 140224 9024 140230 9036
rect 148081 9027 148139 9033
rect 148081 9024 148093 9027
rect 140224 8996 148093 9024
rect 140224 8984 140230 8996
rect 148081 8993 148093 8996
rect 148127 8993 148139 9027
rect 148081 8987 148139 8993
rect 162617 9027 162675 9033
rect 162617 8993 162629 9027
rect 162663 9024 162675 9027
rect 172277 9027 172335 9033
rect 172277 9024 172289 9027
rect 162663 8996 172289 9024
rect 162663 8993 162675 8996
rect 162617 8987 162675 8993
rect 172277 8993 172289 8996
rect 172323 8993 172335 9027
rect 172277 8987 172335 8993
rect 181937 9027 181995 9033
rect 181937 8993 181949 9027
rect 181983 9024 181995 9027
rect 191597 9027 191655 9033
rect 191597 9024 191609 9027
rect 181983 8996 191609 9024
rect 181983 8993 181995 8996
rect 181937 8987 181995 8993
rect 191597 8993 191609 8996
rect 191643 8993 191655 9027
rect 191597 8987 191655 8993
rect 191778 8984 191784 9036
rect 191836 9024 191842 9036
rect 196565 9027 196623 9033
rect 196565 9024 196577 9027
rect 191836 8996 196577 9024
rect 191836 8984 191842 8996
rect 196565 8993 196577 8996
rect 196611 8993 196623 9027
rect 196565 8987 196623 8993
rect 201257 9027 201315 9033
rect 201257 8993 201269 9027
rect 201303 9024 201315 9027
rect 210917 9027 210975 9033
rect 210917 9024 210929 9027
rect 201303 8996 210929 9024
rect 201303 8993 201315 8996
rect 201257 8987 201315 8993
rect 210917 8993 210929 8996
rect 210963 8993 210975 9027
rect 210917 8987 210975 8993
rect 215885 9027 215943 9033
rect 215885 8993 215897 9027
rect 215931 9024 215943 9027
rect 233822 9024 233828 9036
rect 215931 8996 233828 9024
rect 215931 8993 215943 8996
rect 215885 8987 215943 8993
rect 233822 8984 233828 8996
rect 233880 8984 233886 9036
rect 115053 8959 115111 8965
rect 115053 8956 115065 8959
rect 85996 8928 115065 8956
rect 68133 8919 68191 8925
rect 115053 8925 115065 8928
rect 115099 8925 115111 8959
rect 115053 8919 115111 8925
rect 124621 8959 124679 8965
rect 124621 8925 124633 8959
rect 124667 8956 124679 8959
rect 134373 8959 134431 8965
rect 134373 8956 134385 8959
rect 124667 8928 134385 8956
rect 124667 8925 124679 8928
rect 124621 8919 124679 8925
rect 134373 8925 134385 8928
rect 134419 8925 134431 8959
rect 134373 8919 134431 8925
rect 138513 8959 138571 8965
rect 138513 8925 138525 8959
rect 138559 8956 138571 8959
rect 231338 8956 231344 8968
rect 138559 8928 231344 8956
rect 138559 8925 138571 8928
rect 138513 8919 138571 8925
rect 231338 8916 231344 8928
rect 231396 8916 231402 8968
rect 232994 8916 233000 8968
rect 233052 8956 233058 8968
rect 234852 8956 234880 9064
rect 278166 9052 278172 9064
rect 278224 9052 278230 9104
rect 341189 9095 341247 9101
rect 341189 9061 341201 9095
rect 341235 9092 341247 9095
rect 350757 9095 350815 9101
rect 350757 9092 350769 9095
rect 341235 9064 350769 9092
rect 341235 9061 341247 9064
rect 341189 9055 341247 9061
rect 350757 9061 350769 9064
rect 350803 9061 350815 9095
rect 350757 9055 350815 9061
rect 350941 9095 350999 9101
rect 350941 9061 350953 9095
rect 350987 9092 350999 9095
rect 355909 9095 355967 9101
rect 350987 9064 355860 9092
rect 350987 9061 350999 9064
rect 350941 9055 350999 9061
rect 234926 8984 234932 9036
rect 234984 9024 234990 9036
rect 276786 9024 276792 9036
rect 234984 8996 276792 9024
rect 234984 8984 234990 8996
rect 276786 8984 276792 8996
rect 276844 8984 276850 9036
rect 303742 8984 303748 9036
rect 303800 9024 303806 9036
rect 351214 9024 351220 9036
rect 303800 8996 351220 9024
rect 303800 8984 303806 8996
rect 351214 8984 351220 8996
rect 351272 8984 351278 9036
rect 351309 9027 351367 9033
rect 351309 8993 351321 9027
rect 351355 9024 351367 9027
rect 355725 9027 355783 9033
rect 355725 9024 355737 9027
rect 351355 8996 355737 9024
rect 351355 8993 351367 8996
rect 351309 8987 351367 8993
rect 355725 8993 355737 8996
rect 355771 8993 355783 9027
rect 355832 9024 355860 9064
rect 355909 9061 355921 9095
rect 355955 9092 355967 9095
rect 570726 9092 570732 9104
rect 355955 9064 570732 9092
rect 355955 9061 355967 9064
rect 355909 9055 355967 9061
rect 570726 9052 570732 9064
rect 570784 9052 570790 9104
rect 574314 9024 574320 9036
rect 355832 8996 574320 9024
rect 355725 8987 355783 8993
rect 574314 8984 574320 8996
rect 574372 8984 574378 9036
rect 233052 8928 234880 8956
rect 233052 8916 233058 8928
rect 235018 8916 235024 8968
rect 235076 8956 235082 8968
rect 276694 8956 276700 8968
rect 235076 8928 276700 8956
rect 235076 8916 235082 8928
rect 276694 8916 276700 8928
rect 276752 8916 276758 8968
rect 303926 8916 303932 8968
rect 303984 8956 303990 8968
rect 351030 8956 351036 8968
rect 303984 8928 351036 8956
rect 303984 8916 303990 8928
rect 351030 8916 351036 8928
rect 351088 8916 351094 8968
rect 351125 8959 351183 8965
rect 351125 8925 351137 8959
rect 351171 8956 351183 8959
rect 577902 8956 577908 8968
rect 351171 8928 577908 8956
rect 351171 8925 351183 8928
rect 351125 8919 351183 8925
rect 577902 8916 577908 8928
rect 577960 8916 577966 8968
rect 22406 8848 22412 8900
rect 22464 8888 22470 8900
rect 31517 8891 31575 8897
rect 31517 8888 31529 8891
rect 22464 8860 31529 8888
rect 22464 8848 22470 8860
rect 31517 8857 31529 8860
rect 31563 8857 31575 8891
rect 31517 8851 31575 8857
rect 42649 8891 42707 8897
rect 42649 8857 42661 8891
rect 42695 8888 42707 8891
rect 54241 8891 54299 8897
rect 54241 8888 54253 8891
rect 42695 8860 54253 8888
rect 42695 8857 42707 8860
rect 42649 8851 42707 8857
rect 54241 8857 54253 8860
rect 54287 8857 54299 8891
rect 54241 8851 54299 8857
rect 81197 8891 81255 8897
rect 81197 8857 81209 8891
rect 81243 8888 81255 8891
rect 85889 8891 85947 8897
rect 85889 8888 85901 8891
rect 81243 8860 85901 8888
rect 81243 8857 81255 8860
rect 81197 8851 81255 8857
rect 85889 8857 85901 8860
rect 85935 8857 85947 8891
rect 85889 8851 85947 8857
rect 85981 8891 86039 8897
rect 85981 8857 85993 8891
rect 86027 8888 86039 8891
rect 92881 8891 92939 8897
rect 92881 8888 92893 8891
rect 86027 8860 92893 8888
rect 86027 8857 86039 8860
rect 85981 8851 86039 8857
rect 92881 8857 92893 8860
rect 92927 8857 92939 8891
rect 92881 8851 92939 8857
rect 140261 8891 140319 8897
rect 140261 8857 140273 8891
rect 140307 8888 140319 8891
rect 148265 8891 148323 8897
rect 140307 8860 148216 8888
rect 140307 8857 140319 8860
rect 140261 8851 140319 8857
rect 57093 8823 57151 8829
rect 57093 8789 57105 8823
rect 57139 8820 57151 8823
rect 66661 8823 66719 8829
rect 66661 8820 66673 8823
rect 57139 8792 66673 8820
rect 57139 8789 57151 8792
rect 57093 8783 57151 8789
rect 66661 8789 66673 8792
rect 66707 8789 66719 8823
rect 66661 8783 66719 8789
rect 68133 8823 68191 8829
rect 68133 8789 68145 8823
rect 68179 8820 68191 8823
rect 85705 8823 85763 8829
rect 85705 8820 85717 8823
rect 68179 8792 85717 8820
rect 68179 8789 68191 8792
rect 68133 8783 68191 8789
rect 85705 8789 85717 8792
rect 85751 8789 85763 8823
rect 85705 8783 85763 8789
rect 134373 8823 134431 8829
rect 134373 8789 134385 8823
rect 134419 8820 134431 8823
rect 138421 8823 138479 8829
rect 138421 8820 138433 8823
rect 134419 8792 138433 8820
rect 134419 8789 134431 8792
rect 134373 8783 134431 8789
rect 138421 8789 138433 8792
rect 138467 8789 138479 8823
rect 148188 8820 148216 8860
rect 148265 8857 148277 8891
rect 148311 8888 148323 8891
rect 157833 8891 157891 8897
rect 157833 8888 157845 8891
rect 148311 8860 157845 8888
rect 148311 8857 148323 8860
rect 148265 8851 148323 8857
rect 157833 8857 157845 8860
rect 157879 8857 157891 8891
rect 157833 8851 157891 8857
rect 161602 8848 161608 8900
rect 161660 8888 161666 8900
rect 162893 8891 162951 8897
rect 161660 8860 162844 8888
rect 161660 8848 161666 8860
rect 162617 8823 162675 8829
rect 162617 8820 162629 8823
rect 148188 8792 162629 8820
rect 138421 8783 138479 8789
rect 162617 8789 162629 8792
rect 162663 8789 162675 8823
rect 162816 8820 162844 8860
rect 162893 8857 162905 8891
rect 162939 8888 162951 8891
rect 254709 8891 254767 8897
rect 162939 8860 254568 8888
rect 162939 8857 162951 8860
rect 162893 8851 162951 8857
rect 254433 8823 254491 8829
rect 254433 8820 254445 8823
rect 162816 8792 254445 8820
rect 162617 8783 162675 8789
rect 254433 8789 254445 8792
rect 254479 8789 254491 8823
rect 254540 8820 254568 8860
rect 254709 8857 254721 8891
rect 254755 8888 254767 8891
rect 261882 8888 261888 8900
rect 254755 8860 261888 8888
rect 254755 8857 254767 8860
rect 254709 8851 254767 8857
rect 261882 8848 261888 8860
rect 261940 8848 261946 8900
rect 309262 8848 309268 8900
rect 309320 8888 309326 8900
rect 381666 8888 381672 8900
rect 309320 8860 381672 8888
rect 309320 8848 309326 8860
rect 381666 8848 381672 8860
rect 381724 8848 381730 8900
rect 254801 8823 254859 8829
rect 254801 8820 254813 8823
rect 254540 8792 254813 8820
rect 254433 8783 254491 8789
rect 254801 8789 254813 8792
rect 254847 8789 254859 8823
rect 254801 8783 254859 8789
rect 254890 8780 254896 8832
rect 254948 8820 254954 8832
rect 260410 8820 260416 8832
rect 254948 8792 260416 8820
rect 254948 8780 254954 8792
rect 260410 8780 260416 8792
rect 260468 8780 260474 8832
rect 308066 8780 308072 8832
rect 308124 8820 308130 8832
rect 378078 8820 378084 8832
rect 308124 8792 378084 8820
rect 308124 8780 308130 8792
rect 378078 8780 378084 8792
rect 378136 8780 378142 8832
rect 1600 8656 583316 8752
rect 37773 8619 37831 8625
rect 37773 8585 37785 8619
rect 37819 8616 37831 8619
rect 47341 8619 47399 8625
rect 47341 8616 47353 8619
rect 37819 8588 47353 8616
rect 37819 8585 37831 8588
rect 37773 8579 37831 8585
rect 47341 8585 47353 8588
rect 47387 8585 47399 8619
rect 47341 8579 47399 8585
rect 115053 8619 115111 8625
rect 115053 8585 115065 8619
rect 115099 8616 115111 8619
rect 124621 8619 124679 8625
rect 124621 8616 124633 8619
rect 115099 8588 124633 8616
rect 115099 8585 115111 8588
rect 115053 8579 115111 8585
rect 124621 8585 124633 8588
rect 124667 8585 124679 8619
rect 124621 8579 124679 8585
rect 158014 8576 158020 8628
rect 158072 8616 158078 8628
rect 162893 8619 162951 8625
rect 162893 8616 162905 8619
rect 158072 8588 162905 8616
rect 158072 8576 158078 8588
rect 162893 8585 162905 8588
rect 162939 8585 162951 8619
rect 162893 8579 162951 8585
rect 172277 8619 172335 8625
rect 172277 8585 172289 8619
rect 172323 8616 172335 8619
rect 181937 8619 181995 8625
rect 181937 8616 181949 8619
rect 172323 8588 181949 8616
rect 172323 8585 172335 8588
rect 172277 8579 172335 8585
rect 181937 8585 181949 8588
rect 181983 8585 181995 8619
rect 181937 8579 181995 8585
rect 191597 8619 191655 8625
rect 191597 8585 191609 8619
rect 191643 8616 191655 8619
rect 201257 8619 201315 8625
rect 201257 8616 201269 8619
rect 191643 8588 201269 8616
rect 191643 8585 191655 8588
rect 191597 8579 191655 8585
rect 201257 8585 201269 8588
rect 201303 8585 201315 8619
rect 201257 8579 201315 8585
rect 207970 8576 207976 8628
rect 208028 8616 208034 8628
rect 272738 8616 272744 8628
rect 208028 8588 272744 8616
rect 208028 8576 208034 8588
rect 272738 8576 272744 8588
rect 272796 8576 272802 8628
rect 307974 8576 307980 8628
rect 308032 8616 308038 8628
rect 374582 8616 374588 8628
rect 308032 8588 374588 8616
rect 308032 8576 308038 8588
rect 374582 8576 374588 8588
rect 374640 8576 374646 8628
rect 154426 8508 154432 8560
rect 154484 8548 154490 8560
rect 162525 8551 162583 8557
rect 162525 8548 162537 8551
rect 154484 8520 162537 8548
rect 154484 8508 154490 8520
rect 162525 8517 162537 8520
rect 162571 8517 162583 8551
rect 162525 8511 162583 8517
rect 211558 8508 211564 8560
rect 211616 8548 211622 8560
rect 273934 8548 273940 8560
rect 211616 8520 273940 8548
rect 211616 8508 211622 8520
rect 273934 8508 273940 8520
rect 273992 8508 273998 8560
rect 306410 8508 306416 8560
rect 306468 8548 306474 8560
rect 370810 8548 370816 8560
rect 306468 8520 370816 8548
rect 306468 8508 306474 8520
rect 370810 8508 370816 8520
rect 370868 8508 370874 8560
rect 274394 8480 274400 8492
rect 218660 8452 274400 8480
rect 184234 8372 184240 8424
rect 184292 8412 184298 8424
rect 185338 8412 185344 8424
rect 184292 8384 185344 8412
rect 184292 8372 184298 8384
rect 185338 8372 185344 8384
rect 185396 8372 185402 8424
rect 186629 8415 186687 8421
rect 186629 8381 186641 8415
rect 186675 8412 186687 8415
rect 196381 8415 196439 8421
rect 196381 8412 196393 8415
rect 186675 8384 196393 8412
rect 186675 8381 186687 8384
rect 186629 8375 186687 8381
rect 196381 8381 196393 8384
rect 196427 8381 196439 8415
rect 196381 8375 196439 8381
rect 215146 8372 215152 8424
rect 215204 8412 215210 8424
rect 218660 8412 218688 8452
rect 274394 8440 274400 8452
rect 274452 8440 274458 8492
rect 306686 8440 306692 8492
rect 306744 8480 306750 8492
rect 355725 8483 355783 8489
rect 306744 8452 355676 8480
rect 306744 8440 306750 8452
rect 215204 8384 218688 8412
rect 215204 8372 215210 8384
rect 222506 8372 222512 8424
rect 222564 8412 222570 8424
rect 225361 8415 225419 8421
rect 222564 8384 225312 8412
rect 222564 8372 222570 8384
rect 177153 8347 177211 8353
rect 177153 8313 177165 8347
rect 177199 8344 177211 8347
rect 195001 8347 195059 8353
rect 195001 8344 195013 8347
rect 177199 8316 195013 8344
rect 177199 8313 177211 8316
rect 177153 8307 177211 8313
rect 195001 8313 195013 8316
rect 195047 8313 195059 8347
rect 195001 8307 195059 8313
rect 210917 8347 210975 8353
rect 210917 8313 210929 8347
rect 210963 8344 210975 8347
rect 215885 8347 215943 8353
rect 215885 8344 215897 8347
rect 210963 8316 215897 8344
rect 210963 8313 210975 8316
rect 210917 8307 210975 8313
rect 215885 8313 215897 8316
rect 215931 8313 215943 8347
rect 215885 8307 215943 8313
rect 218550 8304 218556 8356
rect 218608 8344 218614 8356
rect 225177 8347 225235 8353
rect 225177 8344 225189 8347
rect 218608 8316 225189 8344
rect 218608 8304 218614 8316
rect 225177 8313 225189 8316
rect 225223 8313 225235 8347
rect 225284 8344 225312 8384
rect 225361 8381 225373 8415
rect 225407 8412 225419 8415
rect 275314 8412 275320 8424
rect 225407 8384 275320 8412
rect 225407 8381 225419 8384
rect 225361 8375 225419 8381
rect 275314 8372 275320 8384
rect 275372 8372 275378 8424
rect 305030 8372 305036 8424
rect 305088 8412 305094 8424
rect 355541 8415 355599 8421
rect 355541 8412 355553 8415
rect 305088 8384 355553 8412
rect 305088 8372 305094 8384
rect 355541 8381 355553 8384
rect 355587 8381 355599 8415
rect 355541 8375 355599 8381
rect 275406 8344 275412 8356
rect 225284 8316 275412 8344
rect 225177 8307 225235 8313
rect 275406 8304 275412 8316
rect 275464 8304 275470 8356
rect 305306 8304 305312 8356
rect 305364 8344 305370 8356
rect 351030 8344 351036 8356
rect 305364 8316 351036 8344
rect 305364 8304 305370 8316
rect 351030 8304 351036 8316
rect 351088 8304 351094 8356
rect 351122 8304 351128 8356
rect 351180 8344 351186 8356
rect 353054 8344 353060 8356
rect 351180 8316 353060 8344
rect 351180 8304 351186 8316
rect 353054 8304 353060 8316
rect 353112 8304 353118 8356
rect 355648 8344 355676 8452
rect 355725 8449 355737 8483
rect 355771 8480 355783 8483
rect 363818 8480 363824 8492
rect 355771 8452 363824 8480
rect 355771 8449 355783 8452
rect 355725 8443 355783 8449
rect 363818 8440 363824 8452
rect 363876 8440 363882 8492
rect 363910 8440 363916 8492
rect 363968 8480 363974 8492
rect 367406 8480 367412 8492
rect 363968 8452 367412 8480
rect 363968 8440 363974 8452
rect 367406 8440 367412 8452
rect 367464 8440 367470 8492
rect 356182 8372 356188 8424
rect 356240 8412 356246 8424
rect 370350 8412 370356 8424
rect 356240 8384 370356 8412
rect 356240 8372 356246 8384
rect 370350 8372 370356 8384
rect 370408 8372 370414 8424
rect 373110 8412 373116 8424
rect 373071 8384 373116 8412
rect 373110 8372 373116 8384
rect 373168 8372 373174 8424
rect 374490 8372 374496 8424
rect 374548 8412 374554 8424
rect 375686 8412 375692 8424
rect 374548 8384 375692 8412
rect 374548 8372 374554 8384
rect 375686 8372 375692 8384
rect 375744 8372 375750 8424
rect 399422 8372 399428 8424
rect 399480 8412 399486 8424
rect 409174 8412 409180 8424
rect 399480 8384 409180 8412
rect 399480 8372 399486 8384
rect 409174 8372 409180 8384
rect 409232 8372 409238 8424
rect 438246 8372 438252 8424
rect 438304 8412 438310 8424
rect 457477 8415 457535 8421
rect 457477 8412 457489 8415
rect 438304 8384 457489 8412
rect 438304 8372 438310 8384
rect 457477 8381 457489 8384
rect 457523 8381 457535 8415
rect 457477 8375 457535 8381
rect 361150 8344 361156 8356
rect 355648 8316 361156 8344
rect 361150 8304 361156 8316
rect 361208 8304 361214 8356
rect 361242 8304 361248 8356
rect 361300 8344 361306 8356
rect 457569 8347 457627 8353
rect 457569 8344 457581 8347
rect 361300 8316 457581 8344
rect 361300 8304 361306 8316
rect 457569 8313 457581 8316
rect 457615 8313 457627 8347
rect 457569 8307 457627 8313
rect 129494 8236 129500 8288
rect 129552 8276 129558 8288
rect 256086 8276 256092 8288
rect 129552 8248 256092 8276
rect 129552 8236 129558 8248
rect 256086 8236 256092 8248
rect 256144 8236 256150 8288
rect 272830 8276 272836 8288
rect 272791 8248 272836 8276
rect 272830 8236 272836 8248
rect 272888 8236 272894 8288
rect 310274 8236 310280 8288
rect 310332 8276 310338 8288
rect 312666 8276 312672 8288
rect 310332 8248 312672 8276
rect 310332 8236 310338 8248
rect 312666 8236 312672 8248
rect 312724 8236 312730 8288
rect 337046 8236 337052 8288
rect 337104 8276 337110 8288
rect 341189 8279 341247 8285
rect 341189 8276 341201 8279
rect 337104 8248 341201 8276
rect 337104 8236 337110 8248
rect 341189 8245 341201 8248
rect 341235 8245 341247 8279
rect 341189 8239 341247 8245
rect 341278 8236 341284 8288
rect 341336 8276 341342 8288
rect 506510 8276 506516 8288
rect 341336 8248 506516 8276
rect 341336 8236 341342 8248
rect 506510 8236 506516 8248
rect 506568 8236 506574 8288
rect 1600 8112 583316 8208
rect 69970 8032 69976 8084
rect 70028 8072 70034 8084
rect 244034 8072 244040 8084
rect 70028 8044 244040 8072
rect 70028 8032 70034 8044
rect 244034 8032 244040 8044
rect 244092 8032 244098 8084
rect 249646 8032 249652 8084
rect 249704 8072 249710 8084
rect 280742 8072 280748 8084
rect 249704 8044 280748 8072
rect 249704 8032 249710 8044
rect 280742 8032 280748 8044
rect 280800 8032 280806 8084
rect 336954 8032 336960 8084
rect 337012 8072 337018 8084
rect 341281 8075 341339 8081
rect 341281 8072 341293 8075
rect 337012 8044 341293 8072
rect 337012 8032 337018 8044
rect 341281 8041 341293 8044
rect 341327 8041 341339 8075
rect 341281 8035 341339 8041
rect 341370 8032 341376 8084
rect 341428 8072 341434 8084
rect 510098 8072 510104 8084
rect 341428 8044 510104 8072
rect 341428 8032 341434 8044
rect 510098 8032 510104 8044
rect 510156 8032 510162 8084
rect 66474 7964 66480 8016
rect 66532 8004 66538 8016
rect 243574 8004 243580 8016
rect 66532 7976 243580 8004
rect 66532 7964 66538 7976
rect 243574 7964 243580 7976
rect 243632 7964 243638 8016
rect 245966 7964 245972 8016
rect 246024 8004 246030 8016
rect 280834 8004 280840 8016
rect 246024 7976 280840 8004
rect 246024 7964 246030 7976
rect 280834 7964 280840 7976
rect 280892 7964 280898 8016
rect 332998 7964 333004 8016
rect 333056 8004 333062 8016
rect 338150 8004 338156 8016
rect 333056 7976 338156 8004
rect 333056 7964 333062 7976
rect 338150 7964 338156 7976
rect 338208 7964 338214 8016
rect 338334 7964 338340 8016
rect 338392 8004 338398 8016
rect 350846 8004 350852 8016
rect 338392 7976 350852 8004
rect 338392 7964 338398 7976
rect 350846 7964 350852 7976
rect 350904 7964 350910 8016
rect 350941 8007 350999 8013
rect 350941 7973 350953 8007
rect 350987 8004 350999 8007
rect 513686 8004 513692 8016
rect 350987 7976 513692 8004
rect 350987 7973 350999 7976
rect 350941 7967 350999 7973
rect 513686 7964 513692 7976
rect 513744 7964 513750 8016
rect 62886 7896 62892 7948
rect 62944 7936 62950 7948
rect 242378 7936 242384 7948
rect 62944 7908 242384 7936
rect 62944 7896 62950 7908
rect 242378 7896 242384 7908
rect 242436 7896 242442 7948
rect 242470 7896 242476 7948
rect 242528 7936 242534 7948
rect 279822 7936 279828 7948
rect 242528 7908 279828 7936
rect 242528 7896 242534 7908
rect 279822 7896 279828 7908
rect 279880 7896 279886 7948
rect 334286 7896 334292 7948
rect 334344 7936 334350 7948
rect 339625 7939 339683 7945
rect 339625 7936 339637 7939
rect 334344 7908 339637 7936
rect 334344 7896 334350 7908
rect 339625 7905 339637 7908
rect 339671 7905 339683 7939
rect 339625 7899 339683 7905
rect 339714 7896 339720 7948
rect 339772 7936 339778 7948
rect 350662 7936 350668 7948
rect 339772 7908 350668 7936
rect 339772 7896 339778 7908
rect 350662 7896 350668 7908
rect 350720 7896 350726 7948
rect 350757 7939 350815 7945
rect 350757 7905 350769 7939
rect 350803 7936 350815 7939
rect 517274 7936 517280 7948
rect 350803 7908 517280 7936
rect 350803 7905 350815 7908
rect 350757 7899 350815 7905
rect 517274 7896 517280 7908
rect 517332 7896 517338 7948
rect 17714 7828 17720 7880
rect 17772 7868 17778 7880
rect 196286 7868 196292 7880
rect 17772 7840 196292 7868
rect 17772 7828 17778 7840
rect 196286 7828 196292 7840
rect 196344 7828 196350 7880
rect 196381 7871 196439 7877
rect 196381 7837 196393 7871
rect 196427 7868 196439 7871
rect 215790 7868 215796 7880
rect 196427 7840 215796 7868
rect 196427 7837 196439 7840
rect 196381 7831 196439 7837
rect 215790 7828 215796 7840
rect 215848 7828 215854 7880
rect 215882 7828 215888 7880
rect 215940 7868 215946 7880
rect 225266 7868 225272 7880
rect 215940 7840 225272 7868
rect 215940 7828 215946 7840
rect 225266 7828 225272 7840
rect 225324 7828 225330 7880
rect 225358 7828 225364 7880
rect 225416 7868 225422 7880
rect 225450 7868 225456 7880
rect 225416 7840 225456 7868
rect 225416 7828 225422 7840
rect 225450 7828 225456 7840
rect 225508 7828 225514 7880
rect 225542 7828 225548 7880
rect 225600 7868 225606 7880
rect 231246 7868 231252 7880
rect 225600 7840 231252 7868
rect 225600 7828 225606 7840
rect 231246 7828 231252 7840
rect 231304 7828 231310 7880
rect 231338 7828 231344 7880
rect 231396 7868 231402 7880
rect 232534 7868 232540 7880
rect 231396 7840 232540 7868
rect 231396 7828 231402 7840
rect 232534 7828 232540 7840
rect 232592 7828 232598 7880
rect 232905 7871 232963 7877
rect 232905 7837 232917 7871
rect 232951 7868 232963 7871
rect 237870 7868 237876 7880
rect 232951 7840 237876 7868
rect 232951 7837 232963 7840
rect 232905 7831 232963 7837
rect 237870 7828 237876 7840
rect 237928 7828 237934 7880
rect 238882 7828 238888 7880
rect 238940 7868 238946 7880
rect 279546 7868 279552 7880
rect 238940 7840 279552 7868
rect 238940 7828 238946 7840
rect 279546 7828 279552 7840
rect 279604 7828 279610 7880
rect 330054 7828 330060 7880
rect 330112 7868 330118 7880
rect 336497 7871 336555 7877
rect 336497 7868 336509 7871
rect 330112 7840 336509 7868
rect 330112 7828 330118 7840
rect 336497 7837 336509 7840
rect 336543 7837 336555 7871
rect 336497 7831 336555 7837
rect 338242 7828 338248 7880
rect 338300 7868 338306 7880
rect 520862 7868 520868 7880
rect 338300 7840 520868 7868
rect 338300 7828 338306 7840
rect 520862 7828 520868 7840
rect 520920 7828 520926 7880
rect 12930 7760 12936 7812
rect 12988 7800 12994 7812
rect 186629 7803 186687 7809
rect 186629 7800 186641 7803
rect 12988 7772 186641 7800
rect 12988 7760 12994 7772
rect 186629 7769 186641 7772
rect 186675 7769 186687 7803
rect 186629 7763 186687 7769
rect 186721 7803 186779 7809
rect 186721 7769 186733 7803
rect 186767 7800 186779 7803
rect 267034 7800 267040 7812
rect 186767 7772 267040 7800
rect 186767 7769 186779 7772
rect 186721 7763 186779 7769
rect 267034 7760 267040 7772
rect 267092 7760 267098 7812
rect 327294 7760 327300 7812
rect 327352 7800 327358 7812
rect 457385 7803 457443 7809
rect 457385 7800 457397 7803
rect 327352 7772 457397 7800
rect 327352 7760 327358 7772
rect 457385 7769 457397 7772
rect 457431 7769 457443 7803
rect 457385 7763 457443 7769
rect 457569 7803 457627 7809
rect 457569 7769 457581 7803
rect 457615 7800 457627 7803
rect 524358 7800 524364 7812
rect 457615 7772 524364 7800
rect 457615 7769 457627 7772
rect 457569 7763 457627 7769
rect 524358 7760 524364 7772
rect 524416 7760 524422 7812
rect 4558 7692 4564 7744
rect 4616 7732 4622 7744
rect 193618 7732 193624 7744
rect 4616 7704 193624 7732
rect 4616 7692 4622 7704
rect 193618 7692 193624 7704
rect 193676 7692 193682 7744
rect 193710 7692 193716 7744
rect 193768 7732 193774 7744
rect 194906 7732 194912 7744
rect 193768 7704 194912 7732
rect 193768 7692 193774 7704
rect 194906 7692 194912 7704
rect 194964 7692 194970 7744
rect 195001 7735 195059 7741
rect 195001 7701 195013 7735
rect 195047 7732 195059 7735
rect 265654 7732 265660 7744
rect 195047 7704 265660 7732
rect 195047 7701 195059 7704
rect 195001 7695 195059 7701
rect 265654 7692 265660 7704
rect 265712 7692 265718 7744
rect 328674 7692 328680 7744
rect 328732 7732 328738 7744
rect 457293 7735 457351 7741
rect 457293 7732 457305 7735
rect 328732 7704 457305 7732
rect 328732 7692 328738 7704
rect 457293 7701 457305 7704
rect 457339 7701 457351 7735
rect 457293 7695 457351 7701
rect 457477 7735 457535 7741
rect 457477 7701 457489 7735
rect 457523 7732 457535 7735
rect 527946 7732 527952 7744
rect 457523 7704 527952 7732
rect 457523 7701 457535 7704
rect 457477 7695 457535 7701
rect 527946 7692 527952 7704
rect 528004 7692 528010 7744
rect 1600 7568 583316 7664
rect 146146 7488 146152 7540
rect 146204 7528 146210 7540
rect 260318 7528 260324 7540
rect 146204 7500 260324 7528
rect 146204 7488 146210 7500
rect 260318 7488 260324 7500
rect 260376 7488 260382 7540
rect 331710 7488 331716 7540
rect 331768 7528 331774 7540
rect 332906 7528 332912 7540
rect 331768 7500 332912 7528
rect 331768 7488 331774 7500
rect 332906 7488 332912 7500
rect 332964 7488 332970 7540
rect 335666 7488 335672 7540
rect 335724 7528 335730 7540
rect 340818 7528 340824 7540
rect 335724 7500 340824 7528
rect 335724 7488 335730 7500
rect 340818 7488 340824 7500
rect 340876 7488 340882 7540
rect 340913 7531 340971 7537
rect 340913 7497 340925 7531
rect 340959 7528 340971 7531
rect 341281 7531 341339 7537
rect 340959 7500 341140 7528
rect 340959 7497 340971 7500
rect 340913 7491 340971 7497
rect 149734 7420 149740 7472
rect 149792 7460 149798 7472
rect 260042 7460 260048 7472
rect 149792 7432 260048 7460
rect 149792 7420 149798 7432
rect 260042 7420 260048 7432
rect 260100 7420 260106 7472
rect 335574 7420 335580 7472
rect 335632 7460 335638 7472
rect 340726 7460 340732 7472
rect 335632 7432 340732 7460
rect 335632 7420 335638 7432
rect 340726 7420 340732 7432
rect 340784 7420 340790 7472
rect 341112 7460 341140 7500
rect 341281 7497 341293 7531
rect 341327 7528 341339 7531
rect 473853 7531 473911 7537
rect 473853 7528 473865 7531
rect 341327 7500 473865 7528
rect 341327 7497 341339 7500
rect 341281 7491 341339 7497
rect 473853 7497 473865 7500
rect 473899 7497 473911 7531
rect 473853 7491 473911 7497
rect 474037 7531 474095 7537
rect 474037 7497 474049 7531
rect 474083 7528 474095 7531
rect 502922 7528 502928 7540
rect 474083 7500 502928 7528
rect 474083 7497 474095 7500
rect 474037 7491 474095 7497
rect 502922 7488 502928 7500
rect 502980 7488 502986 7540
rect 520770 7488 520776 7540
rect 520828 7528 520834 7540
rect 521966 7528 521972 7540
rect 520828 7500 521972 7528
rect 520828 7488 520834 7500
rect 521966 7488 521972 7500
rect 522024 7488 522030 7540
rect 537330 7488 537336 7540
rect 537388 7528 537394 7540
rect 538618 7528 538624 7540
rect 537388 7500 538624 7528
rect 537388 7488 537394 7500
rect 538618 7488 538624 7500
rect 538676 7488 538682 7540
rect 555270 7488 555276 7540
rect 555328 7528 555334 7540
rect 556466 7528 556472 7540
rect 555328 7500 556472 7528
rect 555328 7488 555334 7500
rect 556466 7488 556472 7500
rect 556524 7488 556530 7540
rect 563550 7488 563556 7540
rect 563608 7528 563614 7540
rect 564838 7528 564844 7540
rect 563608 7500 564844 7528
rect 563608 7488 563614 7500
rect 564838 7488 564844 7500
rect 564896 7488 564902 7540
rect 581490 7488 581496 7540
rect 581548 7528 581554 7540
rect 582686 7528 582692 7540
rect 581548 7500 582692 7528
rect 581548 7488 581554 7500
rect 582686 7488 582692 7500
rect 582744 7488 582750 7540
rect 357933 7463 357991 7469
rect 357933 7460 357945 7463
rect 341112 7432 357945 7460
rect 357933 7429 357945 7432
rect 357979 7429 357991 7463
rect 357933 7423 357991 7429
rect 358117 7463 358175 7469
rect 358117 7429 358129 7463
rect 358163 7460 358175 7463
rect 499426 7460 499432 7472
rect 358163 7432 499432 7460
rect 358163 7429 358175 7432
rect 358117 7423 358175 7429
rect 499426 7420 499432 7432
rect 499484 7420 499490 7472
rect 153230 7352 153236 7404
rect 153288 7392 153294 7404
rect 261790 7392 261796 7404
rect 153288 7364 261796 7392
rect 153288 7352 153294 7364
rect 261790 7352 261796 7364
rect 261848 7352 261854 7404
rect 334378 7352 334384 7404
rect 334436 7392 334442 7404
rect 341189 7395 341247 7401
rect 341189 7392 341201 7395
rect 334436 7364 341201 7392
rect 334436 7352 334442 7364
rect 341189 7361 341201 7364
rect 341235 7361 341247 7395
rect 341189 7355 341247 7361
rect 343394 7352 343400 7404
rect 343452 7392 343458 7404
rect 346893 7395 346951 7401
rect 346893 7392 346905 7395
rect 343452 7364 346905 7392
rect 343452 7352 343458 7364
rect 346893 7361 346905 7364
rect 346939 7392 346951 7395
rect 346982 7392 346988 7404
rect 346939 7364 346988 7392
rect 346939 7361 346951 7364
rect 346893 7355 346951 7361
rect 346982 7352 346988 7364
rect 347040 7352 347046 7404
rect 356458 7352 356464 7404
rect 356516 7392 356522 7404
rect 424173 7395 424231 7401
rect 424173 7392 424185 7395
rect 356516 7364 424185 7392
rect 356516 7352 356522 7364
rect 424173 7361 424185 7364
rect 424219 7361 424231 7395
rect 424173 7355 424231 7361
rect 433741 7395 433799 7401
rect 433741 7361 433753 7395
rect 433787 7392 433799 7395
rect 462813 7395 462871 7401
rect 462813 7392 462825 7395
rect 433787 7364 462825 7392
rect 433787 7361 433799 7364
rect 433741 7355 433799 7361
rect 462813 7361 462825 7364
rect 462859 7361 462871 7395
rect 462813 7355 462871 7361
rect 472381 7395 472439 7401
rect 472381 7361 472393 7395
rect 472427 7392 472439 7395
rect 473945 7395 474003 7401
rect 473945 7392 473957 7395
rect 472427 7364 473957 7392
rect 472427 7361 472439 7364
rect 472381 7355 472439 7361
rect 473945 7361 473957 7364
rect 473991 7361 474003 7395
rect 473945 7355 474003 7361
rect 474129 7395 474187 7401
rect 474129 7361 474141 7395
rect 474175 7392 474187 7395
rect 495838 7392 495844 7404
rect 474175 7364 495844 7392
rect 474175 7361 474187 7364
rect 474129 7355 474187 7361
rect 495838 7352 495844 7364
rect 495896 7352 495902 7404
rect 156818 7284 156824 7336
rect 156876 7324 156882 7336
rect 261698 7324 261704 7336
rect 156876 7296 261704 7324
rect 156876 7284 156882 7296
rect 261698 7284 261704 7296
rect 261756 7284 261762 7336
rect 331434 7284 331440 7336
rect 331492 7324 331498 7336
rect 492250 7324 492256 7336
rect 331492 7296 492256 7324
rect 331492 7284 331498 7296
rect 492250 7284 492256 7296
rect 492308 7284 492314 7336
rect 160406 7216 160412 7268
rect 160464 7256 160470 7268
rect 263262 7256 263268 7268
rect 160464 7228 263268 7256
rect 160464 7216 160470 7228
rect 263262 7216 263268 7228
rect 263320 7216 263326 7268
rect 317634 7216 317640 7268
rect 317692 7256 317698 7268
rect 323801 7259 323859 7265
rect 323801 7256 323813 7259
rect 317692 7228 323813 7256
rect 317692 7216 317698 7228
rect 323801 7225 323813 7228
rect 323847 7225 323859 7259
rect 323801 7219 323859 7225
rect 331158 7216 331164 7268
rect 331216 7256 331222 7268
rect 473945 7259 474003 7265
rect 473945 7256 473957 7259
rect 331216 7228 473957 7256
rect 331216 7216 331222 7228
rect 473945 7225 473957 7228
rect 473991 7225 474003 7259
rect 473945 7219 474003 7225
rect 474129 7259 474187 7265
rect 474129 7225 474141 7259
rect 474175 7256 474187 7259
rect 488662 7256 488668 7268
rect 474175 7228 488668 7256
rect 474175 7225 474187 7228
rect 474129 7219 474187 7225
rect 488662 7216 488668 7228
rect 488720 7216 488726 7268
rect 165190 7148 165196 7200
rect 165248 7188 165254 7200
rect 264274 7188 264280 7200
rect 165248 7160 264280 7188
rect 165248 7148 165254 7160
rect 264274 7148 264280 7160
rect 264332 7148 264338 7200
rect 320302 7148 320308 7200
rect 320360 7188 320366 7200
rect 322145 7191 322203 7197
rect 322145 7188 322157 7191
rect 320360 7160 322157 7188
rect 320360 7148 320366 7160
rect 322145 7157 322157 7160
rect 322191 7157 322203 7191
rect 322145 7151 322203 7157
rect 330146 7148 330152 7200
rect 330204 7188 330210 7200
rect 473850 7188 473856 7200
rect 330204 7160 473856 7188
rect 330204 7148 330210 7160
rect 473850 7148 473856 7160
rect 473908 7148 473914 7200
rect 474218 7148 474224 7200
rect 474276 7188 474282 7200
rect 485074 7188 485080 7200
rect 474276 7160 485080 7188
rect 474276 7148 474282 7160
rect 485074 7148 485080 7160
rect 485132 7148 485138 7200
rect 486270 7148 486276 7200
rect 486328 7188 486334 7200
rect 487466 7188 487472 7200
rect 486328 7160 487472 7188
rect 486328 7148 486334 7160
rect 487466 7148 487472 7160
rect 487524 7148 487530 7200
rect 569070 7148 569076 7200
rect 569128 7188 569134 7200
rect 578638 7188 578644 7200
rect 569128 7160 578644 7188
rect 569128 7148 569134 7160
rect 578638 7148 578644 7160
rect 578696 7148 578702 7200
rect 1600 7024 583316 7120
rect 168686 6944 168692 6996
rect 168744 6984 168750 6996
rect 264182 6984 264188 6996
rect 168744 6956 264188 6984
rect 168744 6944 168750 6956
rect 264182 6944 264188 6956
rect 264240 6944 264246 6996
rect 322145 6987 322203 6993
rect 322145 6953 322157 6987
rect 322191 6984 322203 6987
rect 331710 6984 331716 6996
rect 322191 6956 331716 6984
rect 322191 6953 322203 6956
rect 322145 6947 322203 6953
rect 331710 6944 331716 6956
rect 331768 6944 331774 6996
rect 336497 6987 336555 6993
rect 336497 6953 336509 6987
rect 336543 6984 336555 6987
rect 480382 6984 480388 6996
rect 336543 6956 480388 6984
rect 336543 6953 336555 6956
rect 336497 6947 336555 6953
rect 480382 6944 480388 6956
rect 480440 6944 480446 6996
rect 480842 6944 480848 6996
rect 480900 6984 480906 6996
rect 483510 6984 483516 6996
rect 480900 6956 483516 6984
rect 480900 6944 480906 6956
rect 483510 6944 483516 6956
rect 483568 6944 483574 6996
rect 558030 6944 558036 6996
rect 558088 6984 558094 6996
rect 567598 6984 567604 6996
rect 558088 6956 567604 6984
rect 558088 6944 558094 6956
rect 567598 6944 567604 6956
rect 567656 6944 567662 6996
rect 172274 6876 172280 6928
rect 172332 6916 172338 6928
rect 265746 6916 265752 6928
rect 172332 6888 265752 6916
rect 172332 6876 172338 6888
rect 265746 6876 265752 6888
rect 265804 6876 265810 6928
rect 278442 6876 278448 6928
rect 278500 6916 278506 6928
rect 278718 6916 278724 6928
rect 278500 6888 278724 6916
rect 278500 6876 278506 6888
rect 278718 6876 278724 6888
rect 278776 6876 278782 6928
rect 321777 6919 321835 6925
rect 321777 6885 321789 6919
rect 321823 6916 321835 6919
rect 322234 6916 322240 6928
rect 321823 6888 322240 6916
rect 321823 6885 321835 6888
rect 321777 6879 321835 6885
rect 322234 6876 322240 6888
rect 322292 6876 322298 6928
rect 328582 6876 328588 6928
rect 328640 6916 328646 6928
rect 476794 6916 476800 6928
rect 328640 6888 476800 6916
rect 328640 6876 328646 6888
rect 476794 6876 476800 6888
rect 476852 6876 476858 6928
rect 178254 6808 178260 6860
rect 178312 6848 178318 6860
rect 266942 6848 266948 6860
rect 178312 6820 266948 6848
rect 178312 6808 178318 6820
rect 266942 6808 266948 6820
rect 267000 6808 267006 6860
rect 313494 6808 313500 6860
rect 313552 6848 313558 6860
rect 405402 6848 405408 6860
rect 313552 6820 405408 6848
rect 313552 6808 313558 6820
rect 405402 6808 405408 6820
rect 405460 6808 405466 6860
rect 424173 6851 424231 6857
rect 424173 6817 424185 6851
rect 424219 6848 424231 6851
rect 433741 6851 433799 6857
rect 433741 6848 433753 6851
rect 424219 6820 433753 6848
rect 424219 6817 424231 6820
rect 424173 6811 424231 6817
rect 433741 6817 433753 6820
rect 433787 6817 433799 6851
rect 433741 6811 433799 6817
rect 457385 6851 457443 6857
rect 457385 6817 457397 6851
rect 457431 6848 457443 6851
rect 469618 6848 469624 6860
rect 457431 6820 469624 6848
rect 457431 6817 457443 6820
rect 457385 6811 457443 6817
rect 469618 6808 469624 6820
rect 469676 6808 469682 6860
rect 174666 6740 174672 6792
rect 174724 6780 174730 6792
rect 266022 6780 266028 6792
rect 174724 6752 266028 6780
rect 174724 6740 174730 6752
rect 266022 6740 266028 6752
rect 266080 6740 266086 6792
rect 314966 6740 314972 6792
rect 315024 6780 315030 6792
rect 408990 6780 408996 6792
rect 315024 6752 408996 6780
rect 315024 6740 315030 6752
rect 408990 6740 408996 6752
rect 409048 6740 409054 6792
rect 424078 6740 424084 6792
rect 424136 6780 424142 6792
rect 428954 6780 428960 6792
rect 424136 6752 428960 6780
rect 424136 6740 424142 6752
rect 428954 6740 428960 6752
rect 429012 6740 429018 6792
rect 457293 6783 457351 6789
rect 457293 6749 457305 6783
rect 457339 6780 457351 6783
rect 473206 6780 473212 6792
rect 457339 6752 473212 6780
rect 457339 6749 457351 6752
rect 457293 6743 457351 6749
rect 473206 6740 473212 6752
rect 473264 6740 473270 6792
rect 171078 6672 171084 6724
rect 171136 6712 171142 6724
rect 265562 6712 265568 6724
rect 171136 6684 265568 6712
rect 171136 6672 171142 6684
rect 265562 6672 265568 6684
rect 265620 6672 265626 6724
rect 316346 6672 316352 6724
rect 316404 6712 316410 6724
rect 412578 6712 412584 6724
rect 316404 6684 412584 6712
rect 316404 6672 316410 6684
rect 412578 6672 412584 6684
rect 412636 6672 412642 6724
rect 453242 6672 453248 6724
rect 453300 6712 453306 6724
rect 462718 6712 462724 6724
rect 453300 6684 462724 6712
rect 453300 6672 453306 6684
rect 462718 6672 462724 6684
rect 462776 6672 462782 6724
rect 462813 6715 462871 6721
rect 462813 6681 462825 6715
rect 462859 6712 462871 6715
rect 472381 6715 472439 6721
rect 472381 6712 472393 6715
rect 462859 6684 472393 6712
rect 462859 6681 462871 6684
rect 462813 6675 462871 6681
rect 472381 6681 472393 6684
rect 472427 6681 472439 6715
rect 472381 6675 472439 6681
rect 167582 6604 167588 6656
rect 167640 6644 167646 6656
rect 264550 6644 264556 6656
rect 167640 6616 264556 6644
rect 167640 6604 167646 6616
rect 264550 6604 264556 6616
rect 264608 6604 264614 6656
rect 316254 6604 316260 6656
rect 316312 6644 316318 6656
rect 416166 6644 416172 6656
rect 316312 6616 416172 6644
rect 316312 6604 316318 6616
rect 416166 6604 416172 6616
rect 416224 6604 416230 6656
rect 1600 6480 583316 6576
rect 163994 6400 164000 6452
rect 164052 6440 164058 6452
rect 263170 6440 263176 6452
rect 164052 6412 263176 6440
rect 164052 6400 164058 6412
rect 263170 6400 263176 6412
rect 263228 6400 263234 6452
rect 313586 6400 313592 6452
rect 313644 6440 313650 6452
rect 313644 6412 317312 6440
rect 313644 6400 313650 6412
rect 131886 6332 131892 6384
rect 131944 6372 131950 6384
rect 257374 6372 257380 6384
rect 131944 6344 257380 6372
rect 131944 6332 131950 6344
rect 257374 6332 257380 6344
rect 257432 6332 257438 6384
rect 259033 6375 259091 6381
rect 259033 6341 259045 6375
rect 259079 6372 259091 6375
rect 270070 6372 270076 6384
rect 259079 6344 270076 6372
rect 259079 6341 259091 6344
rect 259033 6335 259091 6341
rect 270070 6332 270076 6344
rect 270128 6332 270134 6384
rect 310734 6332 310740 6384
rect 310792 6372 310798 6384
rect 317177 6375 317235 6381
rect 317177 6372 317189 6375
rect 310792 6344 317189 6372
rect 310792 6332 310798 6344
rect 317177 6341 317189 6344
rect 317223 6341 317235 6375
rect 317284 6372 317312 6412
rect 317726 6400 317732 6452
rect 317784 6440 317790 6452
rect 321869 6443 321927 6449
rect 321869 6440 321881 6443
rect 317784 6412 321881 6440
rect 317784 6400 317790 6412
rect 321869 6409 321881 6412
rect 321915 6409 321927 6443
rect 321869 6403 321927 6409
rect 323801 6443 323859 6449
rect 323801 6409 323813 6443
rect 323847 6440 323859 6443
rect 419662 6440 419668 6452
rect 323847 6412 419668 6440
rect 323847 6409 323859 6412
rect 323801 6403 323859 6409
rect 419662 6400 419668 6412
rect 419720 6400 419726 6452
rect 318830 6372 318836 6384
rect 317284 6344 318836 6372
rect 317177 6335 317235 6341
rect 318830 6332 318836 6344
rect 318888 6332 318894 6384
rect 322053 6375 322111 6381
rect 322053 6341 322065 6375
rect 322099 6372 322111 6375
rect 357933 6375 357991 6381
rect 357933 6372 357945 6375
rect 322099 6344 357945 6372
rect 322099 6341 322111 6344
rect 322053 6335 322111 6341
rect 357933 6341 357945 6344
rect 357979 6341 357991 6375
rect 357933 6335 357991 6341
rect 358117 6375 358175 6381
rect 358117 6341 358129 6375
rect 358163 6372 358175 6375
rect 423250 6372 423256 6384
rect 358163 6344 423256 6372
rect 358163 6341 358175 6344
rect 358117 6335 358175 6341
rect 423250 6332 423256 6344
rect 423308 6332 423314 6384
rect 59298 6264 59304 6316
rect 59356 6304 59362 6316
rect 215790 6304 215796 6316
rect 59356 6276 215796 6304
rect 59356 6264 59362 6276
rect 215790 6264 215796 6276
rect 215848 6264 215854 6316
rect 215885 6307 215943 6313
rect 215885 6273 215897 6307
rect 215931 6304 215943 6307
rect 235110 6304 235116 6316
rect 215931 6276 235116 6304
rect 215931 6273 215943 6276
rect 215885 6267 215943 6273
rect 235110 6264 235116 6276
rect 235168 6264 235174 6316
rect 235205 6307 235263 6313
rect 235205 6273 235217 6307
rect 235251 6304 235263 6307
rect 245049 6307 245107 6313
rect 245049 6304 245061 6307
rect 235251 6276 245061 6304
rect 235251 6273 235263 6276
rect 235205 6267 235263 6273
rect 245049 6273 245061 6276
rect 245095 6273 245107 6307
rect 245049 6267 245107 6273
rect 254157 6307 254215 6313
rect 254157 6273 254169 6307
rect 254203 6304 254215 6307
rect 263998 6304 264004 6316
rect 254203 6276 264004 6304
rect 254203 6273 254215 6276
rect 254157 6267 254215 6273
rect 263998 6264 264004 6276
rect 264056 6264 264062 6316
rect 310826 6264 310832 6316
rect 310884 6304 310890 6316
rect 314601 6307 314659 6313
rect 314601 6304 314613 6307
rect 310884 6276 314613 6304
rect 310884 6264 310890 6276
rect 314601 6273 314613 6276
rect 314647 6273 314659 6307
rect 314601 6267 314659 6273
rect 319014 6264 319020 6316
rect 319072 6304 319078 6316
rect 319072 6276 321912 6304
rect 319072 6264 319078 6276
rect 55710 6196 55716 6248
rect 55768 6236 55774 6248
rect 225174 6236 225180 6248
rect 55768 6208 225180 6236
rect 55768 6196 55774 6208
rect 225174 6196 225180 6208
rect 225232 6196 225238 6248
rect 225266 6196 225272 6248
rect 225324 6236 225330 6248
rect 272646 6236 272652 6248
rect 225324 6208 272652 6236
rect 225324 6196 225330 6208
rect 272646 6196 272652 6208
rect 272704 6196 272710 6248
rect 302454 6196 302460 6248
rect 302512 6236 302518 6248
rect 321777 6239 321835 6245
rect 321777 6236 321789 6239
rect 302512 6208 321789 6236
rect 302512 6196 302518 6208
rect 321777 6205 321789 6208
rect 321823 6205 321835 6239
rect 321884 6236 321912 6276
rect 328674 6264 328680 6316
rect 328732 6304 328738 6316
rect 328861 6307 328919 6313
rect 328732 6276 328777 6304
rect 328732 6264 328738 6276
rect 328861 6273 328873 6307
rect 328907 6304 328919 6307
rect 337230 6304 337236 6316
rect 328907 6276 337236 6304
rect 328907 6273 328919 6276
rect 328861 6267 328919 6273
rect 337230 6264 337236 6276
rect 337288 6264 337294 6316
rect 338794 6264 338800 6316
rect 338852 6304 338858 6316
rect 346893 6307 346951 6313
rect 346893 6304 346905 6307
rect 338852 6276 346905 6304
rect 338852 6264 338858 6276
rect 346893 6273 346905 6276
rect 346939 6304 346951 6307
rect 346982 6304 346988 6316
rect 346939 6276 346988 6304
rect 346939 6273 346951 6276
rect 346893 6267 346951 6273
rect 346982 6264 346988 6276
rect 347040 6264 347046 6316
rect 356458 6264 356464 6316
rect 356516 6304 356522 6316
rect 424173 6307 424231 6313
rect 424173 6304 424185 6307
rect 356516 6276 424185 6304
rect 356516 6264 356522 6276
rect 424173 6273 424185 6276
rect 424219 6273 424231 6307
rect 424173 6267 424231 6273
rect 430426 6236 430432 6248
rect 321884 6208 430432 6236
rect 321777 6199 321835 6205
rect 430426 6196 430432 6208
rect 430484 6196 430490 6248
rect 52122 6128 52128 6180
rect 52180 6168 52186 6180
rect 215793 6171 215851 6177
rect 215793 6168 215805 6171
rect 52180 6140 215805 6168
rect 52180 6128 52186 6140
rect 215793 6137 215805 6140
rect 215839 6137 215851 6171
rect 215793 6131 215851 6137
rect 215882 6128 215888 6180
rect 215940 6168 215946 6180
rect 272833 6171 272891 6177
rect 272833 6168 272845 6171
rect 215940 6140 272845 6168
rect 215940 6128 215946 6140
rect 272833 6137 272845 6140
rect 272879 6137 272891 6171
rect 272833 6131 272891 6137
rect 307790 6128 307796 6180
rect 307848 6168 307854 6180
rect 370350 6168 370356 6180
rect 307848 6140 370356 6168
rect 307848 6128 307854 6140
rect 370350 6128 370356 6140
rect 370408 6128 370414 6180
rect 370442 6128 370448 6180
rect 370500 6168 370506 6180
rect 434014 6168 434020 6180
rect 370500 6140 434020 6168
rect 370500 6128 370506 6140
rect 434014 6128 434020 6140
rect 434072 6128 434078 6180
rect 181842 6060 181848 6112
rect 181900 6100 181906 6112
rect 267310 6100 267316 6112
rect 181900 6072 267316 6100
rect 181900 6060 181906 6072
rect 267310 6060 267316 6072
rect 267368 6060 267374 6112
rect 309354 6060 309360 6112
rect 309412 6100 309418 6112
rect 312301 6103 312359 6109
rect 312301 6100 312313 6103
rect 309412 6072 312313 6100
rect 309412 6060 309418 6072
rect 312301 6069 312313 6072
rect 312347 6069 312359 6103
rect 312301 6063 312359 6069
rect 321958 6060 321964 6112
rect 322016 6100 322022 6112
rect 401814 6100 401820 6112
rect 322016 6072 401820 6100
rect 322016 6060 322022 6072
rect 401814 6060 401820 6072
rect 401872 6060 401878 6112
rect 424173 6103 424231 6109
rect 424173 6069 424185 6103
rect 424219 6100 424231 6103
rect 426838 6100 426844 6112
rect 424219 6072 426844 6100
rect 424219 6069 424231 6072
rect 424173 6063 424231 6069
rect 426838 6060 426844 6072
rect 426896 6060 426902 6112
rect 1600 5936 583316 6032
rect 175862 5856 175868 5908
rect 175920 5896 175926 5908
rect 177153 5899 177211 5905
rect 177153 5896 177165 5899
rect 175920 5868 177165 5896
rect 175920 5856 175926 5868
rect 177153 5865 177165 5868
rect 177199 5865 177211 5899
rect 177153 5859 177211 5865
rect 185338 5856 185344 5908
rect 185396 5896 185402 5908
rect 268414 5896 268420 5908
rect 185396 5868 268420 5896
rect 185396 5856 185402 5868
rect 268414 5856 268420 5868
rect 268472 5856 268478 5908
rect 312114 5856 312120 5908
rect 312172 5856 312178 5908
rect 312206 5856 312212 5908
rect 312264 5896 312270 5908
rect 398318 5896 398324 5908
rect 312264 5868 398324 5896
rect 312264 5856 312270 5868
rect 398318 5856 398324 5868
rect 398376 5856 398382 5908
rect 179450 5788 179456 5840
rect 179508 5828 179514 5840
rect 186721 5831 186779 5837
rect 186721 5828 186733 5831
rect 179508 5800 186733 5828
rect 179508 5788 179514 5800
rect 186721 5797 186733 5800
rect 186767 5797 186779 5831
rect 186721 5791 186779 5797
rect 188926 5788 188932 5840
rect 188984 5828 188990 5840
rect 268322 5828 268328 5840
rect 188984 5800 268328 5828
rect 188984 5788 188990 5800
rect 268322 5788 268328 5800
rect 268380 5788 268386 5840
rect 312132 5828 312160 5856
rect 394730 5828 394736 5840
rect 312132 5800 394736 5828
rect 394730 5788 394736 5800
rect 394788 5788 394794 5840
rect 192514 5720 192520 5772
rect 192572 5760 192578 5772
rect 269886 5760 269892 5772
rect 192572 5732 269892 5760
rect 192572 5720 192578 5732
rect 269886 5720 269892 5732
rect 269944 5720 269950 5772
rect 312209 5763 312267 5769
rect 312209 5729 312221 5763
rect 312255 5760 312267 5763
rect 312669 5763 312727 5769
rect 312669 5760 312681 5763
rect 312255 5732 312681 5760
rect 312255 5729 312267 5732
rect 312209 5723 312267 5729
rect 312669 5729 312681 5732
rect 312715 5729 312727 5763
rect 312669 5723 312727 5729
rect 317177 5763 317235 5769
rect 317177 5729 317189 5763
rect 317223 5760 317235 5763
rect 391142 5760 391148 5772
rect 317223 5732 391148 5760
rect 317223 5729 317235 5732
rect 317177 5723 317235 5729
rect 391142 5720 391148 5732
rect 391200 5720 391206 5772
rect 196105 5695 196163 5701
rect 196105 5661 196117 5695
rect 196151 5692 196163 5695
rect 269794 5692 269800 5704
rect 196151 5664 269800 5692
rect 196151 5661 196163 5664
rect 196105 5655 196163 5661
rect 269794 5652 269800 5664
rect 269852 5652 269858 5704
rect 312117 5695 312175 5701
rect 312117 5661 312129 5695
rect 312163 5692 312175 5695
rect 312485 5695 312543 5701
rect 312485 5692 312497 5695
rect 312163 5664 312497 5692
rect 312163 5661 312175 5664
rect 312117 5655 312175 5661
rect 312485 5661 312497 5664
rect 312531 5661 312543 5695
rect 312485 5655 312543 5661
rect 314601 5695 314659 5701
rect 314601 5661 314613 5695
rect 314647 5692 314659 5695
rect 387554 5692 387560 5704
rect 314647 5664 387560 5692
rect 314647 5661 314659 5664
rect 314601 5655 314659 5661
rect 387554 5652 387560 5664
rect 387612 5652 387618 5704
rect 199690 5584 199696 5636
rect 199748 5624 199754 5636
rect 271266 5624 271272 5636
rect 199748 5596 271272 5624
rect 199748 5584 199754 5596
rect 271266 5584 271272 5596
rect 271324 5584 271330 5636
rect 302549 5627 302607 5633
rect 302549 5593 302561 5627
rect 302595 5624 302607 5627
rect 312022 5624 312028 5636
rect 302595 5596 312028 5624
rect 302595 5593 302607 5596
rect 302549 5587 302607 5593
rect 312022 5584 312028 5596
rect 312080 5584 312086 5636
rect 370721 5627 370779 5633
rect 370721 5624 370733 5627
rect 312224 5596 370733 5624
rect 203186 5516 203192 5568
rect 203244 5556 203250 5568
rect 271174 5556 271180 5568
rect 203244 5528 271180 5556
rect 203244 5516 203250 5528
rect 271174 5516 271180 5528
rect 271232 5516 271238 5568
rect 309446 5516 309452 5568
rect 309504 5556 309510 5568
rect 312224 5556 312252 5596
rect 370721 5593 370733 5596
rect 370767 5593 370779 5627
rect 370721 5587 370779 5593
rect 370994 5584 371000 5636
rect 371052 5624 371058 5636
rect 515161 5627 515219 5633
rect 515161 5624 515173 5627
rect 371052 5596 515173 5624
rect 371052 5584 371058 5596
rect 515161 5593 515173 5596
rect 515207 5593 515219 5627
rect 515161 5587 515219 5593
rect 309504 5528 312252 5556
rect 312301 5559 312359 5565
rect 309504 5516 309510 5528
rect 312301 5525 312313 5559
rect 312347 5556 312359 5559
rect 370813 5559 370871 5565
rect 370813 5556 370825 5559
rect 312347 5528 370825 5556
rect 312347 5525 312359 5528
rect 312301 5519 312359 5525
rect 370813 5525 370825 5528
rect 370859 5525 370871 5559
rect 370813 5519 370871 5525
rect 370902 5516 370908 5568
rect 370960 5556 370966 5568
rect 505869 5559 505927 5565
rect 505869 5556 505881 5559
rect 370960 5528 505881 5556
rect 370960 5516 370966 5528
rect 505869 5525 505881 5528
rect 505915 5525 505927 5559
rect 505869 5519 505927 5525
rect 1600 5392 583316 5488
rect 191318 5312 191324 5364
rect 191376 5352 191382 5364
rect 264185 5355 264243 5361
rect 264185 5352 264197 5355
rect 191376 5324 264197 5352
rect 191376 5312 191382 5324
rect 264185 5321 264197 5324
rect 264231 5321 264243 5355
rect 264185 5315 264243 5321
rect 264277 5355 264335 5361
rect 264277 5321 264289 5355
rect 264323 5352 264335 5355
rect 283594 5352 283600 5364
rect 264323 5324 283600 5352
rect 264323 5321 264335 5324
rect 264277 5315 264335 5321
rect 283594 5312 283600 5324
rect 283652 5312 283658 5364
rect 301074 5312 301080 5364
rect 301132 5352 301138 5364
rect 312209 5355 312267 5361
rect 312209 5352 312221 5355
rect 301132 5324 312221 5352
rect 301132 5312 301138 5324
rect 312209 5321 312221 5324
rect 312255 5321 312267 5355
rect 312209 5315 312267 5321
rect 312301 5355 312359 5361
rect 312301 5321 312313 5355
rect 312347 5352 312359 5355
rect 317269 5355 317327 5361
rect 312347 5324 317220 5352
rect 312347 5321 312359 5324
rect 312301 5315 312359 5321
rect 134278 5244 134284 5296
rect 134336 5284 134342 5296
rect 244770 5284 244776 5296
rect 134336 5256 244776 5284
rect 134336 5244 134342 5256
rect 244770 5244 244776 5256
rect 244828 5244 244834 5296
rect 245049 5287 245107 5293
rect 245049 5253 245061 5287
rect 245095 5284 245107 5287
rect 254157 5287 254215 5293
rect 254157 5284 254169 5287
rect 245095 5256 254169 5284
rect 245095 5253 245107 5256
rect 245049 5247 245107 5253
rect 254157 5253 254169 5256
rect 254203 5253 254215 5287
rect 259217 5287 259275 5293
rect 259217 5284 259229 5287
rect 254157 5247 254215 5253
rect 254264 5256 259229 5284
rect 130690 5176 130696 5228
rect 130748 5216 130754 5228
rect 244862 5216 244868 5228
rect 130748 5188 244868 5216
rect 130748 5176 130754 5188
rect 244862 5176 244868 5188
rect 244920 5176 244926 5228
rect 244954 5176 244960 5228
rect 245012 5216 245018 5228
rect 254264 5216 254292 5256
rect 259217 5253 259229 5256
rect 259263 5253 259275 5287
rect 263909 5287 263967 5293
rect 263909 5284 263921 5287
rect 259217 5247 259275 5253
rect 259324 5256 263921 5284
rect 245012 5188 254292 5216
rect 254341 5219 254399 5225
rect 245012 5176 245018 5188
rect 254341 5185 254353 5219
rect 254387 5216 254399 5219
rect 259324 5216 259352 5256
rect 263909 5253 263921 5256
rect 263955 5253 263967 5287
rect 263909 5247 263967 5253
rect 263998 5244 264004 5296
rect 264056 5284 264062 5296
rect 278258 5284 278264 5296
rect 264056 5256 278264 5284
rect 264056 5244 264062 5256
rect 278258 5244 278264 5256
rect 278316 5244 278322 5296
rect 299786 5244 299792 5296
rect 299844 5284 299850 5296
rect 302549 5287 302607 5293
rect 302549 5284 302561 5287
rect 299844 5256 302561 5284
rect 299844 5244 299850 5256
rect 302549 5253 302561 5256
rect 302595 5253 302607 5287
rect 302549 5247 302607 5253
rect 302641 5287 302699 5293
rect 302641 5253 302653 5287
rect 302687 5284 302699 5287
rect 312574 5284 312580 5296
rect 302687 5256 312580 5284
rect 302687 5253 302699 5256
rect 302641 5247 302699 5253
rect 312574 5244 312580 5256
rect 312632 5244 312638 5296
rect 312669 5287 312727 5293
rect 312669 5253 312681 5287
rect 312715 5284 312727 5287
rect 317085 5287 317143 5293
rect 317085 5284 317097 5287
rect 312715 5256 317097 5284
rect 312715 5253 312727 5256
rect 312669 5247 312727 5253
rect 317085 5253 317097 5256
rect 317131 5253 317143 5287
rect 317192 5284 317220 5324
rect 317269 5321 317281 5355
rect 317315 5352 317327 5355
rect 341186 5352 341192 5364
rect 317315 5324 341192 5352
rect 317315 5321 317327 5324
rect 317269 5315 317327 5321
rect 341186 5312 341192 5324
rect 341244 5312 341250 5364
rect 341373 5355 341431 5361
rect 341373 5321 341385 5355
rect 341419 5352 341431 5355
rect 346341 5355 346399 5361
rect 346341 5352 346353 5355
rect 341419 5324 346353 5352
rect 341419 5321 341431 5324
rect 341373 5315 341431 5321
rect 346341 5321 346353 5324
rect 346387 5321 346399 5355
rect 346341 5315 346399 5321
rect 346433 5355 346491 5361
rect 346433 5321 346445 5355
rect 346479 5352 346491 5355
rect 548186 5352 548192 5364
rect 346479 5324 548192 5352
rect 346479 5321 346491 5324
rect 346433 5315 346491 5321
rect 548186 5312 548192 5324
rect 548244 5312 548250 5364
rect 332449 5287 332507 5293
rect 332449 5284 332461 5287
rect 317192 5256 332461 5284
rect 317085 5247 317143 5253
rect 332449 5253 332461 5256
rect 332495 5253 332507 5287
rect 332449 5247 332507 5253
rect 338058 5244 338064 5296
rect 338116 5284 338122 5296
rect 341281 5287 341339 5293
rect 341281 5284 341293 5287
rect 338116 5256 341293 5284
rect 338116 5244 338122 5256
rect 341281 5253 341293 5256
rect 341327 5253 341339 5287
rect 341281 5247 341339 5253
rect 343578 5244 343584 5296
rect 343636 5284 343642 5296
rect 345329 5287 345387 5293
rect 345329 5284 345341 5287
rect 343636 5256 345341 5284
rect 343636 5244 343642 5256
rect 345329 5253 345341 5256
rect 345375 5253 345387 5287
rect 345329 5247 345387 5253
rect 345418 5244 345424 5296
rect 345476 5284 345482 5296
rect 346065 5287 346123 5293
rect 346065 5284 346077 5287
rect 345476 5256 346077 5284
rect 345476 5244 345482 5256
rect 346065 5253 346077 5256
rect 346111 5253 346123 5287
rect 551682 5284 551688 5296
rect 346065 5247 346123 5253
rect 346172 5256 551688 5284
rect 254387 5188 259352 5216
rect 259401 5219 259459 5225
rect 254387 5185 254399 5188
rect 254341 5179 254399 5185
rect 259401 5185 259413 5219
rect 259447 5216 259459 5219
rect 278718 5216 278724 5228
rect 259447 5188 278724 5216
rect 259447 5185 259459 5188
rect 259401 5179 259459 5185
rect 278718 5176 278724 5188
rect 278776 5176 278782 5228
rect 296750 5176 296756 5228
rect 296808 5216 296814 5228
rect 312393 5219 312451 5225
rect 312393 5216 312405 5219
rect 296808 5188 312405 5216
rect 296808 5176 296814 5188
rect 312393 5185 312405 5188
rect 312439 5185 312451 5219
rect 312393 5179 312451 5185
rect 312485 5219 312543 5225
rect 312485 5185 312497 5219
rect 312531 5216 312543 5219
rect 345970 5216 345976 5228
rect 312531 5188 345976 5216
rect 312531 5185 312543 5188
rect 312485 5179 312543 5185
rect 345970 5176 345976 5188
rect 346028 5176 346034 5228
rect 8146 5108 8152 5160
rect 8204 5148 8210 5160
rect 226922 5148 226928 5160
rect 8204 5120 226928 5148
rect 8204 5108 8210 5120
rect 226922 5108 226928 5120
rect 226980 5108 226986 5160
rect 227014 5108 227020 5160
rect 227072 5148 227078 5160
rect 276510 5148 276516 5160
rect 227072 5120 276516 5148
rect 227072 5108 227078 5120
rect 276510 5108 276516 5120
rect 276568 5108 276574 5160
rect 296842 5108 296848 5160
rect 296900 5148 296906 5160
rect 301169 5151 301227 5157
rect 301169 5148 301181 5151
rect 296900 5120 301181 5148
rect 296900 5108 296906 5120
rect 301169 5117 301181 5120
rect 301215 5117 301227 5151
rect 301169 5111 301227 5117
rect 301258 5108 301264 5160
rect 301316 5148 301322 5160
rect 302730 5148 302736 5160
rect 301316 5120 302736 5148
rect 301316 5108 301322 5120
rect 302730 5108 302736 5120
rect 302788 5108 302794 5160
rect 302825 5151 302883 5157
rect 302825 5117 302837 5151
rect 302871 5148 302883 5151
rect 307425 5151 307483 5157
rect 307425 5148 307437 5151
rect 302871 5120 307437 5148
rect 302871 5117 302883 5120
rect 302825 5111 302883 5117
rect 307425 5117 307437 5120
rect 307471 5117 307483 5151
rect 307425 5111 307483 5117
rect 307514 5108 307520 5160
rect 307572 5148 307578 5160
rect 317269 5151 317327 5157
rect 317269 5148 317281 5151
rect 307572 5120 317281 5148
rect 307572 5108 307578 5120
rect 317269 5117 317281 5120
rect 317315 5117 317327 5151
rect 317269 5111 317327 5117
rect 317361 5151 317419 5157
rect 317361 5117 317373 5151
rect 317407 5148 317419 5151
rect 332357 5151 332415 5157
rect 332357 5148 332369 5151
rect 317407 5120 332369 5148
rect 317407 5117 317419 5120
rect 317361 5111 317419 5117
rect 332357 5117 332369 5120
rect 332403 5117 332415 5151
rect 332357 5111 332415 5117
rect 332449 5151 332507 5157
rect 332449 5117 332461 5151
rect 332495 5148 332507 5151
rect 342382 5148 342388 5160
rect 332495 5120 342388 5148
rect 332495 5117 332507 5120
rect 332449 5111 332507 5117
rect 342382 5108 342388 5120
rect 342440 5108 342446 5160
rect 343946 5108 343952 5160
rect 344004 5148 344010 5160
rect 346172 5148 346200 5256
rect 551682 5244 551688 5256
rect 551740 5244 551746 5296
rect 555270 5216 555276 5228
rect 346356 5188 555276 5216
rect 344004 5120 346200 5148
rect 346249 5151 346307 5157
rect 344004 5108 344010 5120
rect 346249 5117 346261 5151
rect 346295 5148 346307 5151
rect 346356 5148 346384 5188
rect 555270 5176 555276 5188
rect 555328 5176 555334 5228
rect 346295 5120 346384 5148
rect 346295 5117 346307 5120
rect 346249 5111 346307 5117
rect 346798 5108 346804 5160
rect 346856 5148 346862 5160
rect 350846 5148 350852 5160
rect 346856 5120 350852 5148
rect 346856 5108 346862 5120
rect 350846 5108 350852 5120
rect 350904 5108 350910 5160
rect 350938 5108 350944 5160
rect 350996 5148 351002 5160
rect 558858 5148 558864 5160
rect 350996 5120 558864 5148
rect 350996 5108 351002 5120
rect 558858 5108 558864 5120
rect 558916 5108 558922 5160
rect 2166 5040 2172 5092
rect 2224 5080 2230 5092
rect 220669 5083 220727 5089
rect 2224 5052 220620 5080
rect 2224 5040 2230 5052
rect 3362 4972 3368 5024
rect 3420 5012 3426 5024
rect 220485 5015 220543 5021
rect 220485 5012 220497 5015
rect 3420 4984 220497 5012
rect 3420 4972 3426 4984
rect 220485 4981 220497 4984
rect 220531 4981 220543 5015
rect 220592 5012 220620 5052
rect 220669 5049 220681 5083
rect 220715 5080 220727 5083
rect 227569 5083 227627 5089
rect 227569 5080 227581 5083
rect 220715 5052 227581 5080
rect 220715 5049 220727 5052
rect 220669 5043 220727 5049
rect 227569 5049 227581 5052
rect 227615 5049 227627 5083
rect 229317 5083 229375 5089
rect 229317 5080 229329 5083
rect 227569 5043 227627 5049
rect 227676 5052 229329 5080
rect 227676 5012 227704 5052
rect 229317 5049 229329 5052
rect 229363 5049 229375 5083
rect 229317 5043 229375 5049
rect 229409 5083 229467 5089
rect 229409 5049 229421 5083
rect 229455 5080 229467 5083
rect 275682 5080 275688 5092
rect 229455 5052 275688 5080
rect 229455 5049 229467 5052
rect 229409 5043 229467 5049
rect 275682 5040 275688 5052
rect 275740 5040 275746 5092
rect 295646 5040 295652 5092
rect 295704 5080 295710 5092
rect 302549 5083 302607 5089
rect 302549 5080 302561 5083
rect 295704 5052 302561 5080
rect 295704 5040 295710 5052
rect 302549 5049 302561 5052
rect 302595 5049 302607 5083
rect 302549 5043 302607 5049
rect 302638 5040 302644 5092
rect 302696 5080 302702 5092
rect 312117 5083 312175 5089
rect 312117 5080 312129 5083
rect 302696 5052 312129 5080
rect 302696 5040 302702 5052
rect 312117 5049 312129 5052
rect 312163 5049 312175 5083
rect 312117 5043 312175 5049
rect 312206 5040 312212 5092
rect 312264 5080 312270 5092
rect 331710 5080 331716 5092
rect 312264 5052 331716 5080
rect 312264 5040 312270 5052
rect 331710 5040 331716 5052
rect 331768 5040 331774 5092
rect 342566 5040 342572 5092
rect 342624 5080 342630 5092
rect 345326 5080 345332 5092
rect 342624 5052 345332 5080
rect 342624 5040 342630 5052
rect 345326 5040 345332 5052
rect 345384 5040 345390 5092
rect 345421 5083 345479 5089
rect 345421 5049 345433 5083
rect 345467 5080 345479 5083
rect 505777 5083 505835 5089
rect 505777 5080 505789 5083
rect 345467 5052 505789 5080
rect 345467 5049 345479 5052
rect 345421 5043 345479 5049
rect 505777 5049 505789 5052
rect 505823 5049 505835 5083
rect 505777 5043 505835 5049
rect 505869 5083 505927 5089
rect 505869 5049 505881 5083
rect 505915 5080 505927 5083
rect 562446 5080 562452 5092
rect 505915 5052 562452 5080
rect 505915 5049 505927 5052
rect 505869 5043 505927 5049
rect 562446 5040 562452 5052
rect 562504 5040 562510 5092
rect 220592 4984 227704 5012
rect 227753 5015 227811 5021
rect 220485 4975 220543 4981
rect 227753 4981 227765 5015
rect 227799 5012 227811 5015
rect 229682 5012 229688 5024
rect 227799 4984 229688 5012
rect 227799 4981 227811 4984
rect 227753 4975 227811 4981
rect 229682 4972 229688 4984
rect 229740 4972 229746 5024
rect 229777 5015 229835 5021
rect 229777 4981 229789 5015
rect 229823 5012 229835 5015
rect 230142 5012 230148 5024
rect 229823 4984 230148 5012
rect 229823 4981 229835 4984
rect 229777 4975 229835 4981
rect 230142 4972 230148 4984
rect 230200 4972 230206 5024
rect 230602 4972 230608 5024
rect 230660 5012 230666 5024
rect 276970 5012 276976 5024
rect 230660 4984 276976 5012
rect 230660 4972 230666 4984
rect 276970 4972 276976 4984
rect 277028 4972 277034 5024
rect 300982 4972 300988 5024
rect 301040 5012 301046 5024
rect 307514 5012 307520 5024
rect 301040 4984 307520 5012
rect 301040 4972 301046 4984
rect 307514 4972 307520 4984
rect 307572 4972 307578 5024
rect 307609 5015 307667 5021
rect 307609 4981 307621 5015
rect 307655 5012 307667 5015
rect 335206 5012 335212 5024
rect 307655 4984 335212 5012
rect 307655 4981 307667 4984
rect 307609 4975 307667 4981
rect 335206 4972 335212 4984
rect 335264 4972 335270 5024
rect 335758 4972 335764 5024
rect 335816 5012 335822 5024
rect 505593 5015 505651 5021
rect 505593 5012 505605 5015
rect 335816 4984 505605 5012
rect 335816 4972 335822 4984
rect 505593 4981 505605 4984
rect 505639 4981 505651 5015
rect 505593 4975 505651 4981
rect 505685 5015 505743 5021
rect 505685 4981 505697 5015
rect 505731 5012 505743 5015
rect 515069 5015 515127 5021
rect 515069 5012 515081 5015
rect 505731 4984 515081 5012
rect 505731 4981 505743 4984
rect 505685 4975 505743 4981
rect 515069 4981 515081 4984
rect 515115 4981 515127 5015
rect 515069 4975 515127 4981
rect 515161 5015 515219 5021
rect 515161 4981 515173 5015
rect 515207 5012 515219 5015
rect 566034 5012 566040 5024
rect 515207 4984 566040 5012
rect 515207 4981 515219 4984
rect 515161 4975 515219 4981
rect 566034 4972 566040 4984
rect 566092 4972 566098 5024
rect 1600 4848 583316 4944
rect 1062 4768 1068 4820
rect 1120 4808 1126 4820
rect 220669 4811 220727 4817
rect 220669 4808 220681 4811
rect 1120 4780 220681 4808
rect 1120 4768 1126 4780
rect 220669 4777 220681 4780
rect 220715 4777 220727 4811
rect 220669 4771 220727 4777
rect 220761 4811 220819 4817
rect 220761 4777 220773 4811
rect 220807 4808 220819 4811
rect 225266 4808 225272 4820
rect 220807 4780 225272 4808
rect 220807 4777 220819 4780
rect 220761 4771 220819 4777
rect 225266 4768 225272 4780
rect 225324 4768 225330 4820
rect 225358 4768 225364 4820
rect 225416 4808 225422 4820
rect 275222 4808 275228 4820
rect 225416 4780 275228 4808
rect 225416 4768 225422 4780
rect 275222 4768 275228 4780
rect 275280 4768 275286 4820
rect 296934 4768 296940 4820
rect 296992 4808 296998 4820
rect 301077 4811 301135 4817
rect 301077 4808 301089 4811
rect 296992 4780 301089 4808
rect 296992 4768 296998 4780
rect 301077 4777 301089 4780
rect 301123 4777 301135 4811
rect 301077 4771 301135 4777
rect 301166 4768 301172 4820
rect 301224 4808 301230 4820
rect 302733 4811 302791 4817
rect 302733 4808 302745 4811
rect 301224 4780 302745 4808
rect 301224 4768 301230 4780
rect 302733 4777 302745 4780
rect 302779 4777 302791 4811
rect 302733 4771 302791 4777
rect 302825 4811 302883 4817
rect 302825 4777 302837 4811
rect 302871 4808 302883 4811
rect 321958 4808 321964 4820
rect 302871 4780 321964 4808
rect 302871 4777 302883 4780
rect 302825 4771 302883 4777
rect 321958 4768 321964 4780
rect 322016 4768 322022 4820
rect 322142 4768 322148 4820
rect 322200 4808 322206 4820
rect 337598 4808 337604 4820
rect 322200 4780 337604 4808
rect 322200 4768 322206 4780
rect 337598 4768 337604 4780
rect 337656 4768 337662 4820
rect 339806 4768 339812 4820
rect 339864 4808 339870 4820
rect 346249 4811 346307 4817
rect 346249 4808 346261 4811
rect 339864 4780 346261 4808
rect 339864 4768 339870 4780
rect 346249 4777 346261 4780
rect 346295 4777 346307 4811
rect 346249 4771 346307 4777
rect 346341 4811 346399 4817
rect 346341 4777 346353 4811
rect 346387 4808 346399 4811
rect 515250 4808 515256 4820
rect 346387 4780 515256 4808
rect 346387 4777 346399 4780
rect 346341 4771 346399 4777
rect 515250 4768 515256 4780
rect 515308 4768 515314 4820
rect 515342 4768 515348 4820
rect 515400 4808 515406 4820
rect 526750 4808 526756 4820
rect 515400 4780 526756 4808
rect 515400 4768 515406 4780
rect 526750 4768 526756 4780
rect 526808 4768 526814 4820
rect 529513 4811 529571 4817
rect 529513 4777 529525 4811
rect 529559 4808 529571 4811
rect 534573 4811 534631 4817
rect 534573 4808 534585 4811
rect 529559 4780 534585 4808
rect 529559 4777 529571 4780
rect 529513 4771 529571 4777
rect 534573 4777 534585 4780
rect 534619 4777 534631 4811
rect 534573 4771 534631 4777
rect 194998 4700 195004 4752
rect 195056 4740 195062 4752
rect 259033 4743 259091 4749
rect 259033 4740 259045 4743
rect 195056 4712 259045 4740
rect 195056 4700 195062 4712
rect 259033 4709 259045 4712
rect 259079 4709 259091 4743
rect 259033 4703 259091 4709
rect 259122 4700 259128 4752
rect 259180 4740 259186 4752
rect 263909 4743 263967 4749
rect 263909 4740 263921 4743
rect 259180 4712 263921 4740
rect 259180 4700 259186 4712
rect 263909 4709 263921 4712
rect 263955 4709 263967 4743
rect 263909 4703 263967 4709
rect 264001 4743 264059 4749
rect 264001 4709 264013 4743
rect 264047 4740 264059 4743
rect 279362 4740 279368 4752
rect 264047 4712 279368 4740
rect 264047 4709 264059 4712
rect 264001 4703 264059 4709
rect 279362 4700 279368 4712
rect 279420 4700 279426 4752
rect 297026 4700 297032 4752
rect 297084 4740 297090 4752
rect 312393 4743 312451 4749
rect 312393 4740 312405 4743
rect 297084 4712 312405 4740
rect 297084 4700 297090 4712
rect 312393 4709 312405 4712
rect 312439 4709 312451 4743
rect 312393 4703 312451 4709
rect 312485 4743 312543 4749
rect 312485 4709 312497 4743
rect 312531 4740 312543 4743
rect 338794 4740 338800 4752
rect 312531 4712 338800 4740
rect 312531 4709 312543 4712
rect 312485 4703 312543 4709
rect 338794 4700 338800 4712
rect 338852 4700 338858 4752
rect 340910 4700 340916 4752
rect 340968 4740 340974 4752
rect 340968 4712 345556 4740
rect 340968 4700 340974 4712
rect 198494 4632 198500 4684
rect 198552 4672 198558 4684
rect 264553 4675 264611 4681
rect 198552 4644 264412 4672
rect 198552 4632 198558 4644
rect 201990 4564 201996 4616
rect 202048 4604 202054 4616
rect 264274 4604 264280 4616
rect 202048 4576 264280 4604
rect 202048 4564 202054 4576
rect 264274 4564 264280 4576
rect 264332 4564 264338 4616
rect 264384 4604 264412 4644
rect 264553 4641 264565 4675
rect 264599 4672 264611 4675
rect 283502 4672 283508 4684
rect 264599 4644 283508 4672
rect 264599 4641 264611 4644
rect 264553 4635 264611 4641
rect 283502 4632 283508 4644
rect 283560 4632 283566 4684
rect 299878 4632 299884 4684
rect 299936 4672 299942 4684
rect 307609 4675 307667 4681
rect 307609 4672 307621 4675
rect 299936 4644 307621 4672
rect 299936 4632 299942 4644
rect 307609 4641 307621 4644
rect 307655 4641 307667 4675
rect 307609 4635 307667 4641
rect 307701 4675 307759 4681
rect 307701 4641 307713 4675
rect 307747 4672 307759 4675
rect 312209 4675 312267 4681
rect 312209 4672 312221 4675
rect 307747 4644 312221 4672
rect 307747 4641 307759 4644
rect 307701 4635 307759 4641
rect 312209 4641 312221 4644
rect 312255 4641 312267 4675
rect 312209 4635 312267 4641
rect 312298 4632 312304 4684
rect 312356 4672 312362 4684
rect 334102 4672 334108 4684
rect 312356 4644 334108 4672
rect 312356 4632 312362 4644
rect 334102 4632 334108 4644
rect 334160 4632 334166 4684
rect 337138 4632 337144 4684
rect 337196 4672 337202 4684
rect 345421 4675 345479 4681
rect 345421 4672 345433 4675
rect 337196 4644 345433 4672
rect 337196 4632 337202 4644
rect 345421 4641 345433 4644
rect 345467 4641 345479 4675
rect 345421 4635 345479 4641
rect 267497 4607 267555 4613
rect 267497 4604 267509 4607
rect 264384 4576 267509 4604
rect 267497 4573 267509 4576
rect 267543 4573 267555 4607
rect 267497 4567 267555 4573
rect 268877 4607 268935 4613
rect 268877 4573 268889 4607
rect 268923 4604 268935 4607
rect 274118 4604 274124 4616
rect 268923 4576 274124 4604
rect 268923 4573 268935 4576
rect 268877 4567 268935 4573
rect 274118 4564 274124 4576
rect 274176 4564 274182 4616
rect 299694 4564 299700 4616
rect 299752 4604 299758 4616
rect 302733 4607 302791 4613
rect 302733 4604 302745 4607
rect 299752 4576 302745 4604
rect 299752 4564 299758 4576
rect 302733 4573 302745 4576
rect 302779 4573 302791 4607
rect 330514 4604 330520 4616
rect 302733 4567 302791 4573
rect 302932 4576 330520 4604
rect 205578 4496 205584 4548
rect 205636 4536 205642 4548
rect 264366 4536 264372 4548
rect 205636 4508 264372 4536
rect 205636 4496 205642 4508
rect 264366 4496 264372 4508
rect 264424 4496 264430 4548
rect 264461 4539 264519 4545
rect 264461 4505 264473 4539
rect 264507 4536 264519 4539
rect 269702 4536 269708 4548
rect 264507 4508 269708 4536
rect 264507 4505 264519 4508
rect 264461 4499 264519 4505
rect 269702 4496 269708 4508
rect 269760 4496 269766 4548
rect 269794 4496 269800 4548
rect 269852 4536 269858 4548
rect 272462 4536 272468 4548
rect 269852 4508 272468 4536
rect 269852 4496 269858 4508
rect 272462 4496 272468 4508
rect 272520 4496 272526 4548
rect 298406 4496 298412 4548
rect 298464 4536 298470 4548
rect 302546 4536 302552 4548
rect 298464 4508 302552 4536
rect 298464 4496 298470 4508
rect 302546 4496 302552 4508
rect 302604 4496 302610 4548
rect 302641 4539 302699 4545
rect 302641 4505 302653 4539
rect 302687 4536 302699 4539
rect 302822 4536 302828 4548
rect 302687 4508 302828 4536
rect 302687 4505 302699 4508
rect 302641 4499 302699 4505
rect 302822 4496 302828 4508
rect 302880 4496 302886 4548
rect 209166 4428 209172 4480
rect 209224 4468 209230 4480
rect 264182 4468 264188 4480
rect 209224 4440 264188 4468
rect 209224 4428 209230 4440
rect 264182 4428 264188 4440
rect 264240 4428 264246 4480
rect 264274 4428 264280 4480
rect 264332 4468 264338 4480
rect 267405 4471 267463 4477
rect 267405 4468 267417 4471
rect 264332 4440 267417 4468
rect 264332 4428 264338 4440
rect 267405 4437 267417 4440
rect 267451 4437 267463 4471
rect 267405 4431 267463 4437
rect 267497 4471 267555 4477
rect 267497 4437 267509 4471
rect 267543 4468 267555 4471
rect 270990 4468 270996 4480
rect 267543 4440 270996 4468
rect 267543 4437 267555 4440
rect 267497 4431 267555 4437
rect 270990 4428 270996 4440
rect 271048 4428 271054 4480
rect 298498 4428 298504 4480
rect 298556 4468 298562 4480
rect 302932 4468 302960 4576
rect 330514 4564 330520 4576
rect 330572 4564 330578 4616
rect 332357 4607 332415 4613
rect 332357 4573 332369 4607
rect 332403 4604 332415 4607
rect 344774 4604 344780 4616
rect 332403 4576 344780 4604
rect 332403 4573 332415 4576
rect 332357 4567 332415 4573
rect 344774 4564 344780 4576
rect 344832 4564 344838 4616
rect 345528 4604 345556 4712
rect 347902 4700 347908 4752
rect 347960 4740 347966 4752
rect 350570 4740 350576 4752
rect 347960 4712 350576 4740
rect 347960 4700 347966 4712
rect 350570 4700 350576 4712
rect 350628 4700 350634 4752
rect 350938 4700 350944 4752
rect 350996 4740 351002 4752
rect 544598 4740 544604 4752
rect 350996 4712 544604 4740
rect 350996 4700 351002 4712
rect 544598 4700 544604 4712
rect 544656 4700 544662 4752
rect 559413 4743 559471 4749
rect 559413 4709 559425 4743
rect 559459 4709 559471 4743
rect 559413 4703 559471 4709
rect 559505 4743 559563 4749
rect 559505 4709 559517 4743
rect 559551 4740 559563 4743
rect 569530 4740 569536 4752
rect 559551 4712 569536 4740
rect 559551 4709 559563 4712
rect 559505 4703 559563 4709
rect 346706 4632 346712 4684
rect 346764 4672 346770 4684
rect 350662 4672 350668 4684
rect 346764 4644 350668 4672
rect 346764 4632 346770 4644
rect 350662 4632 350668 4644
rect 350720 4632 350726 4684
rect 350846 4632 350852 4684
rect 350904 4672 350910 4684
rect 534573 4675 534631 4681
rect 350904 4644 529740 4672
rect 350904 4632 350910 4644
rect 529605 4607 529663 4613
rect 529605 4604 529617 4607
rect 345528 4576 529617 4604
rect 529605 4573 529617 4576
rect 529651 4573 529663 4607
rect 529712 4604 529740 4644
rect 534573 4641 534585 4675
rect 534619 4672 534631 4675
rect 538713 4675 538771 4681
rect 538713 4672 538725 4675
rect 534619 4644 538725 4672
rect 534619 4641 534631 4644
rect 534573 4635 534631 4641
rect 538713 4641 538725 4644
rect 538759 4641 538771 4675
rect 538713 4635 538771 4641
rect 549845 4675 549903 4681
rect 549845 4641 549857 4675
rect 549891 4672 549903 4675
rect 559428 4672 559456 4703
rect 569530 4700 569536 4712
rect 569588 4700 569594 4752
rect 549891 4644 559456 4672
rect 549891 4641 549903 4644
rect 549845 4635 549903 4641
rect 541010 4604 541016 4616
rect 529712 4576 541016 4604
rect 529605 4567 529663 4573
rect 541010 4564 541016 4576
rect 541068 4564 541074 4616
rect 548281 4607 548339 4613
rect 548281 4573 548293 4607
rect 548327 4604 548339 4607
rect 549753 4607 549811 4613
rect 549753 4604 549765 4607
rect 548327 4576 549765 4604
rect 548327 4573 548339 4576
rect 548281 4567 548339 4573
rect 549753 4573 549765 4576
rect 549799 4573 549811 4607
rect 549753 4567 549811 4573
rect 303098 4496 303104 4548
rect 303156 4536 303162 4548
rect 328122 4536 328128 4548
rect 303156 4508 328128 4536
rect 303156 4496 303162 4508
rect 328122 4496 328128 4508
rect 328180 4496 328186 4548
rect 341373 4539 341431 4545
rect 341373 4505 341385 4539
rect 341419 4536 341431 4539
rect 345605 4539 345663 4545
rect 345605 4536 345617 4539
rect 341419 4508 345617 4536
rect 341419 4505 341431 4508
rect 341373 4499 341431 4505
rect 345605 4505 345617 4508
rect 345651 4505 345663 4539
rect 345605 4499 345663 4505
rect 346525 4539 346583 4545
rect 346525 4505 346537 4539
rect 346571 4536 346583 4539
rect 533926 4536 533932 4548
rect 346571 4508 533932 4536
rect 346571 4505 346583 4508
rect 346525 4499 346583 4505
rect 533926 4496 533932 4508
rect 533984 4496 533990 4548
rect 298556 4440 302960 4468
rect 298556 4428 298562 4440
rect 303006 4428 303012 4480
rect 303064 4468 303070 4480
rect 326926 4468 326932 4480
rect 303064 4440 326932 4468
rect 303064 4428 303070 4440
rect 326926 4428 326932 4440
rect 326984 4428 326990 4480
rect 346157 4471 346215 4477
rect 346157 4437 346169 4471
rect 346203 4468 346215 4471
rect 530338 4468 530344 4480
rect 346203 4440 530344 4468
rect 346203 4437 346215 4440
rect 346157 4431 346215 4437
rect 530338 4428 530344 4440
rect 530396 4428 530402 4480
rect 538713 4471 538771 4477
rect 538713 4437 538725 4471
rect 538759 4468 538771 4471
rect 548281 4471 548339 4477
rect 548281 4468 548293 4471
rect 538759 4440 548293 4468
rect 538759 4437 538771 4440
rect 538713 4431 538771 4437
rect 548281 4437 548293 4440
rect 548327 4437 548339 4471
rect 548281 4431 548339 4437
rect 1600 4304 583316 4400
rect 128850 4224 128856 4276
rect 128908 4264 128914 4276
rect 138789 4267 138847 4273
rect 128908 4236 134416 4264
rect 128908 4224 128914 4236
rect 123333 4199 123391 4205
rect 123333 4165 123345 4199
rect 123379 4196 123391 4199
rect 128945 4199 129003 4205
rect 128945 4196 128957 4199
rect 123379 4168 128957 4196
rect 123379 4165 123391 4168
rect 123333 4159 123391 4165
rect 128945 4165 128957 4168
rect 128991 4165 129003 4199
rect 128945 4159 129003 4165
rect 132993 4199 133051 4205
rect 132993 4165 133005 4199
rect 133039 4196 133051 4199
rect 134281 4199 134339 4205
rect 134281 4196 134293 4199
rect 133039 4168 134293 4196
rect 133039 4165 133051 4168
rect 132993 4159 133051 4165
rect 134281 4165 134293 4168
rect 134327 4165 134339 4199
rect 134388 4196 134416 4236
rect 138789 4233 138801 4267
rect 138835 4264 138847 4267
rect 157741 4267 157799 4273
rect 157741 4264 157753 4267
rect 138835 4236 157753 4264
rect 138835 4233 138847 4236
rect 138789 4227 138847 4233
rect 157741 4233 157753 4236
rect 157787 4233 157799 4267
rect 157741 4227 157799 4233
rect 157833 4267 157891 4273
rect 157833 4233 157845 4267
rect 157879 4264 157891 4267
rect 177429 4267 177487 4273
rect 157879 4236 177380 4264
rect 157879 4233 157891 4236
rect 157833 4227 157891 4233
rect 147897 4199 147955 4205
rect 147897 4196 147909 4199
rect 134388 4168 147909 4196
rect 134281 4159 134339 4165
rect 147897 4165 147909 4168
rect 147943 4165 147955 4199
rect 147897 4159 147955 4165
rect 147989 4199 148047 4205
rect 147989 4165 148001 4199
rect 148035 4196 148047 4199
rect 152221 4199 152279 4205
rect 152221 4196 152233 4199
rect 148035 4168 152233 4196
rect 148035 4165 148047 4168
rect 147989 4159 148047 4165
rect 152221 4165 152233 4168
rect 152267 4165 152279 4199
rect 152221 4159 152279 4165
rect 159121 4199 159179 4205
rect 159121 4165 159133 4199
rect 159167 4196 159179 4199
rect 167585 4199 167643 4205
rect 167585 4196 167597 4199
rect 159167 4168 167597 4196
rect 159167 4165 159179 4168
rect 159121 4159 159179 4165
rect 167585 4165 167597 4168
rect 167631 4165 167643 4199
rect 167585 4159 167643 4165
rect 167677 4199 167735 4205
rect 167677 4165 167689 4199
rect 167723 4196 167735 4199
rect 171449 4199 171507 4205
rect 171449 4196 171461 4199
rect 167723 4168 171461 4196
rect 167723 4165 167735 4168
rect 167677 4159 167735 4165
rect 171449 4165 171461 4168
rect 171495 4165 171507 4199
rect 171449 4159 171507 4165
rect 171725 4199 171783 4205
rect 171725 4165 171737 4199
rect 171771 4196 171783 4199
rect 176877 4199 176935 4205
rect 176877 4196 176889 4199
rect 171771 4168 176889 4196
rect 171771 4165 171783 4168
rect 171725 4159 171783 4165
rect 176877 4165 176889 4168
rect 176923 4165 176935 4199
rect 176877 4159 176935 4165
rect 176969 4199 177027 4205
rect 176969 4165 176981 4199
rect 177015 4196 177027 4199
rect 177245 4199 177303 4205
rect 177245 4196 177257 4199
rect 177015 4168 177257 4196
rect 177015 4165 177027 4168
rect 176969 4159 177027 4165
rect 177245 4165 177257 4168
rect 177291 4165 177303 4199
rect 177352 4196 177380 4236
rect 177429 4233 177441 4267
rect 177475 4264 177487 4267
rect 190953 4267 191011 4273
rect 190953 4264 190965 4267
rect 177475 4236 190965 4264
rect 177475 4233 177487 4236
rect 177429 4227 177487 4233
rect 190953 4233 190965 4236
rect 190999 4233 191011 4267
rect 190953 4227 191011 4233
rect 206133 4267 206191 4273
rect 206133 4233 206145 4267
rect 206179 4264 206191 4267
rect 215885 4267 215943 4273
rect 215885 4264 215897 4267
rect 206179 4236 215897 4264
rect 206179 4233 206191 4236
rect 206133 4227 206191 4233
rect 215885 4233 215897 4236
rect 215931 4233 215943 4267
rect 215885 4227 215943 4233
rect 217449 4267 217507 4273
rect 217449 4233 217461 4267
rect 217495 4264 217507 4267
rect 218553 4267 218611 4273
rect 218553 4264 218565 4267
rect 217495 4236 218565 4264
rect 217495 4233 217507 4236
rect 217449 4227 217507 4233
rect 218553 4233 218565 4236
rect 218599 4233 218611 4267
rect 218553 4227 218611 4233
rect 218642 4224 218648 4276
rect 218700 4264 218706 4276
rect 220669 4267 220727 4273
rect 218700 4236 220620 4264
rect 218700 4224 218706 4236
rect 186721 4199 186779 4205
rect 186721 4196 186733 4199
rect 177352 4168 186733 4196
rect 177245 4159 177303 4165
rect 186721 4165 186733 4168
rect 186767 4165 186779 4199
rect 186721 4159 186779 4165
rect 186810 4156 186816 4208
rect 186868 4196 186874 4208
rect 190769 4199 190827 4205
rect 190769 4196 190781 4199
rect 186868 4168 190781 4196
rect 186868 4156 186874 4168
rect 190769 4165 190781 4168
rect 190815 4165 190827 4199
rect 190769 4159 190827 4165
rect 191045 4199 191103 4205
rect 191045 4165 191057 4199
rect 191091 4196 191103 4199
rect 196378 4196 196384 4208
rect 191091 4168 196384 4196
rect 191091 4165 191103 4168
rect 191045 4159 191103 4165
rect 196378 4156 196384 4168
rect 196436 4156 196442 4208
rect 196470 4156 196476 4208
rect 196528 4196 196534 4208
rect 200245 4199 200303 4205
rect 200245 4196 200257 4199
rect 196528 4168 200257 4196
rect 196528 4156 196534 4168
rect 200245 4165 200257 4168
rect 200291 4165 200303 4199
rect 200245 4159 200303 4165
rect 200705 4199 200763 4205
rect 200705 4165 200717 4199
rect 200751 4196 200763 4199
rect 206038 4196 206044 4208
rect 200751 4168 206044 4196
rect 200751 4165 200763 4168
rect 200705 4159 200763 4165
rect 206038 4156 206044 4168
rect 206096 4156 206102 4208
rect 212754 4156 212760 4208
rect 212812 4196 212818 4208
rect 220485 4199 220543 4205
rect 220485 4196 220497 4199
rect 212812 4168 220497 4196
rect 212812 4156 212818 4168
rect 220485 4165 220497 4168
rect 220531 4165 220543 4199
rect 220592 4196 220620 4236
rect 220669 4233 220681 4267
rect 220715 4264 220727 4267
rect 274210 4264 274216 4276
rect 220715 4236 274216 4264
rect 220715 4233 220727 4236
rect 220669 4227 220727 4233
rect 274210 4224 274216 4236
rect 274268 4224 274274 4276
rect 288838 4224 288844 4276
rect 288896 4224 288902 4276
rect 298222 4224 298228 4276
rect 298280 4264 298286 4276
rect 302549 4267 302607 4273
rect 302549 4264 302561 4267
rect 298280 4236 302561 4264
rect 298280 4224 298286 4236
rect 302549 4233 302561 4236
rect 302595 4233 302607 4267
rect 302549 4227 302607 4233
rect 302638 4224 302644 4276
rect 302696 4264 302702 4276
rect 324534 4264 324540 4276
rect 302696 4236 324540 4264
rect 302696 4224 302702 4236
rect 324534 4224 324540 4236
rect 324592 4224 324598 4276
rect 331529 4267 331587 4273
rect 331529 4233 331541 4267
rect 331575 4264 331587 4267
rect 336678 4264 336684 4276
rect 331575 4236 336684 4264
rect 331575 4233 331587 4236
rect 331529 4227 331587 4233
rect 336678 4224 336684 4236
rect 336736 4224 336742 4276
rect 339438 4224 339444 4276
rect 339496 4264 339502 4276
rect 346157 4267 346215 4273
rect 346157 4264 346169 4267
rect 339496 4236 346169 4264
rect 339496 4224 339502 4236
rect 346157 4233 346169 4236
rect 346203 4233 346215 4267
rect 346157 4227 346215 4233
rect 346249 4267 346307 4273
rect 346249 4233 346261 4267
rect 346295 4264 346307 4267
rect 515342 4264 515348 4276
rect 346295 4236 515348 4264
rect 346295 4233 346307 4236
rect 346249 4227 346307 4233
rect 515342 4224 515348 4236
rect 515400 4224 515406 4276
rect 529513 4267 529571 4273
rect 529513 4264 529525 4267
rect 515452 4236 529525 4264
rect 268877 4199 268935 4205
rect 268877 4196 268889 4199
rect 220592 4168 268889 4196
rect 220485 4159 220543 4165
rect 268877 4165 268889 4168
rect 268923 4165 268935 4199
rect 271358 4196 271364 4208
rect 268877 4159 268935 4165
rect 268984 4168 271364 4196
rect 58102 4088 58108 4140
rect 58160 4128 58166 4140
rect 235110 4128 235116 4140
rect 58160 4100 235116 4128
rect 58160 4088 58166 4100
rect 235110 4088 235116 4100
rect 235168 4088 235174 4140
rect 235294 4088 235300 4140
rect 235352 4128 235358 4140
rect 236398 4128 236404 4140
rect 235352 4100 236404 4128
rect 235352 4088 235358 4100
rect 236398 4088 236404 4100
rect 236456 4088 236462 4140
rect 236490 4088 236496 4140
rect 236548 4128 236554 4140
rect 237778 4128 237784 4140
rect 236548 4100 237784 4128
rect 236548 4088 236554 4100
rect 237778 4088 237784 4100
rect 237836 4088 237842 4140
rect 238054 4088 238060 4140
rect 238112 4128 238118 4140
rect 242746 4128 242752 4140
rect 238112 4100 242752 4128
rect 238112 4088 238118 4100
rect 242746 4088 242752 4100
rect 242804 4088 242810 4140
rect 244862 4088 244868 4140
rect 244920 4128 244926 4140
rect 246058 4128 246064 4140
rect 244920 4100 246064 4128
rect 244920 4088 244926 4100
rect 246058 4088 246064 4100
rect 246116 4088 246122 4140
rect 251946 4088 251952 4140
rect 252004 4128 252010 4140
rect 252958 4128 252964 4140
rect 252004 4100 252964 4128
rect 252004 4088 252010 4100
rect 252958 4088 252964 4100
rect 253016 4088 253022 4140
rect 260318 4088 260324 4140
rect 260376 4128 260382 4140
rect 261238 4128 261244 4140
rect 260376 4100 261244 4128
rect 260376 4088 260382 4100
rect 261238 4088 261244 4100
rect 261296 4088 261302 4140
rect 263909 4131 263967 4137
rect 263909 4097 263921 4131
rect 263955 4128 263967 4131
rect 264277 4131 264335 4137
rect 264277 4128 264289 4131
rect 263955 4100 264289 4128
rect 263955 4097 263967 4100
rect 263909 4091 263967 4097
rect 264277 4097 264289 4100
rect 264323 4097 264335 4131
rect 264277 4091 264335 4097
rect 267405 4131 267463 4137
rect 267405 4097 267417 4131
rect 267451 4128 267463 4131
rect 268984 4128 269012 4168
rect 271358 4156 271364 4168
rect 271416 4156 271422 4208
rect 288856 4196 288884 4224
rect 288764 4168 288884 4196
rect 267451 4100 269012 4128
rect 267451 4097 267463 4100
rect 267405 4091 267463 4097
rect 269794 4088 269800 4140
rect 269852 4128 269858 4140
rect 269852 4100 284100 4128
rect 269852 4088 269858 4100
rect 51018 4020 51024 4072
rect 51076 4060 51082 4072
rect 228118 4060 228124 4072
rect 51076 4032 228124 4060
rect 51076 4020 51082 4032
rect 228118 4020 228124 4032
rect 228176 4020 228182 4072
rect 228210 4020 228216 4072
rect 228268 4060 228274 4072
rect 229498 4060 229504 4072
rect 228268 4032 229504 4060
rect 228268 4020 228274 4032
rect 229498 4020 229504 4032
rect 229556 4020 229562 4072
rect 229685 4063 229743 4069
rect 229685 4029 229697 4063
rect 229731 4060 229743 4063
rect 230142 4060 230148 4072
rect 229731 4032 230148 4060
rect 229731 4029 229743 4032
rect 229685 4023 229743 4029
rect 230142 4020 230148 4032
rect 230200 4020 230206 4072
rect 230252 4032 235616 4060
rect 47430 3952 47436 4004
rect 47488 3992 47494 4004
rect 132993 3995 133051 4001
rect 132993 3992 133005 3995
rect 47488 3964 133005 3992
rect 47488 3952 47494 3964
rect 132993 3961 133005 3964
rect 133039 3961 133051 3995
rect 132993 3955 133051 3961
rect 133082 3952 133088 4004
rect 133140 3992 133146 4004
rect 134186 3992 134192 4004
rect 133140 3964 134192 3992
rect 133140 3952 133146 3964
rect 134186 3952 134192 3964
rect 134244 3952 134250 4004
rect 134281 3995 134339 4001
rect 134281 3961 134293 3995
rect 134327 3992 134339 3995
rect 137682 3992 137688 4004
rect 134327 3964 137688 3992
rect 134327 3961 134339 3964
rect 134281 3955 134339 3961
rect 137682 3952 137688 3964
rect 137740 3952 137746 4004
rect 137774 3952 137780 4004
rect 137832 3992 137838 4004
rect 138050 3992 138056 4004
rect 137832 3964 138056 3992
rect 137832 3952 137838 3964
rect 138050 3952 138056 3964
rect 138108 3952 138114 4004
rect 138421 3995 138479 4001
rect 138421 3961 138433 3995
rect 138467 3992 138479 3995
rect 215790 3992 215796 4004
rect 138467 3964 215796 3992
rect 138467 3961 138479 3964
rect 138421 3955 138479 3961
rect 215790 3952 215796 3964
rect 215848 3952 215854 4004
rect 215882 3952 215888 4004
rect 215940 3992 215946 4004
rect 217449 3995 217507 4001
rect 217449 3992 217461 3995
rect 215940 3964 217461 3992
rect 215940 3952 215946 3964
rect 217449 3961 217461 3964
rect 217495 3961 217507 3995
rect 217449 3955 217507 3961
rect 217538 3952 217544 4004
rect 217596 3992 217602 4004
rect 218458 3992 218464 4004
rect 217596 3964 218464 3992
rect 217596 3952 217602 3964
rect 218458 3952 218464 3964
rect 218516 3952 218522 4004
rect 218553 3995 218611 4001
rect 218553 3961 218565 3995
rect 218599 3992 218611 3995
rect 219657 3995 219715 4001
rect 219657 3992 219669 3995
rect 218599 3964 219669 3992
rect 218599 3961 218611 3964
rect 218553 3955 218611 3961
rect 219657 3961 219669 3964
rect 219703 3961 219715 3995
rect 219657 3955 219715 3961
rect 219746 3952 219752 4004
rect 219804 3992 219810 4004
rect 219841 3995 219899 4001
rect 219841 3992 219853 3995
rect 219804 3964 219853 3992
rect 219804 3952 219810 3964
rect 219841 3961 219853 3964
rect 219887 3961 219899 3995
rect 219841 3955 219899 3961
rect 219933 3995 219991 4001
rect 219933 3961 219945 3995
rect 219979 3992 219991 3995
rect 230252 3992 230280 4032
rect 219979 3964 230280 3992
rect 230329 3995 230387 4001
rect 219979 3961 219991 3964
rect 219933 3955 219991 3961
rect 230329 3961 230341 3995
rect 230375 3992 230387 3995
rect 232905 3995 232963 4001
rect 232905 3992 232917 3995
rect 230375 3964 232917 3992
rect 230375 3961 230387 3964
rect 230329 3955 230387 3961
rect 232905 3961 232917 3964
rect 232951 3961 232963 3995
rect 235588 3992 235616 4032
rect 235662 4020 235668 4072
rect 235720 4060 235726 4072
rect 237962 4060 237968 4072
rect 235720 4032 237968 4060
rect 235720 4020 235726 4032
rect 237962 4020 237968 4032
rect 238020 4020 238026 4072
rect 241274 4020 241280 4072
rect 241332 4060 241338 4072
rect 254341 4063 254399 4069
rect 254341 4060 254353 4063
rect 241332 4032 254353 4060
rect 241332 4020 241338 4032
rect 254341 4029 254353 4032
rect 254387 4029 254399 4063
rect 254341 4023 254399 4029
rect 268598 4020 268604 4072
rect 268656 4060 268662 4072
rect 283965 4063 284023 4069
rect 283965 4060 283977 4063
rect 268656 4032 283977 4060
rect 268656 4020 268662 4032
rect 283965 4029 283977 4032
rect 284011 4029 284023 4063
rect 284072 4060 284100 4100
rect 284146 4088 284152 4140
rect 284204 4128 284210 4140
rect 285434 4128 285440 4140
rect 284204 4100 285440 4128
rect 284204 4088 284210 4100
rect 285434 4088 285440 4100
rect 285492 4088 285498 4140
rect 287642 4088 287648 4140
rect 287700 4128 287706 4140
rect 288764 4128 288792 4168
rect 298314 4156 298320 4208
rect 298372 4196 298378 4208
rect 302454 4196 302460 4208
rect 298372 4168 302460 4196
rect 298372 4156 298378 4168
rect 302454 4156 302460 4168
rect 302512 4156 302518 4208
rect 323338 4196 323344 4208
rect 302564 4168 323344 4196
rect 287700 4100 288792 4128
rect 287700 4088 287706 4100
rect 288838 4088 288844 4140
rect 288896 4128 288902 4140
rect 289390 4128 289396 4140
rect 288896 4100 289396 4128
rect 288896 4088 288902 4100
rect 289390 4088 289396 4100
rect 289448 4088 289454 4140
rect 289574 4088 289580 4140
rect 289632 4128 289638 4140
rect 290034 4128 290040 4140
rect 289632 4100 290040 4128
rect 289632 4088 289638 4100
rect 290034 4088 290040 4100
rect 290092 4088 290098 4140
rect 291506 4088 291512 4140
rect 291564 4128 291570 4140
rect 292426 4128 292432 4140
rect 291564 4100 292432 4128
rect 291564 4088 291570 4100
rect 292426 4088 292432 4100
rect 292484 4088 292490 4140
rect 293898 4088 293904 4140
rect 293956 4128 293962 4140
rect 297210 4128 297216 4140
rect 293956 4100 297216 4128
rect 293956 4088 293962 4100
rect 297210 4088 297216 4100
rect 297268 4088 297274 4140
rect 301077 4131 301135 4137
rect 301077 4097 301089 4131
rect 301123 4128 301135 4131
rect 302564 4128 302592 4168
rect 323338 4156 323344 4168
rect 323396 4156 323402 4208
rect 324169 4199 324227 4205
rect 324169 4165 324181 4199
rect 324215 4196 324227 4199
rect 331621 4199 331679 4205
rect 331621 4196 331633 4199
rect 324215 4168 331633 4196
rect 324215 4165 324227 4168
rect 324169 4159 324227 4165
rect 331621 4165 331633 4168
rect 331667 4165 331679 4199
rect 331621 4159 331679 4165
rect 338426 4156 338432 4208
rect 338484 4196 338490 4208
rect 515253 4199 515311 4205
rect 515253 4196 515265 4199
rect 338484 4168 515265 4196
rect 338484 4156 338490 4168
rect 515253 4165 515265 4168
rect 515299 4165 515311 4199
rect 515452 4196 515480 4236
rect 529513 4233 529525 4236
rect 529559 4233 529571 4267
rect 529513 4227 529571 4233
rect 529605 4267 529663 4273
rect 529605 4233 529617 4267
rect 529651 4264 529663 4267
rect 537422 4264 537428 4276
rect 529651 4236 537428 4264
rect 529651 4233 529663 4236
rect 529605 4227 529663 4233
rect 537422 4224 537428 4236
rect 537480 4224 537486 4276
rect 523162 4196 523168 4208
rect 515253 4159 515311 4165
rect 515360 4168 515480 4196
rect 516188 4168 523168 4196
rect 301123 4100 302592 4128
rect 302641 4131 302699 4137
rect 301123 4097 301135 4100
rect 301077 4091 301135 4097
rect 302641 4097 302653 4131
rect 302687 4128 302699 4131
rect 305490 4128 305496 4140
rect 302687 4100 305496 4128
rect 302687 4097 302699 4100
rect 302641 4091 302699 4097
rect 305490 4088 305496 4100
rect 305548 4088 305554 4140
rect 312393 4131 312451 4137
rect 312393 4097 312405 4131
rect 312439 4128 312451 4131
rect 319750 4128 319756 4140
rect 312439 4100 319756 4128
rect 312439 4097 312451 4100
rect 312393 4091 312451 4097
rect 319750 4088 319756 4100
rect 319808 4088 319814 4140
rect 320578 4088 320584 4140
rect 320636 4128 320642 4140
rect 322881 4131 322939 4137
rect 320636 4100 322832 4128
rect 320636 4088 320642 4100
rect 284974 4060 284980 4072
rect 284072 4032 284980 4060
rect 283965 4023 284023 4029
rect 284974 4020 284980 4032
rect 285032 4020 285038 4072
rect 294266 4020 294272 4072
rect 294324 4060 294330 4072
rect 299697 4063 299755 4069
rect 299697 4060 299709 4063
rect 294324 4032 299709 4060
rect 294324 4020 294330 4032
rect 299697 4029 299709 4032
rect 299743 4029 299755 4063
rect 299697 4023 299755 4029
rect 301169 4063 301227 4069
rect 301169 4029 301181 4063
rect 301215 4060 301227 4063
rect 302546 4060 302552 4072
rect 301215 4032 302552 4060
rect 301215 4029 301227 4032
rect 301169 4023 301227 4029
rect 302546 4020 302552 4032
rect 302604 4020 302610 4072
rect 302730 4020 302736 4072
rect 302788 4060 302794 4072
rect 312485 4063 312543 4069
rect 312485 4060 312497 4063
rect 302788 4032 312497 4060
rect 302788 4020 302794 4032
rect 312485 4029 312497 4032
rect 312531 4029 312543 4063
rect 312485 4023 312543 4029
rect 312577 4063 312635 4069
rect 312577 4029 312589 4063
rect 312623 4060 312635 4063
rect 320946 4060 320952 4072
rect 312623 4032 320952 4060
rect 312623 4029 312635 4032
rect 312577 4023 312635 4029
rect 320946 4020 320952 4032
rect 321004 4020 321010 4072
rect 322804 4060 322832 4100
rect 322881 4097 322893 4131
rect 322927 4128 322939 4131
rect 418745 4131 418803 4137
rect 418745 4128 418757 4131
rect 322927 4100 418757 4128
rect 322927 4097 322939 4100
rect 322881 4091 322939 4097
rect 418745 4097 418757 4100
rect 418791 4097 418803 4131
rect 418745 4091 418803 4097
rect 418834 4088 418840 4140
rect 418892 4128 418898 4140
rect 505685 4131 505743 4137
rect 505685 4128 505697 4131
rect 418892 4100 505697 4128
rect 418892 4088 418898 4100
rect 505685 4097 505697 4100
rect 505731 4097 505743 4131
rect 505685 4091 505743 4097
rect 515069 4131 515127 4137
rect 515069 4097 515081 4131
rect 515115 4128 515127 4131
rect 515360 4128 515388 4168
rect 515115 4100 515388 4128
rect 515437 4131 515495 4137
rect 515115 4097 515127 4100
rect 515069 4091 515127 4097
rect 515437 4097 515449 4131
rect 515483 4128 515495 4131
rect 516188 4128 516216 4168
rect 523162 4156 523168 4168
rect 523220 4156 523226 4208
rect 515483 4100 516216 4128
rect 515483 4097 515495 4100
rect 515437 4091 515495 4097
rect 577994 4088 578000 4140
rect 578052 4128 578058 4140
rect 579098 4128 579104 4140
rect 578052 4100 579104 4128
rect 578052 4088 578058 4100
rect 579098 4088 579104 4100
rect 579156 4088 579162 4140
rect 579374 4088 579380 4140
rect 579432 4128 579438 4140
rect 580294 4128 580300 4140
rect 579432 4100 580300 4128
rect 579432 4088 579438 4100
rect 580294 4088 580300 4100
rect 580352 4088 580358 4140
rect 436314 4060 436320 4072
rect 322804 4032 436320 4060
rect 436314 4020 436320 4032
rect 436372 4020 436378 4072
rect 505593 4063 505651 4069
rect 505593 4029 505605 4063
rect 505639 4060 505651 4063
rect 512490 4060 512496 4072
rect 505639 4032 512496 4060
rect 505639 4029 505651 4032
rect 505593 4023 505651 4029
rect 512490 4020 512496 4032
rect 512548 4020 512554 4072
rect 239342 3992 239348 4004
rect 235588 3964 239348 3992
rect 232905 3955 232963 3961
rect 239342 3952 239348 3964
rect 239400 3952 239406 4004
rect 267494 3952 267500 4004
rect 267552 3992 267558 4004
rect 284882 3992 284888 4004
rect 267552 3964 284888 3992
rect 267552 3952 267558 3964
rect 284882 3952 284888 3964
rect 284940 3952 284946 4004
rect 286446 3952 286452 4004
rect 286504 3992 286510 4004
rect 289114 3992 289120 4004
rect 286504 3964 289120 3992
rect 286504 3952 286510 3964
rect 289114 3952 289120 3964
rect 289172 3952 289178 4004
rect 295094 3952 295100 4004
rect 295152 3992 295158 4004
rect 302457 3995 302515 4001
rect 302457 3992 302469 3995
rect 295152 3964 302469 3992
rect 295152 3952 295158 3964
rect 302457 3961 302469 3964
rect 302503 3961 302515 3995
rect 304294 3992 304300 4004
rect 302457 3955 302515 3961
rect 302564 3964 304300 3992
rect 46234 3884 46240 3936
rect 46292 3924 46298 3936
rect 234929 3927 234987 3933
rect 234929 3924 234941 3927
rect 46292 3896 234941 3924
rect 46292 3884 46298 3896
rect 234929 3893 234941 3896
rect 234975 3893 234987 3927
rect 234929 3887 234987 3893
rect 266298 3884 266304 3936
rect 266356 3924 266362 3936
rect 284054 3924 284060 3936
rect 266356 3896 284060 3924
rect 266356 3884 266362 3896
rect 284054 3884 284060 3896
rect 284112 3884 284118 3936
rect 284149 3927 284207 3933
rect 284149 3893 284161 3927
rect 284195 3924 284207 3927
rect 285250 3924 285256 3936
rect 284195 3896 285256 3924
rect 284195 3893 284207 3896
rect 284149 3887 284207 3893
rect 285250 3884 285256 3896
rect 285308 3884 285314 3936
rect 292794 3884 292800 3936
rect 292852 3924 292858 3936
rect 298406 3924 298412 3936
rect 292852 3896 298412 3924
rect 292852 3884 292858 3896
rect 298406 3884 298412 3896
rect 298464 3884 298470 3936
rect 298501 3927 298559 3933
rect 298501 3893 298513 3927
rect 298547 3924 298559 3927
rect 302564 3924 302592 3964
rect 304294 3952 304300 3964
rect 304352 3952 304358 4004
rect 321866 3952 321872 4004
rect 321924 3992 321930 4004
rect 439902 3992 439908 4004
rect 321924 3964 439908 3992
rect 321924 3952 321930 3964
rect 439902 3952 439908 3964
rect 439960 3952 439966 4004
rect 505777 3995 505835 4001
rect 505777 3961 505789 3995
rect 505823 3992 505835 3995
rect 516078 3992 516084 4004
rect 505823 3964 516084 3992
rect 505823 3961 505835 3964
rect 505777 3955 505835 3961
rect 516078 3952 516084 3964
rect 516136 3952 516142 4004
rect 298547 3896 302592 3924
rect 298547 3893 298559 3896
rect 298501 3887 298559 3893
rect 320486 3884 320492 3936
rect 320544 3924 320550 3936
rect 322881 3927 322939 3933
rect 322881 3924 322893 3927
rect 320544 3896 322893 3924
rect 320544 3884 320550 3896
rect 322881 3893 322893 3896
rect 322927 3893 322939 3927
rect 322881 3887 322939 3893
rect 322970 3884 322976 3936
rect 323028 3924 323034 3936
rect 324169 3927 324227 3933
rect 324169 3924 324181 3927
rect 323028 3896 324181 3924
rect 323028 3884 323034 3896
rect 324169 3893 324181 3896
rect 324215 3893 324227 3927
rect 324169 3887 324227 3893
rect 324258 3884 324264 3936
rect 324316 3924 324322 3936
rect 325917 3927 325975 3933
rect 325917 3924 325929 3927
rect 324316 3896 325929 3924
rect 324316 3884 324322 3896
rect 325917 3893 325929 3896
rect 325963 3893 325975 3927
rect 325917 3887 325975 3893
rect 326009 3927 326067 3933
rect 326009 3893 326021 3927
rect 326055 3924 326067 3927
rect 443490 3924 443496 3936
rect 326055 3896 443496 3924
rect 326055 3893 326067 3896
rect 326009 3887 326067 3893
rect 443490 3884 443496 3896
rect 443548 3884 443554 3936
rect 1600 3760 583316 3856
rect 42646 3680 42652 3732
rect 42704 3720 42710 3732
rect 230329 3723 230387 3729
rect 230329 3720 230341 3723
rect 42704 3692 230341 3720
rect 42704 3680 42710 3692
rect 230329 3689 230341 3692
rect 230375 3689 230387 3723
rect 230329 3683 230387 3689
rect 230418 3680 230424 3732
rect 230476 3720 230482 3732
rect 235202 3720 235208 3732
rect 230476 3692 235208 3720
rect 230476 3680 230482 3692
rect 235202 3680 235208 3692
rect 235260 3680 235266 3732
rect 235297 3723 235355 3729
rect 235297 3689 235309 3723
rect 235343 3720 235355 3723
rect 239710 3720 239716 3732
rect 235343 3692 239716 3720
rect 235343 3689 235355 3692
rect 235297 3683 235355 3689
rect 239710 3680 239716 3692
rect 239768 3680 239774 3732
rect 249557 3723 249615 3729
rect 249557 3689 249569 3723
rect 249603 3720 249615 3723
rect 254798 3720 254804 3732
rect 249603 3692 254804 3720
rect 249603 3689 249615 3692
rect 249557 3683 249615 3689
rect 254798 3680 254804 3692
rect 254856 3680 254862 3732
rect 263906 3680 263912 3732
rect 263964 3720 263970 3732
rect 283686 3720 283692 3732
rect 263964 3692 283692 3720
rect 263964 3680 263970 3692
rect 283686 3680 283692 3692
rect 283744 3680 283750 3732
rect 292886 3680 292892 3732
rect 292944 3720 292950 3732
rect 299602 3720 299608 3732
rect 292944 3692 299608 3720
rect 292944 3680 292950 3692
rect 299602 3680 299608 3692
rect 299660 3680 299666 3732
rect 299697 3723 299755 3729
rect 299697 3689 299709 3723
rect 299743 3720 299755 3723
rect 311470 3720 311476 3732
rect 299743 3692 311476 3720
rect 299743 3689 299755 3692
rect 299697 3683 299755 3689
rect 311470 3680 311476 3692
rect 311528 3680 311534 3732
rect 324626 3680 324632 3732
rect 324684 3720 324690 3732
rect 331529 3723 331587 3729
rect 331529 3720 331541 3723
rect 324684 3692 331541 3720
rect 324684 3680 324690 3692
rect 331529 3689 331541 3692
rect 331575 3689 331587 3723
rect 331529 3683 331587 3689
rect 331621 3723 331679 3729
rect 331621 3689 331633 3723
rect 331667 3720 331679 3723
rect 447078 3720 447084 3732
rect 331667 3692 447084 3720
rect 331667 3689 331679 3692
rect 331621 3683 331679 3689
rect 447078 3680 447084 3692
rect 447136 3680 447142 3732
rect 38966 3612 38972 3664
rect 39024 3652 39030 3664
rect 44765 3655 44823 3661
rect 39024 3624 44716 3652
rect 39024 3612 39030 3624
rect 29582 3544 29588 3596
rect 29640 3584 29646 3596
rect 30778 3584 30784 3596
rect 29640 3556 30784 3584
rect 29640 3544 29646 3556
rect 30778 3544 30784 3556
rect 30836 3544 30842 3596
rect 36666 3544 36672 3596
rect 36724 3584 36730 3596
rect 37678 3584 37684 3596
rect 36724 3556 37684 3584
rect 36724 3544 36730 3556
rect 37678 3544 37684 3556
rect 37736 3544 37742 3596
rect 37862 3544 37868 3596
rect 37920 3584 37926 3596
rect 39058 3584 39064 3596
rect 37920 3556 39064 3584
rect 37920 3544 37926 3556
rect 39058 3544 39064 3556
rect 39116 3544 39122 3596
rect 43842 3544 43848 3596
rect 43900 3584 43906 3596
rect 44578 3584 44584 3596
rect 43900 3556 44584 3584
rect 43900 3544 43906 3556
rect 44578 3544 44584 3556
rect 44636 3544 44642 3596
rect 44688 3584 44716 3624
rect 44765 3621 44777 3655
rect 44811 3652 44823 3655
rect 138881 3655 138939 3661
rect 138881 3652 138893 3655
rect 44811 3624 138893 3652
rect 44811 3621 44823 3624
rect 44765 3615 44823 3621
rect 138881 3621 138893 3624
rect 138927 3621 138939 3655
rect 138881 3615 138939 3621
rect 138970 3612 138976 3664
rect 139028 3652 139034 3664
rect 139798 3652 139804 3664
rect 139028 3624 139804 3652
rect 139028 3612 139034 3624
rect 139798 3612 139804 3624
rect 139856 3612 139862 3664
rect 141362 3612 141368 3664
rect 141420 3652 141426 3664
rect 142558 3652 142564 3664
rect 141420 3624 142564 3652
rect 141420 3612 141426 3624
rect 142558 3612 142564 3624
rect 142616 3612 142622 3664
rect 142745 3655 142803 3661
rect 142745 3621 142757 3655
rect 142791 3652 142803 3655
rect 148449 3655 148507 3661
rect 148449 3652 148461 3655
rect 142791 3624 148461 3652
rect 142791 3621 142803 3624
rect 142745 3615 142803 3621
rect 148449 3621 148461 3624
rect 148495 3621 148507 3655
rect 148449 3615 148507 3621
rect 148538 3612 148544 3664
rect 148596 3652 148602 3664
rect 149458 3652 149464 3664
rect 148596 3624 149464 3652
rect 148596 3612 148602 3624
rect 149458 3612 149464 3624
rect 149516 3612 149522 3664
rect 149553 3655 149611 3661
rect 149553 3621 149565 3655
rect 149599 3652 149611 3655
rect 152129 3655 152187 3661
rect 152129 3652 152141 3655
rect 149599 3624 152141 3652
rect 149599 3621 149611 3624
rect 149553 3615 149611 3621
rect 152129 3621 152141 3624
rect 152175 3621 152187 3655
rect 152129 3615 152187 3621
rect 152221 3655 152279 3661
rect 152221 3621 152233 3655
rect 152267 3652 152279 3655
rect 159121 3655 159179 3661
rect 159121 3652 159133 3655
rect 152267 3624 159133 3652
rect 152267 3621 152279 3624
rect 152221 3615 152279 3621
rect 159121 3621 159133 3624
rect 159167 3621 159179 3655
rect 159121 3615 159179 3621
rect 159210 3612 159216 3664
rect 159268 3652 159274 3664
rect 160498 3652 160504 3664
rect 159268 3624 160504 3652
rect 159268 3612 159274 3624
rect 160498 3612 160504 3624
rect 160556 3612 160562 3664
rect 162065 3655 162123 3661
rect 162065 3621 162077 3655
rect 162111 3652 162123 3655
rect 162709 3655 162767 3661
rect 162709 3652 162721 3655
rect 162111 3624 162721 3652
rect 162111 3621 162123 3624
rect 162065 3615 162123 3621
rect 162709 3621 162721 3624
rect 162755 3621 162767 3655
rect 162709 3615 162767 3621
rect 162798 3612 162804 3664
rect 162856 3652 162862 3664
rect 163258 3652 163264 3664
rect 162856 3624 163264 3652
rect 162856 3612 162862 3624
rect 163258 3612 163264 3624
rect 163316 3612 163322 3664
rect 163353 3655 163411 3661
rect 163353 3621 163365 3655
rect 163399 3652 163411 3655
rect 166297 3655 166355 3661
rect 166297 3652 166309 3655
rect 163399 3624 166309 3652
rect 163399 3621 163411 3624
rect 163353 3615 163411 3621
rect 166297 3621 166309 3624
rect 166343 3621 166355 3655
rect 166297 3615 166355 3621
rect 166386 3612 166392 3664
rect 166444 3652 166450 3664
rect 167214 3652 167220 3664
rect 166444 3624 167220 3652
rect 166444 3612 166450 3624
rect 167214 3612 167220 3624
rect 167272 3612 167278 3664
rect 167401 3655 167459 3661
rect 167401 3621 167413 3655
rect 167447 3652 167459 3655
rect 167493 3655 167551 3661
rect 167493 3652 167505 3655
rect 167447 3624 167505 3652
rect 167447 3621 167459 3624
rect 167401 3615 167459 3621
rect 167493 3621 167505 3624
rect 167539 3621 167551 3655
rect 167493 3615 167551 3621
rect 167585 3655 167643 3661
rect 167585 3621 167597 3655
rect 167631 3652 167643 3655
rect 176969 3655 177027 3661
rect 176969 3652 176981 3655
rect 167631 3624 176981 3652
rect 167631 3621 167643 3624
rect 167585 3615 167643 3621
rect 176969 3621 176981 3624
rect 177015 3621 177027 3655
rect 176969 3615 177027 3621
rect 177061 3655 177119 3661
rect 177061 3621 177073 3655
rect 177107 3652 177119 3655
rect 181109 3655 181167 3661
rect 181109 3652 181121 3655
rect 177107 3624 181121 3652
rect 177107 3621 177119 3624
rect 177061 3615 177119 3621
rect 181109 3621 181121 3624
rect 181155 3621 181167 3655
rect 210270 3652 210276 3664
rect 181109 3615 181167 3621
rect 181308 3624 210276 3652
rect 181201 3587 181259 3593
rect 181201 3584 181213 3587
rect 44688 3556 181213 3584
rect 181201 3553 181213 3556
rect 181247 3553 181259 3587
rect 181201 3547 181259 3553
rect 10538 3476 10544 3528
rect 10596 3516 10602 3528
rect 11458 3516 11464 3528
rect 10596 3488 11464 3516
rect 10596 3476 10602 3488
rect 11458 3476 11464 3488
rect 11516 3476 11522 3528
rect 11734 3476 11740 3528
rect 11792 3516 11798 3528
rect 12838 3516 12844 3528
rect 11792 3488 12844 3516
rect 11792 3476 11798 3488
rect 12838 3476 12844 3488
rect 12896 3476 12902 3528
rect 18818 3476 18824 3528
rect 18876 3516 18882 3528
rect 19738 3516 19744 3528
rect 18876 3488 19744 3516
rect 18876 3476 18882 3488
rect 19738 3476 19744 3488
rect 19796 3476 19802 3528
rect 20014 3476 20020 3528
rect 20072 3516 20078 3528
rect 21118 3516 21124 3528
rect 20072 3488 21124 3516
rect 20072 3476 20078 3488
rect 21118 3476 21124 3488
rect 21176 3476 21182 3528
rect 34366 3476 34372 3528
rect 34424 3516 34430 3528
rect 34918 3516 34924 3528
rect 34424 3488 34924 3516
rect 34424 3476 34430 3488
rect 34918 3476 34924 3488
rect 34976 3476 34982 3528
rect 35470 3476 35476 3528
rect 35528 3516 35534 3528
rect 36393 3519 36451 3525
rect 36393 3516 36405 3519
rect 35528 3488 36405 3516
rect 35528 3476 35534 3488
rect 36393 3485 36405 3488
rect 36439 3485 36451 3519
rect 36393 3479 36451 3485
rect 45961 3519 46019 3525
rect 45961 3485 45973 3519
rect 46007 3516 46019 3519
rect 56265 3519 56323 3525
rect 56265 3516 56277 3519
rect 46007 3488 56277 3516
rect 46007 3485 46019 3488
rect 45961 3479 46019 3485
rect 56265 3485 56277 3488
rect 56311 3485 56323 3519
rect 56265 3479 56323 3485
rect 65189 3519 65247 3525
rect 65189 3485 65201 3519
rect 65235 3485 65247 3519
rect 65189 3479 65247 3485
rect 65281 3519 65339 3525
rect 65281 3485 65293 3519
rect 65327 3516 65339 3519
rect 75033 3519 75091 3525
rect 75033 3516 75045 3519
rect 65327 3488 75045 3516
rect 65327 3485 65339 3488
rect 65281 3479 65339 3485
rect 75033 3485 75045 3488
rect 75079 3485 75091 3519
rect 75033 3479 75091 3485
rect 45869 3451 45927 3457
rect 45869 3417 45881 3451
rect 45915 3448 45927 3451
rect 56357 3451 56415 3457
rect 56357 3448 56369 3451
rect 45915 3420 56369 3448
rect 45915 3417 45927 3420
rect 45869 3411 45927 3417
rect 56357 3417 56369 3420
rect 56403 3417 56415 3451
rect 65204 3448 65232 3479
rect 81930 3476 81936 3528
rect 81988 3516 81994 3528
rect 83034 3516 83040 3528
rect 81988 3488 83040 3516
rect 81988 3476 81994 3488
rect 83034 3476 83040 3488
rect 83092 3476 83098 3528
rect 84601 3519 84659 3525
rect 84601 3485 84613 3519
rect 84647 3516 84659 3519
rect 93709 3519 93767 3525
rect 93709 3516 93721 3519
rect 84647 3488 93721 3516
rect 84647 3485 84659 3488
rect 84601 3479 84659 3485
rect 93709 3485 93721 3488
rect 93755 3485 93767 3519
rect 93709 3479 93767 3485
rect 93798 3476 93804 3528
rect 93856 3516 93862 3528
rect 94258 3516 94264 3528
rect 93856 3488 94264 3516
rect 93856 3476 93862 3488
rect 94258 3476 94264 3488
rect 94316 3476 94322 3528
rect 94994 3476 95000 3528
rect 95052 3516 95058 3528
rect 95638 3516 95644 3528
rect 95052 3488 95644 3516
rect 95052 3476 95058 3488
rect 95638 3476 95644 3488
rect 95696 3476 95702 3528
rect 96190 3476 96196 3528
rect 96248 3516 96254 3528
rect 97018 3516 97024 3528
rect 96248 3488 97024 3516
rect 96248 3476 96254 3488
rect 97018 3476 97024 3488
rect 97076 3476 97082 3528
rect 98582 3476 98588 3528
rect 98640 3516 98646 3528
rect 99778 3516 99784 3528
rect 98640 3488 99784 3516
rect 98640 3476 98646 3488
rect 99778 3476 99784 3488
rect 99836 3476 99842 3528
rect 103921 3519 103979 3525
rect 103921 3485 103933 3519
rect 103967 3516 103979 3519
rect 103967 3488 113992 3516
rect 103967 3485 103979 3488
rect 103921 3479 103979 3485
rect 75125 3451 75183 3457
rect 75125 3448 75137 3451
rect 65204 3420 75137 3448
rect 56357 3411 56415 3417
rect 75125 3417 75137 3420
rect 75171 3417 75183 3451
rect 75125 3411 75183 3417
rect 84509 3451 84567 3457
rect 84509 3417 84521 3451
rect 84555 3448 84567 3451
rect 99686 3448 99692 3460
rect 84555 3420 99692 3448
rect 84555 3417 84567 3420
rect 84509 3411 84567 3417
rect 99686 3408 99692 3420
rect 99744 3408 99750 3460
rect 103826 3408 103832 3460
rect 103884 3448 103890 3460
rect 113854 3448 113860 3460
rect 103884 3420 113860 3448
rect 103884 3408 103890 3420
rect 113854 3408 113860 3420
rect 113912 3408 113918 3460
rect 113964 3448 113992 3488
rect 114038 3476 114044 3528
rect 114096 3516 114102 3528
rect 114958 3516 114964 3528
rect 114096 3488 114964 3516
rect 114096 3476 114102 3488
rect 114958 3476 114964 3488
rect 115016 3476 115022 3528
rect 115234 3476 115240 3528
rect 115292 3516 115298 3528
rect 116338 3516 116344 3528
rect 115292 3488 116344 3516
rect 115292 3476 115298 3488
rect 116338 3476 116344 3488
rect 116396 3476 116402 3528
rect 116430 3476 116436 3528
rect 116488 3516 116494 3528
rect 117442 3516 117448 3528
rect 116488 3488 117448 3516
rect 116488 3476 116494 3488
rect 117442 3476 117448 3488
rect 117500 3476 117506 3528
rect 119926 3476 119932 3528
rect 119984 3516 119990 3528
rect 120478 3516 120484 3528
rect 119984 3488 120484 3516
rect 119984 3476 119990 3488
rect 120478 3476 120484 3488
rect 120536 3476 120542 3528
rect 121122 3476 121128 3528
rect 121180 3516 121186 3528
rect 121858 3516 121864 3528
rect 121180 3488 121864 3516
rect 121180 3476 121186 3488
rect 121858 3476 121864 3488
rect 121916 3476 121922 3528
rect 123514 3476 123520 3528
rect 123572 3516 123578 3528
rect 124618 3516 124624 3528
rect 123572 3488 124624 3516
rect 123572 3476 123578 3488
rect 124618 3476 124624 3488
rect 124676 3476 124682 3528
rect 124710 3476 124716 3528
rect 124768 3516 124774 3528
rect 125814 3516 125820 3528
rect 124768 3488 125820 3516
rect 124768 3476 124774 3488
rect 125814 3476 125820 3488
rect 125872 3476 125878 3528
rect 126090 3476 126096 3528
rect 126148 3516 126154 3528
rect 128209 3519 128267 3525
rect 128209 3516 128221 3519
rect 126148 3488 128221 3516
rect 126148 3476 126154 3488
rect 128209 3485 128221 3488
rect 128255 3485 128267 3519
rect 128209 3479 128267 3485
rect 128298 3476 128304 3528
rect 128356 3516 128362 3528
rect 128758 3516 128764 3528
rect 128356 3488 128764 3516
rect 128356 3476 128362 3488
rect 128758 3476 128764 3488
rect 128816 3476 128822 3528
rect 128945 3519 129003 3525
rect 128945 3485 128957 3519
rect 128991 3516 129003 3519
rect 138329 3519 138387 3525
rect 138329 3516 138341 3519
rect 128991 3488 138341 3516
rect 128991 3485 129003 3488
rect 128945 3479 129003 3485
rect 138329 3485 138341 3488
rect 138375 3485 138387 3519
rect 138329 3479 138387 3485
rect 138418 3476 138424 3528
rect 138476 3516 138482 3528
rect 138789 3519 138847 3525
rect 138789 3516 138801 3519
rect 138476 3488 138801 3516
rect 138476 3476 138482 3488
rect 138789 3485 138801 3488
rect 138835 3485 138847 3519
rect 138789 3479 138847 3485
rect 138881 3519 138939 3525
rect 138881 3485 138893 3519
rect 138927 3516 138939 3519
rect 147989 3519 148047 3525
rect 147989 3516 148001 3519
rect 138927 3488 148001 3516
rect 138927 3485 138939 3488
rect 138881 3479 138939 3485
rect 147989 3485 148001 3488
rect 148035 3485 148047 3519
rect 147989 3479 148047 3485
rect 148081 3519 148139 3525
rect 148081 3485 148093 3519
rect 148127 3516 148139 3519
rect 157646 3516 157652 3528
rect 148127 3488 157652 3516
rect 148127 3485 148139 3488
rect 148081 3479 148139 3485
rect 157646 3476 157652 3488
rect 157704 3476 157710 3528
rect 157741 3519 157799 3525
rect 157741 3485 157753 3519
rect 157787 3516 157799 3519
rect 157833 3519 157891 3525
rect 157833 3516 157845 3519
rect 157787 3488 157845 3516
rect 157787 3485 157799 3488
rect 157741 3479 157799 3485
rect 157833 3485 157845 3488
rect 157879 3485 157891 3519
rect 161605 3519 161663 3525
rect 161605 3516 161617 3519
rect 157833 3479 157891 3485
rect 157940 3488 161617 3516
rect 128850 3448 128856 3460
rect 113964 3420 128856 3448
rect 128850 3408 128856 3420
rect 128908 3408 128914 3460
rect 129037 3451 129095 3457
rect 129037 3417 129049 3451
rect 129083 3448 129095 3451
rect 132809 3451 132867 3457
rect 132809 3448 132821 3451
rect 129083 3420 132821 3448
rect 129083 3417 129095 3420
rect 129037 3411 129095 3417
rect 132809 3417 132821 3420
rect 132855 3417 132867 3451
rect 132809 3411 132867 3417
rect 133361 3451 133419 3457
rect 133361 3417 133373 3451
rect 133407 3448 133419 3451
rect 142377 3451 142435 3457
rect 142377 3448 142389 3451
rect 133407 3420 142389 3448
rect 133407 3417 133419 3420
rect 133361 3411 133419 3417
rect 142377 3417 142389 3420
rect 142423 3417 142435 3451
rect 142377 3411 142435 3417
rect 142561 3451 142619 3457
rect 142561 3417 142573 3451
rect 142607 3448 142619 3451
rect 152313 3451 152371 3457
rect 152313 3448 152325 3451
rect 142607 3420 152325 3448
rect 142607 3417 142619 3420
rect 142561 3411 142619 3417
rect 152313 3417 152325 3420
rect 152359 3417 152371 3451
rect 152313 3411 152371 3417
rect 152497 3451 152555 3457
rect 152497 3417 152509 3451
rect 152543 3448 152555 3451
rect 157940 3448 157968 3488
rect 161605 3485 161617 3488
rect 161651 3485 161663 3519
rect 161605 3479 161663 3485
rect 161881 3519 161939 3525
rect 161881 3485 161893 3519
rect 161927 3516 161939 3519
rect 177153 3519 177211 3525
rect 177153 3516 177165 3519
rect 161927 3488 177165 3516
rect 161927 3485 161939 3488
rect 161881 3479 161939 3485
rect 177153 3485 177165 3488
rect 177199 3485 177211 3519
rect 177153 3479 177211 3485
rect 177245 3519 177303 3525
rect 177245 3485 177257 3519
rect 177291 3516 177303 3519
rect 181308 3516 181336 3624
rect 210270 3612 210276 3624
rect 210328 3612 210334 3664
rect 210365 3655 210423 3661
rect 210365 3621 210377 3655
rect 210411 3652 210423 3655
rect 215790 3652 215796 3664
rect 210411 3624 215796 3652
rect 210411 3621 210423 3624
rect 210365 3615 210423 3621
rect 215790 3612 215796 3624
rect 215848 3612 215854 3664
rect 215885 3655 215943 3661
rect 215885 3621 215897 3655
rect 215931 3652 215943 3655
rect 219933 3655 219991 3661
rect 219933 3652 219945 3655
rect 215931 3624 219945 3652
rect 215931 3621 215943 3624
rect 215885 3615 215943 3621
rect 219933 3621 219945 3624
rect 219979 3621 219991 3655
rect 219933 3615 219991 3621
rect 220022 3612 220028 3664
rect 220080 3652 220086 3664
rect 224530 3652 224536 3664
rect 220080 3624 224536 3652
rect 220080 3612 220086 3624
rect 224530 3612 224536 3624
rect 224588 3612 224594 3664
rect 225174 3612 225180 3664
rect 225232 3652 225238 3664
rect 225450 3652 225456 3664
rect 225232 3624 225456 3652
rect 225232 3612 225238 3624
rect 225450 3612 225456 3624
rect 225508 3612 225514 3664
rect 234834 3652 234840 3664
rect 225560 3624 234840 3652
rect 181477 3587 181535 3593
rect 181477 3553 181489 3587
rect 181523 3584 181535 3587
rect 225560 3584 225588 3624
rect 234834 3612 234840 3624
rect 234892 3612 234898 3664
rect 234926 3612 234932 3664
rect 234984 3652 234990 3664
rect 234984 3624 241228 3652
rect 234984 3612 234990 3624
rect 181523 3556 225588 3584
rect 181523 3553 181535 3556
rect 181477 3547 181535 3553
rect 225634 3544 225640 3596
rect 225692 3584 225698 3596
rect 234742 3584 234748 3596
rect 225692 3556 234748 3584
rect 225692 3544 225698 3556
rect 234742 3544 234748 3556
rect 234800 3544 234806 3596
rect 235021 3587 235079 3593
rect 235021 3553 235033 3587
rect 235067 3584 235079 3587
rect 235297 3587 235355 3593
rect 235297 3584 235309 3587
rect 235067 3556 235309 3584
rect 235067 3553 235079 3556
rect 235021 3547 235079 3553
rect 235297 3553 235309 3556
rect 235343 3553 235355 3587
rect 235297 3547 235355 3553
rect 235386 3544 235392 3596
rect 235444 3584 235450 3596
rect 238422 3584 238428 3596
rect 235444 3556 238428 3584
rect 235444 3544 235450 3556
rect 238422 3544 238428 3556
rect 238480 3544 238486 3596
rect 177291 3488 181336 3516
rect 181385 3519 181443 3525
rect 177291 3485 177303 3488
rect 177245 3479 177303 3485
rect 181385 3485 181397 3519
rect 181431 3516 181443 3519
rect 186721 3519 186779 3525
rect 181431 3488 186672 3516
rect 181431 3485 181443 3488
rect 181385 3479 181443 3485
rect 152543 3420 157968 3448
rect 152543 3417 152555 3420
rect 152497 3411 152555 3417
rect 158106 3408 158112 3460
rect 158164 3448 158170 3460
rect 186534 3448 186540 3460
rect 158164 3420 186540 3448
rect 158164 3408 158170 3420
rect 186534 3408 186540 3420
rect 186592 3408 186598 3460
rect 186644 3448 186672 3488
rect 186721 3485 186733 3519
rect 186767 3516 186779 3519
rect 206133 3519 206191 3525
rect 206133 3516 206145 3519
rect 186767 3488 206145 3516
rect 186767 3485 186779 3488
rect 186721 3479 186779 3485
rect 206133 3485 206145 3488
rect 206179 3485 206191 3519
rect 206133 3479 206191 3485
rect 206222 3476 206228 3528
rect 206280 3516 206286 3528
rect 236674 3516 236680 3528
rect 206280 3488 236680 3516
rect 206280 3476 206286 3488
rect 236674 3476 236680 3488
rect 236732 3476 236738 3528
rect 236766 3476 236772 3528
rect 236824 3516 236830 3528
rect 241090 3516 241096 3528
rect 236824 3488 241096 3516
rect 236824 3476 236830 3488
rect 241090 3476 241096 3488
rect 241148 3476 241154 3528
rect 241200 3516 241228 3624
rect 243666 3612 243672 3664
rect 243724 3652 243730 3664
rect 243724 3624 247208 3652
rect 243724 3612 243730 3624
rect 247180 3584 247208 3624
rect 247254 3612 247260 3664
rect 247312 3652 247318 3664
rect 278721 3655 278779 3661
rect 247312 3624 278672 3652
rect 247312 3612 247318 3624
rect 268877 3587 268935 3593
rect 268877 3584 268889 3587
rect 247180 3556 268889 3584
rect 268877 3553 268889 3556
rect 268923 3553 268935 3587
rect 268877 3547 268935 3553
rect 273382 3544 273388 3596
rect 273440 3584 273446 3596
rect 278442 3584 278448 3596
rect 273440 3556 278448 3584
rect 273440 3544 273446 3556
rect 278442 3544 278448 3556
rect 278500 3544 278506 3596
rect 278644 3584 278672 3624
rect 278721 3621 278733 3655
rect 278767 3652 278779 3655
rect 285158 3652 285164 3664
rect 278767 3624 285164 3652
rect 278767 3621 278779 3624
rect 278721 3615 278779 3621
rect 285158 3612 285164 3624
rect 285216 3612 285222 3664
rect 285250 3612 285256 3664
rect 285308 3652 285314 3664
rect 289666 3652 289672 3664
rect 285308 3624 289672 3652
rect 285308 3612 285314 3624
rect 289666 3612 289672 3624
rect 289724 3612 289730 3664
rect 295738 3612 295744 3664
rect 295796 3652 295802 3664
rect 313862 3652 313868 3664
rect 295796 3624 313868 3652
rect 295796 3612 295802 3624
rect 313862 3612 313868 3624
rect 313920 3612 313926 3664
rect 323246 3612 323252 3664
rect 323304 3652 323310 3664
rect 450666 3652 450672 3664
rect 323304 3624 450672 3652
rect 323304 3612 323310 3624
rect 450666 3612 450672 3624
rect 450724 3612 450730 3664
rect 281018 3584 281024 3596
rect 278644 3556 281024 3584
rect 281018 3544 281024 3556
rect 281076 3544 281082 3596
rect 282950 3544 282956 3596
rect 283008 3584 283014 3596
rect 287918 3584 287924 3596
rect 283008 3556 287924 3584
rect 283008 3544 283014 3556
rect 287918 3544 287924 3556
rect 287976 3544 287982 3596
rect 297118 3544 297124 3596
rect 297176 3584 297182 3596
rect 300985 3587 301043 3593
rect 297176 3556 300936 3584
rect 297176 3544 297182 3556
rect 249557 3519 249615 3525
rect 249557 3516 249569 3519
rect 241200 3488 249569 3516
rect 249557 3485 249569 3488
rect 249603 3485 249615 3519
rect 249557 3479 249615 3485
rect 265102 3476 265108 3528
rect 265160 3516 265166 3528
rect 278537 3519 278595 3525
rect 278537 3516 278549 3519
rect 265160 3488 278549 3516
rect 265160 3476 265166 3488
rect 278537 3485 278549 3488
rect 278583 3485 278595 3519
rect 278537 3479 278595 3485
rect 278629 3519 278687 3525
rect 278629 3485 278641 3519
rect 278675 3516 278687 3519
rect 282306 3516 282312 3528
rect 278675 3488 282312 3516
rect 278675 3485 278687 3488
rect 278629 3479 278687 3485
rect 282306 3476 282312 3488
rect 282364 3476 282370 3528
rect 292702 3476 292708 3528
rect 292760 3516 292766 3528
rect 300798 3516 300804 3528
rect 292760 3488 300804 3516
rect 292760 3476 292766 3488
rect 300798 3476 300804 3488
rect 300856 3476 300862 3528
rect 300908 3516 300936 3556
rect 300985 3553 300997 3587
rect 301031 3584 301043 3587
rect 307882 3584 307888 3596
rect 301031 3556 307888 3584
rect 301031 3553 301043 3556
rect 300985 3547 301043 3553
rect 307882 3544 307888 3556
rect 307940 3544 307946 3596
rect 309538 3544 309544 3596
rect 309596 3584 309602 3596
rect 370445 3587 370503 3593
rect 370445 3584 370457 3587
rect 309596 3556 370457 3584
rect 309596 3544 309602 3556
rect 370445 3553 370457 3556
rect 370491 3553 370503 3587
rect 370445 3547 370503 3553
rect 370626 3544 370632 3596
rect 370684 3584 370690 3596
rect 383969 3587 384027 3593
rect 383969 3584 383981 3587
rect 370684 3556 383981 3584
rect 370684 3544 370690 3556
rect 383969 3553 383981 3556
rect 384015 3553 384027 3587
rect 383969 3547 384027 3553
rect 384061 3587 384119 3593
rect 384061 3553 384073 3587
rect 384107 3584 384119 3587
rect 454162 3584 454168 3596
rect 384107 3556 454168 3584
rect 384107 3553 384119 3556
rect 384061 3547 384119 3553
rect 454162 3544 454168 3556
rect 454220 3544 454226 3596
rect 318554 3516 318560 3528
rect 300908 3488 318560 3516
rect 318554 3476 318560 3488
rect 318612 3476 318618 3528
rect 321774 3476 321780 3528
rect 321832 3516 321838 3528
rect 326009 3519 326067 3525
rect 326009 3516 326021 3519
rect 321832 3488 326021 3516
rect 321832 3476 321838 3488
rect 326009 3485 326021 3488
rect 326055 3485 326067 3519
rect 326009 3479 326067 3485
rect 326098 3476 326104 3528
rect 326156 3516 326162 3528
rect 326193 3519 326251 3525
rect 326193 3516 326205 3519
rect 326156 3488 326205 3516
rect 326156 3476 326162 3488
rect 326193 3485 326205 3488
rect 326239 3485 326251 3519
rect 326193 3479 326251 3485
rect 326285 3519 326343 3525
rect 326285 3485 326297 3519
rect 326331 3516 326343 3519
rect 341373 3519 341431 3525
rect 341373 3516 341385 3519
rect 326331 3488 341385 3516
rect 326331 3485 326343 3488
rect 326285 3479 326343 3485
rect 341373 3485 341385 3488
rect 341419 3485 341431 3519
rect 341373 3479 341431 3485
rect 341462 3476 341468 3528
rect 341520 3516 341526 3528
rect 350757 3519 350815 3525
rect 350757 3516 350769 3519
rect 341520 3488 350769 3516
rect 341520 3476 341526 3488
rect 350757 3485 350769 3488
rect 350803 3485 350815 3519
rect 350757 3479 350815 3485
rect 351122 3476 351128 3528
rect 351180 3516 351186 3528
rect 360506 3516 360512 3528
rect 351180 3488 360512 3516
rect 351180 3476 351186 3488
rect 360506 3476 360512 3488
rect 360564 3476 360570 3528
rect 360598 3476 360604 3528
rect 360656 3516 360662 3528
rect 360693 3519 360751 3525
rect 360693 3516 360705 3519
rect 360656 3488 360705 3516
rect 360656 3476 360662 3488
rect 360693 3485 360705 3488
rect 360739 3485 360751 3519
rect 360693 3479 360751 3485
rect 360782 3476 360788 3528
rect 360840 3516 360846 3528
rect 370166 3516 370172 3528
rect 360840 3488 370172 3516
rect 360840 3476 360846 3488
rect 370166 3476 370172 3488
rect 370224 3476 370230 3528
rect 370258 3476 370264 3528
rect 370316 3516 370322 3528
rect 370353 3519 370411 3525
rect 370353 3516 370365 3519
rect 370316 3488 370365 3516
rect 370316 3476 370322 3488
rect 370353 3485 370365 3488
rect 370399 3485 370411 3519
rect 370353 3479 370411 3485
rect 370534 3476 370540 3528
rect 370592 3516 370598 3528
rect 457750 3516 457756 3528
rect 370592 3488 457756 3516
rect 370592 3476 370598 3488
rect 457750 3476 457756 3488
rect 457808 3476 457814 3528
rect 186810 3448 186816 3460
rect 186644 3420 186816 3448
rect 186810 3408 186816 3420
rect 186868 3408 186874 3460
rect 187089 3451 187147 3457
rect 187089 3417 187101 3451
rect 187135 3448 187147 3451
rect 196286 3448 196292 3460
rect 187135 3420 196292 3448
rect 187135 3417 187147 3420
rect 187089 3411 187147 3417
rect 196286 3408 196292 3420
rect 196344 3408 196350 3460
rect 196378 3408 196384 3460
rect 196436 3448 196442 3460
rect 196470 3448 196476 3460
rect 196436 3420 196476 3448
rect 196436 3408 196442 3420
rect 196470 3408 196476 3420
rect 196528 3408 196534 3460
rect 206038 3408 206044 3460
rect 206096 3448 206102 3460
rect 209905 3451 209963 3457
rect 209905 3448 209917 3451
rect 206096 3420 209917 3448
rect 206096 3408 206102 3420
rect 209905 3417 209917 3420
rect 209951 3417 209963 3451
rect 209905 3411 209963 3417
rect 210181 3451 210239 3457
rect 210181 3417 210193 3451
rect 210227 3448 210239 3451
rect 225361 3451 225419 3457
rect 225361 3448 225373 3451
rect 210227 3420 225373 3448
rect 210227 3417 210239 3420
rect 210181 3411 210239 3417
rect 225361 3417 225373 3420
rect 225407 3417 225419 3451
rect 225361 3411 225419 3417
rect 225453 3451 225511 3457
rect 225453 3417 225465 3451
rect 225499 3448 225511 3451
rect 254706 3448 254712 3460
rect 225499 3420 254712 3448
rect 225499 3417 225511 3420
rect 225453 3411 225511 3417
rect 254706 3408 254712 3420
rect 254764 3408 254770 3460
rect 261514 3408 261520 3460
rect 261572 3448 261578 3460
rect 262618 3448 262624 3460
rect 261572 3420 262624 3448
rect 261572 3408 261578 3420
rect 262618 3408 262624 3420
rect 262676 3408 262682 3460
rect 275685 3451 275743 3457
rect 275685 3448 275697 3451
rect 262728 3420 275697 3448
rect 33170 3340 33176 3392
rect 33228 3380 33234 3392
rect 40165 3383 40223 3389
rect 40165 3380 40177 3383
rect 33228 3352 40177 3380
rect 33228 3340 33234 3352
rect 40165 3349 40177 3352
rect 40211 3349 40223 3383
rect 40165 3343 40223 3349
rect 40254 3340 40260 3392
rect 40312 3380 40318 3392
rect 44765 3383 44823 3389
rect 44765 3380 44777 3383
rect 40312 3352 44777 3380
rect 40312 3340 40318 3352
rect 44765 3349 44777 3352
rect 44811 3349 44823 3383
rect 44765 3343 44823 3349
rect 45038 3340 45044 3392
rect 45096 3380 45102 3392
rect 45958 3380 45964 3392
rect 45096 3352 45964 3380
rect 45096 3340 45102 3352
rect 45958 3340 45964 3352
rect 46016 3340 46022 3392
rect 61690 3340 61696 3392
rect 61748 3380 61754 3392
rect 62518 3380 62524 3392
rect 61748 3352 62524 3380
rect 61748 3340 61754 3352
rect 62518 3340 62524 3352
rect 62576 3340 62582 3392
rect 64082 3340 64088 3392
rect 64140 3380 64146 3392
rect 65186 3380 65192 3392
rect 64140 3352 65192 3380
rect 64140 3340 64146 3352
rect 65186 3340 65192 3352
rect 65244 3340 65250 3392
rect 65278 3340 65284 3392
rect 65336 3380 65342 3392
rect 235110 3380 235116 3392
rect 65336 3352 235116 3380
rect 65336 3340 65342 3352
rect 235110 3340 235116 3352
rect 235168 3340 235174 3392
rect 235202 3340 235208 3392
rect 235260 3380 235266 3392
rect 237042 3380 237048 3392
rect 235260 3352 237048 3380
rect 235260 3340 235266 3352
rect 237042 3340 237048 3352
rect 237100 3340 237106 3392
rect 237134 3340 237140 3392
rect 237192 3380 237198 3392
rect 243850 3380 243856 3392
rect 237192 3352 243856 3380
rect 237192 3340 237198 3352
rect 243850 3340 243856 3352
rect 243908 3340 243914 3392
rect 257926 3340 257932 3392
rect 257984 3380 257990 3392
rect 262728 3380 262756 3420
rect 275685 3417 275697 3420
rect 275731 3417 275743 3451
rect 275685 3411 275743 3417
rect 275774 3408 275780 3460
rect 275832 3448 275838 3460
rect 275832 3420 278672 3448
rect 275832 3408 275838 3420
rect 257984 3352 262756 3380
rect 257984 3340 257990 3352
rect 262894 3340 262900 3392
rect 262952 3380 262958 3392
rect 264553 3383 264611 3389
rect 264553 3380 264565 3383
rect 262952 3352 264565 3380
rect 262952 3340 262958 3352
rect 264553 3349 264565 3352
rect 264599 3349 264611 3383
rect 264553 3343 264611 3349
rect 272186 3340 272192 3392
rect 272244 3380 272250 3392
rect 278537 3383 278595 3389
rect 278537 3380 278549 3383
rect 272244 3352 278549 3380
rect 272244 3340 272250 3352
rect 278537 3349 278549 3352
rect 278583 3349 278595 3383
rect 278644 3380 278672 3420
rect 280098 3408 280104 3460
rect 280156 3448 280162 3460
rect 288102 3448 288108 3460
rect 280156 3420 288108 3448
rect 280156 3408 280162 3420
rect 288102 3408 288108 3420
rect 288160 3408 288166 3460
rect 291414 3408 291420 3460
rect 291472 3448 291478 3460
rect 293622 3448 293628 3460
rect 291472 3420 293628 3448
rect 291472 3408 291478 3420
rect 293622 3408 293628 3420
rect 293680 3408 293686 3460
rect 294358 3408 294364 3460
rect 294416 3448 294422 3460
rect 300985 3451 301043 3457
rect 300985 3448 300997 3451
rect 294416 3420 300997 3448
rect 294416 3408 294422 3420
rect 300985 3417 300997 3420
rect 301031 3417 301043 3451
rect 300985 3411 301043 3417
rect 301077 3451 301135 3457
rect 301077 3417 301089 3451
rect 301123 3448 301135 3451
rect 310274 3448 310280 3460
rect 301123 3420 310280 3448
rect 301123 3417 301135 3420
rect 301077 3411 301135 3417
rect 310274 3408 310280 3420
rect 310332 3408 310338 3460
rect 310918 3408 310924 3460
rect 310976 3448 310982 3460
rect 389946 3448 389952 3460
rect 310976 3420 389952 3448
rect 310976 3408 310982 3420
rect 389946 3408 389952 3420
rect 390004 3408 390010 3460
rect 390041 3451 390099 3457
rect 390041 3417 390053 3451
rect 390087 3448 390099 3451
rect 461338 3448 461344 3460
rect 390087 3420 461344 3448
rect 390087 3417 390099 3420
rect 390041 3411 390099 3417
rect 461338 3408 461344 3420
rect 461396 3408 461402 3460
rect 286722 3380 286728 3392
rect 278644 3352 286728 3380
rect 278537 3343 278595 3349
rect 286722 3340 286728 3352
rect 286780 3340 286786 3392
rect 293714 3340 293720 3392
rect 293772 3380 293778 3392
rect 298501 3383 298559 3389
rect 298501 3380 298513 3383
rect 293772 3352 298513 3380
rect 293772 3340 293778 3352
rect 298501 3349 298513 3352
rect 298547 3349 298559 3383
rect 298501 3343 298559 3349
rect 298593 3383 298651 3389
rect 298593 3349 298605 3383
rect 298639 3380 298651 3383
rect 303098 3380 303104 3392
rect 298639 3352 303104 3380
rect 298639 3349 298651 3352
rect 298593 3343 298651 3349
rect 303098 3340 303104 3352
rect 303156 3340 303162 3392
rect 319106 3340 319112 3392
rect 319164 3380 319170 3392
rect 429230 3380 429236 3392
rect 319164 3352 429236 3380
rect 319164 3340 319170 3352
rect 429230 3340 429236 3352
rect 429288 3340 429294 3392
rect 433830 3340 433836 3392
rect 433888 3380 433894 3392
rect 451678 3380 451684 3392
rect 433888 3352 451684 3380
rect 433888 3340 433894 3352
rect 451678 3340 451684 3352
rect 451736 3340 451742 3392
rect 466582 3340 466588 3392
rect 466640 3380 466646 3392
rect 480658 3380 480664 3392
rect 466640 3352 480664 3380
rect 466640 3340 466646 3352
rect 480658 3340 480664 3352
rect 480716 3340 480722 3392
rect 1600 3216 583316 3312
rect 28386 3136 28392 3188
rect 28444 3176 28450 3188
rect 29398 3176 29404 3188
rect 28444 3148 29404 3176
rect 28444 3136 28450 3148
rect 29398 3136 29404 3148
rect 29456 3136 29462 3188
rect 36393 3179 36451 3185
rect 36393 3145 36405 3179
rect 36439 3176 36451 3179
rect 45961 3179 46019 3185
rect 45961 3176 45973 3179
rect 36439 3148 45973 3176
rect 36439 3145 36451 3148
rect 36393 3139 36451 3145
rect 45961 3145 45973 3148
rect 46007 3145 46019 3179
rect 45961 3139 46019 3145
rect 56265 3179 56323 3185
rect 56265 3145 56277 3179
rect 56311 3176 56323 3179
rect 65281 3179 65339 3185
rect 65281 3176 65293 3179
rect 56311 3148 65293 3176
rect 56311 3145 56323 3148
rect 56265 3139 56323 3145
rect 65281 3145 65293 3148
rect 65327 3145 65339 3179
rect 65281 3139 65339 3145
rect 68774 3136 68780 3188
rect 68832 3176 68838 3188
rect 69418 3176 69424 3188
rect 68832 3148 69424 3176
rect 68832 3136 68838 3148
rect 69418 3136 69424 3148
rect 69476 3136 69482 3188
rect 71166 3136 71172 3188
rect 71224 3176 71230 3188
rect 72178 3176 72184 3188
rect 71224 3148 72184 3176
rect 71224 3136 71230 3148
rect 72178 3136 72184 3148
rect 72236 3136 72242 3188
rect 72362 3136 72368 3188
rect 72420 3176 72426 3188
rect 72420 3148 187040 3176
rect 72420 3136 72426 3148
rect 21210 3068 21216 3120
rect 21268 3108 21274 3120
rect 22498 3108 22504 3120
rect 21268 3080 22504 3108
rect 21268 3068 21274 3080
rect 22498 3068 22504 3080
rect 22556 3068 22562 3120
rect 40165 3111 40223 3117
rect 40165 3077 40177 3111
rect 40211 3108 40223 3111
rect 45869 3111 45927 3117
rect 45869 3108 45881 3111
rect 40211 3080 45881 3108
rect 40211 3077 40223 3080
rect 40165 3071 40223 3077
rect 45869 3077 45881 3080
rect 45915 3077 45927 3111
rect 45869 3071 45927 3077
rect 56357 3111 56415 3117
rect 56357 3077 56369 3111
rect 56403 3108 56415 3111
rect 65189 3111 65247 3117
rect 65189 3108 65201 3111
rect 56403 3080 65201 3108
rect 56403 3077 56415 3080
rect 56357 3071 56415 3077
rect 65189 3077 65201 3080
rect 65235 3077 65247 3111
rect 65189 3071 65247 3077
rect 77146 3068 77152 3120
rect 77204 3108 77210 3120
rect 77698 3108 77704 3120
rect 77204 3080 77704 3108
rect 77204 3068 77210 3080
rect 77698 3068 77704 3080
rect 77756 3068 77762 3120
rect 78342 3068 78348 3120
rect 78400 3108 78406 3120
rect 79078 3108 79084 3120
rect 78400 3080 79084 3108
rect 78400 3068 78406 3080
rect 79078 3068 79084 3080
rect 79136 3068 79142 3120
rect 80734 3068 80740 3120
rect 80792 3108 80798 3120
rect 81838 3108 81844 3120
rect 80792 3080 81844 3108
rect 80792 3068 80798 3080
rect 81838 3068 81844 3080
rect 81896 3068 81902 3120
rect 186905 3111 186963 3117
rect 186905 3108 186917 3111
rect 85352 3080 186917 3108
rect 79538 3000 79544 3052
rect 79596 3040 79602 3052
rect 85352 3040 85380 3080
rect 186905 3077 186917 3080
rect 186951 3077 186963 3111
rect 187012 3108 187040 3148
rect 187178 3136 187184 3188
rect 187236 3176 187242 3188
rect 196194 3176 196200 3188
rect 187236 3148 196200 3176
rect 187236 3136 187242 3148
rect 196194 3136 196200 3148
rect 196252 3136 196258 3188
rect 196304 3148 196608 3176
rect 196304 3108 196332 3148
rect 187012 3080 196332 3108
rect 196580 3108 196608 3148
rect 196746 3136 196752 3188
rect 196804 3176 196810 3188
rect 205854 3176 205860 3188
rect 196804 3148 205860 3176
rect 196804 3136 196810 3148
rect 205854 3136 205860 3148
rect 205912 3136 205918 3188
rect 245138 3176 245144 3188
rect 205964 3148 245144 3176
rect 205964 3108 205992 3148
rect 245138 3136 245144 3148
rect 245196 3136 245202 3188
rect 253142 3136 253148 3188
rect 253200 3176 253206 3188
rect 254154 3176 254160 3188
rect 253200 3148 254160 3176
rect 253200 3136 253206 3148
rect 254154 3136 254160 3148
rect 254212 3136 254218 3188
rect 270990 3136 270996 3188
rect 271048 3176 271054 3188
rect 271048 3148 278120 3176
rect 271048 3136 271054 3148
rect 196580 3080 205992 3108
rect 206041 3111 206099 3117
rect 186905 3071 186963 3077
rect 206041 3077 206053 3111
rect 206087 3108 206099 3111
rect 246610 3108 246616 3120
rect 206087 3080 246616 3108
rect 206087 3077 206099 3080
rect 206041 3071 206099 3077
rect 246610 3068 246616 3080
rect 246668 3068 246674 3120
rect 278092 3108 278120 3148
rect 278166 3136 278172 3188
rect 278224 3176 278230 3188
rect 286814 3176 286820 3188
rect 278224 3148 286820 3176
rect 278224 3136 278230 3148
rect 286814 3136 286820 3148
rect 286872 3136 286878 3188
rect 294082 3136 294088 3188
rect 294140 3176 294146 3188
rect 301077 3179 301135 3185
rect 301077 3176 301089 3179
rect 294140 3148 301089 3176
rect 294140 3136 294146 3148
rect 301077 3145 301089 3148
rect 301123 3145 301135 3179
rect 301077 3139 301135 3145
rect 319198 3136 319204 3188
rect 319256 3176 319262 3188
rect 425642 3176 425648 3188
rect 319256 3148 425648 3176
rect 319256 3136 319262 3148
rect 425642 3136 425648 3148
rect 425700 3136 425706 3188
rect 285526 3108 285532 3120
rect 278092 3080 285532 3108
rect 285526 3068 285532 3080
rect 285584 3068 285590 3120
rect 292334 3068 292340 3120
rect 292392 3108 292398 3120
rect 296014 3108 296020 3120
rect 292392 3080 296020 3108
rect 292392 3068 292398 3080
rect 296014 3068 296020 3080
rect 296072 3068 296078 3120
rect 317818 3068 317824 3120
rect 317876 3108 317882 3120
rect 422054 3108 422060 3120
rect 317876 3080 422060 3108
rect 317876 3068 317882 3080
rect 422054 3068 422060 3080
rect 422112 3068 422118 3120
rect 432818 3108 432824 3120
rect 422256 3080 432824 3108
rect 79596 3012 85380 3040
rect 79596 3000 79602 3012
rect 85426 3000 85432 3052
rect 85484 3040 85490 3052
rect 85978 3040 85984 3052
rect 85484 3012 85984 3040
rect 85484 3000 85490 3012
rect 85978 3000 85984 3012
rect 86036 3000 86042 3052
rect 86622 3000 86628 3052
rect 86680 3040 86686 3052
rect 87358 3040 87364 3052
rect 86680 3012 87364 3040
rect 86680 3000 86686 3012
rect 87358 3000 87364 3012
rect 87416 3000 87422 3052
rect 87818 3000 87824 3052
rect 87876 3040 87882 3052
rect 88738 3040 88744 3052
rect 87876 3012 88744 3040
rect 87876 3000 87882 3012
rect 88738 3000 88744 3012
rect 88796 3000 88802 3052
rect 89014 3000 89020 3052
rect 89072 3040 89078 3052
rect 90118 3040 90124 3052
rect 89072 3012 90124 3040
rect 89072 3000 89078 3012
rect 90118 3000 90124 3012
rect 90176 3000 90182 3052
rect 99502 3000 99508 3052
rect 99560 3040 99566 3052
rect 99778 3040 99784 3052
rect 99560 3012 99784 3040
rect 99560 3000 99566 3012
rect 99778 3000 99784 3012
rect 99836 3000 99842 3052
rect 102078 3000 102084 3052
rect 102136 3040 102142 3052
rect 102538 3040 102544 3052
rect 102136 3012 102544 3040
rect 102136 3000 102142 3012
rect 102538 3000 102544 3012
rect 102596 3000 102602 3052
rect 186810 3040 186816 3052
rect 102648 3012 186816 3040
rect 54514 2932 54520 2984
rect 54572 2972 54578 2984
rect 55618 2972 55624 2984
rect 54572 2944 55624 2972
rect 54572 2932 54578 2944
rect 55618 2932 55624 2944
rect 55676 2932 55682 2984
rect 75033 2975 75091 2981
rect 75033 2941 75045 2975
rect 75079 2972 75091 2975
rect 84601 2975 84659 2981
rect 84601 2972 84613 2975
rect 75079 2944 84613 2972
rect 75079 2941 75091 2944
rect 75033 2935 75091 2941
rect 84601 2941 84613 2944
rect 84647 2941 84659 2975
rect 84601 2935 84659 2941
rect 90210 2932 90216 2984
rect 90268 2972 90274 2984
rect 102648 2972 102676 3012
rect 186810 3000 186816 3012
rect 186868 3000 186874 3052
rect 186997 3043 187055 3049
rect 186997 3009 187009 3043
rect 187043 3040 187055 3043
rect 196197 3043 196255 3049
rect 196197 3040 196209 3043
rect 187043 3012 196209 3040
rect 187043 3009 187055 3012
rect 186997 3003 187055 3009
rect 196197 3009 196209 3012
rect 196243 3009 196255 3043
rect 196197 3003 196255 3009
rect 196565 3043 196623 3049
rect 196565 3009 196577 3043
rect 196611 3040 196623 3043
rect 205949 3043 206007 3049
rect 205949 3040 205961 3043
rect 196611 3012 205961 3040
rect 196611 3009 196623 3012
rect 196565 3003 196623 3009
rect 205949 3009 205961 3012
rect 205995 3009 206007 3043
rect 205949 3003 206007 3009
rect 207694 3000 207700 3052
rect 207752 3040 207758 3052
rect 247898 3040 247904 3052
rect 207752 3012 247904 3040
rect 207752 3000 207758 3012
rect 247898 3000 247904 3012
rect 247956 3000 247962 3052
rect 250842 3000 250848 3052
rect 250900 3040 250906 3052
rect 251578 3040 251584 3052
rect 250900 3012 251584 3040
rect 250900 3000 250906 3012
rect 251578 3000 251584 3012
rect 251636 3000 251642 3052
rect 275685 3043 275743 3049
rect 275685 3009 275697 3043
rect 275731 3040 275743 3043
rect 278445 3043 278503 3049
rect 278445 3040 278457 3043
rect 275731 3012 278457 3040
rect 275731 3009 275743 3012
rect 275685 3003 275743 3009
rect 278445 3009 278457 3012
rect 278491 3009 278503 3043
rect 278445 3003 278503 3009
rect 278537 3043 278595 3049
rect 278537 3009 278549 3043
rect 278583 3040 278595 3043
rect 286354 3040 286360 3052
rect 278583 3012 286360 3040
rect 278583 3009 278595 3012
rect 278537 3003 278595 3009
rect 286354 3000 286360 3012
rect 286412 3000 286418 3052
rect 294174 3000 294180 3052
rect 294232 3040 294238 3052
rect 294232 3012 302040 3040
rect 294232 3000 294238 3012
rect 103829 2975 103887 2981
rect 103829 2972 103841 2975
rect 90268 2944 102676 2972
rect 102740 2944 103841 2972
rect 90268 2932 90274 2944
rect 75125 2907 75183 2913
rect 75125 2873 75137 2907
rect 75171 2904 75183 2907
rect 84509 2907 84567 2913
rect 84509 2904 84521 2907
rect 75171 2876 84521 2904
rect 75171 2873 75183 2876
rect 75125 2867 75183 2873
rect 84509 2873 84521 2876
rect 84555 2873 84567 2907
rect 84509 2867 84567 2873
rect 93709 2907 93767 2913
rect 93709 2873 93721 2907
rect 93755 2904 93767 2907
rect 102740 2904 102768 2944
rect 103829 2941 103841 2944
rect 103875 2941 103887 2975
rect 103829 2935 103887 2941
rect 105666 2932 105672 2984
rect 105724 2972 105730 2984
rect 106678 2972 106684 2984
rect 105724 2944 106684 2972
rect 105724 2932 105730 2944
rect 106678 2932 106684 2944
rect 106736 2932 106742 2984
rect 106862 2932 106868 2984
rect 106920 2972 106926 2984
rect 107966 2972 107972 2984
rect 106920 2944 107972 2972
rect 106920 2932 106926 2944
rect 107966 2932 107972 2944
rect 108024 2932 108030 2984
rect 108720 2944 187040 2972
rect 93755 2876 102768 2904
rect 93755 2873 93767 2876
rect 93709 2867 93767 2873
rect 103274 2864 103280 2916
rect 103332 2904 103338 2916
rect 103918 2904 103924 2916
rect 103332 2876 103924 2904
rect 103332 2864 103338 2876
rect 103918 2864 103924 2876
rect 103976 2864 103982 2916
rect 104470 2864 104476 2916
rect 104528 2904 104534 2916
rect 108613 2907 108671 2913
rect 108613 2904 108625 2907
rect 104528 2876 108625 2904
rect 104528 2864 104534 2876
rect 108613 2873 108625 2876
rect 108659 2873 108671 2907
rect 108613 2867 108671 2873
rect 97386 2796 97392 2848
rect 97444 2836 97450 2848
rect 108720 2836 108748 2944
rect 111646 2864 111652 2916
rect 111704 2904 111710 2916
rect 113489 2907 113547 2913
rect 113489 2904 113501 2907
rect 111704 2876 113501 2904
rect 111704 2864 111710 2876
rect 113489 2873 113501 2876
rect 113535 2873 113547 2907
rect 186813 2907 186871 2913
rect 186813 2904 186825 2907
rect 113489 2867 113547 2873
rect 113596 2876 186825 2904
rect 97444 2808 108748 2836
rect 108797 2839 108855 2845
rect 97444 2796 97450 2808
rect 108797 2805 108809 2839
rect 108843 2836 108855 2839
rect 112753 2839 112811 2845
rect 112753 2836 112765 2839
rect 108843 2808 112765 2836
rect 108843 2805 108855 2808
rect 108797 2799 108855 2805
rect 112753 2805 112765 2808
rect 112799 2805 112811 2839
rect 112753 2799 112811 2805
rect 112842 2796 112848 2848
rect 112900 2836 112906 2848
rect 113302 2836 113308 2848
rect 112900 2808 113308 2836
rect 112900 2796 112906 2808
rect 113302 2796 113308 2808
rect 113360 2796 113366 2848
rect 113397 2839 113455 2845
rect 113397 2805 113409 2839
rect 113443 2836 113455 2839
rect 113596 2836 113624 2876
rect 186813 2873 186825 2876
rect 186859 2873 186871 2907
rect 186813 2867 186871 2873
rect 186905 2907 186963 2913
rect 186905 2873 186917 2907
rect 186951 2873 186963 2907
rect 187012 2904 187040 2944
rect 187086 2932 187092 2984
rect 187144 2972 187150 2984
rect 195918 2972 195924 2984
rect 187144 2944 195924 2972
rect 187144 2932 187150 2944
rect 195918 2932 195924 2944
rect 195976 2932 195982 2984
rect 198497 2975 198555 2981
rect 198497 2941 198509 2975
rect 198543 2972 198555 2975
rect 205857 2975 205915 2981
rect 205857 2972 205869 2975
rect 198543 2944 205869 2972
rect 198543 2941 198555 2944
rect 198497 2935 198555 2941
rect 205857 2941 205869 2944
rect 205903 2941 205915 2975
rect 205857 2935 205915 2941
rect 206133 2975 206191 2981
rect 206133 2941 206145 2975
rect 206179 2972 206191 2975
rect 250658 2972 250664 2984
rect 206179 2944 250664 2972
rect 206179 2941 206191 2944
rect 206133 2935 206191 2941
rect 250658 2932 250664 2944
rect 250716 2932 250722 2984
rect 274578 2932 274584 2984
rect 274636 2972 274642 2984
rect 286630 2972 286636 2984
rect 274636 2944 286636 2972
rect 274636 2932 274642 2944
rect 286630 2932 286636 2944
rect 286688 2932 286694 2984
rect 291598 2932 291604 2984
rect 291656 2972 291662 2984
rect 294818 2972 294824 2984
rect 291656 2944 294824 2972
rect 291656 2932 291662 2944
rect 294818 2932 294824 2944
rect 294876 2932 294882 2984
rect 196197 2907 196255 2913
rect 196197 2904 196209 2907
rect 187012 2876 196209 2904
rect 186905 2867 186963 2873
rect 196197 2873 196209 2876
rect 196243 2873 196255 2907
rect 196197 2867 196255 2873
rect 196473 2907 196531 2913
rect 196473 2873 196485 2907
rect 196519 2904 196531 2907
rect 252130 2904 252136 2916
rect 196519 2876 252136 2904
rect 196519 2873 196531 2876
rect 196473 2867 196531 2873
rect 113443 2808 113624 2836
rect 113673 2839 113731 2845
rect 113443 2805 113455 2808
rect 113397 2799 113455 2805
rect 113673 2805 113685 2839
rect 113719 2836 113731 2839
rect 186920 2836 186948 2867
rect 252130 2864 252136 2876
rect 252188 2864 252194 2916
rect 276970 2864 276976 2916
rect 277028 2904 277034 2916
rect 279914 2904 279920 2916
rect 277028 2876 279920 2904
rect 277028 2864 277034 2876
rect 279914 2864 279920 2876
rect 279972 2864 279978 2916
rect 280558 2864 280564 2916
rect 280616 2904 280622 2916
rect 283962 2904 283968 2916
rect 280616 2876 283968 2904
rect 280616 2864 280622 2876
rect 283962 2864 283968 2876
rect 284020 2864 284026 2916
rect 292978 2864 292984 2916
rect 293036 2904 293042 2916
rect 301902 2904 301908 2916
rect 293036 2876 301908 2904
rect 293036 2864 293042 2876
rect 301902 2864 301908 2876
rect 301960 2864 301966 2916
rect 302012 2904 302040 3012
rect 316438 3000 316444 3052
rect 316496 3040 316502 3052
rect 418466 3040 418472 3052
rect 316496 3012 418472 3040
rect 316496 3000 316502 3012
rect 418466 3000 418472 3012
rect 418524 3000 418530 3052
rect 418745 3043 418803 3049
rect 418745 3009 418757 3043
rect 418791 3040 418803 3043
rect 422256 3040 422284 3080
rect 432818 3068 432824 3080
rect 432876 3068 432882 3120
rect 418791 3012 422284 3040
rect 418791 3009 418803 3012
rect 418745 3003 418803 3009
rect 315058 2932 315064 2984
rect 315116 2972 315122 2984
rect 355081 2975 355139 2981
rect 355081 2972 355093 2975
rect 315116 2944 355093 2972
rect 315116 2932 315122 2944
rect 355081 2941 355093 2944
rect 355127 2941 355139 2975
rect 355262 2972 355268 2984
rect 355223 2944 355268 2972
rect 355081 2935 355139 2941
rect 355262 2932 355268 2944
rect 355320 2932 355326 2984
rect 355357 2975 355415 2981
rect 355357 2941 355369 2975
rect 355403 2972 355415 2975
rect 355403 2944 404160 2972
rect 355403 2941 355415 2944
rect 355357 2935 355415 2941
rect 306686 2904 306692 2916
rect 302012 2876 306692 2904
rect 306686 2864 306692 2876
rect 306744 2864 306750 2916
rect 313678 2864 313684 2916
rect 313736 2904 313742 2916
rect 404132 2904 404160 2944
rect 406874 2932 406880 2984
rect 406932 2972 406938 2984
rect 411658 2972 411664 2984
rect 406932 2944 411664 2972
rect 406932 2932 406938 2944
rect 411658 2932 411664 2944
rect 411716 2932 411722 2984
rect 414602 2932 414608 2984
rect 414660 2972 414666 2984
rect 424078 2972 424084 2984
rect 414660 2944 424084 2972
rect 414660 2932 414666 2944
rect 424078 2932 424084 2944
rect 424136 2932 424142 2984
rect 411382 2904 411388 2916
rect 313736 2876 401768 2904
rect 404132 2876 411388 2904
rect 313736 2864 313742 2876
rect 113719 2808 186948 2836
rect 186997 2839 187055 2845
rect 113719 2805 113731 2808
rect 113673 2799 113731 2805
rect 186997 2805 187009 2839
rect 187043 2836 187055 2839
rect 196289 2839 196347 2845
rect 196289 2836 196301 2839
rect 187043 2808 196301 2836
rect 187043 2805 187055 2808
rect 186997 2799 187055 2805
rect 196289 2805 196301 2808
rect 196335 2805 196347 2839
rect 196289 2799 196347 2805
rect 196378 2796 196384 2848
rect 196436 2836 196442 2848
rect 253418 2836 253424 2848
rect 196436 2808 253424 2836
rect 196436 2796 196442 2808
rect 253418 2796 253424 2808
rect 253476 2796 253482 2848
rect 268877 2839 268935 2845
rect 268877 2805 268889 2839
rect 268923 2836 268935 2839
rect 279270 2836 279276 2848
rect 268923 2808 279276 2836
rect 268923 2805 268935 2808
rect 268877 2799 268935 2805
rect 279270 2796 279276 2808
rect 279328 2796 279334 2848
rect 281754 2796 281760 2848
rect 281812 2836 281818 2848
rect 288194 2836 288200 2848
rect 281812 2808 288200 2836
rect 281812 2796 281818 2808
rect 288194 2796 288200 2808
rect 288252 2796 288258 2848
rect 293806 2796 293812 2848
rect 293864 2836 293870 2848
rect 298593 2839 298651 2845
rect 298593 2836 298605 2839
rect 293864 2808 298605 2836
rect 293864 2796 293870 2808
rect 298593 2805 298605 2808
rect 298639 2805 298651 2839
rect 298593 2799 298651 2805
rect 308250 2796 308256 2848
rect 308308 2836 308314 2848
rect 309081 2839 309139 2845
rect 309081 2836 309093 2839
rect 308308 2808 309093 2836
rect 308308 2796 308314 2808
rect 309081 2805 309093 2808
rect 309127 2805 309139 2839
rect 309081 2799 309139 2805
rect 311930 2796 311936 2848
rect 311988 2836 311994 2848
rect 364646 2836 364652 2848
rect 311988 2808 364652 2836
rect 311988 2796 311994 2808
rect 364646 2796 364652 2808
rect 364704 2796 364710 2848
rect 364738 2796 364744 2848
rect 364796 2836 364802 2848
rect 364796 2808 364841 2836
rect 364796 2796 364802 2808
rect 364922 2796 364928 2848
rect 364980 2836 364986 2848
rect 364980 2808 365025 2836
rect 364980 2796 364986 2808
rect 365106 2796 365112 2848
rect 365164 2836 365170 2848
rect 397122 2836 397128 2848
rect 365164 2808 397128 2836
rect 365164 2796 365170 2808
rect 397122 2796 397128 2808
rect 397180 2796 397186 2848
rect 401740 2836 401768 2876
rect 411382 2864 411388 2876
rect 411440 2864 411446 2916
rect 404206 2836 404212 2848
rect 401740 2808 404212 2836
rect 404206 2796 404212 2808
rect 404264 2796 404270 2848
rect 420030 2796 420036 2848
rect 420088 2836 420094 2848
rect 420861 2839 420919 2845
rect 420861 2836 420873 2839
rect 420088 2808 420873 2836
rect 420088 2796 420094 2808
rect 420861 2805 420873 2808
rect 420907 2805 420919 2839
rect 420861 2799 420919 2805
rect 1600 2672 583316 2768
rect 113489 2635 113547 2641
rect 113489 2601 113501 2635
rect 113535 2632 113547 2635
rect 113673 2635 113731 2641
rect 113673 2632 113685 2635
rect 113535 2604 113685 2632
rect 113535 2601 113547 2604
rect 113489 2595 113547 2601
rect 113673 2601 113685 2604
rect 113719 2601 113731 2635
rect 113673 2595 113731 2601
rect 122318 2592 122324 2644
rect 122376 2632 122382 2644
rect 123333 2635 123391 2641
rect 123333 2632 123345 2635
rect 122376 2604 123345 2632
rect 122376 2592 122382 2604
rect 123333 2601 123345 2604
rect 123379 2601 123391 2635
rect 123333 2595 123391 2601
rect 132809 2635 132867 2641
rect 132809 2601 132821 2635
rect 132855 2632 132867 2635
rect 133361 2635 133419 2641
rect 133361 2632 133373 2635
rect 132855 2604 133373 2632
rect 132855 2601 132867 2604
rect 132809 2595 132867 2601
rect 133361 2601 133373 2604
rect 133407 2601 133419 2635
rect 133361 2595 133419 2601
rect 142377 2635 142435 2641
rect 142377 2601 142389 2635
rect 142423 2632 142435 2635
rect 142745 2635 142803 2641
rect 142745 2632 142757 2635
rect 142423 2604 142757 2632
rect 142423 2601 142435 2604
rect 142377 2595 142435 2601
rect 142745 2601 142757 2604
rect 142791 2601 142803 2635
rect 142745 2595 142803 2601
rect 152129 2635 152187 2641
rect 152129 2601 152141 2635
rect 152175 2632 152187 2635
rect 152497 2635 152555 2641
rect 152497 2632 152509 2635
rect 152175 2604 152509 2632
rect 152175 2601 152187 2604
rect 152129 2595 152187 2601
rect 152497 2601 152509 2604
rect 152543 2601 152555 2635
rect 152497 2595 152555 2601
rect 161605 2635 161663 2641
rect 161605 2601 161617 2635
rect 161651 2632 161663 2635
rect 162065 2635 162123 2641
rect 162065 2632 162077 2635
rect 161651 2604 162077 2632
rect 161651 2601 161663 2604
rect 161605 2595 161663 2601
rect 162065 2601 162077 2604
rect 162111 2601 162123 2635
rect 162065 2595 162123 2601
rect 171449 2635 171507 2641
rect 171449 2601 171461 2635
rect 171495 2632 171507 2635
rect 171725 2635 171783 2641
rect 171725 2632 171737 2635
rect 171495 2604 171737 2632
rect 171495 2601 171507 2604
rect 171449 2595 171507 2601
rect 171725 2601 171737 2604
rect 171771 2601 171783 2635
rect 171725 2595 171783 2601
rect 181109 2635 181167 2641
rect 181109 2601 181121 2635
rect 181155 2632 181167 2635
rect 181385 2635 181443 2641
rect 181385 2632 181397 2635
rect 181155 2604 181397 2632
rect 181155 2601 181167 2604
rect 181109 2595 181167 2601
rect 181385 2601 181397 2604
rect 181431 2601 181443 2635
rect 181385 2595 181443 2601
rect 190769 2635 190827 2641
rect 190769 2601 190781 2635
rect 190815 2632 190827 2635
rect 191045 2635 191103 2641
rect 191045 2632 191057 2635
rect 190815 2604 191057 2632
rect 190815 2601 190827 2604
rect 190769 2595 190827 2601
rect 191045 2601 191057 2604
rect 191091 2601 191103 2635
rect 196102 2632 196108 2644
rect 196063 2604 196108 2632
rect 191045 2595 191103 2601
rect 196102 2592 196108 2604
rect 196160 2592 196166 2644
rect 196197 2635 196255 2641
rect 196197 2601 196209 2635
rect 196243 2632 196255 2635
rect 198497 2635 198555 2641
rect 198497 2632 198509 2635
rect 196243 2604 198509 2632
rect 196243 2601 196255 2604
rect 196197 2595 196255 2601
rect 198497 2601 198509 2604
rect 198543 2601 198555 2635
rect 198497 2595 198555 2601
rect 200245 2635 200303 2641
rect 200245 2601 200257 2635
rect 200291 2632 200303 2635
rect 200705 2635 200763 2641
rect 200705 2632 200717 2635
rect 200291 2604 200717 2632
rect 200291 2601 200303 2604
rect 200245 2595 200303 2601
rect 200705 2601 200717 2604
rect 200751 2601 200763 2635
rect 200705 2595 200763 2601
rect 209905 2635 209963 2641
rect 209905 2601 209917 2635
rect 209951 2632 209963 2635
rect 210365 2635 210423 2641
rect 210365 2632 210377 2635
rect 209951 2604 210377 2632
rect 209951 2601 209963 2604
rect 209905 2595 209963 2601
rect 210365 2601 210377 2604
rect 210411 2601 210423 2635
rect 210365 2595 210423 2601
rect 219749 2635 219807 2641
rect 219749 2601 219761 2635
rect 219795 2632 219807 2635
rect 220022 2632 220028 2644
rect 219795 2604 220028 2632
rect 219795 2601 219807 2604
rect 219749 2595 219807 2601
rect 220022 2592 220028 2604
rect 220080 2592 220086 2644
rect 223426 2592 223432 2644
rect 223484 2632 223490 2644
rect 229409 2635 229467 2641
rect 229409 2632 229421 2635
rect 223484 2604 229421 2632
rect 223484 2592 223490 2604
rect 229409 2601 229421 2604
rect 229455 2601 229467 2635
rect 229409 2595 229467 2601
rect 326193 2635 326251 2641
rect 326193 2601 326205 2635
rect 326239 2632 326251 2635
rect 346338 2632 346344 2644
rect 326239 2604 346344 2632
rect 326239 2601 326251 2604
rect 326193 2595 326251 2601
rect 346338 2592 346344 2604
rect 346396 2592 346402 2644
rect 355265 2635 355323 2641
rect 355265 2632 355277 2635
rect 347368 2604 355277 2632
rect 118730 2524 118736 2576
rect 118788 2564 118794 2576
rect 132901 2567 132959 2573
rect 132901 2564 132913 2567
rect 118788 2536 132913 2564
rect 118788 2524 118794 2536
rect 132901 2533 132913 2536
rect 132947 2533 132959 2567
rect 132901 2527 132959 2533
rect 133269 2567 133327 2573
rect 133269 2533 133281 2567
rect 133315 2564 133327 2567
rect 142561 2567 142619 2573
rect 142561 2564 142573 2567
rect 133315 2536 142573 2564
rect 133315 2533 133327 2536
rect 133269 2527 133327 2533
rect 142561 2533 142573 2536
rect 142607 2533 142619 2567
rect 142561 2527 142619 2533
rect 152313 2567 152371 2573
rect 152313 2533 152325 2567
rect 152359 2564 152371 2567
rect 161881 2567 161939 2573
rect 161881 2564 161893 2567
rect 152359 2536 161893 2564
rect 152359 2533 152371 2536
rect 152313 2527 152371 2533
rect 161881 2533 161893 2536
rect 161927 2533 161939 2567
rect 161881 2527 161939 2533
rect 190953 2567 191011 2573
rect 190953 2533 190965 2567
rect 190999 2564 191011 2567
rect 200521 2567 200579 2573
rect 200521 2564 200533 2567
rect 190999 2536 200533 2564
rect 190999 2533 191011 2536
rect 190953 2527 191011 2533
rect 200521 2533 200533 2536
rect 200567 2533 200579 2567
rect 200521 2527 200579 2533
rect 200613 2567 200671 2573
rect 200613 2533 200625 2567
rect 200659 2564 200671 2567
rect 210181 2567 210239 2573
rect 210181 2564 210193 2567
rect 200659 2536 210193 2564
rect 200659 2533 200671 2536
rect 200613 2527 200671 2533
rect 210181 2533 210193 2536
rect 210227 2533 210239 2567
rect 210181 2527 210239 2533
rect 219933 2567 219991 2573
rect 219933 2533 219945 2567
rect 219979 2564 219991 2567
rect 229685 2567 229743 2573
rect 229685 2564 229697 2567
rect 219979 2536 229697 2564
rect 219979 2533 219991 2536
rect 219933 2527 219991 2533
rect 229685 2533 229697 2536
rect 229731 2533 229743 2567
rect 229685 2527 229743 2533
rect 345605 2567 345663 2573
rect 345605 2533 345617 2567
rect 345651 2564 345663 2567
rect 347368 2564 347396 2604
rect 355265 2601 355277 2604
rect 355311 2601 355323 2635
rect 355265 2595 355323 2601
rect 358022 2592 358028 2644
rect 358080 2632 358086 2644
rect 359034 2632 359040 2644
rect 358080 2604 359040 2632
rect 358080 2592 358086 2604
rect 359034 2592 359040 2604
rect 359092 2592 359098 2644
rect 360690 2592 360696 2644
rect 360748 2632 360754 2644
rect 361426 2632 361432 2644
rect 360748 2604 361432 2632
rect 360748 2592 360754 2604
rect 361426 2592 361432 2604
rect 361484 2592 361490 2644
rect 362070 2592 362076 2644
rect 362128 2632 362134 2644
rect 362622 2632 362628 2644
rect 362128 2604 362628 2632
rect 362128 2592 362134 2604
rect 362622 2592 362628 2604
rect 362680 2592 362686 2644
rect 364649 2635 364707 2641
rect 364649 2601 364661 2635
rect 364695 2632 364707 2635
rect 364925 2635 364983 2641
rect 364925 2632 364937 2635
rect 364695 2604 364937 2632
rect 364695 2601 364707 2604
rect 364649 2595 364707 2601
rect 364925 2601 364937 2604
rect 364971 2601 364983 2635
rect 364925 2595 364983 2601
rect 374309 2635 374367 2641
rect 374309 2601 374321 2635
rect 374355 2632 374367 2635
rect 374585 2635 374643 2641
rect 374355 2604 374536 2632
rect 374355 2601 374367 2604
rect 374309 2595 374367 2601
rect 345651 2536 347396 2564
rect 350757 2567 350815 2573
rect 345651 2533 345663 2536
rect 345605 2527 345663 2533
rect 350757 2533 350769 2567
rect 350803 2564 350815 2567
rect 364741 2567 364799 2573
rect 364741 2564 364753 2567
rect 350803 2536 364753 2564
rect 350803 2533 350815 2536
rect 350757 2527 350815 2533
rect 364741 2533 364753 2536
rect 364787 2533 364799 2567
rect 374508 2564 374536 2604
rect 374585 2601 374597 2635
rect 374631 2632 374643 2635
rect 382862 2632 382868 2644
rect 374631 2604 382868 2632
rect 374631 2601 374643 2604
rect 374585 2595 374643 2601
rect 382862 2592 382868 2604
rect 382920 2592 382926 2644
rect 383969 2635 384027 2641
rect 383969 2601 383981 2635
rect 384015 2632 384027 2635
rect 390041 2635 390099 2641
rect 390041 2632 390053 2635
rect 384015 2604 390053 2632
rect 384015 2601 384027 2604
rect 383969 2595 384027 2601
rect 390041 2601 390053 2604
rect 390087 2601 390099 2635
rect 390041 2595 390099 2601
rect 384061 2567 384119 2573
rect 384061 2564 384073 2567
rect 374508 2536 384073 2564
rect 364741 2527 364799 2533
rect 384061 2533 384073 2536
rect 384107 2533 384119 2567
rect 384061 2527 384119 2533
rect 374677 2499 374735 2505
rect 374677 2465 374689 2499
rect 374723 2496 374735 2499
rect 380470 2496 380476 2508
rect 374723 2468 380476 2496
rect 374723 2465 374735 2468
rect 374677 2459 374735 2465
rect 380470 2456 380476 2468
rect 380528 2456 380534 2508
rect 349650 2388 349656 2440
rect 349708 2428 349714 2440
rect 350754 2428 350760 2440
rect 349708 2400 350760 2428
rect 349708 2388 349714 2400
rect 350754 2388 350760 2400
rect 350812 2388 350818 2440
rect 374769 2431 374827 2437
rect 374769 2397 374781 2431
rect 374815 2428 374827 2431
rect 384058 2428 384064 2440
rect 374815 2400 384064 2428
rect 374815 2397 374827 2400
rect 374769 2391 374827 2397
rect 384058 2388 384064 2400
rect 384116 2388 384122 2440
rect 1600 2128 583316 2224
rect 356550 1368 356556 1420
rect 356608 1408 356614 1420
rect 357838 1408 357844 1420
rect 356608 1380 357844 1408
rect 356608 1368 356614 1380
rect 357838 1368 357844 1380
rect 357896 1368 357902 1420
rect 353790 1096 353796 1148
rect 353848 1136 353854 1148
rect 354250 1136 354256 1148
rect 353848 1108 354256 1136
rect 353848 1096 353854 1108
rect 354250 1096 354256 1108
rect 354308 1096 354314 1148
rect 5754 552 5760 604
rect 5812 592 5818 604
rect 5938 592 5944 604
rect 5812 564 5944 592
rect 5812 552 5818 564
rect 5938 552 5944 564
rect 5996 552 6002 604
rect 23602 552 23608 604
rect 23660 592 23666 604
rect 23878 592 23884 604
rect 23660 564 23884 592
rect 23660 552 23666 564
rect 23878 552 23884 564
rect 23936 552 23942 604
rect 74754 552 74760 604
rect 74812 592 74818 604
rect 74938 592 74944 604
rect 74812 564 74944 592
rect 74812 552 74818 564
rect 74938 552 74944 564
rect 74996 552 75002 604
rect 152034 552 152040 604
rect 152092 592 152098 604
rect 152126 592 152132 604
rect 152092 564 152132 592
rect 152092 552 152098 564
rect 152126 552 152132 564
rect 152184 552 152190 604
rect 155622 552 155628 604
rect 155680 592 155686 604
rect 156358 592 156364 604
rect 155680 564 156364 592
rect 155680 552 155686 564
rect 156358 552 156364 564
rect 156416 552 156422 604
rect 169882 552 169888 604
rect 169940 592 169946 604
rect 169974 592 169980 604
rect 169940 564 169980 592
rect 169940 552 169946 564
rect 169974 552 169980 564
rect 170032 552 170038 604
rect 173470 552 173476 604
rect 173528 592 173534 604
rect 174298 592 174304 604
rect 173528 564 174304 592
rect 173528 552 173534 564
rect 174298 552 174304 564
rect 174356 552 174362 604
rect 180646 552 180652 604
rect 180704 592 180710 604
rect 181198 592 181204 604
rect 180704 564 181204 592
rect 180704 552 180710 564
rect 181198 552 181204 564
rect 181256 552 181262 604
rect 183038 552 183044 604
rect 183096 592 183102 604
rect 183958 592 183964 604
rect 183096 564 183964 592
rect 183096 552 183102 564
rect 183958 552 183964 564
rect 184016 552 184022 604
rect 190122 552 190128 604
rect 190180 592 190186 604
rect 190398 592 190404 604
rect 190180 564 190404 592
rect 190180 552 190186 564
rect 190398 552 190404 564
rect 190456 552 190462 604
rect 197298 552 197304 604
rect 197356 592 197362 604
rect 197758 592 197764 604
rect 197356 564 197764 592
rect 197356 552 197362 564
rect 197758 552 197764 564
rect 197816 552 197822 604
rect 200886 552 200892 604
rect 200944 592 200950 604
rect 201898 592 201904 604
rect 200944 564 201904 592
rect 200944 552 200950 564
rect 201898 552 201904 564
rect 201956 552 201962 604
rect 221034 552 221040 604
rect 221092 592 221098 604
rect 221218 592 221224 604
rect 221092 564 221224 592
rect 221092 552 221098 564
rect 221218 552 221224 564
rect 221276 552 221282 604
rect 231798 552 231804 604
rect 231856 592 231862 604
rect 231982 592 231988 604
rect 231856 564 231988 592
rect 231856 552 231862 564
rect 231982 552 231988 564
rect 232040 552 232046 604
rect 234190 552 234196 604
rect 234248 592 234254 604
rect 235205 595 235263 601
rect 235205 592 235217 595
rect 234248 564 235217 592
rect 234248 552 234254 564
rect 235205 561 235217 564
rect 235251 561 235263 595
rect 235205 555 235263 561
rect 248450 552 248456 604
rect 248508 592 248514 604
rect 248818 592 248824 604
rect 248508 564 248824 592
rect 248508 552 248514 564
rect 248818 552 248824 564
rect 248876 552 248882 604
rect 256730 552 256736 604
rect 256788 592 256794 604
rect 257098 592 257104 604
rect 256788 564 257104 592
rect 256788 552 256794 564
rect 257098 552 257104 564
rect 257156 552 257162 604
rect 290586 552 290592 604
rect 290644 592 290650 604
rect 291230 592 291236 604
rect 290644 564 291236 592
rect 290644 552 290650 564
rect 291230 552 291236 564
rect 291288 552 291294 604
rect 309078 592 309084 604
rect 309039 564 309084 592
rect 309078 552 309084 564
rect 309136 552 309142 604
rect 324810 552 324816 604
rect 324868 592 324874 604
rect 325730 592 325736 604
rect 324868 564 325736 592
rect 324868 552 324874 564
rect 325730 552 325736 564
rect 325788 552 325794 604
rect 378630 552 378636 604
rect 378688 592 378694 604
rect 379274 592 379280 604
rect 378688 564 379280 592
rect 378688 552 378694 564
rect 379274 552 379280 564
rect 379332 552 379338 604
rect 395190 552 395196 604
rect 395248 592 395254 604
rect 395926 592 395932 604
rect 395248 564 395932 592
rect 395248 552 395254 564
rect 395926 552 395932 564
rect 395984 552 395990 604
rect 402090 552 402096 604
rect 402148 592 402154 604
rect 403010 592 403016 604
rect 402148 564 403016 592
rect 402148 552 402154 564
rect 403010 552 403016 564
rect 403068 552 403074 604
rect 406230 552 406236 604
rect 406288 592 406294 604
rect 406598 592 406604 604
rect 406288 564 406604 592
rect 406288 552 406294 564
rect 406598 552 406604 564
rect 406656 552 406662 604
rect 420858 592 420864 604
rect 420819 564 420864 592
rect 420858 552 420864 564
rect 420916 552 420922 604
rect 424170 552 424176 604
rect 424228 592 424234 604
rect 424446 592 424452 604
rect 424228 564 424452 592
rect 424228 552 424234 564
rect 424446 552 424452 564
rect 424504 552 424510 604
rect 426930 552 426936 604
rect 426988 592 426994 604
rect 428034 592 428040 604
rect 426988 564 428040 592
rect 426988 552 426994 564
rect 428034 552 428040 564
rect 428092 552 428098 604
rect 431070 552 431076 604
rect 431128 592 431134 604
rect 431622 592 431628 604
rect 431128 564 431628 592
rect 431128 552 431134 564
rect 431622 552 431628 564
rect 431680 552 431686 604
rect 442110 552 442116 604
rect 442168 592 442174 604
rect 442294 592 442300 604
rect 442168 564 442300 592
rect 442168 552 442174 564
rect 442294 552 442300 564
rect 442352 552 442358 604
rect 443582 552 443588 604
rect 443640 592 443646 604
rect 444686 592 444692 604
rect 443640 564 444692 592
rect 443640 552 443646 564
rect 444686 552 444692 564
rect 444744 552 444750 604
rect 444870 552 444876 604
rect 444928 592 444934 604
rect 445882 592 445888 604
rect 444928 564 445888 592
rect 444928 552 444934 564
rect 445882 552 445888 564
rect 445940 552 445946 604
rect 447630 552 447636 604
rect 447688 592 447694 604
rect 448274 592 448280 604
rect 447688 564 448280 592
rect 447688 552 447694 564
rect 448274 552 448280 564
rect 448332 552 448338 604
rect 449010 552 449016 604
rect 449068 592 449074 604
rect 449470 592 449476 604
rect 449068 564 449476 592
rect 449068 552 449074 564
rect 449470 552 449476 564
rect 449528 552 449534 604
rect 451862 552 451868 604
rect 451920 592 451926 604
rect 452966 592 452972 604
rect 451920 564 452972 592
rect 451920 552 451926 564
rect 452966 552 452972 564
rect 453024 552 453030 604
rect 454530 552 454536 604
rect 454588 592 454594 604
rect 455358 592 455364 604
rect 454588 564 455364 592
rect 454588 552 454594 564
rect 455358 552 455364 564
rect 455416 552 455422 604
rect 461430 552 461436 604
rect 461488 592 461494 604
rect 462534 592 462540 604
rect 461488 564 462540 592
rect 461488 552 461494 564
rect 462534 552 462540 564
rect 462592 552 462598 604
rect 462810 552 462816 604
rect 462868 592 462874 604
rect 463730 592 463736 604
rect 462868 564 463736 592
rect 462868 552 462874 564
rect 463730 552 463736 564
rect 463788 552 463794 604
rect 465570 552 465576 604
rect 465628 592 465634 604
rect 466122 592 466128 604
rect 465628 564 466128 592
rect 465628 552 465634 564
rect 466122 552 466128 564
rect 466180 552 466186 604
rect 466950 552 466956 604
rect 467008 592 467014 604
rect 467318 592 467324 604
rect 467008 564 467324 592
rect 467008 552 467014 564
rect 467318 552 467324 564
rect 467376 552 467382 604
rect 469710 552 469716 604
rect 469768 592 469774 604
rect 470814 592 470820 604
rect 469768 564 470820 592
rect 469768 552 469774 564
rect 470814 552 470820 564
rect 470872 552 470878 604
rect 490410 552 490416 604
rect 490468 592 490474 604
rect 491054 592 491060 604
rect 490468 564 491060 592
rect 490468 552 490474 564
rect 491054 552 491060 564
rect 491112 552 491118 604
rect 495930 552 495936 604
rect 495988 592 495994 604
rect 497034 592 497040 604
rect 495988 564 497040 592
rect 495988 552 495994 564
rect 497034 552 497040 564
rect 497092 552 497098 604
rect 497310 552 497316 604
rect 497368 592 497374 604
rect 498230 592 498236 604
rect 497368 564 498236 592
rect 497368 552 497374 564
rect 498230 552 498236 564
rect 498288 552 498294 604
rect 500070 552 500076 604
rect 500128 592 500134 604
rect 500622 592 500628 604
rect 500128 564 500628 592
rect 500128 552 500134 564
rect 500622 552 500628 564
rect 500680 552 500686 604
rect 501450 552 501456 604
rect 501508 592 501514 604
rect 501726 592 501732 604
rect 501508 564 501732 592
rect 501508 552 501514 564
rect 501726 552 501732 564
rect 501784 552 501790 604
rect 504210 552 504216 604
rect 504268 592 504274 604
rect 505314 592 505320 604
rect 504268 564 505320 592
rect 504268 552 504274 564
rect 505314 552 505320 564
rect 505372 552 505378 604
rect 506970 552 506976 604
rect 507028 592 507034 604
rect 507706 592 507712 604
rect 507028 564 507712 592
rect 507028 552 507034 564
rect 507706 552 507712 564
rect 507764 552 507770 604
rect 508350 552 508356 604
rect 508408 592 508414 604
rect 508902 592 508908 604
rect 508408 564 508908 592
rect 508408 552 508414 564
rect 508902 552 508908 564
rect 508960 552 508966 604
rect 529142 552 529148 604
rect 529200 592 529206 604
rect 529234 592 529240 604
rect 529200 564 529240 592
rect 529200 552 529206 564
rect 529234 552 529240 564
rect 529292 552 529298 604
<< via1 >>
rect 119380 700952 119432 701004
rect 249192 700884 249244 700936
rect 250204 700884 250256 700936
rect 284704 700884 284756 700936
rect 299976 700952 300028 701004
rect 184240 700816 184292 700868
rect 185344 700816 185396 700868
rect 286084 700816 286136 700868
rect 288844 700816 288896 700868
rect 465484 700884 465536 700936
rect 487104 700816 487156 700868
rect 97760 700748 97812 700800
rect 301356 700748 301408 700800
rect 76140 700544 76192 700596
rect 301448 700544 301500 700596
rect 54520 700476 54572 700528
rect 302736 700476 302788 700528
rect 280564 700408 280616 700460
rect 530344 700408 530396 700460
rect 280472 700340 280524 700392
rect 551964 700340 552016 700392
rect 32900 700272 32952 700324
rect 305496 700272 305548 700324
rect 141000 700204 141052 700256
rect 298596 700204 298648 700256
rect 162620 700000 162672 700052
rect 270812 699932 270864 699984
rect 287464 699932 287516 699984
rect 422244 699932 422296 699984
rect 283324 699864 283376 699916
rect 205952 699796 206004 699848
rect 294456 699864 294508 699916
rect 400624 699864 400676 699916
rect 290224 699796 290276 699848
rect 292524 699796 292576 699848
rect 227572 699728 227624 699780
rect 291788 699728 291840 699780
rect 295928 699728 295980 699780
rect 335672 699796 335724 699848
rect 297216 699728 297268 699780
rect 291696 699660 291748 699712
rect 292432 699660 292484 699712
rect 292524 699660 292576 699712
rect 357292 699660 357344 699712
rect 276424 695512 276476 695564
rect 580116 695512 580168 695564
rect 378728 695487 378780 695496
rect 378728 695453 378737 695487
rect 378737 695453 378771 695487
rect 378771 695453 378780 695487
rect 378728 695444 378780 695453
rect 508448 695487 508500 695496
rect 508448 695453 508457 695487
rect 508457 695453 508491 695487
rect 508491 695453 508500 695487
rect 508448 695444 508500 695453
rect 3736 694220 3788 694272
rect 305588 694220 305640 694272
rect 314052 688576 314104 688628
rect 314236 688576 314288 688628
rect 443772 688576 443824 688628
rect 443956 688576 444008 688628
rect 573492 688576 573544 688628
rect 573676 688576 573728 688628
rect 378820 685856 378872 685908
rect 508540 685856 508592 685908
rect 277804 680348 277856 680400
rect 580116 680348 580168 680400
rect 3920 677560 3972 677612
rect 308256 677560 308308 677612
rect 314144 676107 314196 676116
rect 314144 676073 314153 676107
rect 314153 676073 314187 676107
rect 314187 676073 314196 676107
rect 314144 676064 314196 676073
rect 378636 676107 378688 676116
rect 378636 676073 378645 676107
rect 378645 676073 378679 676107
rect 378679 676073 378688 676107
rect 378636 676064 378688 676073
rect 443864 676107 443916 676116
rect 443864 676073 443873 676107
rect 443873 676073 443907 676107
rect 443907 676073 443916 676107
rect 443864 676064 443916 676073
rect 508356 676107 508408 676116
rect 508356 676073 508365 676107
rect 508365 676073 508399 676107
rect 508399 676073 508408 676107
rect 508356 676064 508408 676073
rect 573584 676107 573636 676116
rect 573584 676073 573593 676107
rect 573593 676073 573627 676107
rect 573627 676073 573636 676107
rect 573584 676064 573636 676073
rect 314236 666544 314288 666596
rect 378728 666544 378780 666596
rect 443956 666544 444008 666596
rect 508448 666544 508500 666596
rect 573676 666544 573728 666596
rect 275044 663756 275096 663808
rect 580116 663756 580168 663808
rect 3920 661036 3972 661088
rect 306876 661036 306928 661088
rect 378728 659676 378780 659728
rect 378820 659676 378872 659728
rect 508448 659676 508500 659728
rect 508540 659676 508592 659728
rect 378636 654100 378688 654152
rect 378820 654100 378872 654152
rect 508356 654100 508408 654152
rect 508540 654100 508592 654152
rect 273664 648592 273716 648644
rect 580116 648592 580168 648644
rect 313960 647232 314012 647284
rect 314052 647232 314104 647284
rect 443680 647232 443732 647284
rect 443772 647232 443824 647284
rect 573400 647232 573452 647284
rect 573492 647232 573544 647284
rect 3552 644444 3604 644496
rect 309636 644444 309688 644496
rect 314144 637483 314196 637492
rect 314144 637449 314153 637483
rect 314153 637449 314187 637483
rect 314187 637449 314196 637483
rect 314144 637440 314196 637449
rect 443864 637483 443916 637492
rect 443864 637449 443873 637483
rect 443873 637449 443907 637483
rect 443907 637449 443916 637483
rect 443864 637440 443916 637449
rect 573584 637483 573636 637492
rect 573584 637449 573593 637483
rect 573593 637449 573627 637483
rect 573627 637449 573636 637483
rect 573584 637440 573636 637449
rect 274952 633428 275004 633480
rect 580116 633428 580168 633480
rect 3920 627920 3972 627972
rect 311016 627920 311068 627972
rect 314236 627920 314288 627972
rect 443956 627920 444008 627972
rect 573676 627920 573728 627972
rect 314052 618264 314104 618316
rect 314236 618264 314288 618316
rect 443772 618264 443824 618316
rect 443956 618264 444008 618316
rect 573492 618264 573544 618316
rect 573676 618264 573728 618316
rect 573492 618128 573544 618180
rect 573768 618128 573820 618180
rect 272284 616972 272336 617024
rect 580116 616972 580168 617024
rect 378636 615476 378688 615528
rect 378820 615476 378872 615528
rect 508356 615476 508408 615528
rect 508540 615476 508592 615528
rect 3828 611328 3880 611380
rect 309728 611328 309780 611380
rect 313776 608608 313828 608660
rect 313960 608608 314012 608660
rect 443680 608583 443732 608592
rect 443680 608549 443689 608583
rect 443689 608549 443723 608583
rect 443723 608549 443732 608583
rect 443680 608540 443732 608549
rect 573400 608583 573452 608592
rect 573400 608549 573409 608583
rect 573409 608549 573443 608583
rect 573443 608549 573452 608583
rect 573400 608540 573452 608549
rect 270904 601740 270956 601792
rect 580116 601740 580168 601792
rect 443864 601536 443916 601588
rect 573584 601536 573636 601588
rect 313868 598859 313920 598868
rect 313868 598825 313877 598859
rect 313877 598825 313911 598859
rect 313911 598825 313920 598859
rect 313868 598816 313920 598825
rect 443864 598859 443916 598868
rect 443864 598825 443873 598859
rect 443873 598825 443907 598859
rect 443907 598825 443916 598859
rect 443864 598816 443916 598825
rect 573584 598859 573636 598868
rect 573584 598825 573593 598859
rect 573593 598825 573627 598859
rect 573627 598825 573636 598859
rect 573584 598816 573636 598825
rect 3920 594804 3972 594856
rect 312396 594804 312448 594856
rect 314052 589296 314104 589348
rect 443956 589296 444008 589348
rect 573676 589296 573728 589348
rect 378728 589228 378780 589280
rect 508448 589228 508500 589280
rect 270812 586508 270864 586560
rect 580116 586508 580168 586560
rect 314052 582360 314104 582412
rect 443956 582428 444008 582480
rect 573676 582428 573728 582480
rect 314144 582292 314196 582344
rect 443864 582292 443916 582344
rect 573584 582292 573636 582344
rect 378636 579683 378688 579692
rect 378636 579649 378645 579683
rect 378645 579649 378679 579683
rect 378679 579649 378688 579683
rect 378636 579640 378688 579649
rect 508356 579683 508408 579692
rect 508356 579649 508365 579683
rect 508365 579649 508399 579683
rect 508399 579649 508408 579683
rect 508356 579640 508408 579649
rect 314144 579572 314196 579624
rect 3736 576852 3788 576904
rect 313868 576852 313920 576904
rect 313960 570027 314012 570036
rect 313960 569993 313969 570027
rect 313969 569993 314003 570027
rect 314003 569993 314012 570027
rect 313960 569984 314012 569993
rect 269524 569916 269576 569968
rect 580116 569916 580168 569968
rect 378728 569891 378780 569900
rect 378728 569857 378737 569891
rect 378737 569857 378771 569891
rect 378771 569857 378780 569891
rect 378728 569848 378780 569857
rect 508448 569891 508500 569900
rect 508448 569857 508457 569891
rect 508457 569857 508491 569891
rect 508491 569857 508500 569891
rect 508448 569848 508500 569857
rect 378912 562912 378964 562964
rect 508632 562912 508684 562964
rect 3920 560396 3972 560448
rect 313960 560396 314012 560448
rect 266764 554752 266816 554804
rect 580116 554752 580168 554804
rect 443496 553435 443548 553444
rect 443496 553401 443505 553435
rect 443505 553401 443539 553435
rect 443539 553401 443548 553435
rect 443496 553392 443548 553401
rect 573216 553435 573268 553444
rect 573216 553401 573225 553435
rect 573225 553401 573259 553435
rect 573259 553401 573268 553435
rect 573216 553392 573268 553401
rect 313776 552576 313828 552628
rect 314052 552576 314104 552628
rect 378728 550604 378780 550656
rect 379004 550604 379056 550656
rect 443496 550647 443548 550656
rect 443496 550613 443505 550647
rect 443505 550613 443539 550647
rect 443539 550613 443548 550647
rect 443496 550604 443548 550613
rect 508448 550604 508500 550656
rect 508724 550604 508776 550656
rect 573216 550647 573268 550656
rect 573216 550613 573225 550647
rect 573225 550613 573259 550647
rect 573259 550613 573268 550647
rect 573216 550604 573268 550613
rect 3644 543736 3696 543788
rect 315156 543736 315208 543788
rect 379004 543804 379056 543856
rect 443496 543736 443548 543788
rect 378912 543668 378964 543720
rect 508724 543804 508776 543856
rect 573216 543736 573268 543788
rect 508632 543668 508684 543720
rect 443588 543600 443640 543652
rect 573308 543600 573360 543652
rect 268144 539724 268196 539776
rect 580116 539724 580168 539776
rect 313776 538228 313828 538280
rect 314052 538228 314104 538280
rect 378912 534080 378964 534132
rect 443496 534123 443548 534132
rect 443496 534089 443505 534123
rect 443505 534089 443539 534123
rect 443539 534089 443548 534123
rect 443496 534080 443548 534089
rect 508632 534080 508684 534132
rect 573216 534123 573268 534132
rect 573216 534089 573225 534123
rect 573225 534089 573259 534123
rect 573259 534089 573268 534123
rect 573216 534080 573268 534089
rect 379004 533944 379056 533996
rect 508724 533944 508776 533996
rect 443496 531335 443548 531344
rect 443496 531301 443505 531335
rect 443505 531301 443539 531335
rect 443539 531301 443548 531335
rect 443496 531292 443548 531301
rect 573216 531335 573268 531344
rect 573216 531301 573225 531335
rect 573225 531301 573259 531335
rect 573259 531301 573268 531335
rect 573216 531292 573268 531301
rect 443588 531267 443640 531276
rect 443588 531233 443597 531267
rect 443597 531233 443631 531267
rect 443631 531233 443640 531267
rect 443588 531224 443640 531233
rect 573308 531267 573360 531276
rect 573308 531233 573317 531267
rect 573317 531233 573351 531267
rect 573351 531233 573360 531267
rect 573308 531224 573360 531233
rect 313776 528504 313828 528556
rect 314052 528504 314104 528556
rect 3644 527212 3696 527264
rect 317916 527212 317968 527264
rect 443588 524331 443640 524340
rect 443588 524297 443597 524331
rect 443597 524297 443631 524331
rect 443631 524297 443640 524331
rect 443588 524288 443640 524297
rect 573308 524331 573360 524340
rect 573308 524297 573317 524331
rect 573317 524297 573351 524331
rect 573351 524297 573360 524331
rect 573308 524288 573360 524297
rect 266672 522996 266724 523048
rect 580116 522996 580168 523048
rect 379004 514496 379056 514548
rect 379188 514496 379240 514548
rect 508724 514496 508776 514548
rect 508908 514496 508960 514548
rect 313776 513952 313828 514004
rect 314052 513952 314104 514004
rect 4012 510620 4064 510672
rect 316536 510620 316588 510672
rect 264004 507832 264056 507884
rect 580116 507832 580168 507884
rect 378820 502324 378872 502376
rect 379004 502324 379056 502376
rect 443496 502324 443548 502376
rect 443772 502324 443824 502376
rect 508540 502324 508592 502376
rect 508724 502324 508776 502376
rect 573216 502324 573268 502376
rect 573492 502324 573544 502376
rect 313776 499536 313828 499588
rect 314052 499536 314104 499588
rect 3736 494028 3788 494080
rect 318008 494028 318060 494080
rect 265384 492668 265436 492720
rect 580116 492668 580168 492720
rect 313776 489812 313828 489864
rect 314052 489812 314104 489864
rect 443772 485868 443824 485920
rect 573492 485868 573544 485920
rect 443496 485707 443548 485716
rect 443496 485673 443505 485707
rect 443505 485673 443539 485707
rect 443539 485673 443548 485707
rect 443496 485664 443548 485673
rect 573216 485707 573268 485716
rect 573216 485673 573225 485707
rect 573225 485673 573259 485707
rect 573259 485673 573268 485707
rect 573216 485664 573268 485673
rect 313776 480224 313828 480276
rect 314052 480224 314104 480276
rect 378636 480224 378688 480276
rect 378820 480224 378872 480276
rect 508356 480224 508408 480276
rect 508540 480224 508592 480276
rect 3920 477504 3972 477556
rect 320676 477504 320728 477556
rect 262624 476076 262676 476128
rect 580116 476076 580168 476128
rect 313776 475328 313828 475380
rect 314052 475328 314104 475380
rect 443588 471971 443640 471980
rect 443588 471937 443597 471971
rect 443597 471937 443631 471971
rect 443631 471937 443640 471971
rect 443588 471928 443640 471937
rect 573308 471971 573360 471980
rect 573308 471937 573317 471971
rect 573317 471937 573351 471971
rect 573351 471937 573360 471971
rect 573308 471928 573360 471937
rect 314052 463700 314104 463752
rect 359960 463632 360012 463684
rect 257104 463564 257156 463616
rect 355912 463564 355964 463616
rect 258208 463360 258260 463412
rect 358672 463360 358724 463412
rect 253976 463292 254028 463344
rect 354532 463292 354584 463344
rect 185344 463224 185396 463276
rect 283600 463224 283652 463276
rect 250204 463156 250256 463208
rect 293076 463224 293128 463276
rect 293168 463224 293220 463276
rect 378820 463224 378872 463276
rect 261336 463088 261388 463140
rect 278172 463088 278224 463140
rect 282312 463088 282364 463140
rect 282404 463088 282456 463140
rect 283324 463088 283376 463140
rect 283416 463088 283468 463140
rect 264556 463020 264608 463072
rect 265384 463020 265436 463072
rect 265568 463020 265620 463072
rect 266672 463020 266724 463072
rect 268696 463020 268748 463072
rect 269524 463020 269576 463072
rect 269800 463020 269852 463072
rect 270904 463020 270956 463072
rect 272928 463020 272980 463072
rect 273664 463020 273716 463072
rect 273940 463020 273992 463072
rect 274952 463020 275004 463072
rect 279276 463020 279328 463072
rect 280564 463020 280616 463072
rect 281392 463020 281444 463072
rect 283784 463020 283836 463072
rect 284704 463020 284756 463072
rect 286636 463020 286688 463072
rect 287464 463020 287516 463072
rect 288200 463088 288252 463140
rect 291696 463088 291748 463140
rect 292524 463088 292576 463140
rect 301356 463088 301408 463140
rect 302092 463088 302144 463140
rect 508540 463088 508592 463140
rect 255080 462816 255132 462868
rect 357200 462816 357252 462868
rect 4380 462748 4432 462800
rect 330796 462748 330848 462800
rect 4288 462680 4340 462732
rect 333924 462680 333976 462732
rect 4196 462612 4248 462664
rect 337144 462612 337196 462664
rect 4012 462544 4064 462596
rect 339260 462544 339312 462596
rect 4104 462476 4156 462528
rect 340272 462476 340324 462528
rect 291144 462272 291196 462324
rect 313868 462272 313920 462324
rect 314788 462272 314840 462324
rect 284704 462204 284756 462256
rect 296756 462136 296808 462188
rect 228952 461524 229004 461576
rect 328680 461524 328732 461576
rect 220580 461456 220632 461508
rect 324540 461456 324592 461508
rect 240268 461388 240320 461440
rect 351680 461388 351732 461440
rect 235024 461184 235076 461236
rect 361340 461184 361392 461236
rect 259220 461116 259272 461168
rect 411020 461116 411072 461168
rect 179180 461048 179232 461100
rect 332912 461048 332964 461100
rect 6772 460980 6824 461032
rect 322424 460980 322476 461032
rect 260324 460912 260376 460964
rect 580668 460912 580720 460964
rect 228860 460300 228912 460352
rect 335028 460300 335080 460352
rect 243488 460096 243540 460148
rect 353060 460096 353112 460148
rect 3644 459756 3696 459808
rect 227572 460028 227624 460080
rect 325276 460028 325328 460080
rect 223340 459960 223392 460012
rect 326380 459960 326432 460012
rect 252780 459892 252832 459944
rect 355820 459892 355872 459944
rect 248088 459824 248140 459876
rect 358580 459824 358632 459876
rect 224720 459756 224772 459808
rect 335856 459756 335908 459808
rect 234288 459663 234340 459672
rect 234288 459629 234297 459663
rect 234297 459629 234331 459663
rect 234331 459629 234340 459663
rect 234288 459620 234340 459629
rect 250112 459663 250164 459672
rect 250112 459629 250121 459663
rect 250121 459629 250155 459663
rect 250155 459629 250164 459663
rect 250112 459620 250164 459629
rect 256368 459663 256420 459672
rect 256368 459629 256377 459663
rect 256377 459629 256411 459663
rect 256411 459629 256420 459663
rect 256368 459620 256420 459629
rect 319940 459688 319992 459740
rect 323528 459663 323580 459672
rect 323528 459629 323537 459663
rect 323537 459629 323571 459663
rect 323571 459629 323580 459663
rect 323528 459620 323580 459629
rect 327484 459663 327536 459672
rect 327484 459629 327493 459663
rect 327493 459629 327527 459663
rect 327527 459629 327536 459663
rect 327484 459620 327536 459629
rect 329508 459663 329560 459672
rect 329508 459629 329517 459663
rect 329517 459629 329551 459663
rect 329551 459629 329560 459663
rect 329508 459620 329560 459629
rect 331716 459663 331768 459672
rect 331716 459629 331725 459663
rect 331725 459629 331759 459663
rect 331759 459629 331768 459663
rect 331716 459620 331768 459629
rect 337788 459663 337840 459672
rect 337788 459629 337797 459663
rect 337797 459629 337831 459663
rect 337831 459629 337840 459663
rect 337788 459620 337840 459629
rect 341192 459620 341244 459672
rect 345608 459663 345660 459672
rect 345608 459629 345617 459663
rect 345617 459629 345651 459663
rect 345651 459629 345660 459663
rect 345608 459620 345660 459629
rect 227480 458940 227532 458992
rect 354440 458872 354492 458924
rect 226192 458804 226244 458856
rect 226100 458736 226152 458788
rect 221960 458668 222012 458720
rect 219200 458464 219252 458516
rect 406880 458396 406932 458448
rect 6680 458328 6732 458380
rect 9440 458260 9492 458312
rect 580760 458192 580812 458244
rect 359960 447040 360012 447092
rect 580668 447040 580720 447092
rect 3644 444116 3696 444168
rect 6772 444116 6824 444168
rect 411020 430516 411072 430568
rect 580668 430516 580720 430568
rect 3644 427728 3696 427780
rect 220580 427728 220632 427780
rect 355912 415352 355964 415404
rect 580668 415352 580720 415404
rect 3828 411136 3880 411188
rect 226192 411136 226244 411188
rect 358672 400120 358724 400172
rect 580668 400120 580720 400172
rect 3828 394612 3880 394664
rect 227572 394612 227624 394664
rect 406880 383596 406932 383648
rect 580668 383596 580720 383648
rect 3552 377952 3604 378004
rect 221960 377952 222012 378004
rect 354532 368432 354584 368484
rect 580668 368432 580720 368484
rect 3828 361496 3880 361548
rect 223340 361496 223392 361548
rect 357200 353200 357252 353252
rect 580668 353200 580720 353252
rect 3828 343544 3880 343596
rect 228952 343544 229004 343596
rect 240912 339056 240964 339108
rect 241280 339056 241332 339108
rect 242108 339056 242160 339108
rect 242476 339056 242528 339108
rect 268236 339056 268288 339108
rect 268696 339056 268748 339108
rect 254804 338512 254856 338564
rect 255172 338512 255224 338564
rect 272652 338444 272704 338496
rect 273112 338444 273164 338496
rect 278908 338444 278960 338496
rect 279184 338444 279236 338496
rect 234196 338172 234248 338224
rect 129224 338104 129276 338156
rect 142564 338104 142616 338156
rect 152224 338104 152276 338156
rect 161884 338104 161936 338156
rect 171544 338104 171596 338156
rect 181204 338104 181256 338156
rect 190864 338104 190916 338156
rect 200524 338104 200576 338156
rect 210184 338104 210236 338156
rect 219844 338104 219896 338156
rect 232356 338104 232408 338156
rect 308900 338104 308952 338156
rect 309544 338104 309596 338156
rect 62524 338036 62576 338088
rect 242936 338036 242988 338088
rect 259220 338036 259272 338088
rect 283876 338036 283928 338088
rect 303932 338036 303984 338088
rect 356556 338036 356608 338088
rect 45964 337968 46016 338020
rect 55624 337968 55676 338020
rect 236312 337968 236364 338020
rect 44584 337900 44636 337952
rect 142564 337900 142616 337952
rect 152224 337900 152276 337952
rect 161884 337900 161936 337952
rect 171544 337900 171596 337952
rect 181204 337900 181256 337952
rect 190864 337900 190916 337952
rect 200524 337900 200576 337952
rect 210184 337900 210236 337952
rect 219844 337900 219896 337952
rect 237784 337900 237836 337952
rect 292616 337968 292668 338020
rect 293812 337968 293864 338020
rect 297308 337968 297360 338020
rect 304760 337968 304812 338020
rect 305404 337968 305456 338020
rect 364836 337968 364888 338020
rect 298228 337900 298280 337952
rect 298504 337900 298556 337952
rect 300252 337900 300304 337952
rect 303472 337900 303524 337952
rect 304944 337900 304996 337952
rect 305128 337900 305180 337952
rect 309084 337900 309136 337952
rect 309544 337900 309596 337952
rect 22504 337696 22556 337748
rect 37684 337696 37736 337748
rect 30784 337628 30836 337680
rect 45964 337560 46016 337612
rect 65284 337560 65336 337612
rect 84604 337560 84656 337612
rect 126004 337560 126056 337612
rect 12844 337492 12896 337544
rect 116344 337492 116396 337544
rect 128580 337492 128632 337544
rect 128764 337560 128816 337612
rect 129040 337560 129092 337612
rect 138332 337628 138384 337680
rect 138424 337628 138476 337680
rect 232632 337696 232684 337748
rect 232816 337696 232868 337748
rect 234656 337696 234708 337748
rect 241464 337696 241516 337748
rect 264740 337696 264792 337748
rect 280656 337696 280708 337748
rect 284060 337696 284112 337748
rect 293352 337696 293404 337748
rect 294180 337696 294232 337748
rect 294824 337696 294876 337748
rect 295744 337696 295796 337748
rect 296296 337696 296348 337748
rect 296756 337696 296808 337748
rect 296848 337696 296900 337748
rect 297032 337696 297084 337748
rect 297584 337696 297636 337748
rect 298320 337696 298372 337748
rect 298780 337696 298832 337748
rect 299516 337696 299568 337748
rect 300712 337696 300764 337748
rect 301172 337696 301224 337748
rect 302184 337696 302236 337748
rect 302460 337696 302512 337748
rect 302920 337696 302972 337748
rect 303932 337696 303984 337748
rect 304668 337696 304720 337748
rect 305220 337696 305272 337748
rect 306416 337696 306468 337748
rect 306600 337696 306652 337748
rect 307336 337696 307388 337748
rect 307980 337696 308032 337748
rect 310004 337696 310056 337748
rect 310832 337696 310884 337748
rect 312028 337696 312080 337748
rect 312304 337696 312356 337748
rect 378636 337696 378688 337748
rect 230056 337628 230108 337680
rect 292892 337628 292944 337680
rect 293720 337628 293772 337680
rect 293904 337628 293956 337680
rect 295192 337628 295244 337680
rect 295376 337628 295428 337680
rect 295560 337628 295612 337680
rect 296572 337628 296624 337680
rect 142472 337560 142524 337612
rect 142656 337560 142708 337612
rect 142748 337560 142800 337612
rect 152132 337560 152184 337612
rect 152224 337560 152276 337612
rect 152408 337560 152460 337612
rect 161792 337560 161844 337612
rect 161976 337560 162028 337612
rect 162068 337560 162120 337612
rect 171452 337560 171504 337612
rect 171544 337560 171596 337612
rect 171728 337560 171780 337612
rect 181112 337560 181164 337612
rect 181296 337560 181348 337612
rect 181388 337560 181440 337612
rect 190772 337560 190824 337612
rect 190864 337560 190916 337612
rect 191048 337560 191100 337612
rect 200432 337560 200484 337612
rect 200616 337560 200668 337612
rect 200708 337560 200760 337612
rect 210092 337560 210144 337612
rect 210184 337560 210236 337612
rect 210368 337560 210420 337612
rect 219752 337560 219804 337612
rect 219936 337560 219988 337612
rect 220028 337560 220080 337612
rect 239256 337560 239308 337612
rect 251584 337560 251636 337612
rect 281852 337560 281904 337612
rect 293628 337560 293680 337612
rect 294364 337560 294416 337612
rect 296112 337560 296164 337612
rect 297032 337560 297084 337612
rect 297768 337560 297820 337612
rect 298412 337560 298464 337612
rect 128856 337492 128908 337544
rect 129132 337492 129184 337544
rect 253976 337492 254028 337544
rect 254344 337492 254396 337544
rect 282588 337492 282640 337544
rect 295836 337492 295888 337544
rect 297124 337492 297176 337544
rect 299240 337628 299292 337680
rect 299884 337628 299936 337680
rect 299976 337628 300028 337680
rect 301264 337628 301316 337680
rect 302000 337628 302052 337680
rect 302552 337628 302604 337680
rect 304392 337628 304444 337680
rect 305312 337628 305364 337680
rect 305864 337628 305916 337680
rect 306692 337628 306744 337680
rect 310280 337628 310332 337680
rect 310648 337628 310700 337680
rect 311476 337628 311528 337680
rect 312120 337628 312172 337680
rect 385536 337628 385588 337680
rect 299056 337560 299108 337612
rect 299792 337560 299844 337612
rect 301448 337560 301500 337612
rect 302644 337560 302696 337612
rect 306140 337560 306192 337612
rect 306600 337560 306652 337612
rect 311016 337560 311068 337612
rect 312028 337560 312080 337612
rect 392436 337560 392488 337612
rect 303380 337492 303432 337544
rect 306876 337492 306928 337544
rect 21124 337424 21176 337476
rect 142380 337424 142432 337476
rect 152500 337424 152552 337476
rect 161700 337424 161752 337476
rect 171820 337424 171872 337476
rect 181020 337424 181072 337476
rect 191140 337424 191192 337476
rect 200340 337424 200392 337476
rect 210460 337424 210512 337476
rect 219660 337424 219712 337476
rect 11464 337356 11516 337408
rect 26644 337356 26696 337408
rect 36396 337356 36448 337408
rect 45964 337356 46016 337408
rect 55716 337356 55768 337408
rect 65284 337356 65336 337408
rect 75036 337356 75088 337408
rect 84604 337356 84656 337408
rect 94356 337356 94408 337408
rect 103924 337356 103976 337408
rect 123888 337356 123940 337408
rect 138332 337356 138384 337408
rect 142564 337356 142616 337408
rect 152316 337356 152368 337408
rect 161884 337356 161936 337408
rect 171636 337356 171688 337408
rect 181204 337356 181256 337408
rect 190956 337356 191008 337408
rect 200524 337356 200576 337408
rect 210276 337356 210328 337408
rect 219844 337356 219896 337408
rect 226928 337424 226980 337476
rect 230056 337424 230108 337476
rect 256184 337424 256236 337476
rect 257104 337424 257156 337476
rect 283140 337424 283192 337476
rect 294640 337424 294692 337476
rect 310280 337424 310332 337476
rect 310556 337492 310608 337544
rect 310924 337492 310976 337544
rect 311292 337492 311344 337544
rect 314236 337492 314288 337544
rect 400716 337492 400768 337544
rect 407616 337424 407668 337476
rect 252504 337356 252556 337408
rect 254252 337356 254304 337408
rect 282404 337356 282456 337408
rect 295100 337356 295152 337408
rect 308532 337356 308584 337408
rect 309360 337356 309412 337408
rect 312764 337356 312816 337408
rect 313684 337356 313736 337408
rect 315708 337356 315760 337408
rect 414516 337356 414568 337408
rect 26644 337152 26696 337204
rect 65192 337152 65244 337204
rect 69424 337152 69476 337204
rect 244408 337152 244460 337204
rect 251032 337152 251084 337204
rect 280104 337152 280156 337204
rect 287280 337152 287332 337204
rect 293168 337152 293220 337204
rect 295100 337152 295152 337204
rect 301724 337152 301776 337204
rect 313040 337152 313092 337204
rect 313684 337152 313736 337204
rect 342388 337152 342440 337204
rect 342664 337152 342716 337204
rect 342848 337152 342900 337204
rect 343768 337152 343820 337204
rect 344596 337152 344648 337204
rect 345424 337152 345476 337204
rect 346252 337152 346304 337204
rect 346528 337152 346580 337204
rect 347540 337152 347592 337204
rect 348184 337152 348236 337204
rect 348276 337152 348328 337204
rect 349196 337152 349248 337204
rect 349288 337152 349340 337204
rect 349472 337152 349524 337204
rect 349932 337152 349984 337204
rect 350944 337152 350996 337204
rect 76324 337084 76376 337136
rect 245880 337084 245932 337136
rect 278540 337084 278592 337136
rect 286544 337084 286596 337136
rect 291420 337084 291472 337136
rect 293904 337084 293956 337136
rect 314144 337084 314196 337136
rect 341376 337084 341428 337136
rect 342480 337084 342532 337136
rect 344320 337084 344372 337136
rect 345056 337084 345108 337136
rect 346068 337084 346120 337136
rect 346804 337084 346856 337136
rect 346988 337084 347040 337136
rect 348000 337084 348052 337136
rect 348736 337084 348788 337136
rect 351772 337084 351824 337136
rect 36396 337016 36448 337068
rect 45964 337016 46016 337068
rect 55716 337016 55768 337068
rect 65284 337016 65336 337068
rect 83224 337016 83276 337068
rect 247352 337016 247404 337068
rect 261244 337016 261296 337068
rect 283508 337016 283560 337068
rect 284152 337016 284204 337068
rect 291144 337016 291196 337068
rect 292248 337016 292300 337068
rect 300528 337016 300580 337068
rect 300988 337016 301040 337068
rect 309820 337016 309872 337068
rect 318376 337016 318428 337068
rect 318836 337016 318888 337068
rect 321044 337016 321096 337068
rect 321596 337016 321648 337068
rect 326656 337016 326708 337068
rect 327392 337016 327444 337068
rect 332084 337016 332136 337068
rect 332636 337016 332688 337068
rect 336224 337016 336276 337068
rect 336776 337016 336828 337068
rect 341652 337016 341704 337068
rect 342664 337016 342716 337068
rect 343124 337016 343176 337068
rect 343584 337016 343636 337068
rect 343676 337016 343728 337068
rect 344044 337016 344096 337068
rect 345516 337016 345568 337068
rect 346620 337016 346672 337068
rect 347264 337016 347316 337068
rect 347816 337016 347868 337068
rect 348460 337016 348512 337068
rect 349472 337016 349524 337068
rect 84512 336948 84564 337000
rect 87364 336948 87416 337000
rect 248088 336948 248140 337000
rect 94264 336880 94316 336932
rect 249560 336880 249612 336932
rect 288016 336948 288068 337000
rect 290500 336948 290552 337000
rect 291512 336948 291564 337000
rect 291880 336948 291932 337000
rect 292892 336948 292944 337000
rect 298044 336948 298096 337000
rect 306140 336948 306192 337000
rect 308348 336948 308400 337000
rect 315156 336948 315208 337000
rect 316352 336948 316404 337000
rect 316628 336948 316680 337000
rect 317640 336948 317692 337000
rect 318652 336948 318704 337000
rect 319204 336948 319256 337000
rect 320124 336948 320176 337000
rect 320492 336948 320544 337000
rect 320768 336948 320820 337000
rect 321964 336948 322016 337000
rect 326472 336948 326524 337000
rect 327208 336948 327260 337000
rect 328128 336948 328180 337000
rect 328772 336948 328824 337000
rect 330888 336948 330940 337000
rect 331164 336948 331216 337000
rect 331808 336948 331860 337000
rect 332912 336948 332964 337000
rect 333832 336948 333884 337000
rect 334384 336948 334436 337000
rect 334568 336948 334620 337000
rect 335672 336948 335724 337000
rect 335948 336948 336000 337000
rect 336960 336948 337012 337000
rect 338892 336948 338944 337000
rect 339812 336948 339864 337000
rect 340180 336948 340232 337000
rect 341284 336948 341336 337000
rect 345792 336948 345844 337000
rect 346344 336948 346396 337000
rect 347724 336948 347776 337000
rect 348092 336948 348144 337000
rect 349748 336948 349800 337000
rect 350760 336948 350812 337000
rect 290960 336880 291012 336932
rect 291604 336880 291656 336932
rect 291696 336880 291748 336932
rect 292800 336880 292852 336932
rect 307612 336880 307664 336932
rect 307888 336880 307940 336932
rect 313960 336880 314012 336932
rect 314788 336880 314840 336932
rect 315892 336880 315944 336932
rect 316260 336880 316312 336932
rect 317180 336880 317232 336932
rect 317824 336880 317876 336932
rect 319572 336880 319624 336932
rect 320308 336880 320360 336932
rect 321320 336880 321372 336932
rect 321780 336880 321832 336932
rect 322792 336880 322844 336932
rect 323160 336880 323212 336932
rect 323528 336880 323580 336932
rect 324448 336880 324500 336932
rect 325184 336880 325236 336932
rect 326104 336880 326156 336932
rect 326932 336880 326984 336932
rect 327300 336880 327352 336932
rect 329140 336880 329192 336932
rect 330060 336880 330112 336932
rect 330336 336880 330388 336932
rect 331440 336880 331492 336932
rect 332360 336880 332412 336932
rect 333004 336880 333056 336932
rect 333280 336880 333332 336932
rect 334200 336880 334252 336932
rect 335304 336880 335356 336932
rect 335580 336880 335632 336932
rect 336500 336880 336552 336932
rect 337144 336880 337196 336932
rect 337420 336880 337472 336932
rect 338248 336880 338300 336932
rect 339352 336880 339404 336932
rect 339628 336880 339680 336932
rect 340640 336880 340692 336932
rect 341100 336880 341152 336932
rect 342756 336880 342808 336932
rect 343308 336880 343360 336932
rect 75036 336812 75088 336864
rect 84604 336812 84656 336864
rect 101164 336812 101216 336864
rect 245420 336812 245472 336864
rect 247628 336812 247680 336864
rect 249744 336812 249796 336864
rect 250572 336812 250624 336864
rect 256828 336812 256880 336864
rect 258668 336812 258720 336864
rect 276148 336812 276200 336864
rect 278724 336812 278776 336864
rect 284060 336812 284112 336864
rect 284152 336812 284204 336864
rect 285072 336812 285124 336864
rect 287096 336812 287148 336864
rect 287556 336812 287608 336864
rect 288844 336812 288896 336864
rect 289488 336812 289540 336864
rect 290684 336812 290736 336864
rect 291420 336812 291472 336864
rect 292432 336812 292484 336864
rect 292984 336812 293036 336864
rect 312488 336812 312540 336864
rect 313316 336812 313368 336864
rect 313500 336812 313552 336864
rect 313684 336812 313736 336864
rect 314420 336812 314472 336864
rect 314972 336812 315024 336864
rect 315432 336812 315484 336864
rect 316076 336812 316128 336864
rect 316904 336812 316956 336864
rect 317272 336812 317324 336864
rect 317364 336812 317416 336864
rect 317732 336812 317784 336864
rect 318100 336812 318152 336864
rect 318928 336812 318980 336864
rect 319664 336812 319716 336864
rect 320032 336812 320084 336864
rect 320216 336812 320268 336864
rect 320584 336812 320636 336864
rect 321504 336812 321556 336864
rect 321872 336812 321924 336864
rect 322240 336812 322292 336864
rect 322884 336812 322936 336864
rect 322976 336812 323028 336864
rect 323252 336812 323304 336864
rect 323712 336812 323764 336864
rect 324172 336812 324224 336864
rect 324264 336812 324316 336864
rect 324724 336812 324776 336864
rect 325000 336812 325052 336864
rect 325736 336812 325788 336864
rect 326196 336812 326248 336864
rect 327024 336812 327076 336864
rect 327944 336812 327996 336864
rect 328496 336812 328548 336864
rect 329416 336812 329468 336864
rect 329968 336812 330020 336864
rect 331072 336812 331124 336864
rect 331348 336812 331400 336864
rect 332544 336812 332596 336864
rect 332820 336812 332872 336864
rect 334016 336812 334068 336864
rect 334292 336812 334344 336864
rect 334752 336812 334804 336864
rect 335396 336812 335448 336864
rect 336684 336812 336736 336864
rect 337052 336812 337104 336864
rect 337236 336812 337288 336864
rect 338064 336812 338116 336864
rect 338156 336812 338208 336864
rect 338432 336812 338484 336864
rect 339168 336812 339220 336864
rect 339536 336812 339588 336864
rect 340916 336812 340968 336864
rect 341192 336812 341244 336864
rect 108064 336608 108116 336660
rect 355820 336608 355872 336660
rect 580392 336608 580444 336660
rect 119288 336404 119340 336456
rect 284980 336447 285032 336456
rect 284980 336413 284989 336447
rect 284989 336413 285023 336447
rect 285023 336413 285032 336447
rect 284980 336404 285032 336413
rect 225364 336268 225416 336320
rect 276516 336268 276568 336320
rect 302736 336268 302788 336320
rect 351036 336268 351088 336320
rect 181204 336064 181256 336116
rect 267408 336064 267460 336116
rect 304208 336064 304260 336116
rect 357936 336064 357988 336116
rect 127384 335996 127436 336048
rect 256460 335996 256512 336048
rect 323988 335996 324040 336048
rect 454536 335996 454588 336048
rect 275228 335860 275280 335912
rect 275412 335860 275464 335912
rect 275136 335792 275188 335844
rect 275596 335792 275648 335844
rect 231068 335724 231120 335776
rect 231620 335724 231672 335776
rect 235208 335724 235260 335776
rect 235484 335724 235536 335776
rect 237968 335724 238020 335776
rect 238428 335724 238480 335776
rect 239348 335724 239400 335776
rect 239900 335724 239952 335776
rect 245052 335724 245104 335776
rect 245236 335724 245288 335776
rect 247904 335724 247956 335776
rect 248640 335724 248692 335776
rect 253148 335724 253200 335776
rect 254068 335724 254120 335776
rect 254620 335724 254672 335776
rect 255540 335724 255592 335776
rect 260048 335724 260100 335776
rect 260876 335724 260928 335776
rect 264188 335724 264240 335776
rect 264832 335724 264884 335776
rect 265660 335724 265712 335776
rect 266304 335724 266356 335776
rect 268328 335724 268380 335776
rect 268972 335724 269024 335776
rect 269800 335724 269852 335776
rect 270444 335724 270496 335776
rect 271180 335724 271232 335776
rect 271916 335724 271968 335776
rect 273756 335724 273808 335776
rect 274860 335724 274912 335776
rect 276516 335724 276568 335776
rect 276792 335724 276844 335776
rect 328220 335724 328272 335776
rect 328680 335724 328732 335776
rect 229964 335520 230016 335572
rect 230700 335520 230752 335572
rect 231344 335520 231396 335572
rect 231988 335520 232040 335572
rect 233000 335520 233052 335572
rect 233460 335520 233512 335572
rect 233828 335520 233880 335572
rect 234748 335520 234800 335572
rect 235300 335520 235352 335572
rect 235668 335520 235720 335572
rect 236772 335520 236824 335572
rect 237140 335520 237192 335572
rect 238152 335520 238204 335572
rect 238612 335520 238664 335572
rect 239624 335520 239676 335572
rect 240360 335520 240412 335572
rect 240820 335520 240872 335572
rect 241096 335520 241148 335572
rect 242384 335520 242436 335572
rect 242568 335520 242620 335572
rect 244040 335520 244092 335572
rect 244500 335520 244552 335572
rect 244868 335520 244920 335572
rect 245512 335520 245564 335572
rect 247720 335520 247772 335572
rect 248456 335520 248508 335572
rect 249008 335520 249060 335572
rect 249928 335520 249980 335572
rect 253332 335520 253384 335572
rect 253608 335520 253660 335572
rect 254712 335520 254764 335572
rect 255264 335520 255316 335572
rect 257472 335520 257524 335572
rect 258208 335520 258260 335572
rect 258760 335520 258812 335572
rect 259496 335520 259548 335572
rect 260232 335520 260284 335572
rect 260692 335520 260744 335572
rect 261704 335520 261756 335572
rect 262348 335520 262400 335572
rect 262900 335520 262952 335572
rect 263360 335520 263412 335572
rect 264096 335520 264148 335572
rect 264372 335520 264424 335572
rect 265844 335520 265896 335572
rect 266580 335520 266632 335572
rect 267132 335520 267184 335572
rect 267776 335520 267828 335572
rect 268512 335520 268564 335572
rect 269248 335520 269300 335572
rect 269984 335520 270036 335572
rect 270720 335520 270772 335572
rect 274124 335520 274176 335572
rect 274676 335520 274728 335572
rect 276792 335520 276844 335572
rect 277344 335520 277396 335572
rect 278080 335520 278132 335572
rect 278816 335520 278868 335572
rect 279276 335520 279328 335572
rect 280288 335520 280340 335572
rect 280748 335520 280800 335572
rect 281484 335520 281536 335572
rect 327852 335520 327904 335572
rect 328680 335520 328732 335572
rect 333188 335520 333240 335572
rect 334292 335520 334344 335572
rect 337972 335520 338024 335572
rect 338432 335520 338484 335572
rect 231068 335452 231120 335504
rect 231804 335452 231856 335504
rect 232724 335452 232776 335504
rect 233276 335452 233328 335504
rect 237876 335452 237928 335504
rect 238888 335452 238940 335504
rect 239440 335452 239492 335504
rect 240084 335452 240136 335504
rect 242016 335452 242068 335504
rect 242292 335452 242344 335504
rect 243580 335452 243632 335504
rect 243948 335452 244000 335504
rect 270076 335452 270128 335504
rect 270260 335452 270312 335504
rect 272652 335452 272704 335504
rect 273388 335452 273440 335504
rect 284980 335452 285032 335504
rect 285624 335452 285676 335504
rect 289028 335452 289080 335504
rect 289672 335452 289724 335504
rect 313132 335452 313184 335504
rect 313592 335452 313644 335504
rect 318008 335452 318060 335504
rect 319204 335452 319256 335504
rect 319480 335452 319532 335504
rect 320492 335452 320544 335504
rect 322148 335452 322200 335504
rect 323068 335452 323120 335504
rect 240820 335384 240872 335436
rect 241556 335384 241608 335436
rect 264372 335384 264424 335436
rect 265108 335384 265160 335436
rect 250388 335316 250440 335368
rect 251124 335316 251176 335368
rect 251860 335316 251912 335368
rect 252596 335316 252648 335368
rect 338800 335316 338852 335368
rect 339812 335316 339864 335368
rect 250480 335248 250532 335300
rect 250756 335248 250808 335300
rect 251952 335248 252004 335300
rect 252412 335248 252464 335300
rect 277068 335248 277120 335300
rect 277528 335248 277580 335300
rect 319940 335291 319992 335300
rect 319940 335257 319949 335291
rect 319949 335257 319983 335291
rect 319983 335257 319992 335291
rect 319940 335248 319992 335257
rect 263176 334908 263228 334960
rect 263820 334908 263872 334960
rect 305588 334704 305640 334756
rect 366216 334704 366268 334756
rect 261520 334636 261572 334688
rect 342756 334636 342808 334688
rect 548376 334636 548428 334688
rect 280012 334296 280064 334348
rect 276516 333931 276568 333940
rect 276516 333897 276525 333931
rect 276525 333897 276559 333931
rect 276559 333897 276568 333931
rect 276516 333888 276568 333897
rect 236680 333548 236732 333600
rect 237416 333548 237468 333600
rect 204664 333344 204716 333396
rect 272376 333344 272428 333396
rect 303104 333344 303156 333396
rect 353796 333344 353848 333396
rect 163264 333276 163316 333328
rect 263728 333276 263780 333328
rect 284888 333276 284940 333328
rect 285164 333276 285216 333328
rect 329876 333276 329928 333328
rect 483516 333276 483568 333328
rect 145324 333208 145376 333260
rect 260140 333208 260192 333260
rect 262624 333208 262676 333260
rect 348828 333208 348880 333260
rect 575976 333208 576028 333260
rect 279368 332800 279420 332852
rect 279736 332800 279788 332852
rect 274308 331984 274360 332036
rect 287924 331984 287976 332036
rect 288384 331984 288436 332036
rect 307060 331984 307112 332036
rect 373024 331984 373076 332036
rect 117724 331916 117776 331968
rect 254436 331916 254488 331968
rect 278816 331916 278868 331968
rect 337696 331916 337748 331968
rect 520776 331916 520828 331968
rect 282312 331576 282364 331628
rect 283232 331576 283284 331628
rect 285440 331440 285492 331492
rect 259128 331372 259180 331424
rect 254712 331168 254764 331220
rect 254896 331168 254948 331220
rect 259036 331211 259088 331220
rect 259036 331177 259045 331211
rect 259045 331177 259079 331211
rect 259079 331177 259088 331211
rect 259036 331168 259088 331177
rect 340824 331168 340876 331220
rect 341192 331168 341244 331220
rect 259128 331143 259180 331152
rect 259128 331109 259137 331143
rect 259137 331109 259171 331143
rect 259171 331109 259180 331143
rect 259128 331100 259180 331109
rect 285164 331100 285216 331152
rect 285440 331100 285492 331152
rect 288752 331100 288804 331152
rect 371920 331143 371972 331152
rect 371920 331109 371929 331143
rect 371929 331109 371963 331143
rect 371963 331109 371972 331143
rect 371920 331100 371972 331109
rect 246432 331032 246484 331084
rect 246708 331032 246760 331084
rect 271364 331032 271416 331084
rect 271732 331032 271784 331084
rect 167404 330624 167456 330676
rect 264096 330624 264148 330676
rect 303564 330624 303616 330676
rect 355176 330624 355228 330676
rect 156364 330556 156416 330608
rect 262072 330556 262124 330608
rect 330520 330556 330572 330608
rect 486276 330556 486328 330608
rect 23884 330488 23936 330540
rect 235116 330488 235168 330540
rect 342020 330488 342072 330540
rect 342388 330488 342440 330540
rect 339352 330420 339404 330472
rect 530436 330488 530488 330540
rect 221224 329196 221276 329248
rect 275136 329196 275188 329248
rect 322516 329196 322568 329248
rect 447636 329196 447688 329248
rect 252504 328448 252556 328500
rect 252872 328448 252924 328500
rect 259312 328448 259364 328500
rect 259772 328448 259824 328500
rect 285348 328491 285400 328500
rect 285348 328457 285357 328491
rect 285357 328457 285391 328491
rect 285391 328457 285400 328491
rect 285348 328448 285400 328457
rect 285716 328448 285768 328500
rect 285992 328448 286044 328500
rect 333372 328448 333424 328500
rect 333924 328448 333976 328500
rect 229964 328380 230016 328432
rect 235576 328380 235628 328432
rect 268604 328423 268656 328432
rect 268604 328389 268613 328423
rect 268613 328389 268647 328423
rect 268647 328389 268656 328423
rect 268604 328380 268656 328389
rect 318652 328423 318704 328432
rect 318652 328389 318661 328423
rect 318661 328389 318695 328423
rect 318695 328389 318704 328423
rect 318652 328380 318704 328389
rect 328128 328380 328180 328432
rect 328220 328380 328272 328432
rect 371920 328423 371972 328432
rect 371920 328389 371929 328423
rect 371929 328389 371963 328423
rect 371963 328389 371972 328423
rect 371920 328380 371972 328389
rect 218464 327836 218516 327888
rect 273756 327836 273808 327888
rect 305128 327836 305180 327888
rect 362076 327836 362128 327888
rect 264372 327768 264424 327820
rect 331256 327768 331308 327820
rect 490416 327768 490468 327820
rect 77704 327700 77756 327752
rect 246156 327700 246208 327752
rect 341836 327700 341888 327752
rect 541476 327700 541528 327752
rect 152224 327131 152276 327140
rect 152224 327097 152233 327131
rect 152233 327097 152267 327131
rect 152267 327097 152276 327131
rect 152224 327088 152276 327097
rect 170164 327131 170216 327140
rect 170164 327097 170173 327131
rect 170173 327097 170207 327131
rect 170207 327097 170216 327131
rect 170164 327088 170216 327097
rect 214324 327131 214376 327140
rect 214324 327097 214333 327131
rect 214333 327097 214367 327131
rect 214367 327097 214376 327131
rect 214324 327088 214376 327097
rect 246524 327088 246576 327140
rect 246708 327088 246760 327140
rect 279828 327131 279880 327140
rect 279828 327097 279837 327131
rect 279837 327097 279871 327131
rect 279871 327097 279880 327131
rect 279828 327088 279880 327097
rect 392252 327088 392304 327140
rect 392436 327088 392488 327140
rect 328128 327063 328180 327072
rect 328128 327029 328137 327063
rect 328137 327029 328171 327063
rect 328171 327029 328180 327063
rect 328128 327020 328180 327029
rect 373024 327063 373076 327072
rect 373024 327029 373033 327063
rect 373033 327029 373067 327063
rect 373067 327029 373076 327063
rect 373024 327020 373076 327029
rect 278724 326859 278776 326868
rect 278724 326825 278733 326859
rect 278733 326825 278767 326859
rect 278767 326825 278776 326859
rect 278724 326816 278776 326825
rect 186724 326476 186776 326528
rect 268236 326476 268288 326528
rect 327024 326476 327076 326528
rect 465576 326476 465628 326528
rect 229504 325048 229556 325100
rect 276884 325048 276936 325100
rect 306508 325048 306560 325100
rect 368976 325048 369028 325100
rect 174304 324980 174356 325032
rect 265936 324980 265988 325032
rect 332636 324980 332688 325032
rect 494556 324980 494608 325032
rect 73564 324912 73616 324964
rect 245052 324912 245104 324964
rect 345056 324912 345108 324964
rect 553896 324912 553948 324964
rect 275780 324368 275832 324420
rect 276148 324368 276200 324420
rect 276608 324368 276660 324420
rect 272928 324300 272980 324352
rect 273020 324300 273072 324352
rect 275688 324300 275740 324352
rect 275964 324300 276016 324352
rect 194912 323552 194964 323604
rect 270168 323552 270220 323604
rect 313316 323552 313368 323604
rect 399336 323552 399388 323604
rect 177064 322260 177116 322312
rect 265844 322260 265896 322312
rect 332728 322260 332780 322312
rect 497316 322260 497368 322312
rect 135664 322192 135716 322244
rect 257932 322192 257984 322244
rect 299516 322192 299568 322244
rect 331716 322192 331768 322244
rect 343676 322192 343728 322244
rect 552516 322192 552568 322244
rect 235760 321920 235812 321972
rect 239256 321580 239308 321632
rect 239440 321580 239492 321632
rect 258944 321580 258996 321632
rect 259128 321580 259180 321632
rect 272560 321580 272612 321632
rect 272744 321580 272796 321632
rect 340824 321580 340876 321632
rect 341192 321580 341244 321632
rect 229872 321419 229924 321428
rect 229872 321385 229881 321419
rect 229881 321385 229915 321419
rect 229915 321385 229924 321419
rect 229872 321376 229924 321385
rect 268696 321376 268748 321428
rect 318652 321419 318704 321428
rect 318652 321385 318661 321419
rect 318661 321385 318695 321419
rect 318695 321385 318704 321419
rect 318652 321376 318704 321385
rect 340824 321376 340876 321428
rect 341192 321376 341244 321428
rect 371920 321419 371972 321428
rect 371920 321385 371929 321419
rect 371929 321385 371963 321419
rect 371963 321385 371972 321419
rect 371920 321376 371972 321385
rect 110824 320832 110876 320884
rect 252504 320832 252556 320884
rect 261244 320671 261296 320680
rect 261244 320637 261253 320671
rect 261253 320637 261287 320671
rect 261287 320637 261296 320671
rect 261244 320628 261296 320637
rect 254160 320492 254212 320544
rect 261152 320492 261204 320544
rect 488300 320492 488352 320544
rect 493084 320492 493136 320544
rect 418564 320288 418616 320340
rect 425464 320288 425516 320340
rect 437884 320288 437936 320340
rect 444784 320288 444836 320340
rect 457204 320288 457256 320340
rect 464104 320288 464156 320340
rect 476524 320288 476576 320340
rect 483424 320288 483476 320340
rect 541568 320288 541620 320340
rect 544328 320288 544380 320340
rect 261244 320263 261296 320272
rect 261244 320229 261253 320263
rect 261253 320229 261287 320263
rect 261287 320229 261296 320263
rect 261244 320220 261296 320229
rect 290316 320220 290368 320272
rect 294640 320220 294692 320272
rect 311936 319540 311988 319592
rect 395196 319540 395248 319592
rect 185344 319472 185396 319524
rect 267592 319472 267644 319524
rect 333924 319472 333976 319524
rect 501456 319472 501508 319524
rect 134192 319404 134244 319456
rect 257564 319404 257616 319456
rect 346344 319404 346396 319456
rect 560796 319404 560848 319456
rect 235484 318903 235536 318912
rect 235484 318869 235493 318903
rect 235493 318869 235527 318903
rect 235527 318869 235536 318903
rect 235484 318860 235536 318869
rect 235668 318903 235720 318912
rect 235668 318869 235677 318903
rect 235677 318869 235711 318903
rect 235711 318869 235720 318903
rect 235668 318860 235720 318869
rect 277068 318860 277120 318912
rect 235484 318699 235536 318708
rect 235484 318665 235493 318699
rect 235493 318665 235527 318699
rect 235527 318665 235536 318699
rect 235484 318656 235536 318665
rect 235668 318656 235720 318708
rect 235944 318656 235996 318708
rect 276976 318699 277028 318708
rect 276976 318665 276985 318699
rect 276985 318665 277019 318699
rect 277019 318665 277028 318699
rect 276976 318656 277028 318665
rect 285256 318699 285308 318708
rect 285256 318665 285265 318699
rect 285265 318665 285299 318699
rect 285299 318665 285308 318699
rect 285256 318656 285308 318665
rect 285624 318699 285676 318708
rect 285624 318665 285633 318699
rect 285633 318665 285667 318699
rect 285667 318665 285676 318699
rect 285624 318656 285676 318665
rect 318928 318699 318980 318708
rect 318928 318665 318937 318699
rect 318937 318665 318971 318699
rect 318971 318665 318980 318699
rect 318928 318656 318980 318665
rect 319112 318699 319164 318708
rect 319112 318665 319121 318699
rect 319121 318665 319155 318699
rect 319155 318665 319164 318699
rect 319112 318656 319164 318665
rect 373116 318656 373168 318708
rect 319204 318588 319256 318640
rect 319204 318452 319256 318504
rect 197764 318112 197816 318164
rect 269984 318112 270036 318164
rect 314788 318112 314840 318164
rect 406236 318112 406288 318164
rect 138424 318044 138476 318096
rect 256460 318044 256512 318096
rect 334016 318044 334068 318096
rect 504216 318044 504268 318096
rect 320124 317432 320176 317484
rect 328404 317432 328456 317484
rect 135664 317407 135716 317416
rect 135664 317373 135673 317407
rect 135673 317373 135707 317407
rect 135707 317373 135716 317407
rect 135664 317364 135716 317373
rect 152224 317407 152276 317416
rect 152224 317373 152233 317407
rect 152233 317373 152267 317407
rect 152267 317373 152276 317407
rect 152224 317364 152276 317373
rect 170164 317407 170216 317416
rect 170164 317373 170173 317407
rect 170173 317373 170207 317407
rect 170207 317373 170216 317407
rect 170164 317364 170216 317373
rect 214324 317407 214376 317416
rect 214324 317373 214333 317407
rect 214333 317373 214367 317407
rect 214367 317373 214376 317407
rect 214324 317364 214376 317373
rect 385536 317407 385588 317416
rect 385536 317373 385545 317407
rect 385545 317373 385579 317407
rect 385579 317373 385588 317407
rect 392436 317407 392488 317416
rect 385536 317364 385588 317373
rect 392436 317373 392445 317407
rect 392445 317373 392479 317407
rect 392479 317373 392488 317407
rect 392436 317364 392488 317373
rect 342204 316752 342256 316804
rect 342388 316752 342440 316804
rect 121864 316684 121916 316736
rect 254804 316684 254856 316736
rect 317456 316684 317508 316736
rect 420036 316684 420088 316736
rect 201904 315324 201956 315376
rect 271640 315324 271692 315376
rect 316076 315324 316128 315376
rect 413136 315324 413188 315376
rect 142564 315256 142616 315308
rect 258944 315256 258996 315308
rect 335304 315256 335356 315308
rect 508356 315256 508408 315308
rect 275504 314644 275556 314696
rect 275688 314644 275740 314696
rect 318928 314075 318980 314084
rect 318928 314041 318937 314075
rect 318937 314041 318971 314075
rect 318971 314041 318980 314075
rect 318928 314032 318980 314041
rect 242660 313964 242712 314016
rect 242844 313964 242896 314016
rect 305220 313964 305272 314016
rect 360696 313964 360748 314016
rect 149464 312604 149516 312656
rect 260232 312604 260284 312656
rect 313408 312604 313460 312656
rect 402096 312604 402148 312656
rect 14224 312536 14276 312588
rect 233092 312536 233144 312588
rect 350760 312536 350812 312588
rect 579380 312536 579432 312588
rect 268696 311967 268748 311976
rect 268696 311933 268705 311967
rect 268705 311933 268739 311967
rect 268739 311933 268748 311967
rect 268696 311924 268748 311933
rect 318744 311924 318796 311976
rect 331164 311967 331216 311976
rect 331164 311933 331173 311967
rect 331173 311933 331207 311967
rect 331207 311933 331216 311967
rect 331164 311924 331216 311933
rect 372012 311924 372064 311976
rect 235576 311788 235628 311840
rect 249468 311788 249520 311840
rect 249652 311788 249704 311840
rect 309176 311831 309228 311840
rect 309176 311797 309185 311831
rect 309185 311797 309219 311831
rect 309219 311797 309228 311831
rect 309176 311788 309228 311797
rect 318744 311788 318796 311840
rect 371920 311788 371972 311840
rect 268696 311627 268748 311636
rect 268696 311593 268705 311627
rect 268705 311593 268739 311627
rect 268739 311593 268748 311627
rect 268696 311584 268748 311593
rect 306600 311244 306652 311296
rect 367596 311244 367648 311296
rect 3644 310428 3696 310480
rect 226100 310428 226152 310480
rect 319112 309859 319164 309868
rect 319112 309825 319121 309859
rect 319121 309825 319155 309859
rect 319155 309825 319164 309859
rect 319112 309816 319164 309825
rect 321596 309816 321648 309868
rect 440736 309816 440788 309868
rect 268512 309748 268564 309800
rect 345148 309748 345200 309800
rect 555276 309748 555328 309800
rect 285440 309272 285492 309324
rect 331256 309204 331308 309256
rect 242476 309136 242528 309188
rect 242568 309136 242620 309188
rect 285348 309136 285400 309188
rect 285440 309136 285492 309188
rect 285716 309136 285768 309188
rect 309176 309179 309228 309188
rect 309176 309145 309185 309179
rect 309185 309145 309219 309179
rect 309219 309145 309228 309179
rect 309176 309136 309228 309145
rect 340824 309136 340876 309188
rect 341192 309136 341244 309188
rect 225364 309111 225416 309120
rect 225364 309077 225373 309111
rect 225373 309077 225407 309111
rect 225407 309077 225416 309111
rect 225364 309068 225416 309077
rect 259312 309111 259364 309120
rect 259312 309077 259321 309111
rect 259321 309077 259355 309111
rect 259355 309077 259364 309111
rect 259312 309068 259364 309077
rect 357936 309111 357988 309120
rect 357936 309077 357945 309111
rect 357945 309077 357979 309111
rect 357979 309077 357988 309111
rect 357936 309068 357988 309077
rect 371920 309068 371972 309120
rect 373116 309068 373168 309120
rect 373208 309068 373260 309120
rect 552516 309068 552568 309120
rect 552608 309068 552660 309120
rect 135664 307819 135716 307828
rect 135664 307785 135673 307819
rect 135673 307785 135707 307819
rect 135707 307785 135716 307819
rect 135664 307776 135716 307785
rect 152224 307819 152276 307828
rect 152224 307785 152233 307819
rect 152233 307785 152267 307819
rect 152267 307785 152276 307819
rect 152224 307776 152276 307785
rect 170164 307819 170216 307828
rect 170164 307785 170173 307819
rect 170173 307785 170207 307819
rect 170207 307785 170216 307819
rect 170164 307776 170216 307785
rect 190864 307819 190916 307828
rect 190864 307785 190873 307819
rect 190873 307785 190907 307819
rect 190907 307785 190916 307819
rect 190864 307776 190916 307785
rect 214324 307819 214376 307828
rect 214324 307785 214333 307819
rect 214333 307785 214367 307819
rect 214367 307785 214376 307819
rect 214324 307776 214376 307785
rect 319940 307776 319992 307828
rect 320124 307776 320176 307828
rect 385536 307819 385588 307828
rect 385536 307785 385545 307819
rect 385545 307785 385579 307819
rect 385579 307785 385588 307819
rect 392436 307819 392488 307828
rect 385536 307776 385588 307785
rect 392436 307785 392445 307819
rect 392445 307785 392479 307819
rect 392479 307785 392488 307819
rect 392436 307776 392488 307785
rect 229872 307708 229924 307760
rect 229964 307708 230016 307760
rect 372932 307708 372984 307760
rect 373208 307708 373260 307760
rect 160504 307096 160556 307148
rect 263084 307096 263136 307148
rect 321688 307096 321740 307148
rect 443588 307096 443640 307148
rect 103924 307028 103976 307080
rect 250940 307028 250992 307080
rect 339536 307028 339588 307080
rect 529056 307028 529108 307080
rect 342204 306348 342256 306400
rect 342388 306348 342440 306400
rect 272560 304920 272612 304972
rect 272836 304920 272888 304972
rect 273020 304920 273072 304972
rect 273204 304920 273256 304972
rect 276608 304920 276660 304972
rect 276700 304920 276752 304972
rect 276976 304920 277028 304972
rect 277252 304852 277304 304904
rect 322976 304308 323028 304360
rect 451776 304308 451828 304360
rect 128764 304240 128816 304292
rect 256000 304240 256052 304292
rect 343768 304240 343820 304292
rect 546996 304240 547048 304292
rect 235760 302268 235812 302320
rect 239256 302268 239308 302320
rect 239348 302268 239400 302320
rect 285348 302268 285400 302320
rect 285716 302268 285768 302320
rect 235668 302132 235720 302184
rect 239256 302132 239308 302184
rect 239348 302132 239400 302184
rect 285256 302132 285308 302184
rect 331164 302200 331216 302252
rect 331256 302132 331308 302184
rect 340824 302132 340876 302184
rect 341192 302132 341244 302184
rect 371828 302175 371880 302184
rect 371828 302141 371837 302175
rect 371837 302141 371871 302175
rect 371871 302141 371880 302175
rect 371828 302132 371880 302141
rect 285808 302064 285860 302116
rect 324356 301520 324408 301572
rect 458676 301520 458728 301572
rect 139804 301452 139856 301504
rect 258852 301452 258904 301504
rect 346436 301452 346488 301504
rect 563556 301452 563608 301504
rect 325736 300160 325788 300212
rect 461436 300160 461488 300212
rect 142472 300092 142524 300144
rect 258760 300092 258812 300144
rect 347816 300092 347868 300144
rect 567696 300092 567748 300144
rect 225364 299523 225416 299532
rect 225364 299489 225373 299523
rect 225373 299489 225407 299523
rect 225407 299489 225416 299523
rect 225364 299480 225416 299489
rect 242476 299480 242528 299532
rect 242568 299480 242620 299532
rect 259404 299480 259456 299532
rect 271364 299480 271416 299532
rect 275688 299480 275740 299532
rect 357936 299523 357988 299532
rect 357936 299489 357945 299523
rect 357945 299489 357979 299523
rect 357979 299489 357988 299523
rect 357936 299480 357988 299489
rect 235668 299455 235720 299464
rect 235668 299421 235677 299455
rect 235677 299421 235711 299455
rect 235711 299421 235720 299455
rect 235668 299412 235720 299421
rect 239256 299412 239308 299464
rect 239440 299412 239492 299464
rect 309176 299455 309228 299464
rect 309176 299421 309185 299455
rect 309185 299421 309219 299455
rect 309219 299421 309228 299455
rect 309176 299412 309228 299421
rect 553804 299412 553856 299464
rect 553896 299412 553948 299464
rect 271456 299344 271508 299396
rect 272560 298732 272612 298784
rect 272928 298732 272980 298784
rect 229872 297984 229924 298036
rect 230240 297984 230292 298036
rect 319940 298027 319992 298036
rect 319940 297993 319949 298027
rect 319949 297993 319983 298027
rect 319983 297993 319992 298027
rect 319940 297984 319992 297993
rect 183964 297440 184016 297492
rect 267132 297440 267184 297492
rect 307888 297440 307940 297492
rect 374496 297440 374548 297492
rect 29404 297372 29456 297424
rect 340916 297372 340968 297424
rect 534576 297372 534628 297424
rect 275504 296939 275556 296948
rect 275504 296905 275513 296939
rect 275513 296905 275547 296939
rect 275547 296905 275556 296939
rect 275504 296896 275556 296905
rect 278724 296692 278776 296744
rect 278908 296692 278960 296744
rect 342204 296692 342256 296744
rect 342388 296692 342440 296744
rect 272652 295579 272704 295588
rect 272652 295545 272661 295579
rect 272661 295545 272695 295579
rect 272695 295545 272704 295579
rect 272652 295536 272704 295545
rect 272744 295511 272796 295520
rect 272744 295477 272753 295511
rect 272753 295477 272787 295511
rect 272787 295477 272796 295511
rect 272744 295468 272796 295477
rect 249376 295264 249428 295316
rect 249652 295264 249704 295316
rect 272744 295307 272796 295316
rect 272744 295273 272753 295307
rect 272753 295273 272787 295307
rect 272787 295273 272796 295307
rect 272744 295264 272796 295273
rect 276700 295307 276752 295316
rect 276700 295273 276709 295307
rect 276709 295273 276743 295307
rect 276743 295273 276752 295307
rect 276700 295264 276752 295273
rect 278448 295264 278500 295316
rect 278724 295264 278776 295316
rect 272652 295239 272704 295248
rect 272652 295205 272661 295239
rect 272661 295205 272695 295239
rect 272695 295205 272704 295239
rect 272652 295196 272704 295205
rect 276608 295239 276660 295248
rect 276608 295205 276617 295239
rect 276617 295205 276651 295239
rect 276651 295205 276660 295239
rect 276608 295196 276660 295205
rect 340824 294924 340876 294976
rect 341192 294924 341244 294976
rect 81844 294584 81896 294636
rect 246432 294584 246484 294636
rect 303472 294584 303524 294636
rect 339996 294584 340048 294636
rect 341008 294584 341060 294636
rect 537336 294584 537388 294636
rect 3552 293836 3604 293888
rect 6680 293836 6732 293888
rect 331164 292544 331216 292596
rect 268696 292476 268748 292528
rect 331256 292476 331308 292528
rect 320124 292408 320176 292460
rect 268696 292340 268748 292392
rect 84604 291796 84656 291848
rect 245420 291796 245472 291848
rect 342296 291796 342348 291848
rect 545616 291796 545668 291848
rect 235484 289824 235536 289876
rect 235576 289824 235628 289876
rect 309176 289867 309228 289876
rect 309176 289833 309185 289867
rect 309185 289833 309219 289867
rect 309219 289833 309228 289867
rect 309176 289824 309228 289833
rect 259404 289799 259456 289808
rect 259404 289765 259413 289799
rect 259413 289765 259447 289799
rect 259447 289765 259456 289799
rect 259404 289756 259456 289765
rect 341192 289756 341244 289808
rect 354440 289756 354492 289808
rect 580668 289756 580720 289808
rect 357936 289688 357988 289740
rect 371920 289731 371972 289740
rect 371920 289697 371929 289731
rect 371929 289697 371963 289731
rect 371963 289697 371972 289731
rect 371920 289688 371972 289697
rect 553896 289731 553948 289740
rect 553896 289697 553905 289731
rect 553905 289697 553939 289731
rect 553939 289697 553948 289731
rect 553896 289688 553948 289697
rect 88744 289076 88796 289128
rect 248272 289076 248324 289128
rect 135480 288396 135532 288448
rect 135664 288396 135716 288448
rect 152040 288396 152092 288448
rect 152224 288396 152276 288448
rect 170164 288396 170216 288448
rect 170348 288396 170400 288448
rect 190680 288396 190732 288448
rect 190864 288396 190916 288448
rect 214324 288396 214376 288448
rect 214508 288396 214560 288448
rect 385536 288396 385588 288448
rect 385720 288396 385772 288448
rect 392436 288396 392488 288448
rect 392620 288396 392672 288448
rect 528872 288396 528924 288448
rect 529056 288396 529108 288448
rect 372840 288192 372892 288244
rect 373116 288192 373168 288244
rect 229964 287036 230016 287088
rect 230148 287036 230200 287088
rect 314880 286356 314932 286408
rect 408996 286356 409048 286408
rect 249192 286288 249244 286340
rect 347908 286288 347960 286340
rect 571836 286288 571888 286340
rect 276608 285719 276660 285728
rect 276608 285685 276617 285719
rect 276617 285685 276651 285719
rect 276651 285685 276660 285719
rect 276608 285676 276660 285685
rect 276976 285676 277028 285728
rect 235484 285311 235536 285320
rect 235484 285277 235493 285311
rect 235493 285277 235527 285311
rect 235527 285277 235536 285311
rect 235484 285268 235536 285277
rect 276976 285132 277028 285184
rect 268696 284971 268748 284980
rect 268696 284937 268705 284971
rect 268705 284937 268739 284971
rect 268739 284937 268748 284971
rect 268696 284928 268748 284937
rect 272836 284248 272888 284300
rect 272928 284248 272980 284300
rect 316168 283636 316220 283688
rect 417368 283636 417420 283688
rect 95644 283568 95696 283620
rect 249376 283568 249428 283620
rect 349288 283568 349340 283620
rect 578000 283568 578052 283620
rect 271456 283067 271508 283076
rect 271456 283033 271465 283067
rect 271465 283033 271499 283067
rect 271499 283033 271508 283067
rect 271456 283024 271508 283033
rect 341100 282999 341152 283008
rect 341100 282965 341109 282999
rect 341109 282965 341143 282999
rect 341143 282965 341152 282999
rect 341100 282956 341152 282965
rect 235576 282752 235628 282804
rect 268788 282752 268840 282804
rect 271456 282795 271508 282804
rect 271456 282761 271465 282795
rect 271465 282761 271499 282795
rect 271499 282761 271508 282795
rect 271456 282752 271508 282761
rect 341100 282795 341152 282804
rect 341100 282761 341109 282795
rect 341109 282761 341143 282795
rect 341143 282761 341152 282795
rect 341100 282752 341152 282761
rect 371920 282795 371972 282804
rect 371920 282761 371929 282795
rect 371929 282761 371963 282795
rect 371963 282761 371972 282795
rect 371920 282752 371972 282761
rect 276792 280483 276844 280492
rect 276792 280449 276801 280483
rect 276801 280449 276835 280483
rect 276835 280449 276844 280483
rect 276792 280440 276844 280449
rect 357936 280304 357988 280356
rect 91504 280279 91556 280288
rect 91504 280245 91513 280279
rect 91513 280245 91547 280279
rect 91547 280245 91556 280279
rect 91504 280236 91556 280245
rect 259404 280279 259456 280288
rect 259404 280245 259413 280279
rect 259413 280245 259447 280279
rect 259447 280245 259456 280279
rect 259404 280236 259456 280245
rect 340916 280279 340968 280288
rect 340916 280245 340925 280279
rect 340925 280245 340959 280279
rect 340959 280245 340968 280279
rect 340916 280236 340968 280245
rect 373116 280236 373168 280288
rect 553896 280279 553948 280288
rect 553896 280245 553905 280279
rect 553905 280245 553939 280279
rect 553939 280245 553948 280279
rect 553896 280236 553948 280245
rect 276792 280075 276844 280084
rect 276792 280041 276801 280075
rect 276801 280041 276835 280075
rect 276835 280041 276844 280075
rect 276792 280032 276844 280041
rect 309176 280075 309228 280084
rect 309176 280041 309185 280075
rect 309185 280041 309219 280075
rect 309219 280041 309228 280075
rect 309176 280032 309228 280041
rect 331256 280075 331308 280084
rect 331256 280041 331265 280075
rect 331265 280041 331299 280075
rect 331299 280041 331308 280075
rect 331256 280032 331308 280041
rect 276700 280007 276752 280016
rect 276700 279973 276709 280007
rect 276709 279973 276743 280007
rect 276743 279973 276752 280007
rect 276700 279964 276752 279973
rect 285164 279871 285216 279880
rect 285164 279837 285173 279871
rect 285173 279837 285207 279871
rect 285207 279837 285216 279871
rect 285164 279828 285216 279837
rect 285256 279871 285308 279880
rect 285256 279837 285265 279871
rect 285265 279837 285299 279871
rect 285299 279837 285308 279871
rect 285256 279828 285308 279837
rect 99784 279420 99836 279472
rect 249560 279420 249612 279472
rect 335396 279420 335448 279472
rect 506976 279420 507028 279472
rect 242108 278851 242160 278860
rect 242108 278817 242117 278851
rect 242117 278817 242151 278851
rect 242151 278817 242160 278851
rect 242108 278808 242160 278817
rect 246616 278851 246668 278860
rect 246616 278817 246625 278851
rect 246625 278817 246659 278851
rect 246659 278817 246668 278851
rect 246616 278808 246668 278817
rect 229964 278740 230016 278792
rect 230056 278740 230108 278792
rect 372932 278783 372984 278792
rect 372932 278749 372941 278783
rect 372941 278749 372975 278783
rect 372975 278749 372984 278783
rect 372932 278740 372984 278749
rect 552516 278740 552568 278792
rect 552608 278740 552660 278792
rect 285716 278672 285768 278724
rect 285808 278672 285860 278724
rect 242108 277355 242160 277364
rect 242108 277321 242117 277355
rect 242117 277321 242151 277355
rect 242151 277321 242160 277355
rect 242108 277312 242160 277321
rect 246616 277355 246668 277364
rect 246616 277321 246625 277355
rect 246625 277321 246659 277355
rect 246659 277321 246668 277355
rect 246616 277312 246668 277321
rect 90124 276632 90176 276684
rect 247720 276632 247772 276684
rect 336776 276632 336828 276684
rect 513876 276632 513928 276684
rect 273020 275952 273072 276004
rect 273112 275952 273164 276004
rect 328220 275952 328272 276004
rect 328404 275952 328456 276004
rect 272836 274592 272888 274644
rect 273020 274592 273072 274644
rect 358580 274592 358632 274644
rect 580668 274592 580720 274644
rect 19744 273912 19796 273964
rect 234104 273912 234156 273964
rect 239256 273232 239308 273284
rect 239440 273232 239492 273284
rect 246800 273300 246852 273352
rect 259404 273300 259456 273352
rect 372012 273300 372064 273352
rect 246708 273164 246760 273216
rect 371920 273164 371972 273216
rect 125912 271124 125964 271176
rect 255908 271124 255960 271176
rect 341100 271124 341152 271176
rect 259312 270555 259364 270564
rect 259312 270521 259321 270555
rect 259321 270521 259355 270555
rect 259355 270521 259364 270555
rect 259312 270512 259364 270521
rect 285348 270512 285400 270564
rect 309176 270555 309228 270564
rect 309176 270521 309185 270555
rect 309185 270521 309219 270555
rect 309219 270521 309228 270555
rect 309176 270512 309228 270521
rect 331256 270555 331308 270564
rect 331256 270521 331265 270555
rect 331265 270521 331299 270555
rect 331299 270521 331308 270555
rect 331256 270512 331308 270521
rect 91504 270487 91556 270496
rect 91504 270453 91513 270487
rect 91513 270453 91547 270487
rect 91547 270453 91556 270487
rect 91504 270444 91556 270453
rect 225364 270487 225416 270496
rect 225364 270453 225373 270487
rect 225373 270453 225407 270487
rect 225407 270453 225416 270487
rect 225364 270444 225416 270453
rect 357936 270487 357988 270496
rect 357936 270453 357945 270487
rect 357945 270453 357979 270487
rect 357979 270453 357988 270487
rect 553896 270487 553948 270496
rect 357936 270444 357988 270453
rect 553896 270453 553905 270487
rect 553905 270453 553939 270487
rect 553939 270453 553948 270487
rect 553896 270444 553948 270453
rect 278448 270240 278500 270292
rect 278816 270240 278868 270292
rect 242752 269739 242804 269748
rect 242752 269705 242761 269739
rect 242761 269705 242795 269739
rect 242795 269705 242804 269739
rect 242752 269696 242804 269705
rect 135480 269084 135532 269136
rect 135664 269084 135716 269136
rect 152040 269084 152092 269136
rect 152224 269084 152276 269136
rect 170164 269084 170216 269136
rect 170348 269084 170400 269136
rect 190680 269084 190732 269136
rect 190864 269084 190916 269136
rect 214324 269084 214376 269136
rect 214508 269084 214560 269136
rect 229780 269084 229832 269136
rect 229872 269084 229924 269136
rect 235392 269084 235444 269136
rect 235576 269084 235628 269136
rect 268604 269084 268656 269136
rect 268696 269084 268748 269136
rect 279828 269084 279880 269136
rect 280012 269084 280064 269136
rect 285164 269127 285216 269136
rect 285164 269093 285173 269127
rect 285173 269093 285207 269127
rect 285207 269093 285216 269127
rect 285164 269084 285216 269093
rect 372932 269084 372984 269136
rect 373116 269084 373168 269136
rect 385536 269084 385588 269136
rect 385720 269084 385772 269136
rect 392436 269084 392488 269136
rect 392620 269084 392672 269136
rect 528872 269084 528924 269136
rect 529056 269084 529108 269136
rect 535956 269127 536008 269136
rect 535956 269093 535965 269127
rect 535965 269093 535999 269127
rect 535999 269093 536008 269127
rect 535956 269084 536008 269093
rect 552608 269084 552660 269136
rect 552792 269084 552844 269136
rect 571836 269084 571888 269136
rect 572020 269084 572072 269136
rect 342388 268336 342440 268388
rect 542856 268336 542908 268388
rect 242568 267792 242620 267844
rect 242476 267724 242528 267776
rect 242936 267520 242988 267572
rect 300896 265616 300948 265668
rect 342756 265616 342808 265668
rect 343860 265616 343912 265668
rect 549756 265616 549808 265668
rect 242936 264800 242988 264852
rect 235576 263644 235628 263696
rect 239256 263576 239308 263628
rect 239440 263576 239492 263628
rect 285348 263644 285400 263696
rect 320032 263619 320084 263628
rect 320032 263585 320041 263619
rect 320041 263585 320075 263619
rect 320075 263585 320084 263619
rect 320032 263576 320084 263585
rect 328404 263644 328456 263696
rect 341192 263644 341244 263696
rect 285256 263508 285308 263560
rect 328312 263508 328364 263560
rect 341100 263508 341152 263560
rect 235576 263440 235628 263492
rect 345240 262828 345292 262880
rect 556656 262828 556708 262880
rect 351772 261468 351824 261520
rect 574596 261468 574648 261520
rect 553896 260967 553948 260976
rect 553896 260933 553905 260967
rect 553905 260933 553939 260967
rect 553939 260933 553948 260967
rect 553896 260924 553948 260933
rect 91504 260899 91556 260908
rect 91504 260865 91513 260899
rect 91513 260865 91547 260899
rect 91547 260865 91556 260899
rect 91504 260856 91556 260865
rect 225364 260899 225416 260908
rect 225364 260865 225373 260899
rect 225373 260865 225407 260899
rect 225407 260865 225416 260899
rect 225364 260856 225416 260865
rect 279736 260856 279788 260908
rect 279828 260856 279880 260908
rect 357936 260899 357988 260908
rect 357936 260865 357945 260899
rect 357945 260865 357979 260899
rect 357979 260865 357988 260899
rect 357936 260856 357988 260865
rect 3828 260788 3880 260840
rect 179180 260788 179232 260840
rect 235576 260831 235628 260840
rect 235576 260797 235585 260831
rect 235585 260797 235619 260831
rect 235619 260797 235628 260831
rect 235576 260788 235628 260797
rect 285624 260831 285676 260840
rect 285624 260797 285633 260831
rect 285633 260797 285667 260831
rect 285667 260797 285676 260831
rect 285624 260788 285676 260797
rect 331256 260831 331308 260840
rect 331256 260797 331265 260831
rect 331265 260797 331299 260831
rect 331299 260797 331308 260831
rect 331256 260788 331308 260797
rect 341100 260831 341152 260840
rect 341100 260797 341109 260831
rect 341109 260797 341143 260831
rect 341143 260797 341152 260831
rect 341100 260788 341152 260797
rect 553896 260788 553948 260840
rect 285256 260763 285308 260772
rect 285256 260729 285265 260763
rect 285265 260729 285299 260763
rect 285299 260729 285308 260763
rect 285256 260720 285308 260729
rect 553804 260720 553856 260772
rect 305036 259403 305088 259412
rect 305036 259369 305045 259403
rect 305045 259369 305079 259403
rect 305079 259369 305088 259403
rect 305036 259360 305088 259369
rect 320032 258111 320084 258120
rect 320032 258077 320041 258111
rect 320041 258077 320075 258111
rect 320075 258077 320084 258111
rect 320032 258068 320084 258077
rect 273020 256887 273072 256896
rect 273020 256853 273029 256887
rect 273029 256853 273063 256887
rect 273063 256853 273072 256887
rect 273020 256844 273072 256853
rect 328312 256683 328364 256692
rect 328312 256649 328321 256683
rect 328321 256649 328355 256683
rect 328355 256649 328364 256683
rect 328312 256640 328364 256649
rect 279736 256028 279788 256080
rect 279828 255960 279880 256012
rect 242844 255323 242896 255332
rect 242844 255289 242853 255323
rect 242853 255289 242887 255323
rect 242887 255289 242896 255323
rect 242844 255280 242896 255289
rect 273020 255323 273072 255332
rect 273020 255289 273029 255323
rect 273029 255289 273063 255323
rect 273063 255289 273072 255323
rect 273020 255280 273072 255289
rect 242568 255255 242620 255264
rect 242568 255221 242577 255255
rect 242577 255221 242611 255255
rect 242611 255221 242620 255255
rect 242568 255212 242620 255221
rect 275688 255212 275740 255264
rect 246616 254124 246668 254176
rect 308992 253920 309044 253972
rect 371920 253920 371972 253972
rect 372104 253920 372156 253972
rect 273020 253895 273072 253904
rect 273020 253861 273029 253895
rect 273029 253861 273063 253895
rect 273063 253861 273072 253895
rect 273020 253852 273072 253861
rect 309084 253852 309136 253904
rect 328312 253895 328364 253904
rect 328312 253861 328321 253895
rect 328321 253861 328355 253895
rect 328355 253861 328364 253895
rect 328312 253852 328364 253861
rect 235576 253827 235628 253836
rect 235576 253793 235585 253827
rect 235585 253793 235619 253827
rect 235619 253793 235628 253827
rect 235576 253784 235628 253793
rect 302368 253172 302420 253224
rect 349656 253172 349708 253224
rect 350852 253172 350904 253224
rect 581496 253172 581548 253224
rect 278816 251200 278868 251252
rect 285348 251200 285400 251252
rect 285716 251200 285768 251252
rect 331256 251243 331308 251252
rect 331256 251209 331265 251243
rect 331265 251209 331299 251243
rect 331299 251209 331308 251243
rect 331256 251200 331308 251209
rect 341192 251200 341244 251252
rect 91504 251175 91556 251184
rect 91504 251141 91513 251175
rect 91513 251141 91547 251175
rect 91547 251141 91556 251175
rect 91504 251132 91556 251141
rect 225364 251175 225416 251184
rect 225364 251141 225373 251175
rect 225373 251141 225407 251175
rect 225407 251141 225416 251175
rect 225364 251132 225416 251141
rect 229964 251175 230016 251184
rect 229964 251141 229973 251175
rect 229973 251141 230007 251175
rect 230007 251141 230016 251175
rect 229964 251132 230016 251141
rect 357936 251175 357988 251184
rect 357936 251141 357945 251175
rect 357945 251141 357979 251175
rect 357979 251141 357988 251175
rect 553896 251175 553948 251184
rect 357936 251132 357988 251141
rect 553896 251141 553905 251175
rect 553905 251141 553939 251175
rect 553939 251141 553948 251175
rect 553896 251132 553948 251141
rect 278816 251064 278868 251116
rect 135480 249772 135532 249824
rect 135664 249772 135716 249824
rect 152040 249772 152092 249824
rect 152224 249772 152276 249824
rect 170164 249772 170216 249824
rect 170348 249772 170400 249824
rect 190680 249772 190732 249824
rect 190864 249772 190916 249824
rect 214324 249772 214376 249824
rect 214508 249772 214560 249824
rect 246524 249815 246576 249824
rect 246524 249781 246533 249815
rect 246533 249781 246567 249815
rect 246567 249781 246576 249815
rect 246524 249772 246576 249781
rect 305128 249772 305180 249824
rect 372932 249772 372984 249824
rect 373116 249772 373168 249824
rect 385536 249772 385588 249824
rect 385720 249772 385772 249824
rect 392436 249772 392488 249824
rect 392620 249772 392672 249824
rect 528872 249772 528924 249824
rect 529056 249772 529108 249824
rect 535956 249772 536008 249824
rect 536140 249772 536192 249824
rect 571836 249772 571888 249824
rect 572020 249772 572072 249824
rect 242752 246823 242804 246832
rect 242752 246789 242761 246823
rect 242761 246789 242795 246823
rect 242795 246789 242804 246823
rect 242752 246780 242804 246789
rect 242660 245624 242712 245676
rect 275596 245667 275648 245676
rect 275596 245633 275605 245667
rect 275605 245633 275639 245667
rect 275639 245633 275648 245667
rect 275596 245624 275648 245633
rect 239256 244332 239308 244384
rect 239440 244332 239492 244384
rect 285348 244375 285400 244384
rect 285348 244341 285357 244375
rect 285357 244341 285391 244375
rect 285391 244341 285400 244375
rect 285348 244332 285400 244341
rect 3828 244128 3880 244180
rect 228860 244128 228912 244180
rect 229964 244171 230016 244180
rect 229964 244137 229973 244171
rect 229973 244137 230007 244171
rect 230007 244137 230016 244171
rect 229964 244128 230016 244137
rect 239256 244128 239308 244180
rect 239440 244128 239492 244180
rect 285348 244171 285400 244180
rect 285348 244137 285357 244171
rect 285357 244137 285391 244171
rect 285391 244137 285400 244171
rect 285348 244128 285400 244137
rect 328312 243448 328364 243500
rect 328404 243448 328456 243500
rect 242752 241995 242804 242004
rect 242752 241961 242761 241995
rect 242761 241961 242795 241995
rect 242795 241961 242804 241995
rect 242752 241952 242804 241961
rect 251676 241748 251728 241800
rect 261152 241748 261204 241800
rect 91504 241655 91556 241664
rect 91504 241621 91513 241655
rect 91513 241621 91547 241655
rect 91547 241621 91556 241655
rect 91504 241612 91556 241621
rect 225364 241655 225416 241664
rect 225364 241621 225373 241655
rect 225373 241621 225407 241655
rect 225407 241621 225416 241655
rect 225364 241612 225416 241621
rect 290316 241612 290368 241664
rect 294824 241612 294876 241664
rect 357936 241655 357988 241664
rect 357936 241621 357945 241655
rect 357945 241621 357979 241655
rect 357979 241621 357988 241655
rect 553896 241655 553948 241664
rect 357936 241612 357988 241621
rect 553896 241621 553905 241655
rect 553905 241621 553939 241655
rect 553939 241621 553948 241655
rect 553896 241612 553948 241621
rect 246432 241408 246484 241460
rect 246708 241408 246760 241460
rect 309176 241451 309228 241460
rect 309176 241417 309185 241451
rect 309185 241417 309219 241451
rect 309219 241417 309228 241451
rect 309176 241408 309228 241417
rect 279460 240116 279512 240168
rect 279736 240116 279788 240168
rect 235484 240091 235536 240100
rect 235484 240057 235493 240091
rect 235493 240057 235527 240091
rect 235527 240057 235536 240091
rect 235484 240048 235536 240057
rect 242476 237371 242528 237380
rect 242476 237337 242485 237371
rect 242485 237337 242519 237371
rect 242519 237337 242528 237371
rect 242476 237328 242528 237337
rect 276700 237328 276752 237380
rect 276884 237328 276936 237380
rect 285348 236759 285400 236768
rect 285348 236725 285357 236759
rect 285357 236725 285391 236759
rect 285391 236725 285400 236759
rect 285348 236716 285400 236725
rect 273020 236011 273072 236020
rect 273020 235977 273029 236011
rect 273029 235977 273063 236011
rect 273063 235977 273072 236011
rect 273020 235968 273072 235977
rect 272836 235943 272888 235952
rect 272836 235909 272845 235943
rect 272845 235909 272879 235943
rect 272879 235909 272888 235943
rect 272836 235900 272888 235909
rect 328312 235943 328364 235952
rect 328312 235909 328321 235943
rect 328321 235909 328355 235943
rect 328355 235909 328364 235943
rect 328312 235900 328364 235909
rect 371828 234676 371880 234728
rect 275688 234583 275740 234592
rect 275688 234549 275697 234583
rect 275697 234549 275731 234583
rect 275731 234549 275740 234583
rect 275688 234540 275740 234549
rect 371736 234540 371788 234592
rect 309176 234379 309228 234388
rect 309176 234345 309185 234379
rect 309185 234345 309219 234379
rect 309219 234345 309228 234379
rect 309176 234336 309228 234345
rect 319940 234336 319992 234388
rect 320124 234336 320176 234388
rect 276608 232568 276660 232620
rect 277068 232500 277120 232552
rect 277252 232500 277304 232552
rect 285348 231931 285400 231940
rect 285348 231897 285357 231931
rect 285357 231897 285391 231931
rect 285391 231897 285400 231931
rect 285348 231888 285400 231897
rect 242108 231820 242160 231872
rect 242200 231820 242252 231872
rect 246616 231820 246668 231872
rect 246708 231820 246760 231872
rect 285716 231820 285768 231872
rect 285808 231820 285860 231872
rect 331072 231820 331124 231872
rect 331256 231820 331308 231872
rect 341008 231820 341060 231872
rect 341100 231820 341152 231872
rect 272928 231548 272980 231600
rect 135480 230460 135532 230512
rect 135664 230460 135716 230512
rect 152040 230460 152092 230512
rect 152224 230460 152276 230512
rect 170164 230460 170216 230512
rect 170348 230460 170400 230512
rect 190680 230460 190732 230512
rect 190864 230460 190916 230512
rect 214324 230460 214376 230512
rect 214508 230460 214560 230512
rect 235668 230460 235720 230512
rect 385536 230460 385588 230512
rect 385720 230460 385772 230512
rect 392436 230460 392488 230512
rect 392620 230460 392672 230512
rect 528872 230460 528924 230512
rect 529056 230460 529108 230512
rect 535956 230460 536008 230512
rect 536140 230460 536192 230512
rect 552332 230460 552384 230512
rect 552424 230460 552476 230512
rect 571836 230460 571888 230512
rect 572020 230460 572072 230512
rect 242844 227740 242896 227792
rect 276516 227783 276568 227792
rect 276516 227749 276525 227783
rect 276525 227749 276559 227783
rect 276559 227749 276568 227783
rect 276516 227740 276568 227749
rect 268696 227035 268748 227044
rect 268696 227001 268705 227035
rect 268705 227001 268739 227035
rect 268739 227001 268748 227035
rect 268696 226992 268748 227001
rect 300436 226584 300488 226636
rect 308164 226584 308216 226636
rect 360604 226516 360656 226568
rect 362260 226516 362312 226568
rect 239256 225632 239308 225684
rect 239440 225632 239492 225684
rect 229780 224952 229832 225004
rect 229964 224952 230016 225004
rect 275688 224995 275740 225004
rect 275688 224961 275697 224995
rect 275697 224961 275731 224995
rect 275731 224961 275740 224995
rect 275688 224952 275740 224961
rect 285348 224952 285400 225004
rect 285532 224952 285584 225004
rect 285716 224952 285768 225004
rect 304944 224952 304996 225004
rect 320032 224995 320084 225004
rect 320032 224961 320041 224995
rect 320041 224961 320075 224995
rect 320075 224961 320084 224995
rect 320032 224952 320084 224961
rect 271364 224884 271416 224936
rect 271548 224884 271600 224936
rect 272928 224927 272980 224936
rect 272928 224893 272937 224927
rect 272937 224893 272971 224927
rect 272971 224893 272980 224927
rect 272928 224884 272980 224893
rect 341100 225020 341152 225072
rect 341008 224884 341060 224936
rect 275688 224816 275740 224868
rect 304944 224816 304996 224868
rect 239348 222232 239400 222284
rect 91320 222164 91372 222216
rect 91504 222164 91556 222216
rect 242200 222232 242252 222284
rect 246616 222232 246668 222284
rect 246800 222164 246852 222216
rect 268788 222164 268840 222216
rect 276700 222164 276752 222216
rect 276884 222164 276936 222216
rect 357936 222164 357988 222216
rect 358120 222164 358172 222216
rect 371552 222164 371604 222216
rect 371828 222164 371880 222216
rect 553712 222164 553764 222216
rect 553896 222164 553948 222216
rect 239348 222096 239400 222148
rect 242108 222096 242160 222148
rect 246524 222096 246576 222148
rect 246800 222028 246852 222080
rect 320032 220983 320084 220992
rect 320032 220949 320041 220983
rect 320041 220949 320075 220983
rect 320075 220949 320084 220983
rect 320032 220940 320084 220949
rect 276700 220779 276752 220788
rect 276700 220745 276709 220779
rect 276709 220745 276743 220779
rect 276743 220745 276752 220779
rect 276700 220736 276752 220745
rect 341008 220779 341060 220788
rect 341008 220745 341017 220779
rect 341017 220745 341051 220779
rect 341051 220745 341060 220779
rect 341008 220736 341060 220745
rect 373208 220779 373260 220788
rect 373208 220745 373217 220779
rect 373217 220745 373251 220779
rect 373251 220745 373260 220779
rect 373208 220736 373260 220745
rect 279736 219444 279788 219496
rect 279828 219444 279880 219496
rect 285256 219487 285308 219496
rect 285256 219453 285265 219487
rect 285265 219453 285299 219487
rect 285299 219453 285308 219487
rect 285256 219444 285308 219453
rect 272928 217991 272980 218000
rect 272928 217957 272937 217991
rect 272937 217957 272971 217991
rect 272971 217957 272980 217991
rect 272928 217948 272980 217957
rect 242476 216631 242528 216640
rect 242476 216597 242485 216631
rect 242485 216597 242519 216631
rect 242519 216597 242528 216631
rect 242476 216588 242528 216597
rect 275596 215339 275648 215348
rect 275596 215305 275605 215339
rect 275605 215305 275639 215339
rect 275639 215305 275648 215339
rect 275596 215296 275648 215305
rect 272836 215271 272888 215280
rect 272836 215237 272845 215271
rect 272845 215237 272879 215271
rect 272879 215237 272888 215271
rect 272836 215228 272888 215237
rect 341100 215228 341152 215280
rect 331072 212508 331124 212560
rect 331256 212508 331308 212560
rect 553712 212508 553764 212560
rect 553896 212508 553948 212560
rect 279736 212440 279788 212492
rect 279828 212440 279880 212492
rect 357936 212483 357988 212492
rect 357936 212449 357945 212483
rect 357945 212449 357979 212483
rect 357979 212449 357988 212483
rect 373208 212483 373260 212492
rect 357936 212440 357988 212449
rect 373208 212449 373217 212483
rect 373217 212449 373251 212483
rect 373251 212449 373260 212483
rect 373208 212440 373260 212449
rect 275596 211259 275648 211268
rect 275596 211225 275605 211259
rect 275605 211225 275639 211259
rect 275639 211225 275648 211259
rect 275596 211216 275648 211225
rect 235392 211148 235444 211200
rect 235484 211148 235536 211200
rect 276700 211191 276752 211200
rect 276700 211157 276709 211191
rect 276709 211157 276743 211191
rect 276743 211157 276752 211191
rect 276700 211148 276752 211157
rect 328312 211191 328364 211200
rect 328312 211157 328321 211191
rect 328321 211157 328355 211191
rect 328355 211157 328364 211191
rect 328312 211148 328364 211157
rect 385536 211148 385588 211200
rect 385720 211148 385772 211200
rect 392436 211148 392488 211200
rect 392620 211148 392672 211200
rect 528872 211148 528924 211200
rect 529056 211148 529108 211200
rect 535956 211148 536008 211200
rect 536140 211148 536192 211200
rect 552332 211148 552384 211200
rect 552516 211148 552568 211200
rect 571836 211148 571888 211200
rect 572020 211148 572072 211200
rect 272836 210443 272888 210452
rect 272836 210409 272845 210443
rect 272845 210409 272879 210443
rect 272879 210409 272888 210443
rect 272836 210400 272888 210409
rect 275596 210443 275648 210452
rect 275596 210409 275605 210443
rect 275605 210409 275639 210443
rect 275639 210409 275648 210443
rect 275596 210400 275648 210409
rect 3736 209720 3788 209772
rect 224720 209720 224772 209772
rect 328404 209763 328456 209772
rect 328404 209729 328413 209763
rect 328413 209729 328447 209763
rect 328447 209729 328456 209763
rect 328404 209720 328456 209729
rect 285256 208564 285308 208616
rect 285256 208428 285308 208480
rect 285256 208224 285308 208276
rect 268696 207723 268748 207732
rect 268696 207689 268705 207723
rect 268705 207689 268739 207723
rect 268739 207689 268748 207723
rect 268696 207680 268748 207689
rect 242476 207043 242528 207052
rect 242476 207009 242485 207043
rect 242485 207009 242519 207043
rect 242519 207009 242528 207043
rect 242476 207000 242528 207009
rect 273020 206932 273072 206984
rect 273112 206864 273164 206916
rect 230056 205776 230108 205828
rect 341192 205776 341244 205828
rect 235484 205751 235536 205760
rect 235484 205717 235493 205751
rect 235493 205717 235527 205751
rect 235527 205717 235536 205751
rect 235484 205708 235536 205717
rect 271456 205751 271508 205760
rect 271456 205717 271465 205751
rect 271465 205717 271499 205751
rect 271499 205717 271508 205751
rect 271456 205708 271508 205717
rect 309084 205751 309136 205760
rect 309084 205717 309093 205751
rect 309093 205717 309127 205751
rect 309127 205717 309136 205751
rect 309084 205708 309136 205717
rect 229964 205547 230016 205556
rect 229964 205513 229973 205547
rect 229973 205513 230007 205547
rect 230007 205513 230016 205547
rect 229964 205504 230016 205513
rect 239256 205504 239308 205556
rect 239440 205504 239492 205556
rect 268788 205504 268840 205556
rect 271456 205547 271508 205556
rect 271456 205513 271465 205547
rect 271465 205513 271499 205547
rect 271499 205513 271508 205547
rect 271456 205504 271508 205513
rect 309084 205547 309136 205556
rect 309084 205513 309093 205547
rect 309093 205513 309127 205547
rect 309127 205513 309136 205547
rect 309084 205504 309136 205513
rect 341100 205547 341152 205556
rect 341100 205513 341109 205547
rect 341109 205513 341143 205547
rect 341143 205513 341152 205547
rect 341100 205504 341152 205513
rect 328404 204935 328456 204944
rect 328404 204901 328413 204935
rect 328413 204901 328447 204935
rect 328447 204901 328456 204935
rect 328404 204892 328456 204901
rect 91320 202988 91372 203040
rect 91504 202988 91556 203040
rect 225364 202988 225416 203040
rect 225548 202988 225600 203040
rect 235484 203031 235536 203040
rect 235484 202997 235493 203031
rect 235493 202997 235527 203031
rect 235527 202997 235536 203031
rect 235484 202988 235536 202997
rect 357936 203031 357988 203040
rect 357936 202997 357945 203031
rect 357945 202997 357979 203031
rect 357979 202997 357988 203031
rect 357936 202988 357988 202997
rect 235576 202827 235628 202836
rect 235576 202793 235585 202827
rect 235585 202793 235619 202827
rect 235619 202793 235628 202827
rect 235576 202784 235628 202793
rect 341100 202827 341152 202836
rect 341100 202793 341109 202827
rect 341109 202793 341143 202827
rect 341143 202793 341152 202827
rect 341100 202784 341152 202793
rect 242476 201492 242528 201544
rect 285624 201492 285676 201544
rect 285716 201492 285768 201544
rect 135480 201424 135532 201476
rect 135664 201424 135716 201476
rect 152040 201424 152092 201476
rect 152224 201424 152276 201476
rect 170164 201424 170216 201476
rect 170348 201424 170400 201476
rect 190680 201424 190732 201476
rect 190864 201424 190916 201476
rect 214324 201424 214376 201476
rect 214508 201424 214560 201476
rect 268512 201424 268564 201476
rect 268788 201424 268840 201476
rect 385536 201424 385588 201476
rect 385720 201424 385772 201476
rect 392436 201424 392488 201476
rect 392620 201424 392672 201476
rect 528872 201424 528924 201476
rect 529056 201424 529108 201476
rect 535956 201424 536008 201476
rect 536140 201424 536192 201476
rect 552424 201467 552476 201476
rect 552424 201433 552433 201467
rect 552433 201433 552467 201467
rect 552467 201433 552476 201467
rect 552424 201424 552476 201433
rect 571836 201424 571888 201476
rect 572020 201424 572072 201476
rect 242568 201356 242620 201408
rect 279828 200107 279880 200116
rect 279828 200073 279837 200107
rect 279837 200073 279871 200107
rect 279871 200073 279880 200107
rect 279828 200064 279880 200073
rect 320032 200107 320084 200116
rect 320032 200073 320041 200107
rect 320041 200073 320075 200107
rect 320075 200073 320084 200107
rect 320032 200064 320084 200073
rect 372012 200107 372064 200116
rect 372012 200073 372021 200107
rect 372021 200073 372055 200107
rect 372055 200073 372064 200107
rect 372012 200064 372064 200073
rect 373116 200064 373168 200116
rect 328404 200039 328456 200048
rect 328404 200005 328413 200039
rect 328413 200005 328447 200039
rect 328447 200005 328456 200039
rect 328404 199996 328456 200005
rect 285072 198747 285124 198756
rect 285072 198713 285081 198747
rect 285081 198713 285115 198747
rect 285115 198713 285124 198747
rect 285072 198704 285124 198713
rect 242568 198636 242620 198688
rect 276976 198135 277028 198144
rect 276976 198101 276985 198135
rect 276985 198101 277019 198135
rect 277019 198101 277028 198135
rect 276976 198092 277028 198101
rect 275596 197548 275648 197600
rect 275688 197387 275740 197396
rect 275688 197353 275697 197387
rect 275697 197353 275731 197387
rect 275731 197353 275740 197387
rect 275688 197344 275740 197353
rect 552424 196299 552476 196308
rect 552424 196265 552433 196299
rect 552433 196265 552467 196299
rect 552467 196265 552476 196299
rect 552424 196256 552476 196265
rect 320032 195959 320084 195968
rect 320032 195925 320041 195959
rect 320041 195925 320075 195959
rect 320075 195925 320084 195959
rect 320032 195916 320084 195925
rect 353060 195916 353112 195968
rect 580668 195916 580720 195968
rect 235576 195755 235628 195764
rect 235576 195721 235585 195755
rect 235585 195721 235619 195755
rect 235619 195721 235628 195755
rect 235576 195712 235628 195721
rect 328404 195755 328456 195764
rect 328404 195721 328413 195755
rect 328413 195721 328447 195755
rect 328447 195721 328456 195755
rect 328404 195712 328456 195721
rect 246708 193876 246760 193928
rect 246984 193876 247036 193928
rect 341192 193332 341244 193384
rect 331072 193196 331124 193248
rect 331256 193196 331308 193248
rect 553712 193196 553764 193248
rect 553896 193196 553948 193248
rect 3828 192652 3880 192704
rect 9440 192652 9492 192704
rect 235576 191768 235628 191820
rect 235760 191768 235812 191820
rect 552424 191811 552476 191820
rect 552424 191777 552433 191811
rect 552433 191777 552467 191811
rect 552467 191777 552476 191811
rect 552424 191768 552476 191777
rect 372012 191267 372064 191276
rect 372012 191233 372021 191267
rect 372021 191233 372055 191267
rect 372055 191233 372064 191267
rect 372012 191224 372064 191233
rect 373024 190587 373076 190596
rect 373024 190553 373033 190587
rect 373033 190553 373067 190587
rect 373067 190553 373076 190587
rect 373024 190544 373076 190553
rect 279828 190519 279880 190528
rect 279828 190485 279837 190519
rect 279837 190485 279871 190519
rect 279871 190485 279880 190519
rect 279828 190476 279880 190485
rect 242476 189091 242528 189100
rect 242476 189057 242485 189091
rect 242485 189057 242519 189091
rect 242519 189057 242528 189091
rect 242476 189048 242528 189057
rect 246432 189048 246484 189100
rect 246616 189048 246668 189100
rect 272928 189048 272980 189100
rect 276976 189091 277028 189100
rect 276976 189057 276985 189091
rect 276985 189057 277019 189091
rect 277019 189057 277028 189091
rect 276976 189048 277028 189057
rect 242844 189023 242896 189032
rect 242844 188989 242853 189023
rect 242853 188989 242887 189023
rect 242887 188989 242896 189023
rect 242844 188980 242896 188989
rect 272928 188912 272980 188964
rect 229780 186328 229832 186380
rect 229964 186328 230016 186380
rect 285532 186328 285584 186380
rect 305036 186328 305088 186380
rect 305220 186328 305272 186380
rect 309084 186328 309136 186380
rect 341100 186371 341152 186380
rect 341100 186337 341109 186371
rect 341109 186337 341143 186371
rect 341143 186337 341152 186371
rect 341100 186328 341152 186337
rect 285072 186260 285124 186312
rect 285256 186260 285308 186312
rect 285624 186192 285676 186244
rect 91320 183540 91372 183592
rect 91504 183540 91556 183592
rect 279828 183608 279880 183660
rect 341100 183651 341152 183660
rect 341100 183617 341109 183651
rect 341109 183617 341143 183651
rect 341143 183617 341152 183651
rect 341100 183608 341152 183617
rect 308992 183583 309044 183592
rect 308992 183549 309001 183583
rect 309001 183549 309035 183583
rect 309035 183549 309044 183583
rect 308992 183540 309044 183549
rect 357936 183540 357988 183592
rect 358120 183540 358172 183592
rect 553712 183540 553764 183592
rect 553896 183540 553948 183592
rect 279736 183472 279788 183524
rect 341100 183472 341152 183524
rect 341468 183472 341520 183524
rect 552424 183515 552476 183524
rect 552424 183481 552433 183515
rect 552433 183481 552467 183515
rect 552467 183481 552476 183515
rect 552424 183472 552476 183481
rect 135480 182112 135532 182164
rect 135664 182112 135716 182164
rect 152040 182112 152092 182164
rect 152224 182112 152276 182164
rect 170164 182112 170216 182164
rect 170348 182112 170400 182164
rect 190680 182112 190732 182164
rect 190864 182112 190916 182164
rect 214324 182112 214376 182164
rect 214508 182112 214560 182164
rect 229872 182155 229924 182164
rect 229872 182121 229881 182155
rect 229881 182121 229915 182155
rect 229915 182121 229924 182155
rect 229872 182112 229924 182121
rect 242108 182112 242160 182164
rect 242200 182112 242252 182164
rect 246524 182112 246576 182164
rect 246616 182112 246668 182164
rect 285164 182155 285216 182164
rect 285164 182121 285173 182155
rect 285173 182121 285207 182155
rect 285207 182121 285216 182155
rect 285164 182112 285216 182121
rect 285624 182112 285676 182164
rect 285716 182112 285768 182164
rect 328312 182155 328364 182164
rect 328312 182121 328321 182155
rect 328321 182121 328355 182155
rect 328355 182121 328364 182155
rect 328312 182112 328364 182121
rect 385536 182112 385588 182164
rect 385720 182112 385772 182164
rect 392436 182112 392488 182164
rect 392620 182112 392672 182164
rect 528872 182112 528924 182164
rect 529056 182112 529108 182164
rect 535956 182112 536008 182164
rect 536140 182112 536192 182164
rect 571836 182112 571888 182164
rect 572020 182112 572072 182164
rect 242844 182019 242896 182028
rect 242844 181985 242853 182019
rect 242853 181985 242887 182019
rect 242887 181985 242896 182019
rect 242844 181976 242896 181985
rect 295192 181432 295244 181484
rect 308256 181432 308308 181484
rect 273020 180752 273072 180804
rect 273112 180752 273164 180804
rect 278816 180795 278868 180804
rect 278816 180761 278825 180795
rect 278825 180761 278859 180795
rect 278859 180761 278868 180795
rect 278816 180752 278868 180761
rect 371920 180752 371972 180804
rect 372012 180752 372064 180804
rect 251676 179392 251728 179444
rect 259864 179392 259916 179444
rect 371920 179367 371972 179376
rect 371920 179333 371929 179367
rect 371929 179333 371963 179367
rect 371963 179333 371972 179367
rect 371920 179324 371972 179333
rect 304852 178712 304904 178764
rect 305128 178712 305180 178764
rect 319756 177216 319808 177268
rect 320032 177216 320084 177268
rect 235484 176672 235536 176724
rect 229872 176579 229924 176588
rect 229872 176545 229881 176579
rect 229881 176545 229915 176579
rect 229915 176545 229924 176579
rect 229872 176536 229924 176545
rect 235576 176536 235628 176588
rect 328404 176536 328456 176588
rect 268512 173884 268564 173936
rect 268696 173884 268748 173936
rect 308992 173884 309044 173936
rect 309084 173884 309136 173936
rect 331072 173884 331124 173936
rect 331256 173884 331308 173936
rect 275596 173247 275648 173256
rect 275596 173213 275605 173247
rect 275605 173213 275639 173247
rect 275639 173213 275648 173247
rect 275596 173204 275648 173213
rect 285164 172567 285216 172576
rect 285164 172533 285173 172567
rect 285173 172533 285207 172567
rect 285207 172533 285216 172567
rect 285164 172524 285216 172533
rect 278816 171139 278868 171148
rect 278816 171105 278825 171139
rect 278825 171105 278859 171139
rect 278859 171105 278868 171139
rect 278816 171096 278868 171105
rect 246984 169260 247036 169312
rect 273112 168308 273164 168360
rect 235576 167152 235628 167204
rect 239256 167084 239308 167136
rect 239440 167084 239492 167136
rect 235484 166923 235536 166932
rect 235484 166889 235493 166923
rect 235493 166889 235527 166923
rect 235527 166889 235536 166923
rect 235484 166880 235536 166889
rect 239256 166880 239308 166932
rect 239440 166880 239492 166932
rect 285716 166812 285768 166864
rect 285716 166676 285768 166728
rect 272928 166268 272980 166320
rect 272836 166200 272888 166252
rect 284796 164364 284848 164416
rect 285624 164364 285676 164416
rect 382040 164364 382092 164416
rect 385812 164364 385864 164416
rect 391700 164364 391752 164416
rect 392712 164364 392764 164416
rect 526940 164364 526992 164416
rect 529332 164364 529384 164416
rect 535680 164364 535732 164416
rect 536600 164364 536652 164416
rect 552516 164364 552568 164416
rect 552700 164364 552752 164416
rect 571560 164364 571612 164416
rect 572112 164364 572164 164416
rect 242108 164160 242160 164212
rect 242660 164203 242712 164212
rect 242660 164169 242669 164203
rect 242669 164169 242703 164203
rect 242703 164169 242712 164203
rect 242660 164160 242712 164169
rect 246524 164160 246576 164212
rect 259312 164203 259364 164212
rect 259312 164169 259321 164203
rect 259321 164169 259355 164203
rect 259355 164169 259364 164203
rect 259312 164160 259364 164169
rect 305128 164203 305180 164212
rect 305128 164169 305137 164203
rect 305137 164169 305171 164203
rect 305171 164169 305180 164203
rect 305128 164160 305180 164169
rect 308992 164160 309044 164212
rect 309084 164160 309136 164212
rect 331072 164160 331124 164212
rect 331256 164160 331308 164212
rect 341008 164160 341060 164212
rect 341100 164160 341152 164212
rect 553896 164203 553948 164212
rect 553896 164169 553905 164203
rect 553905 164169 553939 164203
rect 553939 164169 553948 164203
rect 553896 164160 553948 164169
rect 242200 164092 242252 164144
rect 246616 164092 246668 164144
rect 320032 164092 320084 164144
rect 320124 164092 320176 164144
rect 273020 163523 273072 163532
rect 273020 163489 273029 163523
rect 273029 163489 273063 163523
rect 273063 163489 273072 163523
rect 273020 163480 273072 163489
rect 275596 163523 275648 163532
rect 275596 163489 275605 163523
rect 275605 163489 275639 163523
rect 275639 163489 275648 163523
rect 275596 163480 275648 163489
rect 135664 162843 135716 162852
rect 135664 162809 135673 162843
rect 135673 162809 135707 162843
rect 135707 162809 135716 162843
rect 135664 162800 135716 162809
rect 152224 162843 152276 162852
rect 152224 162809 152233 162843
rect 152233 162809 152267 162843
rect 152267 162809 152276 162843
rect 152224 162800 152276 162809
rect 170164 162843 170216 162852
rect 170164 162809 170173 162843
rect 170173 162809 170207 162843
rect 170207 162809 170216 162843
rect 170164 162800 170216 162809
rect 190864 162843 190916 162852
rect 190864 162809 190873 162843
rect 190873 162809 190907 162843
rect 190907 162809 190916 162843
rect 190864 162800 190916 162809
rect 214324 162843 214376 162852
rect 214324 162809 214333 162843
rect 214333 162809 214367 162843
rect 214367 162809 214376 162843
rect 214324 162800 214376 162809
rect 230056 162843 230108 162852
rect 230056 162809 230065 162843
rect 230065 162809 230099 162843
rect 230099 162809 230108 162843
rect 230056 162800 230108 162809
rect 242016 162800 242068 162852
rect 242200 162800 242252 162852
rect 242568 162868 242620 162920
rect 246616 162843 246668 162852
rect 246616 162809 246625 162843
rect 246625 162809 246659 162843
rect 246659 162809 246668 162843
rect 246616 162800 246668 162809
rect 385536 162843 385588 162852
rect 385536 162809 385545 162843
rect 385545 162809 385579 162843
rect 385579 162809 385588 162843
rect 392436 162843 392488 162852
rect 385536 162800 385588 162809
rect 392436 162809 392445 162843
rect 392445 162809 392479 162843
rect 392479 162809 392488 162843
rect 392436 162800 392488 162809
rect 529056 162843 529108 162852
rect 529056 162809 529065 162843
rect 529065 162809 529099 162843
rect 529099 162809 529108 162843
rect 529056 162800 529108 162809
rect 535956 162843 536008 162852
rect 535956 162809 535965 162843
rect 535965 162809 535999 162843
rect 535999 162809 536008 162843
rect 535956 162800 536008 162809
rect 552516 162843 552568 162852
rect 552516 162809 552525 162843
rect 552525 162809 552559 162843
rect 552559 162809 552568 162843
rect 552516 162800 552568 162809
rect 571836 162843 571888 162852
rect 571836 162809 571845 162843
rect 571845 162809 571879 162843
rect 571879 162809 571888 162843
rect 571836 162800 571888 162809
rect 246892 161483 246944 161492
rect 246892 161449 246901 161483
rect 246901 161449 246935 161483
rect 246935 161449 246944 161483
rect 246892 161440 246944 161449
rect 285256 161440 285308 161492
rect 285348 161440 285400 161492
rect 372012 161440 372064 161492
rect 268512 161279 268564 161288
rect 268512 161245 268521 161279
rect 268521 161245 268555 161279
rect 268555 161245 268564 161279
rect 268512 161236 268564 161245
rect 246892 159468 246944 159520
rect 235484 159307 235536 159316
rect 235484 159273 235493 159307
rect 235493 159273 235527 159307
rect 235527 159273 235536 159307
rect 235484 159264 235536 159273
rect 273020 158652 273072 158704
rect 273112 158652 273164 158704
rect 319848 157972 319900 158024
rect 320124 157972 320176 158024
rect 242476 157947 242528 157956
rect 242476 157913 242485 157947
rect 242485 157913 242519 157947
rect 242519 157913 242528 157947
rect 242476 157904 242528 157913
rect 285348 157360 285400 157412
rect 259312 157335 259364 157344
rect 259312 157301 259321 157335
rect 259321 157301 259355 157335
rect 259355 157301 259364 157335
rect 259312 157292 259364 157301
rect 273112 157292 273164 157344
rect 275596 157335 275648 157344
rect 275596 157301 275605 157335
rect 275605 157301 275639 157335
rect 275639 157301 275648 157335
rect 275596 157292 275648 157301
rect 305128 157335 305180 157344
rect 305128 157301 305137 157335
rect 305137 157301 305171 157335
rect 305171 157301 305180 157335
rect 305128 157292 305180 157301
rect 230056 157131 230108 157140
rect 230056 157097 230065 157131
rect 230065 157097 230099 157131
rect 230099 157097 230108 157131
rect 230056 157088 230108 157097
rect 235576 157088 235628 157140
rect 242660 157131 242712 157140
rect 242660 157097 242669 157131
rect 242669 157097 242703 157131
rect 242703 157097 242712 157131
rect 242660 157088 242712 157097
rect 246800 157131 246852 157140
rect 246800 157097 246809 157131
rect 246809 157097 246843 157131
rect 246843 157097 246852 157131
rect 246800 157088 246852 157097
rect 268696 157088 268748 157140
rect 285164 156748 285216 156800
rect 553896 154683 553948 154692
rect 553896 154649 553905 154683
rect 553905 154649 553939 154683
rect 553939 154649 553948 154683
rect 553896 154640 553948 154649
rect 268696 154411 268748 154420
rect 268696 154377 268705 154411
rect 268705 154377 268739 154411
rect 268739 154377 268748 154411
rect 268696 154368 268748 154377
rect 135664 153255 135716 153264
rect 135664 153221 135673 153255
rect 135673 153221 135707 153255
rect 135707 153221 135716 153255
rect 135664 153212 135716 153221
rect 152224 153255 152276 153264
rect 152224 153221 152233 153255
rect 152233 153221 152267 153255
rect 152267 153221 152276 153255
rect 152224 153212 152276 153221
rect 170164 153255 170216 153264
rect 170164 153221 170173 153255
rect 170173 153221 170207 153255
rect 170207 153221 170216 153255
rect 170164 153212 170216 153221
rect 190864 153255 190916 153264
rect 190864 153221 190873 153255
rect 190873 153221 190907 153255
rect 190907 153221 190916 153255
rect 190864 153212 190916 153221
rect 214324 153255 214376 153264
rect 214324 153221 214333 153255
rect 214333 153221 214367 153255
rect 214367 153221 214376 153255
rect 214324 153212 214376 153221
rect 246616 153255 246668 153264
rect 246616 153221 246625 153255
rect 246625 153221 246659 153255
rect 246659 153221 246668 153255
rect 246616 153212 246668 153221
rect 372012 153212 372064 153264
rect 385536 153255 385588 153264
rect 385536 153221 385545 153255
rect 385545 153221 385579 153255
rect 385579 153221 385588 153255
rect 392436 153255 392488 153264
rect 385536 153212 385588 153221
rect 392436 153221 392445 153255
rect 392445 153221 392479 153255
rect 392479 153221 392488 153255
rect 392436 153212 392488 153221
rect 529056 153255 529108 153264
rect 529056 153221 529065 153255
rect 529065 153221 529099 153255
rect 529099 153221 529108 153255
rect 529056 153212 529108 153221
rect 535956 153255 536008 153264
rect 535956 153221 535965 153255
rect 535965 153221 535999 153255
rect 535999 153221 536008 153255
rect 535956 153212 536008 153221
rect 552516 153255 552568 153264
rect 552516 153221 552525 153255
rect 552525 153221 552559 153255
rect 552559 153221 552568 153255
rect 552516 153212 552568 153221
rect 571836 153255 571888 153264
rect 571836 153221 571845 153255
rect 571845 153221 571879 153255
rect 571879 153221 571888 153255
rect 571836 153212 571888 153221
rect 371920 153144 371972 153196
rect 373116 153187 373168 153196
rect 373116 153153 373125 153187
rect 373125 153153 373159 153187
rect 373159 153153 373168 153187
rect 373116 153144 373168 153153
rect 278724 149855 278776 149864
rect 278724 149821 278733 149855
rect 278733 149821 278767 149855
rect 278767 149821 278776 149855
rect 278724 149812 278776 149821
rect 271456 149132 271508 149184
rect 271548 149132 271600 149184
rect 351680 148928 351732 148980
rect 580392 148928 580444 148980
rect 246616 147704 246668 147756
rect 273020 147679 273072 147688
rect 273020 147645 273029 147679
rect 273029 147645 273063 147679
rect 273063 147645 273072 147679
rect 273020 147636 273072 147645
rect 275688 147636 275740 147688
rect 285532 147636 285584 147688
rect 285716 147636 285768 147688
rect 305036 147636 305088 147688
rect 305220 147636 305272 147688
rect 341192 147704 341244 147756
rect 246524 147568 246576 147620
rect 268696 147611 268748 147620
rect 268696 147577 268705 147611
rect 268705 147577 268739 147611
rect 268739 147577 268748 147611
rect 268696 147568 268748 147577
rect 341100 147568 341152 147620
rect 373116 145163 373168 145172
rect 373116 145129 373125 145163
rect 373125 145129 373159 145163
rect 373159 145129 373168 145163
rect 373116 145120 373168 145129
rect 320032 144984 320084 145036
rect 320124 144984 320176 145036
rect 328312 144984 328364 145036
rect 328404 144984 328456 145036
rect 225364 144891 225416 144900
rect 225364 144857 225373 144891
rect 225373 144857 225407 144891
rect 225407 144857 225416 144891
rect 225364 144848 225416 144857
rect 242108 144848 242160 144900
rect 242200 144848 242252 144900
rect 285624 144891 285676 144900
rect 285624 144857 285633 144891
rect 285633 144857 285667 144891
rect 285667 144857 285676 144891
rect 285624 144848 285676 144857
rect 331072 144848 331124 144900
rect 331256 144848 331308 144900
rect 341008 144848 341060 144900
rect 341100 144848 341152 144900
rect 553896 144891 553948 144900
rect 553896 144857 553905 144891
rect 553905 144857 553939 144891
rect 553939 144857 553948 144891
rect 553896 144848 553948 144857
rect 242660 144780 242712 144832
rect 242752 144780 242804 144832
rect 273020 143735 273072 143744
rect 273020 143701 273029 143735
rect 273029 143701 273063 143735
rect 273063 143701 273072 143735
rect 273020 143692 273072 143701
rect 4012 143488 4064 143540
rect 227480 143488 227532 143540
rect 242016 143488 242068 143540
rect 242200 143488 242252 143540
rect 242476 143488 242528 143540
rect 242568 143488 242620 143540
rect 276700 143488 276752 143540
rect 276884 143488 276936 143540
rect 320124 143488 320176 143540
rect 328404 143531 328456 143540
rect 328404 143497 328413 143531
rect 328413 143497 328447 143531
rect 328447 143497 328456 143531
rect 328404 143488 328456 143497
rect 373024 143488 373076 143540
rect 373116 143488 373168 143540
rect 385536 143531 385588 143540
rect 385536 143497 385545 143531
rect 385545 143497 385579 143531
rect 385579 143497 385588 143531
rect 392436 143531 392488 143540
rect 385536 143488 385588 143497
rect 392436 143497 392445 143531
rect 392445 143497 392479 143531
rect 392479 143497 392488 143531
rect 392436 143488 392488 143497
rect 529056 143531 529108 143540
rect 529056 143497 529065 143531
rect 529065 143497 529099 143531
rect 529099 143497 529108 143531
rect 529056 143488 529108 143497
rect 535956 143531 536008 143540
rect 535956 143497 535965 143531
rect 535965 143497 535999 143531
rect 535999 143497 536008 143531
rect 535956 143488 536008 143497
rect 552516 143488 552568 143540
rect 571836 143531 571888 143540
rect 571836 143497 571845 143531
rect 571845 143497 571879 143531
rect 571879 143497 571888 143531
rect 571836 143488 571888 143497
rect 135664 143463 135716 143472
rect 135664 143429 135673 143463
rect 135673 143429 135707 143463
rect 135707 143429 135716 143463
rect 135664 143420 135716 143429
rect 152224 143463 152276 143472
rect 152224 143429 152233 143463
rect 152233 143429 152267 143463
rect 152267 143429 152276 143463
rect 152224 143420 152276 143429
rect 170164 143463 170216 143472
rect 170164 143429 170173 143463
rect 170173 143429 170207 143463
rect 170207 143429 170216 143463
rect 170164 143420 170216 143429
rect 190864 143463 190916 143472
rect 190864 143429 190873 143463
rect 190873 143429 190907 143463
rect 190907 143429 190916 143463
rect 190864 143420 190916 143429
rect 214324 143463 214376 143472
rect 214324 143429 214333 143463
rect 214333 143429 214367 143463
rect 214367 143429 214376 143463
rect 214324 143420 214376 143429
rect 278816 142128 278868 142180
rect 309084 140743 309136 140752
rect 309084 140709 309093 140743
rect 309093 140709 309127 140743
rect 309127 140709 309136 140743
rect 309084 140700 309136 140709
rect 275504 139544 275556 139596
rect 275688 139544 275740 139596
rect 271456 139408 271508 139460
rect 271548 139408 271600 139460
rect 273020 139451 273072 139460
rect 273020 139417 273029 139451
rect 273029 139417 273063 139451
rect 273063 139417 273072 139451
rect 273020 139408 273072 139417
rect 279736 139383 279788 139392
rect 279736 139349 279745 139383
rect 279745 139349 279779 139383
rect 279779 139349 279788 139383
rect 279736 139340 279788 139349
rect 229872 137980 229924 138032
rect 235484 137980 235536 138032
rect 229780 137912 229832 137964
rect 246892 138048 246944 138100
rect 285348 138048 285400 138100
rect 259312 137980 259364 138032
rect 235576 137912 235628 137964
rect 246800 137912 246852 137964
rect 268788 137980 268840 138032
rect 305036 137980 305088 138032
rect 371828 137980 371880 138032
rect 268696 137912 268748 137964
rect 271456 137955 271508 137964
rect 271456 137921 271465 137955
rect 271465 137921 271499 137955
rect 271499 137921 271508 137955
rect 271456 137912 271508 137921
rect 285624 137955 285676 137964
rect 285624 137921 285633 137955
rect 285633 137921 285667 137955
rect 285667 137921 285676 137955
rect 285624 137912 285676 137921
rect 305128 137912 305180 137964
rect 371920 137912 371972 137964
rect 285164 137844 285216 137896
rect 259404 137776 259456 137828
rect 285440 135575 285492 135584
rect 285440 135541 285449 135575
rect 285449 135541 285483 135575
rect 285483 135541 285492 135575
rect 285440 135532 285492 135541
rect 225364 135371 225416 135380
rect 225364 135337 225373 135371
rect 225373 135337 225407 135371
rect 225407 135337 225416 135371
rect 225364 135328 225416 135337
rect 553896 135371 553948 135380
rect 553896 135337 553905 135371
rect 553905 135337 553939 135371
rect 553939 135337 553948 135371
rect 553896 135328 553948 135337
rect 246524 135260 246576 135312
rect 285532 135260 285584 135312
rect 91320 135192 91372 135244
rect 91504 135192 91556 135244
rect 235576 135192 235628 135244
rect 235760 135192 235812 135244
rect 259404 135235 259456 135244
rect 259404 135201 259413 135235
rect 259413 135201 259447 135235
rect 259447 135201 259456 135235
rect 259404 135192 259456 135201
rect 268696 135235 268748 135244
rect 268696 135201 268705 135235
rect 268705 135201 268739 135235
rect 268739 135201 268748 135235
rect 268696 135192 268748 135201
rect 341192 135192 341244 135244
rect 341376 135192 341428 135244
rect 371920 135235 371972 135244
rect 371920 135201 371929 135235
rect 371929 135201 371963 135235
rect 371963 135201 371972 135235
rect 371920 135192 371972 135201
rect 553712 135192 553764 135244
rect 553896 135192 553948 135244
rect 246524 135124 246576 135176
rect 309084 134691 309136 134700
rect 309084 134657 309093 134691
rect 309093 134657 309127 134691
rect 309127 134657 309136 134691
rect 309084 134648 309136 134657
rect 135664 133943 135716 133952
rect 135664 133909 135673 133943
rect 135673 133909 135707 133943
rect 135707 133909 135716 133943
rect 135664 133900 135716 133909
rect 152224 133943 152276 133952
rect 152224 133909 152233 133943
rect 152233 133909 152267 133943
rect 152267 133909 152276 133943
rect 152224 133900 152276 133909
rect 170164 133943 170216 133952
rect 170164 133909 170173 133943
rect 170173 133909 170207 133943
rect 170207 133909 170216 133943
rect 170164 133900 170216 133909
rect 190864 133943 190916 133952
rect 190864 133909 190873 133943
rect 190873 133909 190907 133943
rect 190907 133909 190916 133943
rect 190864 133900 190916 133909
rect 214324 133943 214376 133952
rect 214324 133909 214333 133943
rect 214333 133909 214367 133943
rect 214367 133909 214376 133943
rect 214324 133900 214376 133909
rect 319940 133943 319992 133952
rect 319940 133909 319949 133943
rect 319949 133909 319983 133943
rect 319983 133909 319992 133943
rect 319940 133900 319992 133909
rect 328404 133943 328456 133952
rect 328404 133909 328413 133943
rect 328413 133909 328447 133943
rect 328447 133909 328456 133943
rect 328404 133900 328456 133909
rect 385536 133943 385588 133952
rect 385536 133909 385545 133943
rect 385545 133909 385579 133943
rect 385579 133909 385588 133943
rect 392436 133943 392488 133952
rect 385536 133900 385588 133909
rect 392436 133909 392445 133943
rect 392445 133909 392479 133943
rect 392479 133909 392488 133943
rect 392436 133900 392488 133909
rect 529056 133943 529108 133952
rect 529056 133909 529065 133943
rect 529065 133909 529099 133943
rect 529099 133909 529108 133943
rect 529056 133900 529108 133909
rect 535956 133943 536008 133952
rect 535956 133909 535965 133943
rect 535965 133909 535999 133943
rect 535999 133909 536008 133943
rect 535956 133900 536008 133909
rect 552240 133943 552292 133952
rect 552240 133909 552249 133943
rect 552249 133909 552283 133943
rect 552283 133909 552292 133943
rect 552240 133900 552292 133909
rect 571836 133943 571888 133952
rect 571836 133909 571845 133943
rect 571845 133909 571879 133943
rect 571879 133909 571888 133943
rect 571836 133900 571888 133909
rect 552240 133739 552292 133748
rect 552240 133705 552249 133739
rect 552249 133705 552283 133739
rect 552283 133705 552292 133739
rect 552240 133696 552292 133705
rect 290316 132812 290368 132864
rect 293260 132812 293312 132864
rect 399244 132812 399296 132864
rect 406144 132812 406196 132864
rect 375876 132540 375928 132592
rect 385444 132540 385496 132592
rect 275504 129820 275556 129872
rect 275688 129820 275740 129872
rect 279828 129752 279880 129804
rect 275596 129684 275648 129736
rect 275688 129684 275740 129736
rect 239256 128460 239308 128512
rect 239440 128460 239492 128512
rect 271456 128503 271508 128512
rect 271456 128469 271465 128503
rect 271465 128469 271499 128503
rect 271499 128469 271508 128503
rect 271456 128460 271508 128469
rect 239256 128256 239308 128308
rect 239440 128256 239492 128308
rect 259404 128299 259456 128308
rect 259404 128265 259413 128299
rect 259413 128265 259447 128299
rect 259447 128265 259456 128299
rect 259404 128256 259456 128265
rect 268696 128299 268748 128308
rect 268696 128265 268705 128299
rect 268705 128265 268739 128299
rect 268739 128265 268748 128299
rect 268696 128256 268748 128265
rect 371920 128299 371972 128308
rect 371920 128265 371929 128299
rect 371929 128265 371963 128299
rect 371963 128265 371972 128299
rect 371920 128256 371972 128265
rect 242844 125579 242896 125588
rect 242844 125545 242853 125579
rect 242853 125545 242887 125579
rect 242887 125545 242896 125579
rect 242844 125536 242896 125545
rect 246524 125536 246576 125588
rect 305128 125579 305180 125588
rect 305128 125545 305137 125579
rect 305137 125545 305171 125579
rect 305171 125545 305180 125579
rect 305128 125536 305180 125545
rect 308992 125579 309044 125588
rect 308992 125545 309001 125579
rect 309001 125545 309035 125579
rect 309035 125545 309044 125579
rect 308992 125536 309044 125545
rect 331072 125536 331124 125588
rect 331256 125536 331308 125588
rect 341100 125579 341152 125588
rect 341100 125545 341109 125579
rect 341109 125545 341143 125579
rect 341143 125545 341152 125579
rect 341100 125536 341152 125545
rect 246616 125468 246668 125520
rect 552516 125400 552568 125452
rect 135664 124151 135716 124160
rect 135664 124117 135673 124151
rect 135673 124117 135707 124151
rect 135707 124117 135716 124151
rect 135664 124108 135716 124117
rect 152224 124151 152276 124160
rect 152224 124117 152233 124151
rect 152233 124117 152267 124151
rect 152267 124117 152276 124151
rect 152224 124108 152276 124117
rect 170164 124151 170216 124160
rect 170164 124117 170173 124151
rect 170173 124117 170207 124151
rect 170207 124117 170216 124151
rect 170164 124108 170216 124117
rect 190864 124151 190916 124160
rect 190864 124117 190873 124151
rect 190873 124117 190907 124151
rect 190907 124117 190916 124151
rect 190864 124108 190916 124117
rect 214324 124151 214376 124160
rect 214324 124117 214333 124151
rect 214333 124117 214367 124151
rect 214367 124117 214376 124151
rect 214324 124108 214376 124117
rect 373116 124151 373168 124160
rect 373116 124117 373125 124151
rect 373125 124117 373159 124151
rect 373159 124117 373168 124151
rect 373116 124108 373168 124117
rect 385536 124151 385588 124160
rect 385536 124117 385545 124151
rect 385545 124117 385579 124151
rect 385579 124117 385588 124151
rect 392436 124151 392488 124160
rect 385536 124108 385588 124117
rect 392436 124117 392445 124151
rect 392445 124117 392479 124151
rect 392479 124117 392488 124151
rect 392436 124108 392488 124117
rect 529056 124151 529108 124160
rect 529056 124117 529065 124151
rect 529065 124117 529099 124151
rect 529099 124117 529108 124151
rect 529056 124108 529108 124117
rect 535956 124151 536008 124160
rect 535956 124117 535965 124151
rect 535965 124117 535999 124151
rect 535999 124117 536008 124151
rect 535956 124108 536008 124117
rect 571836 124151 571888 124160
rect 571836 124117 571845 124151
rect 571845 124117 571879 124151
rect 571879 124117 571888 124151
rect 571836 124108 571888 124117
rect 553436 122748 553488 122800
rect 553896 122748 553948 122800
rect 272836 121431 272888 121440
rect 272836 121397 272845 121431
rect 272845 121397 272879 121431
rect 272879 121397 272888 121431
rect 272836 121388 272888 121397
rect 273020 121388 273072 121440
rect 273112 121388 273164 121440
rect 279736 121388 279788 121440
rect 279828 121388 279880 121440
rect 285624 120071 285676 120080
rect 285624 120037 285633 120071
rect 285633 120037 285667 120071
rect 285667 120037 285676 120071
rect 285624 120028 285676 120037
rect 242568 119348 242620 119400
rect 242936 119348 242988 119400
rect 309176 119348 309228 119400
rect 229872 118736 229924 118788
rect 305128 118507 305180 118516
rect 305128 118473 305137 118507
rect 305137 118473 305171 118507
rect 305171 118473 305180 118507
rect 305128 118464 305180 118473
rect 242844 116739 242896 116748
rect 242844 116705 242853 116739
rect 242853 116705 242887 116739
rect 242887 116705 242896 116739
rect 242844 116696 242896 116705
rect 341192 116016 341244 116068
rect 259312 115948 259364 116000
rect 259496 115948 259548 116000
rect 91504 115787 91556 115796
rect 91504 115753 91513 115787
rect 91513 115753 91547 115787
rect 91547 115753 91556 115787
rect 91504 115744 91556 115753
rect 235576 115787 235628 115796
rect 235576 115753 235585 115787
rect 235585 115753 235619 115787
rect 235619 115753 235628 115787
rect 235576 115744 235628 115753
rect 357936 115787 357988 115796
rect 357936 115753 357945 115787
rect 357945 115753 357979 115787
rect 357979 115753 357988 115787
rect 357936 115744 357988 115753
rect 229780 114699 229832 114708
rect 229780 114665 229789 114699
rect 229789 114665 229823 114699
rect 229823 114665 229832 114699
rect 229780 114656 229832 114665
rect 135664 114563 135716 114572
rect 135664 114529 135673 114563
rect 135673 114529 135707 114563
rect 135707 114529 135716 114563
rect 135664 114520 135716 114529
rect 152224 114563 152276 114572
rect 152224 114529 152233 114563
rect 152233 114529 152267 114563
rect 152267 114529 152276 114563
rect 152224 114520 152276 114529
rect 170164 114563 170216 114572
rect 170164 114529 170173 114563
rect 170173 114529 170207 114563
rect 170207 114529 170216 114563
rect 170164 114520 170216 114529
rect 190864 114563 190916 114572
rect 190864 114529 190873 114563
rect 190873 114529 190907 114563
rect 190907 114529 190916 114563
rect 190864 114520 190916 114529
rect 214324 114563 214376 114572
rect 214324 114529 214333 114563
rect 214333 114529 214367 114563
rect 214367 114529 214376 114563
rect 214324 114520 214376 114529
rect 319940 114520 319992 114572
rect 320124 114520 320176 114572
rect 373116 114563 373168 114572
rect 373116 114529 373125 114563
rect 373125 114529 373159 114563
rect 373159 114529 373168 114563
rect 373116 114520 373168 114529
rect 385536 114563 385588 114572
rect 385536 114529 385545 114563
rect 385545 114529 385579 114563
rect 385579 114529 385588 114563
rect 392436 114563 392488 114572
rect 385536 114520 385588 114529
rect 392436 114529 392445 114563
rect 392445 114529 392479 114563
rect 392479 114529 392488 114563
rect 392436 114520 392488 114529
rect 529056 114563 529108 114572
rect 529056 114529 529065 114563
rect 529065 114529 529099 114563
rect 529099 114529 529108 114563
rect 529056 114520 529108 114529
rect 535956 114563 536008 114572
rect 535956 114529 535965 114563
rect 535965 114529 535999 114563
rect 535999 114529 536008 114563
rect 535956 114520 536008 114529
rect 571836 114563 571888 114572
rect 571836 114529 571845 114563
rect 571845 114529 571879 114563
rect 571879 114529 571888 114563
rect 571836 114520 571888 114529
rect 242844 114495 242896 114504
rect 242844 114461 242853 114495
rect 242853 114461 242887 114495
rect 242887 114461 242896 114495
rect 242844 114452 242896 114461
rect 552516 114452 552568 114504
rect 552608 114452 552660 114504
rect 272836 111843 272888 111852
rect 272836 111809 272845 111843
rect 272845 111809 272879 111843
rect 272879 111809 272888 111843
rect 272836 111800 272888 111809
rect 285256 111800 285308 111852
rect 285348 111800 285400 111852
rect 285624 111299 285676 111308
rect 285624 111265 285633 111299
rect 285633 111265 285667 111299
rect 285667 111265 285676 111299
rect 285624 111256 285676 111265
rect 242936 111120 242988 111172
rect 242936 110508 242988 110560
rect 553620 109692 553672 109744
rect 229780 109012 229832 109064
rect 275504 109012 275556 109064
rect 275596 109012 275648 109064
rect 305036 109012 305088 109064
rect 305220 109012 305272 109064
rect 320124 109055 320176 109064
rect 320124 109021 320133 109055
rect 320133 109021 320167 109055
rect 320167 109021 320176 109055
rect 320124 109012 320176 109021
rect 328404 109055 328456 109064
rect 328404 109021 328413 109055
rect 328413 109021 328447 109055
rect 328447 109021 328456 109055
rect 328404 109012 328456 109021
rect 229872 108944 229924 108996
rect 235576 108987 235628 108996
rect 235576 108953 235585 108987
rect 235585 108953 235619 108987
rect 235619 108953 235628 108987
rect 235576 108944 235628 108953
rect 91504 106335 91556 106344
rect 91504 106301 91513 106335
rect 91513 106301 91547 106335
rect 91547 106301 91556 106335
rect 91504 106292 91556 106301
rect 275596 106292 275648 106344
rect 309176 106292 309228 106344
rect 357936 106335 357988 106344
rect 357936 106301 357945 106335
rect 357945 106301 357979 106335
rect 357979 106301 357988 106335
rect 357936 106292 357988 106301
rect 235484 106267 235536 106276
rect 235484 106233 235493 106267
rect 235493 106233 235527 106267
rect 235527 106233 235536 106267
rect 235484 106224 235536 106233
rect 239256 106224 239308 106276
rect 239440 106224 239492 106276
rect 309084 106224 309136 106276
rect 331072 106224 331124 106276
rect 331256 106224 331308 106276
rect 341008 106224 341060 106276
rect 341100 106224 341152 106276
rect 242660 104907 242712 104916
rect 242660 104873 242669 104907
rect 242669 104873 242703 104907
rect 242703 104873 242712 104907
rect 242660 104864 242712 104873
rect 320124 104907 320176 104916
rect 320124 104873 320133 104907
rect 320133 104873 320167 104907
rect 320167 104873 320176 104907
rect 320124 104864 320176 104873
rect 328404 104907 328456 104916
rect 328404 104873 328413 104907
rect 328413 104873 328447 104907
rect 328447 104873 328456 104907
rect 328404 104864 328456 104873
rect 371828 104864 371880 104916
rect 371920 104864 371972 104916
rect 135664 104839 135716 104848
rect 135664 104805 135673 104839
rect 135673 104805 135707 104839
rect 135707 104805 135716 104839
rect 135664 104796 135716 104805
rect 152224 104839 152276 104848
rect 152224 104805 152233 104839
rect 152233 104805 152267 104839
rect 152267 104805 152276 104839
rect 152224 104796 152276 104805
rect 170164 104839 170216 104848
rect 170164 104805 170173 104839
rect 170173 104805 170207 104839
rect 170207 104805 170216 104839
rect 170164 104796 170216 104805
rect 190864 104839 190916 104848
rect 190864 104805 190873 104839
rect 190873 104805 190907 104839
rect 190907 104805 190916 104839
rect 190864 104796 190916 104805
rect 214324 104839 214376 104848
rect 214324 104805 214333 104839
rect 214333 104805 214367 104839
rect 214367 104805 214376 104839
rect 214324 104796 214376 104805
rect 305036 104839 305088 104848
rect 305036 104805 305045 104839
rect 305045 104805 305079 104839
rect 305079 104805 305088 104839
rect 305036 104796 305088 104805
rect 373116 104839 373168 104848
rect 373116 104805 373125 104839
rect 373125 104805 373159 104839
rect 373159 104805 373168 104839
rect 373116 104796 373168 104805
rect 385536 104839 385588 104848
rect 385536 104805 385545 104839
rect 385545 104805 385579 104839
rect 385579 104805 385588 104839
rect 392436 104839 392488 104848
rect 385536 104796 385588 104805
rect 392436 104805 392445 104839
rect 392445 104805 392479 104839
rect 392479 104805 392488 104839
rect 392436 104796 392488 104805
rect 529056 104839 529108 104848
rect 529056 104805 529065 104839
rect 529065 104805 529099 104839
rect 529099 104805 529108 104839
rect 529056 104796 529108 104805
rect 535956 104839 536008 104848
rect 535956 104805 535965 104839
rect 535965 104805 535999 104839
rect 535999 104805 536008 104839
rect 535956 104796 536008 104805
rect 571836 104839 571888 104848
rect 571836 104805 571845 104839
rect 571845 104805 571879 104839
rect 571879 104805 571888 104839
rect 571836 104796 571888 104805
rect 229872 103436 229924 103488
rect 309084 103436 309136 103488
rect 320124 103436 320176 103488
rect 552424 103436 552476 103488
rect 285348 102348 285400 102400
rect 285256 102187 285308 102196
rect 285256 102153 285265 102187
rect 285265 102153 285299 102187
rect 285299 102153 285308 102187
rect 285256 102144 285308 102153
rect 242108 101396 242160 101448
rect 360420 100920 360472 100972
rect 366124 100920 366176 100972
rect 251676 100852 251728 100904
rect 261152 100852 261204 100904
rect 275504 100759 275556 100768
rect 275504 100725 275513 100759
rect 275513 100725 275547 100759
rect 275547 100725 275556 100759
rect 275504 100716 275556 100725
rect 279736 100716 279788 100768
rect 280012 100716 280064 100768
rect 246616 99424 246668 99476
rect 268696 99356 268748 99408
rect 271456 99356 271508 99408
rect 271640 99356 271692 99408
rect 246616 99288 246668 99340
rect 305128 99288 305180 99340
rect 268696 99220 268748 99272
rect 553896 96747 553948 96756
rect 553896 96713 553905 96747
rect 553905 96713 553939 96747
rect 553939 96713 553948 96747
rect 553896 96704 553948 96713
rect 235484 96679 235536 96688
rect 235484 96645 235493 96679
rect 235493 96645 235527 96679
rect 235527 96645 235536 96679
rect 235484 96636 235536 96645
rect 91320 96568 91372 96620
rect 91504 96568 91556 96620
rect 235576 96611 235628 96620
rect 235576 96577 235585 96611
rect 235585 96577 235619 96611
rect 235619 96577 235628 96611
rect 235576 96568 235628 96577
rect 268696 96611 268748 96620
rect 268696 96577 268705 96611
rect 268705 96577 268739 96611
rect 268739 96577 268748 96611
rect 268696 96568 268748 96577
rect 307888 96568 307940 96620
rect 308256 96568 308308 96620
rect 341192 96568 341244 96620
rect 341376 96568 341428 96620
rect 357936 96568 357988 96620
rect 358212 96568 358264 96620
rect 553712 96568 553764 96620
rect 553896 96568 553948 96620
rect 135664 95319 135716 95328
rect 135664 95285 135673 95319
rect 135673 95285 135707 95319
rect 135707 95285 135716 95319
rect 135664 95276 135716 95285
rect 152224 95319 152276 95328
rect 152224 95285 152233 95319
rect 152233 95285 152267 95319
rect 152267 95285 152276 95319
rect 152224 95276 152276 95285
rect 170164 95319 170216 95328
rect 170164 95285 170173 95319
rect 170173 95285 170207 95319
rect 170207 95285 170216 95319
rect 170164 95276 170216 95285
rect 190864 95319 190916 95328
rect 190864 95285 190873 95319
rect 190873 95285 190907 95319
rect 190907 95285 190916 95319
rect 190864 95276 190916 95285
rect 214324 95319 214376 95328
rect 214324 95285 214333 95319
rect 214333 95285 214367 95319
rect 214367 95285 214376 95319
rect 214324 95276 214376 95285
rect 371920 95276 371972 95328
rect 372012 95276 372064 95328
rect 373116 95319 373168 95328
rect 373116 95285 373125 95319
rect 373125 95285 373159 95319
rect 373159 95285 373168 95319
rect 373116 95276 373168 95285
rect 385536 95319 385588 95328
rect 385536 95285 385545 95319
rect 385545 95285 385579 95319
rect 385579 95285 385588 95319
rect 392436 95319 392488 95328
rect 385536 95276 385588 95285
rect 392436 95285 392445 95319
rect 392445 95285 392479 95319
rect 392479 95285 392488 95319
rect 392436 95276 392488 95285
rect 529056 95319 529108 95328
rect 529056 95285 529065 95319
rect 529065 95285 529099 95319
rect 529099 95285 529108 95319
rect 529056 95276 529108 95285
rect 535956 95319 536008 95328
rect 535956 95285 535965 95319
rect 535965 95285 535999 95319
rect 535999 95285 536008 95319
rect 535956 95276 536008 95285
rect 571836 95319 571888 95328
rect 571836 95285 571845 95319
rect 571845 95285 571879 95319
rect 571879 95285 571888 95319
rect 571836 95276 571888 95285
rect 328588 95072 328640 95124
rect 371920 95115 371972 95124
rect 371920 95081 371929 95115
rect 371929 95081 371963 95115
rect 371963 95081 371972 95115
rect 371920 95072 371972 95081
rect 328588 94936 328640 94988
rect 278816 93916 278868 93968
rect 242016 93891 242068 93900
rect 242016 93857 242025 93891
rect 242025 93857 242059 93891
rect 242059 93857 242068 93891
rect 242016 93848 242068 93857
rect 276516 93848 276568 93900
rect 278724 93848 278776 93900
rect 285256 93848 285308 93900
rect 285348 93848 285400 93900
rect 308900 93891 308952 93900
rect 308900 93857 308909 93891
rect 308909 93857 308943 93891
rect 308943 93857 308952 93891
rect 308900 93848 308952 93857
rect 319940 93891 319992 93900
rect 319940 93857 319949 93891
rect 319949 93857 319983 93891
rect 319983 93857 319992 93891
rect 319940 93848 319992 93857
rect 552424 93848 552476 93900
rect 276608 93780 276660 93832
rect 275504 91060 275556 91112
rect 275688 91060 275740 91112
rect 279828 91060 279880 91112
rect 280012 91060 280064 91112
rect 246616 90040 246668 90092
rect 235576 89675 235628 89684
rect 235576 89641 235585 89675
rect 235585 89641 235619 89675
rect 235619 89641 235628 89675
rect 235576 89632 235628 89641
rect 268696 89675 268748 89684
rect 268696 89641 268705 89675
rect 268705 89641 268739 89675
rect 268739 89641 268748 89675
rect 268696 89632 268748 89641
rect 97024 88952 97076 89004
rect 249008 88952 249060 89004
rect 246524 88451 246576 88460
rect 246524 88417 246533 88451
rect 246533 88417 246567 88451
rect 246567 88417 246576 88451
rect 246524 88408 246576 88417
rect 242476 87227 242528 87236
rect 242476 87193 242485 87227
rect 242485 87193 242519 87227
rect 242519 87193 242528 87227
rect 242476 87184 242528 87193
rect 552424 87159 552476 87168
rect 552424 87125 552433 87159
rect 552433 87125 552467 87159
rect 552467 87125 552476 87159
rect 552424 87116 552476 87125
rect 242844 86912 242896 86964
rect 242936 86912 242988 86964
rect 305128 86955 305180 86964
rect 305128 86921 305137 86955
rect 305137 86921 305171 86955
rect 305171 86921 305180 86955
rect 305128 86912 305180 86921
rect 331072 86912 331124 86964
rect 331256 86912 331308 86964
rect 341100 86955 341152 86964
rect 341100 86921 341109 86955
rect 341109 86921 341143 86955
rect 341143 86921 341152 86955
rect 341100 86912 341152 86921
rect 361340 86912 361392 86964
rect 580668 86912 580720 86964
rect 242476 86887 242528 86896
rect 242476 86853 242485 86887
rect 242485 86853 242519 86887
rect 242519 86853 242528 86887
rect 242476 86844 242528 86853
rect 552424 86887 552476 86896
rect 552424 86853 552433 86887
rect 552433 86853 552467 86887
rect 552467 86853 552476 86887
rect 552424 86844 552476 86853
rect 279828 86776 279880 86828
rect 280012 86776 280064 86828
rect 230056 85552 230108 85604
rect 372012 85552 372064 85604
rect 135664 85527 135716 85536
rect 135664 85493 135673 85527
rect 135673 85493 135707 85527
rect 135707 85493 135716 85527
rect 135664 85484 135716 85493
rect 152224 85527 152276 85536
rect 152224 85493 152233 85527
rect 152233 85493 152267 85527
rect 152267 85493 152276 85527
rect 152224 85484 152276 85493
rect 170164 85527 170216 85536
rect 170164 85493 170173 85527
rect 170173 85493 170207 85527
rect 170207 85493 170216 85527
rect 170164 85484 170216 85493
rect 190864 85527 190916 85536
rect 190864 85493 190873 85527
rect 190873 85493 190907 85527
rect 190907 85493 190916 85527
rect 190864 85484 190916 85493
rect 214324 85527 214376 85536
rect 214324 85493 214333 85527
rect 214333 85493 214367 85527
rect 214367 85493 214376 85527
rect 214324 85484 214376 85493
rect 242476 85527 242528 85536
rect 242476 85493 242485 85527
rect 242485 85493 242519 85527
rect 242519 85493 242528 85527
rect 242476 85484 242528 85493
rect 319940 85527 319992 85536
rect 319940 85493 319949 85527
rect 319949 85493 319983 85527
rect 319983 85493 319992 85527
rect 319940 85484 319992 85493
rect 373116 85527 373168 85536
rect 373116 85493 373125 85527
rect 373125 85493 373159 85527
rect 373159 85493 373168 85527
rect 373116 85484 373168 85493
rect 385536 85527 385588 85536
rect 385536 85493 385545 85527
rect 385545 85493 385579 85527
rect 385579 85493 385588 85527
rect 392436 85527 392488 85536
rect 385536 85484 385588 85493
rect 392436 85493 392445 85527
rect 392445 85493 392479 85527
rect 392479 85493 392488 85527
rect 392436 85484 392488 85493
rect 529056 85527 529108 85536
rect 529056 85493 529065 85527
rect 529065 85493 529099 85527
rect 529099 85493 529108 85527
rect 529056 85484 529108 85493
rect 535956 85527 536008 85536
rect 535956 85493 535965 85527
rect 535965 85493 535999 85527
rect 535999 85493 536008 85527
rect 535956 85484 536008 85493
rect 552424 85484 552476 85536
rect 571836 85527 571888 85536
rect 571836 85493 571845 85527
rect 571845 85493 571879 85527
rect 571879 85493 571888 85527
rect 571836 85484 571888 85493
rect 242568 85280 242620 85332
rect 280012 84192 280064 84244
rect 279920 84124 279972 84176
rect 276976 82900 277028 82952
rect 277068 82832 277120 82884
rect 276608 82807 276660 82816
rect 276608 82773 276617 82807
rect 276617 82773 276651 82807
rect 276651 82773 276660 82807
rect 276608 82764 276660 82773
rect 279828 82764 279880 82816
rect 280104 82764 280156 82816
rect 285256 82807 285308 82816
rect 285256 82773 285265 82807
rect 285265 82773 285299 82807
rect 285299 82773 285308 82807
rect 285256 82764 285308 82773
rect 271456 81472 271508 81524
rect 230056 80112 230108 80164
rect 271364 80087 271416 80096
rect 271364 80053 271373 80087
rect 271373 80053 271407 80087
rect 271407 80053 271416 80087
rect 271364 80044 271416 80053
rect 229964 79883 230016 79892
rect 229964 79849 229973 79883
rect 229973 79849 230007 79883
rect 230007 79849 230016 79883
rect 229964 79840 230016 79849
rect 305128 79883 305180 79892
rect 305128 79849 305137 79883
rect 305137 79849 305171 79883
rect 305171 79849 305180 79883
rect 305128 79840 305180 79849
rect 285256 77979 285308 77988
rect 285256 77945 285265 77979
rect 285265 77945 285299 77979
rect 285299 77945 285308 77979
rect 285256 77936 285308 77945
rect 341192 77392 341244 77444
rect 91504 77163 91556 77172
rect 91504 77129 91513 77163
rect 91513 77129 91547 77163
rect 91547 77129 91556 77163
rect 91504 77120 91556 77129
rect 235576 77120 235628 77172
rect 341192 77120 341244 77172
rect 357936 77163 357988 77172
rect 357936 77129 357945 77163
rect 357945 77129 357979 77163
rect 357979 77129 357988 77163
rect 552332 77163 552384 77172
rect 357936 77120 357988 77129
rect 552332 77129 552341 77163
rect 552341 77129 552375 77163
rect 552375 77129 552384 77163
rect 552332 77120 552384 77129
rect 271364 76576 271416 76628
rect 135664 75939 135716 75948
rect 135664 75905 135673 75939
rect 135673 75905 135707 75939
rect 135707 75905 135716 75939
rect 135664 75896 135716 75905
rect 152224 75939 152276 75948
rect 152224 75905 152233 75939
rect 152233 75905 152267 75939
rect 152267 75905 152276 75939
rect 152224 75896 152276 75905
rect 170164 75939 170216 75948
rect 170164 75905 170173 75939
rect 170173 75905 170207 75939
rect 170207 75905 170216 75939
rect 170164 75896 170216 75905
rect 190864 75939 190916 75948
rect 190864 75905 190873 75939
rect 190873 75905 190907 75939
rect 190907 75905 190916 75939
rect 190864 75896 190916 75905
rect 214324 75939 214376 75948
rect 214324 75905 214333 75939
rect 214333 75905 214367 75939
rect 214367 75905 214376 75939
rect 214324 75896 214376 75905
rect 320124 75896 320176 75948
rect 373116 75939 373168 75948
rect 373116 75905 373125 75939
rect 373125 75905 373159 75939
rect 373159 75905 373168 75939
rect 373116 75896 373168 75905
rect 385536 75939 385588 75948
rect 385536 75905 385545 75939
rect 385545 75905 385579 75939
rect 385579 75905 385588 75939
rect 392436 75939 392488 75948
rect 385536 75896 385588 75905
rect 392436 75905 392445 75939
rect 392445 75905 392479 75939
rect 392479 75905 392488 75939
rect 392436 75896 392488 75905
rect 529056 75939 529108 75948
rect 529056 75905 529065 75939
rect 529065 75905 529099 75939
rect 529099 75905 529108 75939
rect 529056 75896 529108 75905
rect 535956 75939 536008 75948
rect 535956 75905 535965 75939
rect 535965 75905 535999 75939
rect 535999 75905 536008 75939
rect 535956 75896 536008 75905
rect 571836 75939 571888 75948
rect 571836 75905 571845 75939
rect 571845 75905 571879 75939
rect 571879 75905 571888 75939
rect 571836 75896 571888 75905
rect 279920 74647 279972 74656
rect 279920 74613 279929 74647
rect 279929 74613 279963 74647
rect 279963 74613 279972 74647
rect 279920 74604 279972 74613
rect 279920 74443 279972 74452
rect 279920 74409 279929 74443
rect 279929 74409 279963 74443
rect 279963 74409 279972 74443
rect 279920 74400 279972 74409
rect 276608 73219 276660 73228
rect 276608 73185 276617 73219
rect 276617 73185 276651 73219
rect 276651 73185 276660 73219
rect 276608 73176 276660 73185
rect 275688 73108 275740 73160
rect 371920 72156 371972 72208
rect 372104 72156 372156 72208
rect 246708 70499 246760 70508
rect 246708 70465 246717 70499
rect 246717 70465 246751 70499
rect 246751 70465 246760 70499
rect 246708 70456 246760 70465
rect 91504 67643 91556 67652
rect 91504 67609 91513 67643
rect 91513 67609 91547 67643
rect 91547 67609 91556 67643
rect 91504 67600 91556 67609
rect 235484 67643 235536 67652
rect 235484 67609 235493 67643
rect 235493 67609 235527 67643
rect 235527 67609 235536 67643
rect 235484 67600 235536 67609
rect 242016 67600 242068 67652
rect 242108 67600 242160 67652
rect 276976 67600 277028 67652
rect 278724 67668 278776 67720
rect 341100 67643 341152 67652
rect 341100 67609 341109 67643
rect 341109 67609 341143 67643
rect 341143 67609 341152 67643
rect 341100 67600 341152 67609
rect 357936 67643 357988 67652
rect 357936 67609 357945 67643
rect 357945 67609 357979 67643
rect 357979 67609 357988 67643
rect 357936 67600 357988 67609
rect 553896 67600 553948 67652
rect 553988 67600 554040 67652
rect 278632 67532 278684 67584
rect 331256 67575 331308 67584
rect 331256 67541 331265 67575
rect 331265 67541 331299 67575
rect 331299 67541 331308 67575
rect 331256 67532 331308 67541
rect 229872 66240 229924 66292
rect 229964 66240 230016 66292
rect 246708 66283 246760 66292
rect 246708 66249 246717 66283
rect 246717 66249 246751 66283
rect 246751 66249 246760 66283
rect 246708 66240 246760 66249
rect 285624 66240 285676 66292
rect 285808 66240 285860 66292
rect 373208 66240 373260 66292
rect 373300 66240 373352 66292
rect 135664 66215 135716 66224
rect 135664 66181 135673 66215
rect 135673 66181 135707 66215
rect 135707 66181 135716 66215
rect 135664 66172 135716 66181
rect 152224 66215 152276 66224
rect 152224 66181 152233 66215
rect 152233 66181 152267 66215
rect 152267 66181 152276 66215
rect 152224 66172 152276 66181
rect 170164 66215 170216 66224
rect 170164 66181 170173 66215
rect 170173 66181 170207 66215
rect 170207 66181 170216 66215
rect 170164 66172 170216 66181
rect 190864 66215 190916 66224
rect 190864 66181 190873 66215
rect 190873 66181 190907 66215
rect 190907 66181 190916 66215
rect 190864 66172 190916 66181
rect 214324 66215 214376 66224
rect 214324 66181 214333 66215
rect 214333 66181 214367 66215
rect 214367 66181 214376 66215
rect 214324 66172 214376 66181
rect 309084 66172 309136 66224
rect 320124 66215 320176 66224
rect 320124 66181 320133 66215
rect 320133 66181 320167 66215
rect 320167 66181 320176 66215
rect 320124 66172 320176 66181
rect 385536 66215 385588 66224
rect 385536 66181 385545 66215
rect 385545 66181 385579 66215
rect 385579 66181 385588 66215
rect 392436 66215 392488 66224
rect 385536 66172 385588 66181
rect 392436 66181 392445 66215
rect 392445 66181 392479 66215
rect 392479 66181 392488 66215
rect 392436 66172 392488 66181
rect 529056 66215 529108 66224
rect 529056 66181 529065 66215
rect 529065 66181 529099 66215
rect 529099 66181 529108 66215
rect 529056 66172 529108 66181
rect 535956 66215 536008 66224
rect 535956 66181 535965 66215
rect 535965 66181 535999 66215
rect 535999 66181 536008 66215
rect 535956 66172 536008 66181
rect 552516 66215 552568 66224
rect 552516 66181 552525 66215
rect 552525 66181 552559 66215
rect 552559 66181 552568 66215
rect 552516 66172 552568 66181
rect 571836 66215 571888 66224
rect 571836 66181 571845 66215
rect 571845 66181 571879 66215
rect 571879 66181 571888 66215
rect 571836 66172 571888 66181
rect 242568 64948 242620 65000
rect 242476 64880 242528 64932
rect 278632 64855 278684 64864
rect 278632 64821 278641 64855
rect 278641 64821 278675 64855
rect 278675 64821 278684 64855
rect 278632 64812 278684 64821
rect 279736 64855 279788 64864
rect 279736 64821 279745 64855
rect 279745 64821 279779 64855
rect 279779 64821 279788 64855
rect 279736 64812 279788 64821
rect 285256 64855 285308 64864
rect 285256 64821 285265 64855
rect 285265 64821 285299 64855
rect 285299 64821 285308 64855
rect 285256 64812 285308 64821
rect 372012 64812 372064 64864
rect 271456 63563 271508 63572
rect 271456 63529 271465 63563
rect 271465 63529 271499 63563
rect 271499 63529 271508 63563
rect 271456 63520 271508 63529
rect 275596 63563 275648 63572
rect 275596 63529 275605 63563
rect 275605 63529 275639 63563
rect 275639 63529 275648 63563
rect 275596 63520 275648 63529
rect 242476 63495 242528 63504
rect 242476 63461 242485 63495
rect 242485 63461 242519 63495
rect 242519 63461 242528 63495
rect 242476 63452 242528 63461
rect 331256 62815 331308 62824
rect 331256 62781 331265 62815
rect 331265 62781 331299 62815
rect 331299 62781 331308 62815
rect 331256 62772 331308 62781
rect 277068 62747 277120 62756
rect 277068 62713 277077 62747
rect 277077 62713 277111 62747
rect 277111 62713 277120 62747
rect 277068 62704 277120 62713
rect 273020 62092 273072 62144
rect 273112 62092 273164 62144
rect 229872 60800 229924 60852
rect 235484 60732 235536 60784
rect 229780 60664 229832 60716
rect 341192 60732 341244 60784
rect 341100 60664 341152 60716
rect 235576 60596 235628 60648
rect 3644 59168 3696 59220
rect 219200 59168 219252 59220
rect 553896 58012 553948 58064
rect 275596 57987 275648 57996
rect 275596 57953 275605 57987
rect 275605 57953 275639 57987
rect 275639 57953 275648 57987
rect 275596 57944 275648 57953
rect 91504 57919 91556 57928
rect 91504 57885 91513 57919
rect 91513 57885 91547 57919
rect 91547 57885 91556 57919
rect 91504 57876 91556 57885
rect 225180 57876 225232 57928
rect 225364 57876 225416 57928
rect 235576 57876 235628 57928
rect 272836 57919 272888 57928
rect 272836 57885 272845 57919
rect 272845 57885 272879 57919
rect 272879 57885 272888 57919
rect 272836 57876 272888 57885
rect 340916 57876 340968 57928
rect 341192 57876 341244 57928
rect 357936 57919 357988 57928
rect 357936 57885 357945 57919
rect 357945 57885 357979 57919
rect 357979 57885 357988 57919
rect 357936 57876 357988 57885
rect 553988 57876 554040 57928
rect 276424 57264 276476 57316
rect 135664 56695 135716 56704
rect 135664 56661 135673 56695
rect 135673 56661 135707 56695
rect 135707 56661 135716 56695
rect 135664 56652 135716 56661
rect 152224 56695 152276 56704
rect 152224 56661 152233 56695
rect 152233 56661 152267 56695
rect 152267 56661 152276 56695
rect 152224 56652 152276 56661
rect 170164 56695 170216 56704
rect 170164 56661 170173 56695
rect 170173 56661 170207 56695
rect 170207 56661 170216 56695
rect 170164 56652 170216 56661
rect 190864 56695 190916 56704
rect 190864 56661 190873 56695
rect 190873 56661 190907 56695
rect 190907 56661 190916 56695
rect 190864 56652 190916 56661
rect 214324 56695 214376 56704
rect 214324 56661 214333 56695
rect 214333 56661 214367 56695
rect 214367 56661 214376 56695
rect 214324 56652 214376 56661
rect 308900 56695 308952 56704
rect 308900 56661 308909 56695
rect 308909 56661 308943 56695
rect 308943 56661 308952 56695
rect 308900 56652 308952 56661
rect 320124 56695 320176 56704
rect 320124 56661 320133 56695
rect 320133 56661 320167 56695
rect 320167 56661 320176 56695
rect 320124 56652 320176 56661
rect 373116 56652 373168 56704
rect 373300 56652 373352 56704
rect 385536 56695 385588 56704
rect 385536 56661 385545 56695
rect 385545 56661 385579 56695
rect 385579 56661 385588 56695
rect 392436 56695 392488 56704
rect 385536 56652 385588 56661
rect 392436 56661 392445 56695
rect 392445 56661 392479 56695
rect 392479 56661 392488 56695
rect 392436 56652 392488 56661
rect 529056 56695 529108 56704
rect 529056 56661 529065 56695
rect 529065 56661 529099 56695
rect 529099 56661 529108 56695
rect 529056 56652 529108 56661
rect 535956 56695 536008 56704
rect 535956 56661 535965 56695
rect 535965 56661 535999 56695
rect 535999 56661 536008 56695
rect 535956 56652 536008 56661
rect 552516 56695 552568 56704
rect 552516 56661 552525 56695
rect 552525 56661 552559 56695
rect 552559 56661 552568 56695
rect 552516 56652 552568 56661
rect 571836 56695 571888 56704
rect 571836 56661 571845 56695
rect 571845 56661 571879 56695
rect 571879 56661 571888 56695
rect 571836 56652 571888 56661
rect 285256 56491 285308 56500
rect 285256 56457 285265 56491
rect 285265 56457 285299 56491
rect 285299 56457 285308 56491
rect 285256 56448 285308 56457
rect 278724 55224 278776 55276
rect 279736 55267 279788 55276
rect 279736 55233 279745 55267
rect 279745 55233 279779 55267
rect 279779 55233 279788 55267
rect 279736 55224 279788 55233
rect 371920 55267 371972 55276
rect 371920 55233 371929 55267
rect 371929 55233 371963 55267
rect 371963 55233 371972 55267
rect 371920 55224 371972 55233
rect 246892 55199 246944 55208
rect 246892 55165 246901 55199
rect 246901 55165 246935 55199
rect 246935 55165 246944 55199
rect 246892 55156 246944 55165
rect 268604 52504 268656 52556
rect 268696 52504 268748 52556
rect 275596 52479 275648 52488
rect 275596 52445 275605 52479
rect 275605 52445 275639 52479
rect 275639 52445 275648 52479
rect 275596 52436 275648 52445
rect 279736 51756 279788 51808
rect 280012 51756 280064 51808
rect 239256 51008 239308 51060
rect 239440 51008 239492 51060
rect 259220 51008 259272 51060
rect 259404 51008 259456 51060
rect 271364 51008 271416 51060
rect 271548 51008 271600 51060
rect 91504 48331 91556 48340
rect 91504 48297 91513 48331
rect 91513 48297 91547 48331
rect 91547 48297 91556 48331
rect 91504 48288 91556 48297
rect 235392 48331 235444 48340
rect 235392 48297 235401 48331
rect 235401 48297 235435 48331
rect 235435 48297 235444 48331
rect 235392 48288 235444 48297
rect 242752 48288 242804 48340
rect 242844 48288 242896 48340
rect 272836 48331 272888 48340
rect 272836 48297 272845 48331
rect 272845 48297 272879 48331
rect 272879 48297 272888 48331
rect 272836 48288 272888 48297
rect 278816 48288 278868 48340
rect 357936 48331 357988 48340
rect 357936 48297 357945 48331
rect 357945 48297 357979 48331
rect 357979 48297 357988 48331
rect 357936 48288 357988 48297
rect 259404 48220 259456 48272
rect 341008 48220 341060 48272
rect 341100 48220 341152 48272
rect 553804 48220 553856 48272
rect 553896 48220 553948 48272
rect 319848 46996 319900 47048
rect 320032 46996 320084 47048
rect 275596 46971 275648 46980
rect 275596 46937 275605 46971
rect 275605 46937 275639 46971
rect 275639 46937 275648 46971
rect 275596 46928 275648 46937
rect 135664 46903 135716 46912
rect 135664 46869 135673 46903
rect 135673 46869 135707 46903
rect 135707 46869 135716 46903
rect 135664 46860 135716 46869
rect 152224 46903 152276 46912
rect 152224 46869 152233 46903
rect 152233 46869 152267 46903
rect 152267 46869 152276 46903
rect 152224 46860 152276 46869
rect 170164 46903 170216 46912
rect 170164 46869 170173 46903
rect 170173 46869 170207 46903
rect 170207 46869 170216 46903
rect 170164 46860 170216 46869
rect 190864 46903 190916 46912
rect 190864 46869 190873 46903
rect 190873 46869 190907 46903
rect 190907 46869 190916 46903
rect 190864 46860 190916 46869
rect 214324 46903 214376 46912
rect 214324 46869 214333 46903
rect 214333 46869 214367 46903
rect 214367 46869 214376 46903
rect 214324 46860 214376 46869
rect 225364 46903 225416 46912
rect 225364 46869 225373 46903
rect 225373 46869 225407 46903
rect 225407 46869 225416 46903
rect 225364 46860 225416 46869
rect 242016 46860 242068 46912
rect 242108 46860 242160 46912
rect 272836 46903 272888 46912
rect 272836 46869 272845 46903
rect 272845 46869 272879 46903
rect 272879 46869 272888 46903
rect 272836 46860 272888 46869
rect 285072 46860 285124 46912
rect 285256 46860 285308 46912
rect 308992 46860 309044 46912
rect 309176 46860 309228 46912
rect 320032 46860 320084 46912
rect 328404 46860 328456 46912
rect 385536 46903 385588 46912
rect 385536 46869 385545 46903
rect 385545 46869 385579 46903
rect 385579 46869 385588 46903
rect 392436 46903 392488 46912
rect 385536 46860 385588 46869
rect 392436 46869 392445 46903
rect 392445 46869 392479 46903
rect 392479 46869 392488 46903
rect 392436 46860 392488 46869
rect 529056 46903 529108 46912
rect 529056 46869 529065 46903
rect 529065 46869 529099 46903
rect 529099 46869 529108 46903
rect 529056 46860 529108 46869
rect 535956 46903 536008 46912
rect 535956 46869 535965 46903
rect 535965 46869 535999 46903
rect 535999 46869 536008 46903
rect 535956 46860 536008 46869
rect 552516 46903 552568 46912
rect 552516 46869 552525 46903
rect 552525 46869 552559 46903
rect 552559 46869 552568 46903
rect 552516 46860 552568 46869
rect 553804 46903 553856 46912
rect 553804 46869 553813 46903
rect 553813 46869 553847 46903
rect 553847 46869 553856 46903
rect 553804 46860 553856 46869
rect 571836 46903 571888 46912
rect 571836 46869 571845 46903
rect 571845 46869 571879 46903
rect 571879 46869 571888 46903
rect 571836 46860 571888 46869
rect 392528 46656 392580 46708
rect 242568 45568 242620 45620
rect 246892 45611 246944 45620
rect 246892 45577 246901 45611
rect 246901 45577 246935 45611
rect 246935 45577 246944 45611
rect 246892 45568 246944 45577
rect 278724 45611 278776 45620
rect 278724 45577 278733 45611
rect 278733 45577 278767 45611
rect 278767 45577 278776 45611
rect 278724 45568 278776 45577
rect 276608 44140 276660 44192
rect 273112 42780 273164 42832
rect 273296 42780 273348 42832
rect 275596 42823 275648 42832
rect 275596 42789 275605 42823
rect 275605 42789 275639 42823
rect 275639 42789 275648 42823
rect 275596 42780 275648 42789
rect 273112 42644 273164 42696
rect 273020 42576 273072 42628
rect 285624 42032 285676 42084
rect 399244 38836 399296 38888
rect 406144 38836 406196 38888
rect 298596 38768 298648 38820
rect 308164 38768 308216 38820
rect 259312 38743 259364 38752
rect 259312 38709 259321 38743
rect 259321 38709 259355 38743
rect 259355 38709 259364 38743
rect 259312 38700 259364 38709
rect 261060 38700 261112 38752
rect 268144 38700 268196 38752
rect 377348 38700 377400 38752
rect 382040 38700 382092 38752
rect 91504 38539 91556 38548
rect 91504 38505 91513 38539
rect 91513 38505 91547 38539
rect 91547 38505 91556 38539
rect 91504 38496 91556 38505
rect 320308 38539 320360 38548
rect 320308 38505 320317 38539
rect 320317 38505 320351 38539
rect 320351 38505 320360 38539
rect 320308 38496 320360 38505
rect 357936 38539 357988 38548
rect 357936 38505 357945 38539
rect 357945 38505 357979 38539
rect 357979 38505 357988 38539
rect 357936 38496 357988 38505
rect 553804 38403 553856 38412
rect 553804 38369 553813 38403
rect 553813 38369 553847 38403
rect 553847 38369 553856 38403
rect 553804 38360 553856 38369
rect 275504 37952 275556 38004
rect 276240 37952 276292 38004
rect 276608 37952 276660 38004
rect 135664 37315 135716 37324
rect 135664 37281 135673 37315
rect 135673 37281 135707 37315
rect 135707 37281 135716 37315
rect 135664 37272 135716 37281
rect 152224 37315 152276 37324
rect 152224 37281 152233 37315
rect 152233 37281 152267 37315
rect 152267 37281 152276 37315
rect 152224 37272 152276 37281
rect 170164 37315 170216 37324
rect 170164 37281 170173 37315
rect 170173 37281 170207 37315
rect 170207 37281 170216 37315
rect 170164 37272 170216 37281
rect 190864 37315 190916 37324
rect 190864 37281 190873 37315
rect 190873 37281 190907 37315
rect 190907 37281 190916 37315
rect 190864 37272 190916 37281
rect 214324 37315 214376 37324
rect 214324 37281 214333 37315
rect 214333 37281 214367 37315
rect 214367 37281 214376 37315
rect 214324 37272 214376 37281
rect 225456 37272 225508 37324
rect 271456 37272 271508 37324
rect 271548 37272 271600 37324
rect 272836 37315 272888 37324
rect 272836 37281 272845 37315
rect 272845 37281 272879 37315
rect 272879 37281 272888 37315
rect 272836 37272 272888 37281
rect 276976 37272 277028 37324
rect 277068 37272 277120 37324
rect 280012 37272 280064 37324
rect 319940 37315 319992 37324
rect 319940 37281 319949 37315
rect 319949 37281 319983 37315
rect 319983 37281 319992 37315
rect 319940 37272 319992 37281
rect 328220 37315 328272 37324
rect 328220 37281 328229 37315
rect 328229 37281 328263 37315
rect 328263 37281 328272 37315
rect 328220 37272 328272 37281
rect 371920 37272 371972 37324
rect 372012 37272 372064 37324
rect 373024 37272 373076 37324
rect 373116 37272 373168 37324
rect 385536 37315 385588 37324
rect 385536 37281 385545 37315
rect 385545 37281 385579 37315
rect 385579 37281 385588 37315
rect 529056 37315 529108 37324
rect 385536 37272 385588 37281
rect 529056 37281 529065 37315
rect 529065 37281 529099 37315
rect 529099 37281 529108 37315
rect 529056 37272 529108 37281
rect 535956 37315 536008 37324
rect 535956 37281 535965 37315
rect 535965 37281 535999 37315
rect 535999 37281 536008 37315
rect 535956 37272 536008 37281
rect 552608 37272 552660 37324
rect 571836 37315 571888 37324
rect 571836 37281 571845 37315
rect 571845 37281 571879 37315
rect 571879 37281 571888 37315
rect 571836 37272 571888 37281
rect 242016 37204 242068 37256
rect 242108 37204 242160 37256
rect 278724 37204 278776 37256
rect 278908 37204 278960 37256
rect 279828 37204 279880 37256
rect 320308 31875 320360 31884
rect 320308 31841 320317 31875
rect 320317 31841 320351 31875
rect 320351 31841 320360 31875
rect 320308 31832 320360 31841
rect 341100 31832 341152 31884
rect 229964 31764 230016 31816
rect 235484 31807 235536 31816
rect 235484 31773 235493 31807
rect 235493 31773 235527 31807
rect 235527 31773 235536 31807
rect 235484 31764 235536 31773
rect 229964 31628 230016 31680
rect 91504 29019 91556 29028
rect 91504 28985 91513 29019
rect 91513 28985 91547 29019
rect 91547 28985 91556 29019
rect 91504 28976 91556 28985
rect 235484 29019 235536 29028
rect 235484 28985 235493 29019
rect 235493 28985 235527 29019
rect 235527 28985 235536 29019
rect 235484 28976 235536 28985
rect 242660 29044 242712 29096
rect 246892 29044 246944 29096
rect 242752 28976 242804 29028
rect 242844 28976 242896 29028
rect 246524 28976 246576 29028
rect 246616 28976 246668 29028
rect 246708 28976 246760 29028
rect 285072 28976 285124 29028
rect 285256 28976 285308 29028
rect 285808 28976 285860 29028
rect 308992 28976 309044 29028
rect 309176 28976 309228 29028
rect 341008 29019 341060 29028
rect 341008 28985 341017 29019
rect 341017 28985 341051 29019
rect 341051 28985 341060 29019
rect 341008 28976 341060 28985
rect 357936 29019 357988 29028
rect 357936 28985 357945 29019
rect 357945 28985 357979 29019
rect 357979 28985 357988 29019
rect 357936 28976 357988 28985
rect 553804 28976 553856 29028
rect 553896 28976 553948 29028
rect 242568 28908 242620 28960
rect 254896 28908 254948 28960
rect 285164 28951 285216 28960
rect 285164 28917 285173 28951
rect 285173 28917 285207 28951
rect 285207 28917 285216 28951
rect 285164 28908 285216 28917
rect 276240 27616 276292 27668
rect 276516 27616 276568 27668
rect 278816 27659 278868 27668
rect 278816 27625 278825 27659
rect 278825 27625 278859 27659
rect 278859 27625 278868 27659
rect 278816 27616 278868 27625
rect 135664 27548 135716 27600
rect 152224 27548 152276 27600
rect 170164 27548 170216 27600
rect 190220 27548 190272 27600
rect 190864 27548 190916 27600
rect 214324 27548 214376 27600
rect 214508 27548 214560 27600
rect 225364 27548 225416 27600
rect 242568 27591 242620 27600
rect 242568 27557 242577 27591
rect 242577 27557 242611 27591
rect 242611 27557 242620 27591
rect 242568 27548 242620 27557
rect 246524 27548 246576 27600
rect 246616 27548 246668 27600
rect 272836 27591 272888 27600
rect 272836 27557 272845 27591
rect 272845 27557 272879 27591
rect 272879 27557 272888 27591
rect 272836 27548 272888 27557
rect 305128 27591 305180 27600
rect 305128 27557 305137 27591
rect 305137 27557 305171 27591
rect 305171 27557 305180 27591
rect 305128 27548 305180 27557
rect 385536 27548 385588 27600
rect 385996 27548 386048 27600
rect 392436 27548 392488 27600
rect 392620 27548 392672 27600
rect 529056 27591 529108 27600
rect 529056 27557 529065 27591
rect 529065 27557 529099 27591
rect 529099 27557 529108 27591
rect 529056 27548 529108 27557
rect 535956 27591 536008 27600
rect 535956 27557 535965 27591
rect 535965 27557 535999 27591
rect 535999 27557 536008 27591
rect 535956 27548 536008 27557
rect 552516 27591 552568 27600
rect 552516 27557 552525 27591
rect 552525 27557 552559 27591
rect 552559 27557 552568 27591
rect 552516 27548 552568 27557
rect 571836 27591 571888 27600
rect 571836 27557 571845 27591
rect 571845 27557 571879 27591
rect 571879 27557 571888 27591
rect 571836 27548 571888 27557
rect 278816 26299 278868 26308
rect 278816 26265 278825 26299
rect 278825 26265 278859 26299
rect 278859 26265 278868 26299
rect 278816 26256 278868 26265
rect 3920 26188 3972 26240
rect 350024 26188 350076 26240
rect 275688 24828 275740 24880
rect 229964 24148 230016 24200
rect 230148 24148 230200 24200
rect 285808 24148 285860 24200
rect 319940 24148 319992 24200
rect 320124 24148 320176 24200
rect 242568 22695 242620 22704
rect 242568 22661 242577 22695
rect 242577 22661 242611 22695
rect 242611 22661 242620 22695
rect 242568 22652 242620 22661
rect 235484 22108 235536 22160
rect 277068 22108 277120 22160
rect 276976 22040 277028 22092
rect 367596 22040 367648 22092
rect 368332 22040 368384 22092
rect 368976 22040 369028 22092
rect 369528 22040 369580 22092
rect 235576 21972 235628 22024
rect 254804 21403 254856 21412
rect 254804 21369 254813 21403
rect 254813 21369 254847 21403
rect 254847 21369 254856 21403
rect 254804 21360 254856 21369
rect 313040 21360 313092 21412
rect 346896 21360 346948 21412
rect 285072 19388 285124 19440
rect 285164 19363 285216 19372
rect 285164 19329 285173 19363
rect 285173 19329 285207 19363
rect 285207 19329 285216 19363
rect 285164 19320 285216 19329
rect 285348 19320 285400 19372
rect 285716 19363 285768 19372
rect 285716 19329 285725 19363
rect 285725 19329 285759 19363
rect 285759 19329 285768 19363
rect 285716 19320 285768 19329
rect 91504 19295 91556 19304
rect 91504 19261 91513 19295
rect 91513 19261 91547 19295
rect 91547 19261 91556 19295
rect 91504 19252 91556 19261
rect 145324 19252 145376 19304
rect 308256 19295 308308 19304
rect 308256 19261 308265 19295
rect 308265 19261 308299 19295
rect 308299 19261 308308 19295
rect 308256 19252 308308 19261
rect 340732 19252 340784 19304
rect 341008 19252 341060 19304
rect 346896 19252 346948 19304
rect 347080 19252 347132 19304
rect 351036 19252 351088 19304
rect 351312 19252 351364 19304
rect 414516 19252 414568 19304
rect 414884 19252 414936 19304
rect 541476 19295 541528 19304
rect 541476 19261 541485 19295
rect 541485 19261 541519 19295
rect 541519 19261 541528 19295
rect 541476 19252 541528 19261
rect 560796 19295 560848 19304
rect 560796 19261 560805 19295
rect 560805 19261 560839 19295
rect 560839 19261 560848 19295
rect 560796 19252 560848 19261
rect 145232 19184 145284 19236
rect 273020 18776 273072 18828
rect 273204 18776 273256 18828
rect 236404 18572 236456 18624
rect 275780 18572 275832 18624
rect 299608 18572 299660 18624
rect 336132 18572 336184 18624
rect 242752 18096 242804 18148
rect 135296 18071 135348 18080
rect 135296 18037 135305 18071
rect 135305 18037 135339 18071
rect 135339 18037 135348 18071
rect 135296 18028 135348 18037
rect 151856 18071 151908 18080
rect 151856 18037 151865 18071
rect 151865 18037 151899 18071
rect 151899 18037 151908 18071
rect 151856 18028 151908 18037
rect 169704 18071 169756 18080
rect 169704 18037 169713 18071
rect 169713 18037 169747 18071
rect 169747 18037 169756 18071
rect 169704 18028 169756 18037
rect 225088 18071 225140 18080
rect 225088 18037 225097 18071
rect 225097 18037 225131 18071
rect 225131 18037 225140 18071
rect 225088 18028 225140 18037
rect 242660 18028 242712 18080
rect 272836 18071 272888 18080
rect 272836 18037 272845 18071
rect 272845 18037 272879 18071
rect 272879 18037 272888 18071
rect 272836 18028 272888 18037
rect 305128 18071 305180 18080
rect 305128 18037 305137 18071
rect 305137 18037 305171 18071
rect 305171 18037 305180 18071
rect 305128 18028 305180 18037
rect 373116 17867 373168 17876
rect 373116 17833 373125 17867
rect 373125 17833 373159 17867
rect 373159 17833 373168 17867
rect 373116 17824 373168 17833
rect 239256 17280 239308 17332
rect 239532 17280 239584 17332
rect 242476 17280 242528 17332
rect 242660 17280 242712 17332
rect 232172 17212 232224 17264
rect 277160 17212 277212 17264
rect 306140 17212 306192 17264
rect 328956 17212 329008 17264
rect 278632 16600 278684 16652
rect 278816 16600 278868 16652
rect 347908 16532 347960 16584
rect 348184 16532 348236 16584
rect 392344 15444 392396 15496
rect 393540 15444 393592 15496
rect 483516 14560 483568 14612
rect 483976 14560 484028 14612
rect 246064 14492 246116 14544
rect 264740 14492 264792 14544
rect 252964 14424 253016 14476
rect 282220 14424 282272 14476
rect 303380 14424 303432 14476
rect 322056 14424 322108 14476
rect 114964 12384 115016 12436
rect 253332 12384 253384 12436
rect 332912 12384 332964 12436
rect 493176 12384 493228 12436
rect 513876 12384 513928 12436
rect 514888 12384 514940 12436
rect 530436 12384 530488 12436
rect 531540 12384 531592 12436
rect 534576 12384 534628 12436
rect 535036 12384 535088 12436
rect 542856 12384 542908 12436
rect 543408 12384 543460 12436
rect 548376 12384 548428 12436
rect 549388 12384 549440 12436
rect 549756 12384 549808 12436
rect 550584 12384 550636 12436
rect 556656 12384 556708 12436
rect 557668 12384 557720 12436
rect 567696 12384 567748 12436
rect 568340 12384 568392 12436
rect 574596 12384 574648 12436
rect 575516 12384 575568 12436
rect 575976 12384 576028 12436
rect 576712 12384 576764 12436
rect 107972 12316 108024 12368
rect 251952 12316 252004 12368
rect 332820 12316 332872 12368
rect 495936 12316 495988 12368
rect 99508 12248 99560 12300
rect 250480 12248 250532 12300
rect 334200 12248 334252 12300
rect 500076 12248 500128 12300
rect 92608 12180 92660 12232
rect 249284 12180 249336 12232
rect 334108 12180 334160 12232
rect 504124 12180 504176 12232
rect 85984 12112 86036 12164
rect 248180 12112 248232 12164
rect 335488 12112 335540 12164
rect 511300 12112 511352 12164
rect 83132 12044 83184 12096
rect 246708 12044 246760 12096
rect 336868 12044 336920 12096
rect 518384 12044 518436 12096
rect 79084 11840 79136 11892
rect 246248 11840 246300 11892
rect 338156 11840 338208 11892
rect 525560 11840 525612 11892
rect 74944 11772 74996 11824
rect 244868 11772 244920 11824
rect 295560 11772 295612 11824
rect 316168 11772 316220 11824
rect 339628 11772 339680 11824
rect 532736 11772 532788 11824
rect 72184 11704 72236 11756
rect 244960 11704 245012 11756
rect 248824 11704 248876 11756
rect 281300 11704 281352 11756
rect 304760 11704 304812 11756
rect 324816 11704 324868 11756
rect 342480 11704 342532 11756
rect 539820 11704 539872 11756
rect 331348 11636 331400 11688
rect 489864 11636 489916 11688
rect 235300 11228 235352 11280
rect 117632 11092 117684 11144
rect 167588 11160 167640 11212
rect 215980 11160 216032 11212
rect 177248 11092 177300 11144
rect 56912 10956 56964 11008
rect 167496 11024 167548 11076
rect 215796 11024 215848 11076
rect 234932 11024 234984 11076
rect 236772 10956 236824 11008
rect 242292 10956 242344 11008
rect 323160 10956 323212 11008
rect 331348 11024 331400 11076
rect 328404 10956 328456 11008
rect 341468 11160 341520 11212
rect 348092 11228 348144 11280
rect 346528 11160 346580 11212
rect 408996 11160 409048 11212
rect 410192 11160 410244 11212
rect 460148 10956 460200 11008
rect 53324 10752 53376 10804
rect 147808 10752 147860 10804
rect 148452 10752 148504 10804
rect 153052 10752 153104 10804
rect 187092 10752 187144 10804
rect 191692 10752 191744 10804
rect 234656 10752 234708 10804
rect 235024 10752 235076 10804
rect 238152 10752 238204 10804
rect 238520 10752 238572 10804
rect 244132 10752 244184 10804
rect 327208 10752 327260 10804
rect 462816 10752 462868 10804
rect 50104 10684 50156 10736
rect 45964 10616 46016 10668
rect 153052 10616 153104 10668
rect 186816 10684 186868 10736
rect 191692 10616 191744 10668
rect 234840 10684 234892 10736
rect 239256 10684 239308 10736
rect 323068 10684 323120 10736
rect 328404 10684 328456 10736
rect 328496 10684 328548 10736
rect 235392 10616 235444 10668
rect 238244 10616 238296 10668
rect 243764 10616 243816 10668
rect 324448 10616 324500 10668
rect 329876 10616 329928 10668
rect 329968 10616 330020 10668
rect 466956 10684 467008 10736
rect 469716 10616 469768 10668
rect 41824 10548 41876 10600
rect 39064 10480 39116 10532
rect 123520 10548 123572 10600
rect 254988 10548 255040 10600
rect 318836 10548 318888 10600
rect 138424 10480 138476 10532
rect 254620 10480 254672 10532
rect 317548 10480 317600 10532
rect 408996 10480 409048 10532
rect 474408 10548 474460 10600
rect 477996 10480 478048 10532
rect 34924 10412 34976 10464
rect 253148 10412 253200 10464
rect 255724 10412 255776 10464
rect 282496 10412 282548 10464
rect 318652 10412 318704 10464
rect 418748 10412 418800 10464
rect 481584 10412 481636 10464
rect 60500 10208 60552 10260
rect 65284 10140 65336 10192
rect 128856 10140 128908 10192
rect 143300 10208 143352 10260
rect 138608 10140 138660 10192
rect 157468 10140 157520 10192
rect 68044 10072 68096 10124
rect 138240 10072 138292 10124
rect 143300 10072 143352 10124
rect 157560 10072 157612 10124
rect 167588 10140 167640 10192
rect 167864 10140 167916 10192
rect 195924 10140 195976 10192
rect 167772 10072 167824 10124
rect 196016 10072 196068 10124
rect 196384 10208 196436 10260
rect 225456 10140 225508 10192
rect 225640 10208 225692 10260
rect 232448 10251 232500 10260
rect 232448 10217 232457 10251
rect 232457 10217 232491 10251
rect 232491 10217 232500 10251
rect 232448 10208 232500 10217
rect 239624 10208 239676 10260
rect 327116 10208 327168 10260
rect 240912 10140 240964 10192
rect 253516 10140 253568 10192
rect 325828 10140 325880 10192
rect 455916 10208 455968 10260
rect 331624 10140 331676 10192
rect 451868 10140 451920 10192
rect 225640 10072 225692 10124
rect 235024 10072 235076 10124
rect 241924 10072 241976 10124
rect 242384 10072 242436 10124
rect 244776 10072 244828 10124
rect 325920 10072 325972 10124
rect 102544 10004 102596 10056
rect 250388 10004 250440 10056
rect 324540 10004 324592 10056
rect 331348 10072 331400 10124
rect 449016 10072 449068 10124
rect 331624 10004 331676 10056
rect 444876 10004 444928 10056
rect 106684 9936 106736 9988
rect 252320 9936 252372 9988
rect 321780 9936 321832 9988
rect 442116 9936 442168 9988
rect 109444 9868 109496 9920
rect 251860 9868 251912 9920
rect 320216 9868 320268 9920
rect 437976 9868 438028 9920
rect 91504 9707 91556 9716
rect 91504 9673 91513 9707
rect 91513 9673 91547 9707
rect 91547 9673 91556 9707
rect 91504 9664 91556 9673
rect 113584 9664 113636 9716
rect 124624 9596 124676 9648
rect 138240 9596 138292 9648
rect 128856 9528 128908 9580
rect 169520 9596 169572 9648
rect 170164 9596 170216 9648
rect 257472 9596 257524 9648
rect 285072 9664 285124 9716
rect 285256 9664 285308 9716
rect 305036 9664 305088 9716
rect 305128 9664 305180 9716
rect 308256 9707 308308 9716
rect 308256 9673 308265 9707
rect 308265 9673 308299 9707
rect 308299 9673 308308 9707
rect 308256 9664 308308 9673
rect 320124 9664 320176 9716
rect 262808 9596 262860 9648
rect 309176 9596 309228 9648
rect 385168 9596 385220 9648
rect 431076 9596 431128 9648
rect 150936 9528 150988 9580
rect 261612 9528 261664 9580
rect 310648 9528 310700 9580
rect 388756 9528 388808 9580
rect 426936 9528 426988 9580
rect 147348 9460 147400 9512
rect 259036 9460 259088 9512
rect 262900 9460 262952 9512
rect 312028 9460 312080 9512
rect 392344 9460 392396 9512
rect 435124 9664 435176 9716
rect 529148 9664 529200 9716
rect 536232 9664 536284 9716
rect 542212 9664 542264 9716
rect 545524 9664 545576 9716
rect 545800 9664 545852 9716
rect 552884 9664 552936 9716
rect 561256 9664 561308 9716
rect 571928 9664 571980 9716
rect 143760 9324 143812 9376
rect 259220 9392 259272 9444
rect 349380 9392 349432 9444
rect 350852 9392 350904 9444
rect 351128 9392 351180 9444
rect 560060 9392 560112 9444
rect 244868 9324 244920 9376
rect 279644 9324 279696 9376
rect 341284 9324 341336 9376
rect 346620 9324 346672 9376
rect 349288 9324 349340 9376
rect 349472 9324 349524 9376
rect 563648 9324 563700 9376
rect 136584 9120 136636 9172
rect 244776 9120 244828 9172
rect 244868 9120 244920 9172
rect 254252 9120 254304 9172
rect 254436 9120 254488 9172
rect 254528 9120 254580 9172
rect 278080 9120 278132 9172
rect 567236 9120 567288 9172
rect 27196 9052 27248 9104
rect 9348 8916 9400 8968
rect 140172 8984 140224 9036
rect 191784 8984 191836 9036
rect 233828 8984 233880 9036
rect 231344 8916 231396 8968
rect 233000 8916 233052 8968
rect 278172 9052 278224 9104
rect 234932 8984 234984 9036
rect 276792 8984 276844 9036
rect 303748 8984 303800 9036
rect 351220 8984 351272 9036
rect 570732 9052 570784 9104
rect 574320 8984 574372 9036
rect 235024 8916 235076 8968
rect 276700 8916 276752 8968
rect 303932 8916 303984 8968
rect 351036 8916 351088 8968
rect 577908 8916 577960 8968
rect 22412 8848 22464 8900
rect 161608 8848 161660 8900
rect 261888 8848 261940 8900
rect 309268 8848 309320 8900
rect 381672 8848 381724 8900
rect 254896 8780 254948 8832
rect 260416 8780 260468 8832
rect 308072 8780 308124 8832
rect 378084 8780 378136 8832
rect 158020 8576 158072 8628
rect 207976 8576 208028 8628
rect 272744 8576 272796 8628
rect 307980 8576 308032 8628
rect 374588 8576 374640 8628
rect 154432 8508 154484 8560
rect 211564 8508 211616 8560
rect 273940 8508 273992 8560
rect 306416 8508 306468 8560
rect 370816 8508 370868 8560
rect 184240 8372 184292 8424
rect 185344 8372 185396 8424
rect 215152 8372 215204 8424
rect 274400 8440 274452 8492
rect 306692 8440 306744 8492
rect 222512 8372 222564 8424
rect 218556 8304 218608 8356
rect 275320 8372 275372 8424
rect 305036 8372 305088 8424
rect 275412 8304 275464 8356
rect 305312 8304 305364 8356
rect 351036 8304 351088 8356
rect 351128 8304 351180 8356
rect 353060 8304 353112 8356
rect 363824 8440 363876 8492
rect 363916 8440 363968 8492
rect 367412 8440 367464 8492
rect 356188 8372 356240 8424
rect 370356 8372 370408 8424
rect 373116 8415 373168 8424
rect 373116 8381 373125 8415
rect 373125 8381 373159 8415
rect 373159 8381 373168 8415
rect 373116 8372 373168 8381
rect 374496 8372 374548 8424
rect 375692 8372 375744 8424
rect 399428 8372 399480 8424
rect 409180 8372 409232 8424
rect 438252 8372 438304 8424
rect 361156 8304 361208 8356
rect 361248 8304 361300 8356
rect 129500 8236 129552 8288
rect 256092 8236 256144 8288
rect 272836 8279 272888 8288
rect 272836 8245 272845 8279
rect 272845 8245 272879 8279
rect 272879 8245 272888 8279
rect 272836 8236 272888 8245
rect 310280 8236 310332 8288
rect 312672 8236 312724 8288
rect 337052 8236 337104 8288
rect 341284 8236 341336 8288
rect 506516 8236 506568 8288
rect 69976 8032 70028 8084
rect 244040 8032 244092 8084
rect 249652 8032 249704 8084
rect 280748 8032 280800 8084
rect 336960 8032 337012 8084
rect 341376 8032 341428 8084
rect 510104 8032 510156 8084
rect 66480 7964 66532 8016
rect 243580 7964 243632 8016
rect 245972 7964 246024 8016
rect 280840 7964 280892 8016
rect 333004 7964 333056 8016
rect 338156 7964 338208 8016
rect 338340 7964 338392 8016
rect 350852 7964 350904 8016
rect 513692 7964 513744 8016
rect 62892 7896 62944 7948
rect 242384 7896 242436 7948
rect 242476 7896 242528 7948
rect 279828 7896 279880 7948
rect 334292 7896 334344 7948
rect 339720 7896 339772 7948
rect 350668 7896 350720 7948
rect 517280 7896 517332 7948
rect 17720 7828 17772 7880
rect 196292 7828 196344 7880
rect 215796 7828 215848 7880
rect 215888 7828 215940 7880
rect 225272 7828 225324 7880
rect 225364 7828 225416 7880
rect 225456 7828 225508 7880
rect 225548 7828 225600 7880
rect 231252 7828 231304 7880
rect 231344 7828 231396 7880
rect 232540 7828 232592 7880
rect 237876 7828 237928 7880
rect 238888 7828 238940 7880
rect 279552 7828 279604 7880
rect 330060 7828 330112 7880
rect 338248 7828 338300 7880
rect 520868 7828 520920 7880
rect 12936 7760 12988 7812
rect 267040 7760 267092 7812
rect 327300 7760 327352 7812
rect 524364 7760 524416 7812
rect 4564 7692 4616 7744
rect 193624 7692 193676 7744
rect 193716 7692 193768 7744
rect 194912 7692 194964 7744
rect 265660 7692 265712 7744
rect 328680 7692 328732 7744
rect 527952 7692 528004 7744
rect 146152 7488 146204 7540
rect 260324 7488 260376 7540
rect 331716 7488 331768 7540
rect 332912 7488 332964 7540
rect 335672 7488 335724 7540
rect 340824 7488 340876 7540
rect 149740 7420 149792 7472
rect 260048 7420 260100 7472
rect 335580 7420 335632 7472
rect 340732 7420 340784 7472
rect 502928 7488 502980 7540
rect 520776 7488 520828 7540
rect 521972 7488 522024 7540
rect 537336 7488 537388 7540
rect 538624 7488 538676 7540
rect 555276 7488 555328 7540
rect 556472 7488 556524 7540
rect 563556 7488 563608 7540
rect 564844 7488 564896 7540
rect 581496 7488 581548 7540
rect 582692 7488 582744 7540
rect 499432 7420 499484 7472
rect 153236 7352 153288 7404
rect 261796 7352 261848 7404
rect 334384 7352 334436 7404
rect 343400 7352 343452 7404
rect 346988 7395 347040 7404
rect 346988 7361 346997 7395
rect 346997 7361 347031 7395
rect 347031 7361 347040 7395
rect 346988 7352 347040 7361
rect 356464 7352 356516 7404
rect 495844 7352 495896 7404
rect 156824 7284 156876 7336
rect 261704 7284 261756 7336
rect 331440 7284 331492 7336
rect 492256 7284 492308 7336
rect 160412 7216 160464 7268
rect 263268 7216 263320 7268
rect 317640 7216 317692 7268
rect 331164 7216 331216 7268
rect 488668 7216 488720 7268
rect 165196 7148 165248 7200
rect 264280 7148 264332 7200
rect 320308 7148 320360 7200
rect 330152 7148 330204 7200
rect 473856 7148 473908 7200
rect 474224 7148 474276 7200
rect 485080 7148 485132 7200
rect 486276 7148 486328 7200
rect 487472 7148 487524 7200
rect 569076 7148 569128 7200
rect 578644 7148 578696 7200
rect 168692 6944 168744 6996
rect 264188 6944 264240 6996
rect 331716 6944 331768 6996
rect 480388 6944 480440 6996
rect 480848 6944 480900 6996
rect 483516 6944 483568 6996
rect 558036 6944 558088 6996
rect 567604 6944 567656 6996
rect 172280 6876 172332 6928
rect 265752 6876 265804 6928
rect 278448 6876 278500 6928
rect 278724 6876 278776 6928
rect 322240 6876 322292 6928
rect 328588 6876 328640 6928
rect 476800 6876 476852 6928
rect 178260 6808 178312 6860
rect 266948 6808 267000 6860
rect 313500 6808 313552 6860
rect 405408 6808 405460 6860
rect 469624 6808 469676 6860
rect 174672 6740 174724 6792
rect 266028 6740 266080 6792
rect 314972 6740 315024 6792
rect 408996 6740 409048 6792
rect 424084 6740 424136 6792
rect 428960 6740 429012 6792
rect 473212 6740 473264 6792
rect 171084 6672 171136 6724
rect 265568 6672 265620 6724
rect 316352 6672 316404 6724
rect 412584 6672 412636 6724
rect 453248 6672 453300 6724
rect 462724 6672 462776 6724
rect 167588 6604 167640 6656
rect 264556 6604 264608 6656
rect 316260 6604 316312 6656
rect 416172 6604 416224 6656
rect 164000 6400 164052 6452
rect 263176 6400 263228 6452
rect 313592 6400 313644 6452
rect 131892 6332 131944 6384
rect 257380 6332 257432 6384
rect 270076 6332 270128 6384
rect 310740 6332 310792 6384
rect 317732 6400 317784 6452
rect 419668 6400 419720 6452
rect 318836 6332 318888 6384
rect 423256 6332 423308 6384
rect 59304 6264 59356 6316
rect 215796 6264 215848 6316
rect 235116 6264 235168 6316
rect 264004 6264 264056 6316
rect 310832 6264 310884 6316
rect 319020 6264 319072 6316
rect 55716 6196 55768 6248
rect 225180 6196 225232 6248
rect 225272 6196 225324 6248
rect 272652 6196 272704 6248
rect 302460 6196 302512 6248
rect 328680 6307 328732 6316
rect 328680 6273 328689 6307
rect 328689 6273 328723 6307
rect 328723 6273 328732 6307
rect 328680 6264 328732 6273
rect 337236 6264 337288 6316
rect 338800 6264 338852 6316
rect 346988 6307 347040 6316
rect 346988 6273 346997 6307
rect 346997 6273 347031 6307
rect 347031 6273 347040 6307
rect 346988 6264 347040 6273
rect 356464 6264 356516 6316
rect 430432 6196 430484 6248
rect 52128 6128 52180 6180
rect 215888 6128 215940 6180
rect 307796 6128 307848 6180
rect 370356 6128 370408 6180
rect 370448 6128 370500 6180
rect 434020 6128 434072 6180
rect 181848 6060 181900 6112
rect 267316 6060 267368 6112
rect 309360 6060 309412 6112
rect 321964 6060 322016 6112
rect 401820 6060 401872 6112
rect 426844 6060 426896 6112
rect 175868 5856 175920 5908
rect 185344 5856 185396 5908
rect 268420 5856 268472 5908
rect 312120 5856 312172 5908
rect 312212 5856 312264 5908
rect 398324 5856 398376 5908
rect 179456 5788 179508 5840
rect 188932 5788 188984 5840
rect 268328 5788 268380 5840
rect 394736 5788 394788 5840
rect 192520 5720 192572 5772
rect 269892 5720 269944 5772
rect 391148 5720 391200 5772
rect 269800 5652 269852 5704
rect 387560 5652 387612 5704
rect 199696 5584 199748 5636
rect 271272 5584 271324 5636
rect 312028 5584 312080 5636
rect 203192 5516 203244 5568
rect 271180 5516 271232 5568
rect 309452 5516 309504 5568
rect 371000 5584 371052 5636
rect 370908 5516 370960 5568
rect 191324 5312 191376 5364
rect 283600 5312 283652 5364
rect 301080 5312 301132 5364
rect 134284 5244 134336 5296
rect 244776 5244 244828 5296
rect 130696 5176 130748 5228
rect 244868 5176 244920 5228
rect 244960 5176 245012 5228
rect 264004 5244 264056 5296
rect 278264 5244 278316 5296
rect 299792 5244 299844 5296
rect 312580 5244 312632 5296
rect 341192 5312 341244 5364
rect 548192 5312 548244 5364
rect 338064 5244 338116 5296
rect 343584 5244 343636 5296
rect 345424 5244 345476 5296
rect 278724 5176 278776 5228
rect 296756 5176 296808 5228
rect 345976 5176 346028 5228
rect 8152 5108 8204 5160
rect 226928 5108 226980 5160
rect 227020 5108 227072 5160
rect 276516 5108 276568 5160
rect 296848 5108 296900 5160
rect 301264 5108 301316 5160
rect 302736 5108 302788 5160
rect 307520 5108 307572 5160
rect 342388 5108 342440 5160
rect 343952 5108 344004 5160
rect 551688 5244 551740 5296
rect 555276 5176 555328 5228
rect 346804 5108 346856 5160
rect 350852 5108 350904 5160
rect 350944 5108 350996 5160
rect 558864 5108 558916 5160
rect 2172 5040 2224 5092
rect 3368 4972 3420 5024
rect 275688 5040 275740 5092
rect 295652 5040 295704 5092
rect 302644 5040 302696 5092
rect 312212 5040 312264 5092
rect 331716 5040 331768 5092
rect 342572 5040 342624 5092
rect 345332 5040 345384 5092
rect 562452 5040 562504 5092
rect 229688 4972 229740 5024
rect 230148 4972 230200 5024
rect 230608 4972 230660 5024
rect 276976 4972 277028 5024
rect 300988 4972 301040 5024
rect 307520 4972 307572 5024
rect 335212 4972 335264 5024
rect 335764 4972 335816 5024
rect 566040 4972 566092 5024
rect 1068 4768 1120 4820
rect 225272 4768 225324 4820
rect 225364 4768 225416 4820
rect 275228 4768 275280 4820
rect 296940 4768 296992 4820
rect 301172 4768 301224 4820
rect 321964 4768 322016 4820
rect 322148 4768 322200 4820
rect 337604 4768 337656 4820
rect 339812 4768 339864 4820
rect 515256 4768 515308 4820
rect 515348 4768 515400 4820
rect 526756 4768 526808 4820
rect 195004 4700 195056 4752
rect 259128 4700 259180 4752
rect 279368 4700 279420 4752
rect 297032 4700 297084 4752
rect 338800 4700 338852 4752
rect 340916 4700 340968 4752
rect 198500 4632 198552 4684
rect 201996 4564 202048 4616
rect 264280 4564 264332 4616
rect 283508 4632 283560 4684
rect 299884 4632 299936 4684
rect 312304 4632 312356 4684
rect 334108 4632 334160 4684
rect 337144 4632 337196 4684
rect 274124 4564 274176 4616
rect 299700 4564 299752 4616
rect 205584 4496 205636 4548
rect 264372 4496 264424 4548
rect 269708 4496 269760 4548
rect 269800 4496 269852 4548
rect 272468 4496 272520 4548
rect 298412 4496 298464 4548
rect 302552 4496 302604 4548
rect 302828 4496 302880 4548
rect 209172 4428 209224 4480
rect 264188 4428 264240 4480
rect 264280 4428 264332 4480
rect 270996 4428 271048 4480
rect 298504 4428 298556 4480
rect 330520 4564 330572 4616
rect 344780 4564 344832 4616
rect 347908 4700 347960 4752
rect 350576 4700 350628 4752
rect 350944 4700 350996 4752
rect 544604 4700 544656 4752
rect 346712 4632 346764 4684
rect 350668 4632 350720 4684
rect 350852 4632 350904 4684
rect 569536 4700 569588 4752
rect 541016 4564 541068 4616
rect 303104 4496 303156 4548
rect 328128 4496 328180 4548
rect 533932 4496 533984 4548
rect 303012 4428 303064 4480
rect 326932 4428 326984 4480
rect 530344 4428 530396 4480
rect 128856 4224 128908 4276
rect 218648 4224 218700 4276
rect 186816 4156 186868 4208
rect 196384 4156 196436 4208
rect 196476 4156 196528 4208
rect 206044 4156 206096 4208
rect 212760 4156 212812 4208
rect 274216 4224 274268 4276
rect 288844 4224 288896 4276
rect 298228 4224 298280 4276
rect 302644 4224 302696 4276
rect 324540 4224 324592 4276
rect 336684 4224 336736 4276
rect 339444 4224 339496 4276
rect 515348 4224 515400 4276
rect 58108 4088 58160 4140
rect 235116 4088 235168 4140
rect 235300 4088 235352 4140
rect 236404 4088 236456 4140
rect 236496 4088 236548 4140
rect 237784 4088 237836 4140
rect 238060 4088 238112 4140
rect 242752 4088 242804 4140
rect 244868 4088 244920 4140
rect 246064 4088 246116 4140
rect 251952 4088 252004 4140
rect 252964 4088 253016 4140
rect 260324 4088 260376 4140
rect 261244 4088 261296 4140
rect 271364 4156 271416 4208
rect 269800 4088 269852 4140
rect 51024 4020 51076 4072
rect 228124 4020 228176 4072
rect 228216 4020 228268 4072
rect 229504 4020 229556 4072
rect 230148 4020 230200 4072
rect 47436 3952 47488 4004
rect 133088 3952 133140 4004
rect 134192 3952 134244 4004
rect 137688 3952 137740 4004
rect 137780 3952 137832 4004
rect 138056 3952 138108 4004
rect 215796 3952 215848 4004
rect 215888 3952 215940 4004
rect 217544 3952 217596 4004
rect 218464 3952 218516 4004
rect 219752 3952 219804 4004
rect 235668 4020 235720 4072
rect 237968 4020 238020 4072
rect 241280 4020 241332 4072
rect 268604 4020 268656 4072
rect 284152 4088 284204 4140
rect 285440 4088 285492 4140
rect 287648 4088 287700 4140
rect 298320 4156 298372 4208
rect 302460 4156 302512 4208
rect 288844 4088 288896 4140
rect 289396 4088 289448 4140
rect 289580 4088 289632 4140
rect 290040 4088 290092 4140
rect 291512 4088 291564 4140
rect 292432 4088 292484 4140
rect 293904 4088 293956 4140
rect 297216 4088 297268 4140
rect 323344 4156 323396 4208
rect 338432 4156 338484 4208
rect 537428 4224 537480 4276
rect 305496 4088 305548 4140
rect 319756 4088 319808 4140
rect 320584 4088 320636 4140
rect 284980 4020 285032 4072
rect 294272 4020 294324 4072
rect 302552 4020 302604 4072
rect 302736 4020 302788 4072
rect 320952 4020 321004 4072
rect 418840 4088 418892 4140
rect 523168 4156 523220 4208
rect 578000 4088 578052 4140
rect 579104 4088 579156 4140
rect 579380 4088 579432 4140
rect 580300 4088 580352 4140
rect 436320 4020 436372 4072
rect 512496 4020 512548 4072
rect 239348 3952 239400 4004
rect 267500 3952 267552 4004
rect 284888 3952 284940 4004
rect 286452 3952 286504 4004
rect 289120 3952 289172 4004
rect 295100 3952 295152 4004
rect 46240 3884 46292 3936
rect 266304 3884 266356 3936
rect 284060 3884 284112 3936
rect 285256 3884 285308 3936
rect 292800 3884 292852 3936
rect 298412 3884 298464 3936
rect 304300 3952 304352 4004
rect 321872 3952 321924 4004
rect 439908 3952 439960 4004
rect 516084 3952 516136 4004
rect 320492 3884 320544 3936
rect 322976 3884 323028 3936
rect 324264 3884 324316 3936
rect 443496 3884 443548 3936
rect 42652 3680 42704 3732
rect 230424 3680 230476 3732
rect 235208 3680 235260 3732
rect 239716 3680 239768 3732
rect 254804 3680 254856 3732
rect 263912 3680 263964 3732
rect 283692 3680 283744 3732
rect 292892 3680 292944 3732
rect 299608 3680 299660 3732
rect 311476 3680 311528 3732
rect 324632 3680 324684 3732
rect 447084 3680 447136 3732
rect 38972 3612 39024 3664
rect 29588 3544 29640 3596
rect 30784 3544 30836 3596
rect 36672 3544 36724 3596
rect 37684 3544 37736 3596
rect 37868 3544 37920 3596
rect 39064 3544 39116 3596
rect 43848 3544 43900 3596
rect 44584 3544 44636 3596
rect 138976 3612 139028 3664
rect 139804 3612 139856 3664
rect 141368 3612 141420 3664
rect 142564 3612 142616 3664
rect 148544 3612 148596 3664
rect 149464 3612 149516 3664
rect 159216 3612 159268 3664
rect 160504 3612 160556 3664
rect 162804 3612 162856 3664
rect 163264 3612 163316 3664
rect 166392 3612 166444 3664
rect 167220 3612 167272 3664
rect 10544 3476 10596 3528
rect 11464 3476 11516 3528
rect 11740 3476 11792 3528
rect 12844 3476 12896 3528
rect 18824 3476 18876 3528
rect 19744 3476 19796 3528
rect 20020 3476 20072 3528
rect 21124 3476 21176 3528
rect 34372 3476 34424 3528
rect 34924 3476 34976 3528
rect 35476 3476 35528 3528
rect 81936 3476 81988 3528
rect 83040 3476 83092 3528
rect 93804 3476 93856 3528
rect 94264 3476 94316 3528
rect 95000 3476 95052 3528
rect 95644 3476 95696 3528
rect 96196 3476 96248 3528
rect 97024 3476 97076 3528
rect 98588 3476 98640 3528
rect 99784 3476 99836 3528
rect 99692 3408 99744 3460
rect 103832 3408 103884 3460
rect 113860 3408 113912 3460
rect 114044 3476 114096 3528
rect 114964 3476 115016 3528
rect 115240 3476 115292 3528
rect 116344 3476 116396 3528
rect 116436 3476 116488 3528
rect 117448 3476 117500 3528
rect 119932 3476 119984 3528
rect 120484 3476 120536 3528
rect 121128 3476 121180 3528
rect 121864 3476 121916 3528
rect 123520 3476 123572 3528
rect 124624 3476 124676 3528
rect 124716 3476 124768 3528
rect 125820 3476 125872 3528
rect 126096 3476 126148 3528
rect 128304 3476 128356 3528
rect 128764 3476 128816 3528
rect 138424 3476 138476 3528
rect 157652 3476 157704 3528
rect 128856 3408 128908 3460
rect 210276 3612 210328 3664
rect 215796 3612 215848 3664
rect 220028 3612 220080 3664
rect 224536 3612 224588 3664
rect 225180 3612 225232 3664
rect 225456 3612 225508 3664
rect 234840 3612 234892 3664
rect 234932 3612 234984 3664
rect 225640 3544 225692 3596
rect 234748 3544 234800 3596
rect 235392 3544 235444 3596
rect 238428 3544 238480 3596
rect 158112 3408 158164 3460
rect 186540 3408 186592 3460
rect 206228 3476 206280 3528
rect 236680 3476 236732 3528
rect 236772 3476 236824 3528
rect 241096 3476 241148 3528
rect 243672 3612 243724 3664
rect 247260 3612 247312 3664
rect 273388 3544 273440 3596
rect 278448 3544 278500 3596
rect 285164 3612 285216 3664
rect 285256 3612 285308 3664
rect 289672 3612 289724 3664
rect 295744 3612 295796 3664
rect 313868 3612 313920 3664
rect 323252 3612 323304 3664
rect 450672 3612 450724 3664
rect 281024 3544 281076 3596
rect 282956 3544 283008 3596
rect 287924 3544 287976 3596
rect 297124 3544 297176 3596
rect 265108 3476 265160 3528
rect 282312 3476 282364 3528
rect 292708 3476 292760 3528
rect 300804 3476 300856 3528
rect 307888 3544 307940 3596
rect 309544 3544 309596 3596
rect 370632 3544 370684 3596
rect 454168 3544 454220 3596
rect 318560 3476 318612 3528
rect 321780 3476 321832 3528
rect 326104 3476 326156 3528
rect 341468 3476 341520 3528
rect 351128 3476 351180 3528
rect 360512 3476 360564 3528
rect 360604 3476 360656 3528
rect 360788 3476 360840 3528
rect 370172 3476 370224 3528
rect 370264 3476 370316 3528
rect 370540 3476 370592 3528
rect 457756 3476 457808 3528
rect 186816 3408 186868 3460
rect 196292 3408 196344 3460
rect 196384 3408 196436 3460
rect 196476 3408 196528 3460
rect 206044 3408 206096 3460
rect 254712 3408 254764 3460
rect 261520 3408 261572 3460
rect 262624 3408 262676 3460
rect 33176 3340 33228 3392
rect 40260 3340 40312 3392
rect 45044 3340 45096 3392
rect 45964 3340 46016 3392
rect 61696 3340 61748 3392
rect 62524 3340 62576 3392
rect 64088 3340 64140 3392
rect 65192 3340 65244 3392
rect 65284 3340 65336 3392
rect 235116 3340 235168 3392
rect 235208 3340 235260 3392
rect 237048 3340 237100 3392
rect 237140 3340 237192 3392
rect 243856 3340 243908 3392
rect 257932 3340 257984 3392
rect 275780 3408 275832 3460
rect 262900 3340 262952 3392
rect 272192 3340 272244 3392
rect 280104 3408 280156 3460
rect 288108 3408 288160 3460
rect 291420 3408 291472 3460
rect 293628 3408 293680 3460
rect 294364 3408 294416 3460
rect 310280 3408 310332 3460
rect 310924 3408 310976 3460
rect 389952 3408 390004 3460
rect 461344 3408 461396 3460
rect 286728 3340 286780 3392
rect 293720 3340 293772 3392
rect 303104 3340 303156 3392
rect 319112 3340 319164 3392
rect 429236 3340 429288 3392
rect 433836 3340 433888 3392
rect 451684 3340 451736 3392
rect 466588 3340 466640 3392
rect 480664 3340 480716 3392
rect 28392 3136 28444 3188
rect 29404 3136 29456 3188
rect 68780 3136 68832 3188
rect 69424 3136 69476 3188
rect 71172 3136 71224 3188
rect 72184 3136 72236 3188
rect 72368 3136 72420 3188
rect 21216 3068 21268 3120
rect 22504 3068 22556 3120
rect 77152 3068 77204 3120
rect 77704 3068 77756 3120
rect 78348 3068 78400 3120
rect 79084 3068 79136 3120
rect 80740 3068 80792 3120
rect 81844 3068 81896 3120
rect 79544 3000 79596 3052
rect 187184 3136 187236 3188
rect 196200 3136 196252 3188
rect 196752 3136 196804 3188
rect 205860 3136 205912 3188
rect 245144 3136 245196 3188
rect 253148 3136 253200 3188
rect 254160 3136 254212 3188
rect 270996 3136 271048 3188
rect 246616 3068 246668 3120
rect 278172 3136 278224 3188
rect 286820 3136 286872 3188
rect 294088 3136 294140 3188
rect 319204 3136 319256 3188
rect 425648 3136 425700 3188
rect 285532 3068 285584 3120
rect 292340 3068 292392 3120
rect 296020 3068 296072 3120
rect 317824 3068 317876 3120
rect 422060 3068 422112 3120
rect 85432 3000 85484 3052
rect 85984 3000 86036 3052
rect 86628 3000 86680 3052
rect 87364 3000 87416 3052
rect 87824 3000 87876 3052
rect 88744 3000 88796 3052
rect 89020 3000 89072 3052
rect 90124 3000 90176 3052
rect 99508 3000 99560 3052
rect 99784 3000 99836 3052
rect 102084 3000 102136 3052
rect 102544 3000 102596 3052
rect 54520 2932 54572 2984
rect 55624 2932 55676 2984
rect 90216 2932 90268 2984
rect 186816 3000 186868 3052
rect 207700 3000 207752 3052
rect 247904 3000 247956 3052
rect 250848 3000 250900 3052
rect 251584 3000 251636 3052
rect 286360 3000 286412 3052
rect 294180 3000 294232 3052
rect 105672 2932 105724 2984
rect 106684 2932 106736 2984
rect 106868 2932 106920 2984
rect 107972 2932 108024 2984
rect 103280 2864 103332 2916
rect 103924 2864 103976 2916
rect 104476 2864 104528 2916
rect 97392 2796 97444 2848
rect 111652 2864 111704 2916
rect 112848 2796 112900 2848
rect 113308 2796 113360 2848
rect 187092 2932 187144 2984
rect 195924 2932 195976 2984
rect 250664 2932 250716 2984
rect 274584 2932 274636 2984
rect 286636 2932 286688 2984
rect 291604 2932 291656 2984
rect 294824 2932 294876 2984
rect 252136 2864 252188 2916
rect 276976 2864 277028 2916
rect 279920 2864 279972 2916
rect 280564 2864 280616 2916
rect 283968 2864 284020 2916
rect 292984 2864 293036 2916
rect 301908 2864 301960 2916
rect 316444 3000 316496 3052
rect 418472 3000 418524 3052
rect 432824 3068 432876 3120
rect 315064 2932 315116 2984
rect 355268 2975 355320 2984
rect 355268 2941 355277 2975
rect 355277 2941 355311 2975
rect 355311 2941 355320 2975
rect 355268 2932 355320 2941
rect 306692 2864 306744 2916
rect 313684 2864 313736 2916
rect 406880 2932 406932 2984
rect 411664 2932 411716 2984
rect 414608 2932 414660 2984
rect 424084 2932 424136 2984
rect 196384 2796 196436 2848
rect 253424 2796 253476 2848
rect 279276 2796 279328 2848
rect 281760 2796 281812 2848
rect 288200 2796 288252 2848
rect 293812 2796 293864 2848
rect 308256 2796 308308 2848
rect 311936 2796 311988 2848
rect 364652 2796 364704 2848
rect 364744 2839 364796 2848
rect 364744 2805 364753 2839
rect 364753 2805 364787 2839
rect 364787 2805 364796 2839
rect 364744 2796 364796 2805
rect 364928 2839 364980 2848
rect 364928 2805 364937 2839
rect 364937 2805 364971 2839
rect 364971 2805 364980 2839
rect 364928 2796 364980 2805
rect 365112 2796 365164 2848
rect 397128 2796 397180 2848
rect 411388 2864 411440 2916
rect 404212 2796 404264 2848
rect 420036 2796 420088 2848
rect 122324 2592 122376 2644
rect 196108 2635 196160 2644
rect 196108 2601 196117 2635
rect 196117 2601 196151 2635
rect 196151 2601 196160 2635
rect 196108 2592 196160 2601
rect 220028 2592 220080 2644
rect 223432 2592 223484 2644
rect 346344 2592 346396 2644
rect 118736 2524 118788 2576
rect 358028 2592 358080 2644
rect 359040 2592 359092 2644
rect 360696 2592 360748 2644
rect 361432 2592 361484 2644
rect 362076 2592 362128 2644
rect 362628 2592 362680 2644
rect 382868 2592 382920 2644
rect 380476 2456 380528 2508
rect 349656 2388 349708 2440
rect 350760 2388 350812 2440
rect 384064 2388 384116 2440
rect 356556 1368 356608 1420
rect 357844 1368 357896 1420
rect 353796 1096 353848 1148
rect 354256 1096 354308 1148
rect 5760 552 5812 604
rect 5944 552 5996 604
rect 23608 552 23660 604
rect 23884 552 23936 604
rect 74760 552 74812 604
rect 74944 552 74996 604
rect 152040 552 152092 604
rect 152132 552 152184 604
rect 155628 552 155680 604
rect 156364 552 156416 604
rect 169888 552 169940 604
rect 169980 552 170032 604
rect 173476 552 173528 604
rect 174304 552 174356 604
rect 180652 552 180704 604
rect 181204 552 181256 604
rect 183044 552 183096 604
rect 183964 552 184016 604
rect 190128 552 190180 604
rect 190404 552 190456 604
rect 197304 552 197356 604
rect 197764 552 197816 604
rect 200892 552 200944 604
rect 201904 552 201956 604
rect 221040 552 221092 604
rect 221224 552 221276 604
rect 231804 552 231856 604
rect 231988 552 232040 604
rect 234196 552 234248 604
rect 248456 552 248508 604
rect 248824 552 248876 604
rect 256736 552 256788 604
rect 257104 552 257156 604
rect 290592 552 290644 604
rect 291236 552 291288 604
rect 309084 595 309136 604
rect 309084 561 309093 595
rect 309093 561 309127 595
rect 309127 561 309136 595
rect 309084 552 309136 561
rect 324816 552 324868 604
rect 325736 552 325788 604
rect 378636 552 378688 604
rect 379280 552 379332 604
rect 395196 552 395248 604
rect 395932 552 395984 604
rect 402096 552 402148 604
rect 403016 552 403068 604
rect 406236 552 406288 604
rect 406604 552 406656 604
rect 420864 595 420916 604
rect 420864 561 420873 595
rect 420873 561 420907 595
rect 420907 561 420916 595
rect 420864 552 420916 561
rect 424176 552 424228 604
rect 424452 552 424504 604
rect 426936 552 426988 604
rect 428040 552 428092 604
rect 431076 552 431128 604
rect 431628 552 431680 604
rect 442116 552 442168 604
rect 442300 552 442352 604
rect 443588 552 443640 604
rect 444692 552 444744 604
rect 444876 552 444928 604
rect 445888 552 445940 604
rect 447636 552 447688 604
rect 448280 552 448332 604
rect 449016 552 449068 604
rect 449476 552 449528 604
rect 451868 552 451920 604
rect 452972 552 453024 604
rect 454536 552 454588 604
rect 455364 552 455416 604
rect 461436 552 461488 604
rect 462540 552 462592 604
rect 462816 552 462868 604
rect 463736 552 463788 604
rect 465576 552 465628 604
rect 466128 552 466180 604
rect 466956 552 467008 604
rect 467324 552 467376 604
rect 469716 552 469768 604
rect 470820 552 470872 604
rect 490416 552 490468 604
rect 491060 552 491112 604
rect 495936 552 495988 604
rect 497040 552 497092 604
rect 497316 552 497368 604
rect 498236 552 498288 604
rect 500076 552 500128 604
rect 500628 552 500680 604
rect 501456 552 501508 604
rect 501732 552 501784 604
rect 504216 552 504268 604
rect 505320 552 505372 604
rect 506976 552 507028 604
rect 507712 552 507764 604
rect 508356 552 508408 604
rect 508908 552 508960 604
rect 529148 552 529200 604
rect 529240 552 529292 604
<< metal2 >>
rect 11278 703520 11334 704000
rect 32898 703520 32954 704000
rect 54518 703520 54574 704000
rect 76138 703520 76194 704000
rect 97758 703520 97814 704000
rect 119378 703520 119434 704000
rect 140998 703520 141054 704000
rect 162618 703520 162674 704000
rect 184238 703520 184294 704000
rect 205950 703520 206006 704000
rect 227570 703520 227626 704000
rect 249190 703520 249246 704000
rect 270810 703520 270866 704000
rect 292430 703520 292486 704000
rect 314050 703520 314106 704000
rect 335670 703520 335726 704000
rect 357290 703520 357346 704000
rect 378910 703520 378966 704000
rect 400622 703520 400678 704000
rect 422242 703520 422298 704000
rect 443862 703520 443918 704000
rect 465482 703520 465538 704000
rect 487102 703520 487158 704000
rect 508722 703520 508778 704000
rect 530342 703520 530398 704000
rect 551962 703520 552018 704000
rect 573582 703520 573638 704000
rect 11292 700369 11320 703520
rect 11278 700360 11334 700369
rect 32912 700330 32940 703520
rect 54532 700534 54560 703520
rect 76152 700602 76180 703520
rect 97772 700806 97800 703520
rect 119392 701010 119420 703520
rect 119380 701004 119432 701010
rect 119380 700946 119432 700952
rect 97760 700800 97812 700806
rect 97760 700742 97812 700748
rect 76140 700596 76192 700602
rect 76140 700538 76192 700544
rect 54520 700528 54572 700534
rect 54520 700470 54572 700476
rect 11278 700295 11334 700304
rect 32900 700324 32952 700330
rect 32900 700266 32952 700272
rect 141012 700262 141040 703520
rect 141000 700256 141052 700262
rect 141000 700198 141052 700204
rect 162632 700058 162660 703520
rect 184252 700874 184280 703520
rect 184240 700868 184292 700874
rect 184240 700810 184292 700816
rect 185344 700868 185396 700874
rect 185344 700810 185396 700816
rect 162620 700052 162672 700058
rect 162620 699994 162672 700000
rect 3734 695464 3790 695473
rect 3734 695399 3790 695408
rect 3748 694278 3776 695399
rect 3736 694272 3788 694278
rect 3736 694214 3788 694220
rect 3918 678736 3974 678745
rect 3918 678671 3974 678680
rect 3932 677618 3960 678671
rect 3920 677612 3972 677618
rect 3920 677554 3972 677560
rect 3918 662008 3974 662017
rect 3918 661943 3974 661952
rect 3932 661094 3960 661943
rect 3920 661088 3972 661094
rect 3920 661030 3972 661036
rect 3550 645280 3606 645289
rect 3550 645215 3606 645224
rect 3564 644502 3592 645215
rect 3552 644496 3604 644502
rect 3552 644438 3604 644444
rect 3918 628416 3974 628425
rect 3918 628351 3974 628360
rect 3932 627978 3960 628351
rect 3920 627972 3972 627978
rect 3920 627914 3972 627920
rect 3826 611688 3882 611697
rect 3826 611623 3882 611632
rect 3840 611386 3868 611623
rect 3828 611380 3880 611386
rect 3828 611322 3880 611328
rect 3918 594960 3974 594969
rect 3918 594895 3974 594904
rect 3932 594862 3960 594895
rect 3920 594856 3972 594862
rect 3920 594798 3972 594804
rect 3734 578232 3790 578241
rect 3734 578167 3790 578176
rect 3748 576910 3776 578167
rect 3736 576904 3788 576910
rect 3736 576846 3788 576852
rect 3918 561368 3974 561377
rect 3918 561303 3974 561312
rect 3932 560454 3960 561303
rect 3920 560448 3972 560454
rect 3920 560390 3972 560396
rect 3642 544640 3698 544649
rect 3642 544575 3698 544584
rect 3656 543794 3684 544575
rect 3644 543788 3696 543794
rect 3644 543730 3696 543736
rect 3642 527912 3698 527921
rect 3642 527847 3698 527856
rect 3656 527270 3684 527847
rect 3644 527264 3696 527270
rect 3644 527206 3696 527212
rect 4010 511184 4066 511193
rect 4010 511119 4066 511128
rect 4024 510678 4052 511119
rect 4012 510672 4064 510678
rect 4012 510614 4064 510620
rect 3734 494320 3790 494329
rect 3734 494255 3790 494264
rect 3748 494086 3776 494255
rect 3736 494080 3788 494086
rect 3736 494022 3788 494028
rect 3918 477592 3974 477601
rect 3918 477527 3920 477536
rect 3972 477527 3974 477536
rect 3920 477498 3972 477504
rect 185356 463282 185384 700810
rect 205964 699854 205992 703520
rect 205952 699848 206004 699854
rect 205952 699790 206004 699796
rect 227584 699786 227612 703520
rect 249204 700942 249232 703520
rect 249192 700936 249244 700942
rect 249192 700878 249244 700884
rect 250204 700936 250256 700942
rect 250204 700878 250256 700884
rect 227572 699780 227624 699786
rect 227572 699722 227624 699728
rect 185344 463276 185396 463282
rect 185344 463218 185396 463224
rect 250216 463214 250244 700878
rect 270824 699990 270852 703520
rect 284704 700936 284756 700942
rect 284704 700878 284756 700884
rect 280564 700460 280616 700466
rect 280564 700402 280616 700408
rect 280472 700392 280524 700398
rect 280472 700334 280524 700340
rect 270812 699984 270864 699990
rect 270812 699926 270864 699932
rect 276424 695564 276476 695570
rect 276424 695506 276476 695512
rect 275044 663808 275096 663814
rect 275044 663750 275096 663756
rect 273664 648644 273716 648650
rect 273664 648586 273716 648592
rect 272284 617024 272336 617030
rect 272284 616966 272336 616972
rect 270904 601792 270956 601798
rect 270904 601734 270956 601740
rect 270812 586560 270864 586566
rect 270812 586502 270864 586508
rect 269524 569968 269576 569974
rect 269524 569910 269576 569916
rect 266764 554804 266816 554810
rect 266764 554746 266816 554752
rect 266672 523048 266724 523054
rect 266672 522990 266724 522996
rect 264004 507884 264056 507890
rect 264004 507826 264056 507832
rect 262624 476128 262676 476134
rect 262624 476070 262676 476076
rect 257104 463616 257156 463622
rect 257104 463558 257156 463564
rect 253976 463344 254028 463350
rect 253976 463286 254028 463292
rect 250204 463208 250256 463214
rect 250204 463150 250256 463156
rect 4380 462800 4432 462806
rect 4380 462742 4432 462748
rect 4288 462732 4340 462738
rect 4288 462674 4340 462680
rect 4196 462664 4248 462670
rect 4196 462606 4248 462612
rect 4012 462596 4064 462602
rect 4012 462538 4064 462544
rect 3918 462496 3974 462505
rect 3918 462431 3974 462440
rect 3642 460864 3698 460873
rect 3642 460799 3698 460808
rect 3656 459814 3684 460799
rect 3644 459808 3696 459814
rect 3644 459750 3696 459756
rect 3644 444168 3696 444174
rect 3642 444136 3644 444145
rect 3696 444136 3698 444145
rect 3642 444071 3698 444080
rect 3644 427780 3696 427786
rect 3644 427722 3696 427728
rect 3656 427281 3684 427722
rect 3642 427272 3698 427281
rect 3642 427207 3698 427216
rect 3828 411188 3880 411194
rect 3828 411130 3880 411136
rect 3840 410553 3868 411130
rect 3826 410544 3882 410553
rect 3826 410479 3882 410488
rect 3828 394664 3880 394670
rect 3828 394606 3880 394612
rect 3840 393825 3868 394606
rect 3826 393816 3882 393825
rect 3826 393751 3882 393760
rect 3552 378004 3604 378010
rect 3552 377946 3604 377952
rect 3564 377097 3592 377946
rect 3550 377088 3606 377097
rect 3550 377023 3606 377032
rect 3828 361548 3880 361554
rect 3828 361490 3880 361496
rect 3840 360369 3868 361490
rect 3826 360360 3882 360369
rect 3826 360295 3882 360304
rect 3828 343596 3880 343602
rect 3828 343538 3880 343544
rect 3840 343505 3868 343538
rect 3826 343496 3882 343505
rect 3826 343431 3882 343440
rect 3644 310480 3696 310486
rect 3644 310422 3696 310428
rect 3656 310049 3684 310422
rect 3642 310040 3698 310049
rect 3642 309975 3698 309984
rect 3552 293888 3604 293894
rect 3552 293830 3604 293836
rect 3564 293321 3592 293830
rect 3550 293312 3606 293321
rect 3550 293247 3606 293256
rect 3828 260840 3880 260846
rect 3828 260782 3880 260788
rect 3840 259729 3868 260782
rect 3826 259720 3882 259729
rect 3826 259655 3882 259664
rect 3828 244180 3880 244186
rect 3828 244122 3880 244128
rect 3840 243001 3868 244122
rect 3826 242992 3882 243001
rect 3826 242927 3882 242936
rect 3736 209772 3788 209778
rect 3736 209714 3788 209720
rect 3748 209409 3776 209714
rect 3734 209400 3790 209409
rect 3734 209335 3790 209344
rect 3828 192704 3880 192710
rect 3826 192672 3828 192681
rect 3880 192672 3882 192681
rect 3826 192607 3882 192616
rect 3932 108905 3960 462431
rect 4024 159225 4052 462538
rect 4104 462528 4156 462534
rect 4104 462470 4156 462476
rect 4116 175953 4144 462470
rect 4208 226273 4236 462606
rect 4300 276457 4328 462674
rect 4392 326777 4420 462742
rect 228952 461576 229004 461582
rect 228952 461518 229004 461524
rect 220580 461508 220632 461514
rect 220580 461450 220632 461456
rect 179180 461100 179232 461106
rect 179180 461042 179232 461048
rect 6772 461032 6824 461038
rect 6772 460974 6824 460980
rect 6680 458380 6732 458386
rect 6680 458322 6732 458328
rect 5942 337376 5998 337385
rect 5942 337311 5998 337320
rect 4378 326768 4434 326777
rect 4378 326703 4434 326712
rect 4286 276448 4342 276457
rect 4286 276383 4342 276392
rect 4194 226264 4250 226273
rect 4194 226199 4250 226208
rect 4102 175944 4158 175953
rect 4102 175879 4158 175888
rect 4010 159216 4066 159225
rect 4010 159151 4066 159160
rect 4012 143540 4064 143546
rect 4012 143482 4064 143488
rect 4024 142361 4052 143482
rect 4010 142352 4066 142361
rect 4010 142287 4066 142296
rect 4010 126984 4066 126993
rect 4010 126919 4066 126928
rect 4024 125633 4052 126919
rect 4010 125624 4066 125633
rect 4010 125559 4066 125568
rect 3918 108896 3974 108905
rect 3918 108831 3974 108840
rect 3644 59220 3696 59226
rect 3644 59162 3696 59168
rect 3656 58585 3684 59162
rect 3642 58576 3698 58585
rect 3642 58511 3698 58520
rect 3918 42800 3974 42809
rect 3918 42735 3974 42744
rect 3932 41857 3960 42735
rect 3918 41848 3974 41857
rect 3918 41783 3974 41792
rect 3920 26240 3972 26246
rect 3920 26182 3972 26188
rect 3932 25129 3960 26182
rect 3918 25120 3974 25129
rect 3918 25055 3974 25064
rect 3918 9616 3974 9625
rect 3918 9551 3974 9560
rect 3932 8401 3960 9551
rect 3918 8392 3974 8401
rect 3918 8327 3974 8336
rect 4564 7744 4616 7750
rect 4564 7686 4616 7692
rect 2172 5092 2224 5098
rect 2172 5034 2224 5040
rect 1068 4820 1120 4826
rect 1068 4762 1120 4768
rect 1080 480 1108 4762
rect 2184 480 2212 5034
rect 3368 5024 3420 5030
rect 3368 4966 3420 4972
rect 3380 480 3408 4966
rect 4576 480 4604 7686
rect 5956 610 5984 337311
rect 6692 293894 6720 458322
rect 6784 444174 6812 460974
rect 9440 458312 9492 458318
rect 9440 458254 9492 458260
rect 6772 444168 6824 444174
rect 6772 444110 6824 444116
rect 6680 293888 6732 293894
rect 6680 293830 6732 293836
rect 9452 192710 9480 458254
rect 129224 338156 129276 338162
rect 129224 338098 129276 338104
rect 142564 338156 142616 338162
rect 142564 338098 142616 338104
rect 152224 338156 152276 338162
rect 152224 338098 152276 338104
rect 161884 338156 161936 338162
rect 161884 338098 161936 338104
rect 171544 338156 171596 338162
rect 171544 338098 171596 338104
rect 62524 338088 62576 338094
rect 62524 338030 62576 338036
rect 45964 338020 46016 338026
rect 45964 337962 46016 337968
rect 55624 338020 55676 338026
rect 55624 337962 55676 337968
rect 44584 337952 44636 337958
rect 44584 337894 44636 337900
rect 22504 337748 22556 337754
rect 22504 337690 22556 337696
rect 37684 337748 37736 337754
rect 37684 337690 37736 337696
rect 12844 337544 12896 337550
rect 12844 337486 12896 337492
rect 11464 337408 11516 337414
rect 11464 337350 11516 337356
rect 9440 192704 9492 192710
rect 9440 192646 9492 192652
rect 9348 8968 9400 8974
rect 9348 8910 9400 8916
rect 8152 5160 8204 5166
rect 8152 5102 8204 5108
rect 6954 3360 7010 3369
rect 6954 3295 7010 3304
rect 5760 604 5812 610
rect 5760 546 5812 552
rect 5944 604 5996 610
rect 5944 546 5996 552
rect 5772 480 5800 546
rect 6968 480 6996 3295
rect 8164 480 8192 5102
rect 9360 480 9388 8910
rect 11476 3534 11504 337350
rect 12856 3534 12884 337486
rect 21124 337476 21176 337482
rect 21124 337418 21176 337424
rect 14224 312588 14276 312594
rect 14224 312530 14276 312536
rect 12936 7812 12988 7818
rect 12936 7754 12988 7760
rect 10544 3528 10596 3534
rect 10544 3470 10596 3476
rect 11464 3528 11516 3534
rect 11464 3470 11516 3476
rect 11740 3528 11792 3534
rect 11740 3470 11792 3476
rect 12844 3528 12896 3534
rect 12844 3470 12896 3476
rect 10556 480 10584 3470
rect 11752 480 11780 3470
rect 12948 480 12976 7754
rect 14236 626 14264 312530
rect 19744 273964 19796 273970
rect 19744 273906 19796 273912
rect 17720 7880 17772 7886
rect 17720 7822 17772 7828
rect 16522 3632 16578 3641
rect 16522 3567 16578 3576
rect 15326 3496 15382 3505
rect 15326 3431 15382 3440
rect 14144 598 14264 626
rect 14144 480 14172 598
rect 15340 480 15368 3431
rect 16536 480 16564 3567
rect 17732 480 17760 7822
rect 19756 3534 19784 273906
rect 21136 3534 21164 337418
rect 22412 8900 22464 8906
rect 22412 8842 22464 8848
rect 18824 3528 18876 3534
rect 18824 3470 18876 3476
rect 19744 3528 19796 3534
rect 19744 3470 19796 3476
rect 20020 3528 20072 3534
rect 20020 3470 20072 3476
rect 21124 3528 21176 3534
rect 21124 3470 21176 3476
rect 18836 480 18864 3470
rect 20032 480 20060 3470
rect 21216 3120 21268 3126
rect 21216 3062 21268 3068
rect 21228 480 21256 3062
rect 22424 480 22452 8842
rect 22516 3126 22544 337690
rect 30784 337680 30836 337686
rect 30784 337622 30836 337628
rect 26644 337408 26696 337414
rect 26644 337350 26696 337356
rect 26656 337210 26684 337350
rect 26644 337204 26696 337210
rect 26644 337146 26696 337152
rect 23884 330540 23936 330546
rect 23884 330482 23936 330488
rect 22504 3120 22556 3126
rect 22504 3062 22556 3068
rect 23896 610 23924 330482
rect 29404 297424 29456 297430
rect 29404 297366 29456 297372
rect 27196 9104 27248 9110
rect 27196 9046 27248 9052
rect 25998 3904 26054 3913
rect 25998 3839 26054 3848
rect 24802 3768 24858 3777
rect 24802 3703 24858 3712
rect 23608 604 23660 610
rect 23608 546 23660 552
rect 23884 604 23936 610
rect 23884 546 23936 552
rect 23620 480 23648 546
rect 24816 480 24844 3703
rect 26012 480 26040 3839
rect 27208 480 27236 9046
rect 29416 3194 29444 297366
rect 30690 10296 30746 10305
rect 30690 10231 30746 10240
rect 29588 3596 29640 3602
rect 29588 3538 29640 3544
rect 28392 3188 28444 3194
rect 28392 3130 28444 3136
rect 29404 3188 29456 3194
rect 29404 3130 29456 3136
rect 28404 480 28432 3130
rect 29600 480 29628 3538
rect 30704 3482 30732 10231
rect 30796 3602 30824 337622
rect 36396 337408 36448 337414
rect 36396 337350 36448 337356
rect 36408 337074 36436 337350
rect 36396 337068 36448 337074
rect 36396 337010 36448 337016
rect 34924 10464 34976 10470
rect 34924 10406 34976 10412
rect 31978 4040 32034 4049
rect 31978 3975 32034 3984
rect 30784 3596 30836 3602
rect 30784 3538 30836 3544
rect 30704 3454 30824 3482
rect 30796 480 30824 3454
rect 31992 480 32020 3975
rect 34936 3534 34964 10406
rect 37696 3602 37724 337690
rect 41824 10600 41876 10606
rect 41824 10542 41876 10548
rect 39064 10532 39116 10538
rect 39064 10474 39116 10480
rect 38972 3664 39024 3670
rect 38972 3606 39024 3612
rect 36672 3596 36724 3602
rect 36672 3538 36724 3544
rect 37684 3596 37736 3602
rect 37684 3538 37736 3544
rect 37868 3596 37920 3602
rect 37868 3538 37920 3544
rect 34372 3528 34424 3534
rect 34372 3470 34424 3476
rect 34924 3528 34976 3534
rect 34924 3470 34976 3476
rect 35476 3528 35528 3534
rect 35476 3470 35528 3476
rect 33176 3392 33228 3398
rect 33176 3334 33228 3340
rect 33188 480 33216 3334
rect 34384 480 34412 3470
rect 35488 480 35516 3470
rect 36684 480 36712 3538
rect 37880 480 37908 3538
rect 38984 1850 39012 3606
rect 39076 3602 39104 10474
rect 39064 3596 39116 3602
rect 39064 3538 39116 3544
rect 40260 3392 40312 3398
rect 41836 3346 41864 10542
rect 42652 3732 42704 3738
rect 42652 3674 42704 3680
rect 40260 3334 40312 3340
rect 38984 1822 39104 1850
rect 39076 480 39104 1822
rect 40272 480 40300 3334
rect 41468 3318 41864 3346
rect 41468 480 41496 3318
rect 42664 480 42692 3674
rect 44596 3602 44624 337894
rect 45976 337618 46004 337962
rect 45964 337612 46016 337618
rect 45964 337554 46016 337560
rect 45964 337408 46016 337414
rect 45964 337350 46016 337356
rect 45976 337074 46004 337350
rect 45964 337068 46016 337074
rect 45964 337010 46016 337016
rect 53324 10804 53376 10810
rect 53324 10746 53376 10752
rect 50104 10736 50156 10742
rect 50104 10678 50156 10684
rect 45964 10668 46016 10674
rect 45964 10610 46016 10616
rect 43848 3596 43900 3602
rect 43848 3538 43900 3544
rect 44584 3596 44636 3602
rect 44584 3538 44636 3544
rect 43860 480 43888 3538
rect 45976 3398 46004 10610
rect 48630 6216 48686 6225
rect 48630 6151 48686 6160
rect 47436 4004 47488 4010
rect 47436 3946 47488 3952
rect 46240 3936 46292 3942
rect 46240 3878 46292 3884
rect 45044 3392 45096 3398
rect 45044 3334 45096 3340
rect 45964 3392 46016 3398
rect 45964 3334 46016 3340
rect 45056 480 45084 3334
rect 46252 480 46280 3878
rect 47448 480 47476 3946
rect 48644 480 48672 6151
rect 50116 3380 50144 10678
rect 52128 6180 52180 6186
rect 52128 6122 52180 6128
rect 51024 4072 51076 4078
rect 51024 4014 51076 4020
rect 49840 3352 50144 3380
rect 49840 480 49868 3352
rect 51036 480 51064 4014
rect 52140 480 52168 6122
rect 53336 480 53364 10746
rect 55636 2990 55664 337962
rect 55716 337408 55768 337414
rect 55716 337350 55768 337356
rect 55728 337074 55756 337350
rect 55716 337068 55768 337074
rect 55716 337010 55768 337016
rect 56912 11008 56964 11014
rect 56912 10950 56964 10956
rect 55716 6248 55768 6254
rect 55716 6190 55768 6196
rect 54520 2984 54572 2990
rect 54520 2926 54572 2932
rect 55624 2984 55676 2990
rect 55624 2926 55676 2932
rect 54532 480 54560 2926
rect 55728 480 55756 6190
rect 56924 480 56952 10950
rect 60500 10260 60552 10266
rect 60500 10202 60552 10208
rect 59304 6316 59356 6322
rect 59304 6258 59356 6264
rect 58108 4140 58160 4146
rect 58108 4082 58160 4088
rect 58120 480 58148 4082
rect 58212 3590 58424 3618
rect 58212 3505 58240 3590
rect 58396 3505 58424 3590
rect 58198 3496 58254 3505
rect 58198 3431 58254 3440
rect 58382 3496 58438 3505
rect 58382 3431 58438 3440
rect 58198 3360 58254 3369
rect 58198 3295 58254 3304
rect 58382 3360 58438 3369
rect 58382 3295 58438 3304
rect 58212 3210 58240 3295
rect 58396 3210 58424 3295
rect 58212 3182 58424 3210
rect 59316 480 59344 6258
rect 60512 480 60540 10202
rect 62536 3398 62564 338030
rect 128854 337920 128910 337929
rect 128854 337855 128910 337864
rect 119286 337784 119342 337793
rect 119286 337719 119342 337728
rect 65284 337612 65336 337618
rect 65284 337554 65336 337560
rect 84604 337612 84656 337618
rect 84604 337554 84656 337560
rect 65296 337498 65324 337554
rect 84616 337498 84644 337554
rect 116344 337544 116396 337550
rect 65204 337470 65324 337498
rect 84524 337470 84644 337498
rect 94354 337512 94410 337521
rect 65204 337210 65232 337470
rect 65284 337408 65336 337414
rect 65284 337350 65336 337356
rect 75036 337408 75088 337414
rect 75036 337350 75088 337356
rect 65192 337204 65244 337210
rect 65192 337146 65244 337152
rect 65296 337074 65324 337350
rect 69424 337204 69476 337210
rect 69424 337146 69476 337152
rect 65284 337068 65336 337074
rect 65284 337010 65336 337016
rect 65284 10192 65336 10198
rect 65284 10134 65336 10140
rect 62892 7948 62944 7954
rect 62892 7890 62944 7896
rect 61696 3392 61748 3398
rect 61696 3334 61748 3340
rect 62524 3392 62576 3398
rect 62524 3334 62576 3340
rect 61708 480 61736 3334
rect 62904 480 62932 7890
rect 65296 3482 65324 10134
rect 68044 10124 68096 10130
rect 68044 10066 68096 10072
rect 66480 8016 66532 8022
rect 66480 7958 66532 7964
rect 65204 3454 65324 3482
rect 65204 3398 65232 3454
rect 64088 3392 64140 3398
rect 64088 3334 64140 3340
rect 65192 3392 65244 3398
rect 65192 3334 65244 3340
rect 65284 3392 65336 3398
rect 65284 3334 65336 3340
rect 64100 480 64128 3334
rect 65296 480 65324 3334
rect 66492 480 66520 7958
rect 68056 626 68084 10066
rect 69436 3194 69464 337146
rect 75048 336870 75076 337350
rect 76324 337136 76376 337142
rect 76324 337078 76376 337084
rect 75036 336864 75088 336870
rect 75036 336806 75088 336812
rect 73564 324964 73616 324970
rect 73564 324906 73616 324912
rect 72184 11756 72236 11762
rect 72184 11698 72236 11704
rect 69976 8084 70028 8090
rect 69976 8026 70028 8032
rect 68780 3188 68832 3194
rect 68780 3130 68832 3136
rect 69424 3188 69476 3194
rect 69424 3130 69476 3136
rect 67688 598 68084 626
rect 67688 480 67716 598
rect 68792 480 68820 3130
rect 69988 480 70016 8026
rect 72196 3194 72224 11698
rect 71172 3188 71224 3194
rect 71172 3130 71224 3136
rect 72184 3188 72236 3194
rect 72184 3130 72236 3136
rect 72368 3188 72420 3194
rect 72368 3130 72420 3136
rect 71184 480 71212 3130
rect 72380 480 72408 3130
rect 73576 480 73604 324906
rect 74944 11824 74996 11830
rect 74944 11766 74996 11772
rect 74956 610 74984 11766
rect 76336 3346 76364 337078
rect 83224 337068 83276 337074
rect 83224 337010 83276 337016
rect 77704 327752 77756 327758
rect 77704 327694 77756 327700
rect 75968 3318 76364 3346
rect 74760 604 74812 610
rect 74760 546 74812 552
rect 74944 604 74996 610
rect 74944 546 74996 552
rect 74772 480 74800 546
rect 75968 480 75996 3318
rect 77716 3126 77744 327694
rect 81844 294636 81896 294642
rect 81844 294578 81896 294584
rect 79084 11892 79136 11898
rect 79084 11834 79136 11840
rect 79096 3126 79124 11834
rect 81856 3126 81884 294578
rect 83132 12096 83184 12102
rect 83132 12038 83184 12044
rect 83144 3618 83172 12038
rect 83052 3590 83172 3618
rect 83052 3534 83080 3590
rect 81936 3528 81988 3534
rect 81936 3470 81988 3476
rect 83040 3528 83092 3534
rect 83236 3482 83264 337010
rect 84524 337006 84552 337470
rect 94354 337447 94410 337456
rect 103922 337512 103978 337521
rect 116344 337486 116396 337492
rect 103922 337447 103978 337456
rect 94368 337414 94396 337447
rect 103936 337414 103964 337447
rect 84604 337408 84656 337414
rect 84604 337350 84656 337356
rect 94356 337408 94408 337414
rect 94356 337350 94408 337356
rect 103924 337408 103976 337414
rect 103924 337350 103976 337356
rect 84512 337000 84564 337006
rect 84512 336942 84564 336948
rect 84616 336870 84644 337350
rect 87364 337000 87416 337006
rect 87364 336942 87416 336948
rect 84604 336864 84656 336870
rect 84604 336806 84656 336812
rect 84604 291848 84656 291854
rect 84604 291790 84656 291796
rect 83040 3470 83092 3476
rect 77152 3120 77204 3126
rect 77152 3062 77204 3068
rect 77704 3120 77756 3126
rect 77704 3062 77756 3068
rect 78348 3120 78400 3126
rect 78348 3062 78400 3068
rect 79084 3120 79136 3126
rect 79084 3062 79136 3068
rect 80740 3120 80792 3126
rect 80740 3062 80792 3068
rect 81844 3120 81896 3126
rect 81844 3062 81896 3068
rect 77164 480 77192 3062
rect 78360 480 78388 3062
rect 79544 3052 79596 3058
rect 79544 2994 79596 3000
rect 79556 480 79584 2994
rect 80752 480 80780 3062
rect 81948 480 81976 3470
rect 83144 3454 83264 3482
rect 83144 480 83172 3454
rect 84616 3346 84644 291790
rect 85984 12164 86036 12170
rect 85984 12106 86036 12112
rect 84340 3318 84644 3346
rect 84340 480 84368 3318
rect 85996 3058 86024 12106
rect 87376 3058 87404 336942
rect 94264 336932 94316 336938
rect 94264 336874 94316 336880
rect 88744 289128 88796 289134
rect 88744 289070 88796 289076
rect 88756 3058 88784 289070
rect 91504 280288 91556 280294
rect 91504 280230 91556 280236
rect 90124 276684 90176 276690
rect 90124 276626 90176 276632
rect 90136 3058 90164 276626
rect 91516 270502 91544 280230
rect 91504 270496 91556 270502
rect 91504 270438 91556 270444
rect 91504 260908 91556 260914
rect 91504 260850 91556 260856
rect 91516 251190 91544 260850
rect 91504 251184 91556 251190
rect 91504 251126 91556 251132
rect 91504 241664 91556 241670
rect 91504 241606 91556 241612
rect 91516 231849 91544 241606
rect 91318 231840 91374 231849
rect 91318 231775 91374 231784
rect 91502 231840 91558 231849
rect 91502 231775 91558 231784
rect 91332 222222 91360 231775
rect 91320 222216 91372 222222
rect 91320 222158 91372 222164
rect 91504 222216 91556 222222
rect 91504 222158 91556 222164
rect 91516 212537 91544 222158
rect 91318 212528 91374 212537
rect 91318 212463 91374 212472
rect 91502 212528 91558 212537
rect 91502 212463 91558 212472
rect 91332 203046 91360 212463
rect 91320 203040 91372 203046
rect 91320 202982 91372 202988
rect 91504 203040 91556 203046
rect 91504 202982 91556 202988
rect 91516 193225 91544 202982
rect 91318 193216 91374 193225
rect 91318 193151 91374 193160
rect 91502 193216 91558 193225
rect 91502 193151 91558 193160
rect 91332 183598 91360 193151
rect 91320 183592 91372 183598
rect 91320 183534 91372 183540
rect 91504 183592 91556 183598
rect 91504 183534 91556 183540
rect 91516 173913 91544 183534
rect 91502 173904 91558 173913
rect 91502 173839 91558 173848
rect 91502 164248 91558 164257
rect 91502 164183 91558 164192
rect 91516 154465 91544 164183
rect 91502 154456 91558 154465
rect 91502 154391 91558 154400
rect 91778 154456 91834 154465
rect 91778 154391 91834 154400
rect 91792 144945 91820 154391
rect 91502 144936 91558 144945
rect 91502 144871 91558 144880
rect 91778 144936 91834 144945
rect 91778 144871 91834 144880
rect 91516 135250 91544 144871
rect 91320 135244 91372 135250
rect 91320 135186 91372 135192
rect 91504 135244 91556 135250
rect 91504 135186 91556 135192
rect 91332 125769 91360 135186
rect 91318 125760 91374 125769
rect 91318 125695 91374 125704
rect 91502 125624 91558 125633
rect 91502 125559 91558 125568
rect 91516 115802 91544 125559
rect 91504 115796 91556 115802
rect 91504 115738 91556 115744
rect 91504 106344 91556 106350
rect 91504 106286 91556 106292
rect 91516 96626 91544 106286
rect 91320 96620 91372 96626
rect 91320 96562 91372 96568
rect 91504 96620 91556 96626
rect 91504 96562 91556 96568
rect 91332 87145 91360 96562
rect 91318 87136 91374 87145
rect 91318 87071 91374 87080
rect 91502 87000 91558 87009
rect 91502 86935 91558 86944
rect 91516 77178 91544 86935
rect 91504 77172 91556 77178
rect 91504 77114 91556 77120
rect 91504 67652 91556 67658
rect 91504 67594 91556 67600
rect 91516 57934 91544 67594
rect 91504 57928 91556 57934
rect 91504 57870 91556 57876
rect 91504 48340 91556 48346
rect 91504 48282 91556 48288
rect 91516 38554 91544 48282
rect 91504 38548 91556 38554
rect 91504 38490 91556 38496
rect 91504 29028 91556 29034
rect 91504 28970 91556 28976
rect 91516 19310 91544 28970
rect 91504 19304 91556 19310
rect 91504 19246 91556 19252
rect 92608 12232 92660 12238
rect 92608 12174 92660 12180
rect 91504 9716 91556 9722
rect 91504 9658 91556 9664
rect 91516 4842 91544 9658
rect 91424 4814 91544 4842
rect 85432 3052 85484 3058
rect 85432 2994 85484 3000
rect 85984 3052 86036 3058
rect 85984 2994 86036 3000
rect 86628 3052 86680 3058
rect 86628 2994 86680 3000
rect 87364 3052 87416 3058
rect 87364 2994 87416 3000
rect 87824 3052 87876 3058
rect 87824 2994 87876 3000
rect 88744 3052 88796 3058
rect 88744 2994 88796 3000
rect 89020 3052 89072 3058
rect 89020 2994 89072 3000
rect 90124 3052 90176 3058
rect 90124 2994 90176 3000
rect 85444 480 85472 2994
rect 86640 480 86668 2994
rect 87836 480 87864 2994
rect 89032 480 89060 2994
rect 90216 2984 90268 2990
rect 90216 2926 90268 2932
rect 90228 480 90256 2926
rect 91424 480 91452 4814
rect 92620 480 92648 12174
rect 94276 3534 94304 336874
rect 101164 336864 101216 336870
rect 101164 336806 101216 336812
rect 95644 283620 95696 283626
rect 95644 283562 95696 283568
rect 95656 3534 95684 283562
rect 99784 279472 99836 279478
rect 99784 279414 99836 279420
rect 97024 89004 97076 89010
rect 97024 88946 97076 88952
rect 97036 3534 97064 88946
rect 99508 12300 99560 12306
rect 99508 12242 99560 12248
rect 93804 3528 93856 3534
rect 93804 3470 93856 3476
rect 94264 3528 94316 3534
rect 94264 3470 94316 3476
rect 95000 3528 95052 3534
rect 95000 3470 95052 3476
rect 95644 3528 95696 3534
rect 95644 3470 95696 3476
rect 96196 3528 96248 3534
rect 96196 3470 96248 3476
rect 97024 3528 97076 3534
rect 97024 3470 97076 3476
rect 98588 3528 98640 3534
rect 98588 3470 98640 3476
rect 93816 480 93844 3470
rect 95012 480 95040 3470
rect 96208 480 96236 3470
rect 97392 2848 97444 2854
rect 97392 2790 97444 2796
rect 97404 480 97432 2790
rect 98600 480 98628 3470
rect 99520 3058 99548 12242
rect 99796 3534 99824 279414
rect 99784 3528 99836 3534
rect 99784 3470 99836 3476
rect 99692 3460 99744 3466
rect 99692 3402 99744 3408
rect 99704 3233 99732 3402
rect 101176 3346 101204 336806
rect 108064 336660 108116 336666
rect 108064 336602 108116 336608
rect 103924 307080 103976 307086
rect 103924 307022 103976 307028
rect 102544 10056 102596 10062
rect 102544 9998 102596 10004
rect 100992 3318 101204 3346
rect 99690 3224 99746 3233
rect 99690 3159 99746 3168
rect 99508 3052 99560 3058
rect 99508 2994 99560 3000
rect 99784 3052 99836 3058
rect 99784 2994 99836 3000
rect 99796 480 99824 2994
rect 100992 480 101020 3318
rect 102556 3058 102584 9998
rect 103832 3460 103884 3466
rect 103832 3402 103884 3408
rect 103844 3233 103872 3402
rect 103830 3224 103886 3233
rect 103830 3159 103886 3168
rect 102084 3052 102136 3058
rect 102084 2994 102136 3000
rect 102544 3052 102596 3058
rect 102544 2994 102596 3000
rect 102096 480 102124 2994
rect 103936 2922 103964 307022
rect 107972 12368 108024 12374
rect 107972 12310 108024 12316
rect 106684 9988 106736 9994
rect 106684 9930 106736 9936
rect 106696 2990 106724 9930
rect 107984 2990 108012 12310
rect 105672 2984 105724 2990
rect 105672 2926 105724 2932
rect 106684 2984 106736 2990
rect 106684 2926 106736 2932
rect 106868 2984 106920 2990
rect 106868 2926 106920 2932
rect 107972 2984 108024 2990
rect 107972 2926 108024 2932
rect 103280 2916 103332 2922
rect 103280 2858 103332 2864
rect 103924 2916 103976 2922
rect 103924 2858 103976 2864
rect 104476 2916 104528 2922
rect 104476 2858 104528 2864
rect 103292 480 103320 2858
rect 104488 480 104516 2858
rect 105684 480 105712 2926
rect 106880 480 106908 2926
rect 108076 480 108104 336602
rect 110824 320884 110876 320890
rect 110824 320826 110876 320832
rect 109444 9920 109496 9926
rect 109444 9862 109496 9868
rect 109456 3482 109484 9862
rect 110836 3482 110864 320826
rect 114964 12436 115016 12442
rect 114964 12378 115016 12384
rect 113584 9716 113636 9722
rect 113584 9658 113636 9664
rect 109272 3454 109484 3482
rect 110468 3454 110864 3482
rect 109272 480 109300 3454
rect 110468 480 110496 3454
rect 111652 2916 111704 2922
rect 111652 2858 111704 2864
rect 111664 480 111692 2858
rect 112848 2848 112900 2854
rect 112848 2790 112900 2796
rect 113308 2848 113360 2854
rect 113596 2802 113624 9658
rect 114976 3534 115004 12378
rect 116356 3534 116384 337486
rect 119300 336462 119328 337719
rect 128578 337648 128634 337657
rect 126004 337612 126056 337618
rect 128578 337583 128634 337592
rect 128764 337612 128816 337618
rect 126004 337554 126056 337560
rect 123886 337512 123942 337521
rect 123886 337447 123942 337456
rect 123900 337414 123928 337447
rect 123888 337408 123940 337414
rect 123888 337350 123940 337356
rect 119288 336456 119340 336462
rect 119288 336398 119340 336404
rect 117724 331968 117776 331974
rect 117724 331910 117776 331916
rect 117632 11144 117684 11150
rect 117632 11086 117684 11092
rect 117644 3618 117672 11086
rect 117460 3590 117672 3618
rect 117460 3534 117488 3590
rect 114044 3528 114096 3534
rect 114044 3470 114096 3476
rect 114964 3528 115016 3534
rect 114964 3470 115016 3476
rect 115240 3528 115292 3534
rect 115240 3470 115292 3476
rect 116344 3528 116396 3534
rect 116344 3470 116396 3476
rect 116436 3528 116488 3534
rect 116436 3470 116488 3476
rect 117448 3528 117500 3534
rect 117736 3482 117764 331910
rect 121864 316736 121916 316742
rect 121864 316678 121916 316684
rect 120482 10568 120538 10577
rect 120482 10503 120538 10512
rect 120496 3534 120524 10503
rect 121876 3534 121904 316678
rect 125912 271176 125964 271182
rect 125912 271118 125964 271124
rect 123520 10600 123572 10606
rect 123518 10568 123520 10577
rect 123572 10568 123574 10577
rect 123518 10503 123574 10512
rect 124624 9648 124676 9654
rect 124624 9590 124676 9596
rect 124636 3534 124664 9590
rect 125924 3618 125952 271118
rect 125832 3590 125952 3618
rect 125832 3534 125860 3590
rect 117448 3470 117500 3476
rect 113860 3460 113912 3466
rect 113860 3402 113912 3408
rect 113872 3233 113900 3402
rect 113858 3224 113914 3233
rect 113858 3159 113914 3168
rect 113360 2796 113624 2802
rect 113308 2790 113624 2796
rect 112860 480 112888 2790
rect 113320 2774 113624 2790
rect 114056 480 114084 3470
rect 115252 480 115280 3470
rect 116448 480 116476 3470
rect 117644 3454 117764 3482
rect 119932 3528 119984 3534
rect 119932 3470 119984 3476
rect 120484 3528 120536 3534
rect 120484 3470 120536 3476
rect 121128 3528 121180 3534
rect 121128 3470 121180 3476
rect 121864 3528 121916 3534
rect 121864 3470 121916 3476
rect 123520 3528 123572 3534
rect 123520 3470 123572 3476
rect 124624 3528 124676 3534
rect 124624 3470 124676 3476
rect 124716 3528 124768 3534
rect 124716 3470 124768 3476
rect 125820 3528 125872 3534
rect 126016 3482 126044 337554
rect 128592 337550 128620 337583
rect 128764 337554 128816 337560
rect 128580 337544 128632 337550
rect 128776 337521 128804 337554
rect 128868 337550 128896 337855
rect 129038 337784 129094 337793
rect 129038 337719 129094 337728
rect 128946 337648 129002 337657
rect 129052 337618 129080 337719
rect 129236 337657 129264 338098
rect 142576 337958 142604 338098
rect 152236 337958 152264 338098
rect 161896 337958 161924 338098
rect 171556 337958 171584 338098
rect 142564 337952 142616 337958
rect 138422 337920 138478 337929
rect 142564 337894 142616 337900
rect 152224 337952 152276 337958
rect 152224 337894 152276 337900
rect 161884 337952 161936 337958
rect 161884 337894 161936 337900
rect 171544 337952 171596 337958
rect 171544 337894 171596 337900
rect 138422 337855 138478 337864
rect 138436 337686 138464 337855
rect 142654 337784 142710 337793
rect 142654 337719 142710 337728
rect 152222 337784 152278 337793
rect 152222 337719 152278 337728
rect 161974 337784 162030 337793
rect 161974 337719 162030 337728
rect 171542 337784 171598 337793
rect 171542 337719 171598 337728
rect 138332 337680 138384 337686
rect 129222 337648 129278 337657
rect 128946 337583 129002 337592
rect 129040 337612 129092 337618
rect 128856 337544 128908 337550
rect 128580 337486 128632 337492
rect 128762 337512 128818 337521
rect 128856 337486 128908 337492
rect 128960 337498 128988 337583
rect 129222 337583 129278 337592
rect 138330 337648 138332 337657
rect 138424 337680 138476 337686
rect 138384 337648 138386 337657
rect 138424 337622 138476 337628
rect 142668 337618 142696 337719
rect 152236 337618 152264 337719
rect 161988 337618 162016 337719
rect 171556 337618 171584 337719
rect 138330 337583 138386 337592
rect 142472 337612 142524 337618
rect 129040 337554 129092 337560
rect 142472 337554 142524 337560
rect 142656 337612 142708 337618
rect 142656 337554 142708 337560
rect 142748 337612 142800 337618
rect 142748 337554 142800 337560
rect 152132 337612 152184 337618
rect 152132 337554 152184 337560
rect 152224 337612 152276 337618
rect 152224 337554 152276 337560
rect 152408 337612 152460 337618
rect 152408 337554 152460 337560
rect 161792 337612 161844 337618
rect 161792 337554 161844 337560
rect 161976 337612 162028 337618
rect 161976 337554 162028 337560
rect 162068 337612 162120 337618
rect 162068 337554 162120 337560
rect 171452 337612 171504 337618
rect 171452 337554 171504 337560
rect 171544 337612 171596 337618
rect 171544 337554 171596 337560
rect 171728 337612 171780 337618
rect 171728 337554 171780 337560
rect 129132 337544 129184 337550
rect 128960 337492 129132 337498
rect 142484 337521 142512 337554
rect 142760 337521 142788 337554
rect 152144 337521 152172 337554
rect 152420 337521 152448 337554
rect 161804 337521 161832 337554
rect 162080 337521 162108 337554
rect 171464 337521 171492 337554
rect 171740 337521 171768 337554
rect 128960 337486 129184 337492
rect 142286 337512 142342 337521
rect 128960 337470 129172 337486
rect 128762 337447 128818 337456
rect 142470 337512 142526 337521
rect 142342 337482 142420 337498
rect 142342 337476 142432 337482
rect 142342 337470 142380 337476
rect 142286 337447 142342 337456
rect 142470 337447 142526 337456
rect 142746 337512 142802 337521
rect 142746 337447 142802 337456
rect 152130 337512 152186 337521
rect 152130 337447 152186 337456
rect 152406 337512 152462 337521
rect 152590 337512 152646 337521
rect 152512 337482 152590 337498
rect 152406 337447 152462 337456
rect 152500 337476 152590 337482
rect 142380 337418 142432 337424
rect 152552 337470 152590 337476
rect 152590 337447 152646 337456
rect 161606 337512 161662 337521
rect 161790 337512 161846 337521
rect 161662 337482 161740 337498
rect 161662 337476 161752 337482
rect 161662 337470 161700 337476
rect 161606 337447 161662 337456
rect 152500 337418 152552 337424
rect 161790 337447 161846 337456
rect 162066 337512 162122 337521
rect 162066 337447 162122 337456
rect 171450 337512 171506 337521
rect 171450 337447 171506 337456
rect 171726 337512 171782 337521
rect 171910 337512 171966 337521
rect 171832 337482 171910 337498
rect 171726 337447 171782 337456
rect 171820 337476 171910 337482
rect 161700 337418 161752 337424
rect 171872 337470 171910 337476
rect 171910 337447 171966 337456
rect 171820 337418 171872 337424
rect 138332 337408 138384 337414
rect 138332 337350 138384 337356
rect 142564 337408 142616 337414
rect 142564 337350 142616 337356
rect 152316 337408 152368 337414
rect 152316 337350 152368 337356
rect 161884 337408 161936 337414
rect 161884 337350 161936 337356
rect 171636 337408 171688 337414
rect 171636 337350 171688 337356
rect 138344 337249 138372 337350
rect 142576 337249 142604 337350
rect 152328 337249 152356 337350
rect 161896 337249 161924 337350
rect 171648 337249 171676 337350
rect 138330 337240 138386 337249
rect 138330 337175 138386 337184
rect 142562 337240 142618 337249
rect 142562 337175 142618 337184
rect 152314 337240 152370 337249
rect 152314 337175 152370 337184
rect 161882 337240 161938 337249
rect 161882 337175 161938 337184
rect 171634 337240 171690 337249
rect 171634 337175 171690 337184
rect 127384 336048 127436 336054
rect 127384 335990 127436 335996
rect 125820 3470 125872 3476
rect 117644 480 117672 3454
rect 118736 2576 118788 2582
rect 118736 2518 118788 2524
rect 118748 480 118776 2518
rect 119944 480 119972 3470
rect 121140 480 121168 3470
rect 122324 2644 122376 2650
rect 122324 2586 122376 2592
rect 122336 480 122364 2586
rect 123532 480 123560 3470
rect 124728 480 124756 3470
rect 125924 3454 126044 3482
rect 126096 3528 126148 3534
rect 126096 3470 126148 3476
rect 125924 480 125952 3454
rect 126108 3233 126136 3470
rect 127396 3346 127424 335990
rect 163264 333328 163316 333334
rect 163264 333270 163316 333276
rect 145324 333260 145376 333266
rect 145324 333202 145376 333208
rect 135664 322244 135716 322250
rect 135664 322186 135716 322192
rect 134192 319456 134244 319462
rect 134192 319398 134244 319404
rect 128764 304292 128816 304298
rect 128764 304234 128816 304240
rect 128776 3534 128804 304234
rect 128856 10192 128908 10198
rect 128856 10134 128908 10140
rect 128868 9586 128896 10134
rect 128856 9580 128908 9586
rect 128856 9522 128908 9528
rect 129500 8288 129552 8294
rect 129500 8230 129552 8236
rect 128856 4276 128908 4282
rect 128856 4218 128908 4224
rect 128304 3528 128356 3534
rect 128304 3470 128356 3476
rect 128764 3528 128816 3534
rect 128764 3470 128816 3476
rect 127120 3318 127424 3346
rect 126094 3224 126150 3233
rect 126094 3159 126150 3168
rect 127120 480 127148 3318
rect 128316 480 128344 3470
rect 128868 3466 128896 4218
rect 128856 3460 128908 3466
rect 128856 3402 128908 3408
rect 129512 480 129540 8230
rect 131892 6384 131944 6390
rect 131892 6326 131944 6332
rect 130696 5228 130748 5234
rect 130696 5170 130748 5176
rect 130708 480 130736 5170
rect 131904 480 131932 6326
rect 134204 4010 134232 319398
rect 135676 317422 135704 322186
rect 138424 318096 138476 318102
rect 138424 318038 138476 318044
rect 135664 317416 135716 317422
rect 135664 317358 135716 317364
rect 135664 307828 135716 307834
rect 135664 307770 135716 307776
rect 135676 298081 135704 307770
rect 135478 298072 135534 298081
rect 135478 298007 135534 298016
rect 135662 298072 135718 298081
rect 135662 298007 135718 298016
rect 135492 288454 135520 298007
rect 135480 288448 135532 288454
rect 135480 288390 135532 288396
rect 135664 288448 135716 288454
rect 135664 288390 135716 288396
rect 135676 278769 135704 288390
rect 135478 278760 135534 278769
rect 135478 278695 135534 278704
rect 135662 278760 135718 278769
rect 135662 278695 135718 278704
rect 135492 269142 135520 278695
rect 135480 269136 135532 269142
rect 135480 269078 135532 269084
rect 135664 269136 135716 269142
rect 135664 269078 135716 269084
rect 135676 259457 135704 269078
rect 135478 259448 135534 259457
rect 135478 259383 135534 259392
rect 135662 259448 135718 259457
rect 135662 259383 135718 259392
rect 135492 249830 135520 259383
rect 135480 249824 135532 249830
rect 135480 249766 135532 249772
rect 135664 249824 135716 249830
rect 135664 249766 135716 249772
rect 135676 240145 135704 249766
rect 135478 240136 135534 240145
rect 135478 240071 135534 240080
rect 135662 240136 135718 240145
rect 135662 240071 135718 240080
rect 135492 230518 135520 240071
rect 135480 230512 135532 230518
rect 135480 230454 135532 230460
rect 135664 230512 135716 230518
rect 135664 230454 135716 230460
rect 135676 220833 135704 230454
rect 135478 220824 135534 220833
rect 135478 220759 135534 220768
rect 135662 220824 135718 220833
rect 135662 220759 135718 220768
rect 135492 211177 135520 220759
rect 135478 211168 135534 211177
rect 135478 211103 135534 211112
rect 135662 211168 135718 211177
rect 135662 211103 135718 211112
rect 135676 201482 135704 211103
rect 135480 201476 135532 201482
rect 135480 201418 135532 201424
rect 135664 201476 135716 201482
rect 135664 201418 135716 201424
rect 135492 191865 135520 201418
rect 135478 191856 135534 191865
rect 135478 191791 135534 191800
rect 135662 191856 135718 191865
rect 135662 191791 135718 191800
rect 135676 182170 135704 191791
rect 135480 182164 135532 182170
rect 135480 182106 135532 182112
rect 135664 182164 135716 182170
rect 135664 182106 135716 182112
rect 135492 172553 135520 182106
rect 135478 172544 135534 172553
rect 135478 172479 135534 172488
rect 135662 172544 135718 172553
rect 135662 172479 135718 172488
rect 135676 164529 135704 172479
rect 135662 164520 135718 164529
rect 135662 164455 135718 164464
rect 135570 164384 135626 164393
rect 135626 164342 135704 164370
rect 135570 164319 135626 164328
rect 135676 162858 135704 164342
rect 135664 162852 135716 162858
rect 135664 162794 135716 162800
rect 135664 153264 135716 153270
rect 135664 153206 135716 153212
rect 135676 143478 135704 153206
rect 135664 143472 135716 143478
rect 135664 143414 135716 143420
rect 135664 133952 135716 133958
rect 135664 133894 135716 133900
rect 135676 124166 135704 133894
rect 135664 124160 135716 124166
rect 135664 124102 135716 124108
rect 135664 114572 135716 114578
rect 135664 114514 135716 114520
rect 135676 104854 135704 114514
rect 135664 104848 135716 104854
rect 135664 104790 135716 104796
rect 135664 95328 135716 95334
rect 135664 95270 135716 95276
rect 135676 85542 135704 95270
rect 135664 85536 135716 85542
rect 135664 85478 135716 85484
rect 135664 75948 135716 75954
rect 135664 75890 135716 75896
rect 135676 66230 135704 75890
rect 135664 66224 135716 66230
rect 135664 66166 135716 66172
rect 135664 56704 135716 56710
rect 135664 56646 135716 56652
rect 135676 48657 135704 56646
rect 135662 48648 135718 48657
rect 135662 48583 135718 48592
rect 135662 48512 135718 48521
rect 135662 48447 135718 48456
rect 135676 46918 135704 48447
rect 135664 46912 135716 46918
rect 135664 46854 135716 46860
rect 135664 37324 135716 37330
rect 135664 37266 135716 37272
rect 135676 27606 135704 37266
rect 135664 27600 135716 27606
rect 135664 27542 135716 27548
rect 135296 18080 135348 18086
rect 135296 18022 135348 18028
rect 135308 9761 135336 18022
rect 138436 10690 138464 318038
rect 142564 315308 142616 315314
rect 142564 315250 142616 315256
rect 139804 301504 139856 301510
rect 139804 301446 139856 301452
rect 138068 10662 138464 10690
rect 135294 9752 135350 9761
rect 135294 9687 135350 9696
rect 135478 9752 135534 9761
rect 135478 9687 135534 9696
rect 134284 5296 134336 5302
rect 134284 5238 134336 5244
rect 133088 4004 133140 4010
rect 133088 3946 133140 3952
rect 134192 4004 134244 4010
rect 134192 3946 134244 3952
rect 133100 480 133128 3946
rect 134296 480 134324 5238
rect 135492 626 135520 9687
rect 136584 9172 136636 9178
rect 136584 9114 136636 9120
rect 135400 598 135520 626
rect 135400 480 135428 598
rect 136596 480 136624 9114
rect 137700 4134 137912 4162
rect 137700 4010 137728 4134
rect 137688 4004 137740 4010
rect 137688 3946 137740 3952
rect 137780 4004 137832 4010
rect 137780 3946 137832 3952
rect 137792 480 137820 3946
rect 137884 3516 137912 4134
rect 138068 4010 138096 10662
rect 138424 10532 138476 10538
rect 138424 10474 138476 10480
rect 138238 10160 138294 10169
rect 138238 10095 138240 10104
rect 138292 10095 138294 10104
rect 138240 10066 138292 10072
rect 138436 9874 138464 10474
rect 138608 10192 138660 10198
rect 138606 10160 138608 10169
rect 138660 10160 138662 10169
rect 138606 10095 138662 10104
rect 138252 9846 138464 9874
rect 138252 9654 138280 9846
rect 138240 9648 138292 9654
rect 138240 9590 138292 9596
rect 138056 4004 138108 4010
rect 138056 3946 138108 3952
rect 139816 3670 139844 301446
rect 142472 300144 142524 300150
rect 142472 300086 142524 300092
rect 140172 9036 140224 9042
rect 140172 8978 140224 8984
rect 138976 3664 139028 3670
rect 138976 3606 139028 3612
rect 139804 3664 139856 3670
rect 139804 3606 139856 3612
rect 138424 3528 138476 3534
rect 137884 3488 138424 3516
rect 138424 3470 138476 3476
rect 138988 480 139016 3606
rect 140184 480 140212 8978
rect 141368 3664 141420 3670
rect 141368 3606 141420 3612
rect 141380 480 141408 3606
rect 142484 3516 142512 300086
rect 142576 3670 142604 315250
rect 145336 19310 145364 333202
rect 156364 330608 156416 330614
rect 156364 330550 156416 330556
rect 152224 327140 152276 327146
rect 152224 327082 152276 327088
rect 152236 317422 152264 327082
rect 152224 317416 152276 317422
rect 152224 317358 152276 317364
rect 149464 312656 149516 312662
rect 149464 312598 149516 312604
rect 145324 19304 145376 19310
rect 145324 19246 145376 19252
rect 145232 19236 145284 19242
rect 145232 19178 145284 19184
rect 145244 12186 145272 19178
rect 145060 12158 145272 12186
rect 143300 10260 143352 10266
rect 143300 10202 143352 10208
rect 143312 10130 143340 10202
rect 143300 10124 143352 10130
rect 143300 10066 143352 10072
rect 143760 9376 143812 9382
rect 143760 9318 143812 9324
rect 142564 3664 142616 3670
rect 142564 3606 142616 3612
rect 142484 3488 142604 3516
rect 142576 480 142604 3488
rect 143772 480 143800 9318
rect 145060 626 145088 12158
rect 147808 10804 147860 10810
rect 147808 10746 147860 10752
rect 148452 10804 148504 10810
rect 148452 10746 148504 10752
rect 147820 10577 147848 10746
rect 148464 10577 148492 10746
rect 147806 10568 147862 10577
rect 147806 10503 147862 10512
rect 148450 10568 148506 10577
rect 148450 10503 148506 10512
rect 147348 9512 147400 9518
rect 147348 9454 147400 9460
rect 146152 7540 146204 7546
rect 146152 7482 146204 7488
rect 144968 598 145088 626
rect 144968 480 144996 598
rect 146164 480 146192 7482
rect 147360 480 147388 9454
rect 149476 3670 149504 312598
rect 152224 307828 152276 307834
rect 152224 307770 152276 307776
rect 152236 298081 152264 307770
rect 152038 298072 152094 298081
rect 152038 298007 152094 298016
rect 152222 298072 152278 298081
rect 152222 298007 152278 298016
rect 152052 288454 152080 298007
rect 152040 288448 152092 288454
rect 152040 288390 152092 288396
rect 152224 288448 152276 288454
rect 152224 288390 152276 288396
rect 152236 278769 152264 288390
rect 152038 278760 152094 278769
rect 152038 278695 152094 278704
rect 152222 278760 152278 278769
rect 152222 278695 152278 278704
rect 152052 269142 152080 278695
rect 152040 269136 152092 269142
rect 152040 269078 152092 269084
rect 152224 269136 152276 269142
rect 152224 269078 152276 269084
rect 152236 259457 152264 269078
rect 152038 259448 152094 259457
rect 152038 259383 152094 259392
rect 152222 259448 152278 259457
rect 152222 259383 152278 259392
rect 152052 249830 152080 259383
rect 152040 249824 152092 249830
rect 152040 249766 152092 249772
rect 152224 249824 152276 249830
rect 152224 249766 152276 249772
rect 152236 240145 152264 249766
rect 152038 240136 152094 240145
rect 152038 240071 152094 240080
rect 152222 240136 152278 240145
rect 152222 240071 152278 240080
rect 152052 230518 152080 240071
rect 152040 230512 152092 230518
rect 152040 230454 152092 230460
rect 152224 230512 152276 230518
rect 152224 230454 152276 230460
rect 152236 220833 152264 230454
rect 152038 220824 152094 220833
rect 152038 220759 152094 220768
rect 152222 220824 152278 220833
rect 152222 220759 152278 220768
rect 152052 211177 152080 220759
rect 152038 211168 152094 211177
rect 152038 211103 152094 211112
rect 152222 211168 152278 211177
rect 152222 211103 152278 211112
rect 152236 201482 152264 211103
rect 152040 201476 152092 201482
rect 152040 201418 152092 201424
rect 152224 201476 152276 201482
rect 152224 201418 152276 201424
rect 152052 191865 152080 201418
rect 152038 191856 152094 191865
rect 152038 191791 152094 191800
rect 152222 191856 152278 191865
rect 152222 191791 152278 191800
rect 152236 182170 152264 191791
rect 152040 182164 152092 182170
rect 152040 182106 152092 182112
rect 152224 182164 152276 182170
rect 152224 182106 152276 182112
rect 152052 172553 152080 182106
rect 152038 172544 152094 172553
rect 152038 172479 152094 172488
rect 152222 172544 152278 172553
rect 152222 172479 152278 172488
rect 152236 162858 152264 172479
rect 152224 162852 152276 162858
rect 152224 162794 152276 162800
rect 152224 153264 152276 153270
rect 152224 153206 152276 153212
rect 152236 143478 152264 153206
rect 152224 143472 152276 143478
rect 152224 143414 152276 143420
rect 152224 133952 152276 133958
rect 152224 133894 152276 133900
rect 152236 124166 152264 133894
rect 152224 124160 152276 124166
rect 152224 124102 152276 124108
rect 152224 114572 152276 114578
rect 152224 114514 152276 114520
rect 152236 104854 152264 114514
rect 152224 104848 152276 104854
rect 152224 104790 152276 104796
rect 152224 95328 152276 95334
rect 152224 95270 152276 95276
rect 152236 85542 152264 95270
rect 152224 85536 152276 85542
rect 152224 85478 152276 85484
rect 152224 75948 152276 75954
rect 152224 75890 152276 75896
rect 152236 66230 152264 75890
rect 152224 66224 152276 66230
rect 152224 66166 152276 66172
rect 152224 56704 152276 56710
rect 152224 56646 152276 56652
rect 152236 46918 152264 56646
rect 152224 46912 152276 46918
rect 152224 46854 152276 46860
rect 152224 37324 152276 37330
rect 152224 37266 152276 37272
rect 152236 27606 152264 37266
rect 152224 27600 152276 27606
rect 152224 27542 152276 27548
rect 151856 18080 151908 18086
rect 151856 18022 151908 18028
rect 151868 9761 151896 18022
rect 153052 10804 153104 10810
rect 153052 10746 153104 10752
rect 153064 10674 153092 10746
rect 153052 10668 153104 10674
rect 153052 10610 153104 10616
rect 151854 9752 151910 9761
rect 151854 9687 151910 9696
rect 152038 9752 152094 9761
rect 152038 9687 152094 9696
rect 150936 9580 150988 9586
rect 152052 9568 152080 9687
rect 152052 9540 152172 9568
rect 150936 9522 150988 9528
rect 149740 7472 149792 7478
rect 149740 7414 149792 7420
rect 148544 3664 148596 3670
rect 148544 3606 148596 3612
rect 149464 3664 149516 3670
rect 149464 3606 149516 3612
rect 148174 3360 148230 3369
rect 148174 3295 148230 3304
rect 148082 3088 148138 3097
rect 148188 3074 148216 3295
rect 148138 3046 148216 3074
rect 148082 3023 148138 3032
rect 148556 480 148584 3606
rect 149752 480 149780 7414
rect 150948 480 150976 9522
rect 152144 610 152172 9540
rect 154432 8560 154484 8566
rect 154432 8502 154484 8508
rect 153236 7404 153288 7410
rect 153236 7346 153288 7352
rect 152040 604 152092 610
rect 152040 546 152092 552
rect 152132 604 152184 610
rect 152132 546 152184 552
rect 152052 480 152080 546
rect 153248 480 153276 7346
rect 154444 480 154472 8502
rect 156376 610 156404 330550
rect 160504 307148 160556 307154
rect 160504 307090 160556 307096
rect 157834 10432 157890 10441
rect 157834 10367 157890 10376
rect 157468 10192 157520 10198
rect 157466 10160 157468 10169
rect 157848 10169 157876 10367
rect 157520 10160 157522 10169
rect 157834 10160 157890 10169
rect 157466 10095 157522 10104
rect 157560 10124 157612 10130
rect 157834 10095 157890 10104
rect 157560 10066 157612 10072
rect 157572 10033 157600 10066
rect 157558 10024 157614 10033
rect 157558 9959 157614 9968
rect 158020 8628 158072 8634
rect 158020 8570 158072 8576
rect 156824 7336 156876 7342
rect 156824 7278 156876 7284
rect 155628 604 155680 610
rect 155628 546 155680 552
rect 156364 604 156416 610
rect 156364 546 156416 552
rect 155640 480 155668 546
rect 156836 480 156864 7278
rect 157652 3528 157704 3534
rect 157652 3470 157704 3476
rect 157664 3233 157692 3470
rect 157650 3224 157706 3233
rect 157650 3159 157706 3168
rect 158032 480 158060 8570
rect 160412 7268 160464 7274
rect 160412 7210 160464 7216
rect 159216 3664 159268 3670
rect 159216 3606 159268 3612
rect 158112 3460 158164 3466
rect 158112 3402 158164 3408
rect 158124 3233 158152 3402
rect 158110 3224 158166 3233
rect 158110 3159 158166 3168
rect 159228 480 159256 3606
rect 160424 480 160452 7210
rect 160516 3670 160544 307090
rect 161608 8900 161660 8906
rect 161608 8842 161660 8848
rect 160504 3664 160556 3670
rect 160504 3606 160556 3612
rect 161620 480 161648 8842
rect 163276 3670 163304 333270
rect 167404 330676 167456 330682
rect 167404 330618 167456 330624
rect 165196 7200 165248 7206
rect 165196 7142 165248 7148
rect 164000 6452 164052 6458
rect 164000 6394 164052 6400
rect 162804 3664 162856 3670
rect 162804 3606 162856 3612
rect 163264 3664 163316 3670
rect 163264 3606 163316 3612
rect 162816 480 162844 3606
rect 164012 480 164040 6394
rect 165208 480 165236 7142
rect 166392 3664 166444 3670
rect 166392 3606 166444 3612
rect 167220 3664 167272 3670
rect 167416 3618 167444 330618
rect 170164 327140 170216 327146
rect 170164 327082 170216 327088
rect 170176 317422 170204 327082
rect 174304 325032 174356 325038
rect 174304 324974 174356 324980
rect 170164 317416 170216 317422
rect 170164 317358 170216 317364
rect 170164 307828 170216 307834
rect 170164 307770 170216 307776
rect 170176 298081 170204 307770
rect 170162 298072 170218 298081
rect 170162 298007 170218 298016
rect 170346 298072 170402 298081
rect 170346 298007 170402 298016
rect 170360 288454 170388 298007
rect 170164 288448 170216 288454
rect 170164 288390 170216 288396
rect 170348 288448 170400 288454
rect 170348 288390 170400 288396
rect 170176 278769 170204 288390
rect 170162 278760 170218 278769
rect 170162 278695 170218 278704
rect 170346 278760 170402 278769
rect 170346 278695 170402 278704
rect 170360 269142 170388 278695
rect 170164 269136 170216 269142
rect 170164 269078 170216 269084
rect 170348 269136 170400 269142
rect 170348 269078 170400 269084
rect 170176 259457 170204 269078
rect 170162 259448 170218 259457
rect 170162 259383 170218 259392
rect 170346 259448 170402 259457
rect 170346 259383 170402 259392
rect 170360 249830 170388 259383
rect 170164 249824 170216 249830
rect 170164 249766 170216 249772
rect 170348 249824 170400 249830
rect 170348 249766 170400 249772
rect 170176 240145 170204 249766
rect 170162 240136 170218 240145
rect 170162 240071 170218 240080
rect 170346 240136 170402 240145
rect 170346 240071 170402 240080
rect 170360 230518 170388 240071
rect 170164 230512 170216 230518
rect 170164 230454 170216 230460
rect 170348 230512 170400 230518
rect 170348 230454 170400 230460
rect 170176 220833 170204 230454
rect 170162 220824 170218 220833
rect 170162 220759 170218 220768
rect 170346 220824 170402 220833
rect 170346 220759 170402 220768
rect 170360 211177 170388 220759
rect 170162 211168 170218 211177
rect 170162 211103 170218 211112
rect 170346 211168 170402 211177
rect 170346 211103 170402 211112
rect 170176 201482 170204 211103
rect 170164 201476 170216 201482
rect 170164 201418 170216 201424
rect 170348 201476 170400 201482
rect 170348 201418 170400 201424
rect 170360 191865 170388 201418
rect 170162 191856 170218 191865
rect 170162 191791 170218 191800
rect 170346 191856 170402 191865
rect 170346 191791 170402 191800
rect 170176 182170 170204 191791
rect 170164 182164 170216 182170
rect 170164 182106 170216 182112
rect 170348 182164 170400 182170
rect 170348 182106 170400 182112
rect 170360 172553 170388 182106
rect 170162 172544 170218 172553
rect 170162 172479 170218 172488
rect 170346 172544 170402 172553
rect 170346 172479 170402 172488
rect 170176 162858 170204 172479
rect 170164 162852 170216 162858
rect 170164 162794 170216 162800
rect 170164 153264 170216 153270
rect 170164 153206 170216 153212
rect 170176 143478 170204 153206
rect 170164 143472 170216 143478
rect 170164 143414 170216 143420
rect 170164 133952 170216 133958
rect 170164 133894 170216 133900
rect 170176 124166 170204 133894
rect 170164 124160 170216 124166
rect 170164 124102 170216 124108
rect 170164 114572 170216 114578
rect 170164 114514 170216 114520
rect 170176 104854 170204 114514
rect 170164 104848 170216 104854
rect 170164 104790 170216 104796
rect 170164 95328 170216 95334
rect 170164 95270 170216 95276
rect 170176 85542 170204 95270
rect 170164 85536 170216 85542
rect 170164 85478 170216 85484
rect 170164 75948 170216 75954
rect 170164 75890 170216 75896
rect 170176 66230 170204 75890
rect 170164 66224 170216 66230
rect 170164 66166 170216 66172
rect 170164 56704 170216 56710
rect 170164 56646 170216 56652
rect 170176 46918 170204 56646
rect 170164 46912 170216 46918
rect 170164 46854 170216 46860
rect 170164 37324 170216 37330
rect 170164 37266 170216 37272
rect 170176 27606 170204 37266
rect 170164 27600 170216 27606
rect 170164 27542 170216 27548
rect 169704 18080 169756 18086
rect 169704 18022 169756 18028
rect 167588 11212 167640 11218
rect 167588 11154 167640 11160
rect 167496 11076 167548 11082
rect 167496 11018 167548 11024
rect 167508 10033 167536 11018
rect 167600 10198 167628 11154
rect 167862 10432 167918 10441
rect 167862 10367 167918 10376
rect 167876 10198 167904 10367
rect 167588 10192 167640 10198
rect 167864 10192 167916 10198
rect 167588 10134 167640 10140
rect 167770 10160 167826 10169
rect 167864 10134 167916 10140
rect 167770 10095 167772 10104
rect 167824 10095 167826 10104
rect 167772 10066 167824 10072
rect 167494 10024 167550 10033
rect 167494 9959 167550 9968
rect 169716 9761 169744 18022
rect 169702 9752 169758 9761
rect 169702 9687 169758 9696
rect 169886 9752 169942 9761
rect 169886 9687 169942 9696
rect 169520 9648 169572 9654
rect 169520 9590 169572 9596
rect 169900 9602 169928 9687
rect 170164 9648 170216 9654
rect 169532 9489 169560 9590
rect 169900 9574 170020 9602
rect 170164 9590 170216 9596
rect 169518 9480 169574 9489
rect 169518 9415 169574 9424
rect 168692 6996 168744 7002
rect 168692 6938 168744 6944
rect 167588 6656 167640 6662
rect 167588 6598 167640 6604
rect 167272 3612 167444 3618
rect 167220 3606 167444 3612
rect 166404 480 166432 3606
rect 167232 3590 167444 3606
rect 167600 480 167628 6598
rect 168704 480 168732 6938
rect 169992 610 170020 9574
rect 170176 9489 170204 9590
rect 170162 9480 170218 9489
rect 170162 9415 170218 9424
rect 172280 6928 172332 6934
rect 172280 6870 172332 6876
rect 171084 6724 171136 6730
rect 171084 6666 171136 6672
rect 169888 604 169940 610
rect 169888 546 169940 552
rect 169980 604 170032 610
rect 169980 546 170032 552
rect 169900 480 169928 546
rect 171096 480 171124 6666
rect 172292 480 172320 6870
rect 174316 610 174344 324974
rect 177064 322312 177116 322318
rect 177064 322254 177116 322260
rect 174672 6792 174724 6798
rect 174672 6734 174724 6740
rect 173476 604 173528 610
rect 173476 546 173528 552
rect 174304 604 174356 610
rect 174304 546 174356 552
rect 173488 480 173516 546
rect 174684 480 174712 6734
rect 175868 5908 175920 5914
rect 175868 5850 175920 5856
rect 175880 480 175908 5850
rect 177076 480 177104 322254
rect 179192 260846 179220 461042
rect 219200 458516 219252 458522
rect 219200 458458 219252 458464
rect 181204 338156 181256 338162
rect 181204 338098 181256 338104
rect 190864 338156 190916 338162
rect 190864 338098 190916 338104
rect 200524 338156 200576 338162
rect 200524 338098 200576 338104
rect 210184 338156 210236 338162
rect 210184 338098 210236 338104
rect 181216 337958 181244 338098
rect 190876 337958 190904 338098
rect 200536 337958 200564 338098
rect 210196 337958 210224 338098
rect 181204 337952 181256 337958
rect 181204 337894 181256 337900
rect 190864 337952 190916 337958
rect 190864 337894 190916 337900
rect 200524 337952 200576 337958
rect 200524 337894 200576 337900
rect 210184 337952 210236 337958
rect 210184 337894 210236 337900
rect 181294 337784 181350 337793
rect 181294 337719 181350 337728
rect 190862 337784 190918 337793
rect 190862 337719 190918 337728
rect 200614 337784 200670 337793
rect 200614 337719 200670 337728
rect 210182 337784 210238 337793
rect 210182 337719 210238 337728
rect 181308 337618 181336 337719
rect 190876 337618 190904 337719
rect 200628 337618 200656 337719
rect 210196 337618 210224 337719
rect 181112 337612 181164 337618
rect 181112 337554 181164 337560
rect 181296 337612 181348 337618
rect 181296 337554 181348 337560
rect 181388 337612 181440 337618
rect 181388 337554 181440 337560
rect 190772 337612 190824 337618
rect 190772 337554 190824 337560
rect 190864 337612 190916 337618
rect 190864 337554 190916 337560
rect 191048 337612 191100 337618
rect 191048 337554 191100 337560
rect 200432 337612 200484 337618
rect 200432 337554 200484 337560
rect 200616 337612 200668 337618
rect 200616 337554 200668 337560
rect 200708 337612 200760 337618
rect 200708 337554 200760 337560
rect 210092 337612 210144 337618
rect 210092 337554 210144 337560
rect 210184 337612 210236 337618
rect 210184 337554 210236 337560
rect 210368 337612 210420 337618
rect 210368 337554 210420 337560
rect 181124 337521 181152 337554
rect 181400 337521 181428 337554
rect 190784 337521 190812 337554
rect 191060 337521 191088 337554
rect 200444 337521 200472 337554
rect 200720 337521 200748 337554
rect 210104 337521 210132 337554
rect 210380 337521 210408 337554
rect 180926 337512 180982 337521
rect 181110 337512 181166 337521
rect 180982 337482 181060 337498
rect 180982 337476 181072 337482
rect 180982 337470 181020 337476
rect 180926 337447 180982 337456
rect 181110 337447 181166 337456
rect 181386 337512 181442 337521
rect 181386 337447 181442 337456
rect 190770 337512 190826 337521
rect 190770 337447 190826 337456
rect 191046 337512 191102 337521
rect 191230 337512 191286 337521
rect 191152 337482 191230 337498
rect 191046 337447 191102 337456
rect 191140 337476 191230 337482
rect 181020 337418 181072 337424
rect 191192 337470 191230 337476
rect 191230 337447 191286 337456
rect 200246 337512 200302 337521
rect 200430 337512 200486 337521
rect 200302 337482 200380 337498
rect 200302 337476 200392 337482
rect 200302 337470 200340 337476
rect 200246 337447 200302 337456
rect 191140 337418 191192 337424
rect 200430 337447 200486 337456
rect 200706 337512 200762 337521
rect 200706 337447 200762 337456
rect 210090 337512 210146 337521
rect 210090 337447 210146 337456
rect 210366 337512 210422 337521
rect 210550 337512 210606 337521
rect 210472 337482 210550 337498
rect 210366 337447 210422 337456
rect 210460 337476 210550 337482
rect 200340 337418 200392 337424
rect 210512 337470 210550 337476
rect 210550 337447 210606 337456
rect 210460 337418 210512 337424
rect 181204 337408 181256 337414
rect 181204 337350 181256 337356
rect 190956 337408 191008 337414
rect 190956 337350 191008 337356
rect 200524 337408 200576 337414
rect 200524 337350 200576 337356
rect 210276 337408 210328 337414
rect 210276 337350 210328 337356
rect 181216 337249 181244 337350
rect 190968 337249 190996 337350
rect 200536 337249 200564 337350
rect 210288 337249 210316 337350
rect 181202 337240 181258 337249
rect 181202 337175 181258 337184
rect 190954 337240 191010 337249
rect 190954 337175 191010 337184
rect 200522 337240 200578 337249
rect 200522 337175 200578 337184
rect 210274 337240 210330 337249
rect 210274 337175 210330 337184
rect 181204 336116 181256 336122
rect 181204 336058 181256 336064
rect 179180 260840 179232 260846
rect 179180 260782 179232 260788
rect 177248 11144 177300 11150
rect 177248 11086 177300 11092
rect 177260 10577 177288 11086
rect 177246 10568 177302 10577
rect 177246 10503 177302 10512
rect 178260 6860 178312 6866
rect 178260 6802 178312 6808
rect 178272 480 178300 6802
rect 179456 5840 179508 5846
rect 179456 5782 179508 5788
rect 179468 480 179496 5782
rect 181216 610 181244 336058
rect 204664 333396 204716 333402
rect 204664 333338 204716 333344
rect 186724 326528 186776 326534
rect 186724 326470 186776 326476
rect 185344 319524 185396 319530
rect 185344 319466 185396 319472
rect 183964 297492 184016 297498
rect 183964 297434 184016 297440
rect 181848 6112 181900 6118
rect 181848 6054 181900 6060
rect 180652 604 180704 610
rect 180652 546 180704 552
rect 181204 604 181256 610
rect 181204 546 181256 552
rect 180664 480 180692 546
rect 181860 480 181888 6054
rect 183976 610 184004 297434
rect 185356 8430 185384 319466
rect 184240 8424 184292 8430
rect 184240 8366 184292 8372
rect 185344 8424 185396 8430
rect 185344 8366 185396 8372
rect 183044 604 183096 610
rect 183044 546 183096 552
rect 183964 604 184016 610
rect 183964 546 184016 552
rect 183056 480 183084 546
rect 184252 480 184280 8366
rect 185344 5908 185396 5914
rect 185344 5850 185396 5856
rect 185356 480 185384 5850
rect 186540 3460 186592 3466
rect 186540 3402 186592 3408
rect 186552 3233 186580 3402
rect 186538 3224 186594 3233
rect 186538 3159 186594 3168
rect 186736 626 186764 326470
rect 194912 323604 194964 323610
rect 194912 323546 194964 323552
rect 190864 307828 190916 307834
rect 190864 307770 190916 307776
rect 190876 298081 190904 307770
rect 190678 298072 190734 298081
rect 190678 298007 190734 298016
rect 190862 298072 190918 298081
rect 190862 298007 190918 298016
rect 190692 288454 190720 298007
rect 190680 288448 190732 288454
rect 190680 288390 190732 288396
rect 190864 288448 190916 288454
rect 190864 288390 190916 288396
rect 190876 278769 190904 288390
rect 190678 278760 190734 278769
rect 190678 278695 190734 278704
rect 190862 278760 190918 278769
rect 190862 278695 190918 278704
rect 190692 269142 190720 278695
rect 190680 269136 190732 269142
rect 190680 269078 190732 269084
rect 190864 269136 190916 269142
rect 190864 269078 190916 269084
rect 190876 259457 190904 269078
rect 190678 259448 190734 259457
rect 190678 259383 190734 259392
rect 190862 259448 190918 259457
rect 190862 259383 190918 259392
rect 190692 249830 190720 259383
rect 190680 249824 190732 249830
rect 190680 249766 190732 249772
rect 190864 249824 190916 249830
rect 190864 249766 190916 249772
rect 190876 240145 190904 249766
rect 190678 240136 190734 240145
rect 190678 240071 190734 240080
rect 190862 240136 190918 240145
rect 190862 240071 190918 240080
rect 190692 230518 190720 240071
rect 190680 230512 190732 230518
rect 190680 230454 190732 230460
rect 190864 230512 190916 230518
rect 190864 230454 190916 230460
rect 190876 220833 190904 230454
rect 190678 220824 190734 220833
rect 190678 220759 190734 220768
rect 190862 220824 190918 220833
rect 190862 220759 190918 220768
rect 190692 211177 190720 220759
rect 190678 211168 190734 211177
rect 190678 211103 190734 211112
rect 190862 211168 190918 211177
rect 190862 211103 190918 211112
rect 190876 201482 190904 211103
rect 190680 201476 190732 201482
rect 190680 201418 190732 201424
rect 190864 201476 190916 201482
rect 190864 201418 190916 201424
rect 190692 191865 190720 201418
rect 190678 191856 190734 191865
rect 190678 191791 190734 191800
rect 190862 191856 190918 191865
rect 190862 191791 190918 191800
rect 190876 182170 190904 191791
rect 190680 182164 190732 182170
rect 190680 182106 190732 182112
rect 190864 182164 190916 182170
rect 190864 182106 190916 182112
rect 190692 172553 190720 182106
rect 190678 172544 190734 172553
rect 190678 172479 190734 172488
rect 190862 172544 190918 172553
rect 190862 172479 190918 172488
rect 190876 162858 190904 172479
rect 190864 162852 190916 162858
rect 190864 162794 190916 162800
rect 190864 153264 190916 153270
rect 190864 153206 190916 153212
rect 190876 143478 190904 153206
rect 190864 143472 190916 143478
rect 190864 143414 190916 143420
rect 190864 133952 190916 133958
rect 190864 133894 190916 133900
rect 190876 124166 190904 133894
rect 190864 124160 190916 124166
rect 190864 124102 190916 124108
rect 190864 114572 190916 114578
rect 190864 114514 190916 114520
rect 190876 104854 190904 114514
rect 190864 104848 190916 104854
rect 190864 104790 190916 104796
rect 190864 95328 190916 95334
rect 190864 95270 190916 95276
rect 190876 85542 190904 95270
rect 190864 85536 190916 85542
rect 190864 85478 190916 85484
rect 190864 75948 190916 75954
rect 190864 75890 190916 75896
rect 190876 66230 190904 75890
rect 190864 66224 190916 66230
rect 190864 66166 190916 66172
rect 190864 56704 190916 56710
rect 190864 56646 190916 56652
rect 190876 46918 190904 56646
rect 190864 46912 190916 46918
rect 190864 46854 190916 46860
rect 190864 37324 190916 37330
rect 190864 37266 190916 37272
rect 190876 27606 190904 37266
rect 190220 27600 190272 27606
rect 190220 27542 190272 27548
rect 190864 27600 190916 27606
rect 190864 27542 190916 27548
rect 190232 18057 190260 27542
rect 190218 18048 190274 18057
rect 190218 17983 190274 17992
rect 190402 18048 190458 18057
rect 190402 17983 190458 17992
rect 187092 10804 187144 10810
rect 187092 10746 187144 10752
rect 186816 10736 186868 10742
rect 186814 10704 186816 10713
rect 186868 10704 186870 10713
rect 186814 10639 186870 10648
rect 187104 10577 187132 10746
rect 187090 10568 187146 10577
rect 187090 10503 187146 10512
rect 190416 9761 190444 17983
rect 191692 10804 191744 10810
rect 191692 10746 191744 10752
rect 191704 10674 191732 10746
rect 191692 10668 191744 10674
rect 191692 10610 191744 10616
rect 191782 10160 191838 10169
rect 191782 10095 191838 10104
rect 190402 9752 190458 9761
rect 190402 9687 190458 9696
rect 190586 9752 190642 9761
rect 190586 9687 190642 9696
rect 190600 9602 190628 9687
rect 190416 9574 190628 9602
rect 188932 5840 188984 5846
rect 188932 5782 188984 5788
rect 187734 4856 187790 4865
rect 187734 4791 187790 4800
rect 186816 4208 186868 4214
rect 186816 4150 186868 4156
rect 186828 3466 186856 4150
rect 186816 3460 186868 3466
rect 186816 3402 186868 3408
rect 187182 3224 187238 3233
rect 187182 3159 187184 3168
rect 187236 3159 187238 3168
rect 187184 3130 187236 3136
rect 186828 3058 187132 3074
rect 186816 3052 187132 3058
rect 186868 3046 187132 3052
rect 186816 2994 186868 3000
rect 187104 2990 187132 3046
rect 187092 2984 187144 2990
rect 187092 2926 187144 2932
rect 186644 598 186764 626
rect 186644 592 186672 598
rect 186552 564 186672 592
rect 186552 480 186580 564
rect 187748 480 187776 4791
rect 188944 480 188972 5782
rect 190416 610 190444 9574
rect 191796 9042 191824 10095
rect 191784 9036 191836 9042
rect 191784 8978 191836 8984
rect 194924 7750 194952 323546
rect 197764 318164 197816 318170
rect 197764 318106 197816 318112
rect 196382 10704 196438 10713
rect 196382 10639 196438 10648
rect 196396 10266 196424 10639
rect 196474 10432 196530 10441
rect 196474 10367 196530 10376
rect 196384 10260 196436 10266
rect 196384 10202 196436 10208
rect 195924 10192 195976 10198
rect 195922 10160 195924 10169
rect 196488 10169 196516 10367
rect 195976 10160 195978 10169
rect 196474 10160 196530 10169
rect 195922 10095 195978 10104
rect 196016 10124 196068 10130
rect 196474 10095 196530 10104
rect 196016 10066 196068 10072
rect 196028 10033 196056 10066
rect 196014 10024 196070 10033
rect 196014 9959 196070 9968
rect 196292 7880 196344 7886
rect 196290 7848 196292 7857
rect 196344 7848 196346 7857
rect 196290 7783 196346 7792
rect 193624 7744 193676 7750
rect 193622 7712 193624 7721
rect 193716 7744 193768 7750
rect 193676 7712 193678 7721
rect 193716 7686 193768 7692
rect 194912 7744 194964 7750
rect 194912 7686 194964 7692
rect 193622 7647 193678 7656
rect 192520 5772 192572 5778
rect 192520 5714 192572 5720
rect 191324 5364 191376 5370
rect 191324 5306 191376 5312
rect 190128 604 190180 610
rect 190128 546 190180 552
rect 190404 604 190456 610
rect 190404 546 190456 552
rect 190140 480 190168 546
rect 191336 480 191364 5306
rect 192532 480 192560 5714
rect 193728 480 193756 7686
rect 195004 4752 195056 4758
rect 195004 4694 195056 4700
rect 195016 2394 195044 4694
rect 196384 4208 196436 4214
rect 196384 4150 196436 4156
rect 196476 4208 196528 4214
rect 196476 4150 196528 4156
rect 196396 3466 196424 4150
rect 196488 3466 196516 4150
rect 196292 3460 196344 3466
rect 196292 3402 196344 3408
rect 196384 3460 196436 3466
rect 196384 3402 196436 3408
rect 196476 3460 196528 3466
rect 196476 3402 196528 3408
rect 196198 3224 196254 3233
rect 196198 3159 196200 3168
rect 196252 3159 196254 3168
rect 196200 3130 196252 3136
rect 195924 2984 195976 2990
rect 195922 2952 195924 2961
rect 195976 2952 195978 2961
rect 195922 2887 195978 2896
rect 196304 2836 196332 3402
rect 196750 3224 196806 3233
rect 196750 3159 196752 3168
rect 196804 3159 196806 3168
rect 196752 3130 196804 3136
rect 196384 2848 196436 2854
rect 196304 2808 196384 2836
rect 196384 2790 196436 2796
rect 196108 2644 196160 2650
rect 196108 2586 196160 2592
rect 194924 2366 195044 2394
rect 194924 480 194952 2366
rect 196120 480 196148 2586
rect 197776 610 197804 318106
rect 201904 315376 201956 315382
rect 201904 315318 201956 315324
rect 199696 5636 199748 5642
rect 199696 5578 199748 5584
rect 198500 4684 198552 4690
rect 198500 4626 198552 4632
rect 197304 604 197356 610
rect 197304 546 197356 552
rect 197764 604 197816 610
rect 197764 546 197816 552
rect 197316 480 197344 546
rect 198512 480 198540 4626
rect 199708 480 199736 5578
rect 201916 610 201944 315318
rect 203192 5568 203244 5574
rect 203192 5510 203244 5516
rect 201996 4616 202048 4622
rect 201996 4558 202048 4564
rect 200892 604 200944 610
rect 200892 546 200944 552
rect 201904 604 201956 610
rect 201904 546 201956 552
rect 200904 480 200932 546
rect 202008 480 202036 4558
rect 203204 480 203232 5510
rect 204676 626 204704 333338
rect 218464 327888 218516 327894
rect 218464 327830 218516 327836
rect 214324 327140 214376 327146
rect 214324 327082 214376 327088
rect 214336 317422 214364 327082
rect 214324 317416 214376 317422
rect 214324 317358 214376 317364
rect 214324 307828 214376 307834
rect 214324 307770 214376 307776
rect 214336 298081 214364 307770
rect 214322 298072 214378 298081
rect 214322 298007 214378 298016
rect 214506 298072 214562 298081
rect 214506 298007 214562 298016
rect 214520 288454 214548 298007
rect 214324 288448 214376 288454
rect 214324 288390 214376 288396
rect 214508 288448 214560 288454
rect 214508 288390 214560 288396
rect 214336 278769 214364 288390
rect 214322 278760 214378 278769
rect 214322 278695 214378 278704
rect 214506 278760 214562 278769
rect 214506 278695 214562 278704
rect 214520 269142 214548 278695
rect 214324 269136 214376 269142
rect 214324 269078 214376 269084
rect 214508 269136 214560 269142
rect 214508 269078 214560 269084
rect 214336 259457 214364 269078
rect 214322 259448 214378 259457
rect 214322 259383 214378 259392
rect 214506 259448 214562 259457
rect 214506 259383 214562 259392
rect 214520 249830 214548 259383
rect 214324 249824 214376 249830
rect 214324 249766 214376 249772
rect 214508 249824 214560 249830
rect 214508 249766 214560 249772
rect 214336 240145 214364 249766
rect 214322 240136 214378 240145
rect 214322 240071 214378 240080
rect 214506 240136 214562 240145
rect 214506 240071 214562 240080
rect 214520 230518 214548 240071
rect 214324 230512 214376 230518
rect 214324 230454 214376 230460
rect 214508 230512 214560 230518
rect 214508 230454 214560 230460
rect 214336 220833 214364 230454
rect 214322 220824 214378 220833
rect 214322 220759 214378 220768
rect 214506 220824 214562 220833
rect 214506 220759 214562 220768
rect 214520 211177 214548 220759
rect 214322 211168 214378 211177
rect 214322 211103 214378 211112
rect 214506 211168 214562 211177
rect 214506 211103 214562 211112
rect 214336 201482 214364 211103
rect 214324 201476 214376 201482
rect 214324 201418 214376 201424
rect 214508 201476 214560 201482
rect 214508 201418 214560 201424
rect 214520 191865 214548 201418
rect 214322 191856 214378 191865
rect 214322 191791 214378 191800
rect 214506 191856 214562 191865
rect 214506 191791 214562 191800
rect 214336 182170 214364 191791
rect 214324 182164 214376 182170
rect 214324 182106 214376 182112
rect 214508 182164 214560 182170
rect 214508 182106 214560 182112
rect 214520 172553 214548 182106
rect 214322 172544 214378 172553
rect 214322 172479 214378 172488
rect 214506 172544 214562 172553
rect 214506 172479 214562 172488
rect 214336 162858 214364 172479
rect 214324 162852 214376 162858
rect 214324 162794 214376 162800
rect 214324 153264 214376 153270
rect 214324 153206 214376 153212
rect 214336 143478 214364 153206
rect 214324 143472 214376 143478
rect 214324 143414 214376 143420
rect 214324 133952 214376 133958
rect 214324 133894 214376 133900
rect 214336 124166 214364 133894
rect 214324 124160 214376 124166
rect 214324 124102 214376 124108
rect 214324 114572 214376 114578
rect 214324 114514 214376 114520
rect 214336 104854 214364 114514
rect 214324 104848 214376 104854
rect 214324 104790 214376 104796
rect 214324 95328 214376 95334
rect 214324 95270 214376 95276
rect 214336 85542 214364 95270
rect 214324 85536 214376 85542
rect 214324 85478 214376 85484
rect 214324 75948 214376 75954
rect 214324 75890 214376 75896
rect 214336 66230 214364 75890
rect 214324 66224 214376 66230
rect 214324 66166 214376 66172
rect 214324 56704 214376 56710
rect 214324 56646 214376 56652
rect 214336 46918 214364 56646
rect 214324 46912 214376 46918
rect 214324 46854 214376 46860
rect 214324 37324 214376 37330
rect 214324 37266 214376 37272
rect 214336 27606 214364 37266
rect 214324 27600 214376 27606
rect 214324 27542 214376 27548
rect 214508 27600 214560 27606
rect 214508 27542 214560 27548
rect 206318 10432 206374 10441
rect 206318 10367 206374 10376
rect 206332 10169 206360 10367
rect 206318 10160 206374 10169
rect 206318 10095 206374 10104
rect 214520 9761 214548 27542
rect 215980 11212 216032 11218
rect 215980 11154 216032 11160
rect 215796 11076 215848 11082
rect 215796 11018 215848 11024
rect 215808 10033 215836 11018
rect 215794 10024 215850 10033
rect 215794 9959 215850 9968
rect 215992 9897 216020 11154
rect 216162 10432 216218 10441
rect 216162 10367 216218 10376
rect 216176 10169 216204 10367
rect 216162 10160 216218 10169
rect 216162 10095 216218 10104
rect 215978 9888 216034 9897
rect 215978 9823 216034 9832
rect 213954 9752 214010 9761
rect 213954 9687 214010 9696
rect 214506 9752 214562 9761
rect 214506 9687 214562 9696
rect 207976 8628 208028 8634
rect 207976 8570 208028 8576
rect 206778 5944 206834 5953
rect 206778 5879 206834 5888
rect 205584 4548 205636 4554
rect 205584 4490 205636 4496
rect 204400 598 204704 626
rect 204400 480 204428 598
rect 205596 480 205624 4490
rect 206044 4208 206096 4214
rect 206044 4150 206096 4156
rect 206056 3466 206084 4150
rect 206228 3528 206280 3534
rect 206228 3470 206280 3476
rect 206044 3460 206096 3466
rect 206044 3402 206096 3408
rect 206240 3233 206268 3470
rect 205858 3224 205914 3233
rect 205858 3159 205860 3168
rect 205912 3159 205914 3168
rect 206226 3224 206282 3233
rect 206226 3159 206282 3168
rect 205860 3130 205912 3136
rect 206792 480 206820 5879
rect 207700 3052 207752 3058
rect 207700 2994 207752 3000
rect 207712 2961 207740 2994
rect 207698 2952 207754 2961
rect 207698 2887 207754 2896
rect 207988 480 208016 8570
rect 211564 8560 211616 8566
rect 211564 8502 211616 8508
rect 210366 5808 210422 5817
rect 210366 5743 210422 5752
rect 209172 4480 209224 4486
rect 209172 4422 209224 4428
rect 208158 3360 208214 3369
rect 208158 3295 208214 3304
rect 208172 2553 208200 3295
rect 208158 2544 208214 2553
rect 208158 2479 208214 2488
rect 209184 480 209212 4422
rect 210276 3664 210328 3670
rect 210276 3606 210328 3612
rect 210288 3097 210316 3606
rect 210274 3088 210330 3097
rect 210274 3023 210330 3032
rect 210380 480 210408 5743
rect 211576 480 211604 8502
rect 212760 4208 212812 4214
rect 212760 4150 212812 4156
rect 212772 480 212800 4150
rect 213968 480 213996 9687
rect 215152 8424 215204 8430
rect 215152 8366 215204 8372
rect 215164 480 215192 8366
rect 215794 7984 215850 7993
rect 215794 7919 215850 7928
rect 215808 7886 215836 7919
rect 215796 7880 215848 7886
rect 215796 7822 215848 7828
rect 215888 7880 215940 7886
rect 215888 7822 215940 7828
rect 215900 7721 215928 7822
rect 215886 7712 215942 7721
rect 215886 7647 215942 7656
rect 215796 6316 215848 6322
rect 215796 6258 215848 6264
rect 215808 6089 215836 6258
rect 215888 6180 215940 6186
rect 215888 6122 215940 6128
rect 215794 6080 215850 6089
rect 215794 6015 215850 6024
rect 215900 5953 215928 6122
rect 215886 5944 215942 5953
rect 215886 5879 215942 5888
rect 216346 4312 216402 4321
rect 216346 4247 216402 4256
rect 215794 4176 215850 4185
rect 215794 4111 215850 4120
rect 215808 4010 215836 4111
rect 215796 4004 215848 4010
rect 215796 3946 215848 3952
rect 215888 4004 215940 4010
rect 215888 3946 215940 3952
rect 215796 3664 215848 3670
rect 215900 3652 215928 3946
rect 215848 3624 215928 3652
rect 215796 3606 215848 3612
rect 216360 480 216388 4247
rect 218476 4010 218504 327830
rect 219212 59226 219240 458458
rect 220592 427786 220620 461450
rect 228860 460352 228912 460358
rect 228860 460294 228912 460300
rect 227572 460080 227624 460086
rect 227572 460022 227624 460028
rect 223340 460012 223392 460018
rect 223340 459954 223392 459960
rect 221960 458720 222012 458726
rect 221960 458662 222012 458668
rect 220580 427780 220632 427786
rect 220580 427722 220632 427728
rect 221972 378010 222000 458662
rect 221960 378004 222012 378010
rect 221960 377946 222012 377952
rect 223352 361554 223380 459954
rect 224720 459808 224772 459814
rect 224720 459750 224772 459756
rect 223340 361548 223392 361554
rect 223340 361490 223392 361496
rect 219844 338156 219896 338162
rect 219844 338098 219896 338104
rect 219856 337958 219884 338098
rect 219844 337952 219896 337958
rect 219844 337894 219896 337900
rect 219934 337784 219990 337793
rect 219934 337719 219990 337728
rect 219948 337618 219976 337719
rect 219752 337612 219804 337618
rect 219752 337554 219804 337560
rect 219936 337612 219988 337618
rect 219936 337554 219988 337560
rect 220028 337612 220080 337618
rect 220028 337554 220080 337560
rect 219764 337521 219792 337554
rect 220040 337521 220068 337554
rect 219566 337512 219622 337521
rect 219750 337512 219806 337521
rect 219622 337482 219700 337498
rect 219622 337476 219712 337482
rect 219622 337470 219660 337476
rect 219566 337447 219622 337456
rect 219750 337447 219806 337456
rect 220026 337512 220082 337521
rect 220026 337447 220082 337456
rect 219660 337418 219712 337424
rect 219844 337408 219896 337414
rect 219844 337350 219896 337356
rect 219856 337249 219884 337350
rect 219842 337240 219898 337249
rect 219842 337175 219898 337184
rect 221224 329248 221276 329254
rect 221224 329190 221276 329196
rect 219200 59220 219252 59226
rect 219200 59162 219252 59168
rect 218556 8356 218608 8362
rect 218556 8298 218608 8304
rect 217544 4004 217596 4010
rect 217544 3946 217596 3952
rect 218464 4004 218516 4010
rect 218464 3946 218516 3952
rect 217556 480 217584 3946
rect 218568 2802 218596 8298
rect 219658 4720 219714 4729
rect 219658 4655 219714 4664
rect 218646 4312 218702 4321
rect 218646 4247 218648 4256
rect 218700 4247 218702 4256
rect 218648 4218 218700 4224
rect 218568 2774 218688 2802
rect 218660 480 218688 2774
rect 219672 1306 219700 4655
rect 219750 4176 219806 4185
rect 219750 4111 219806 4120
rect 219764 4010 219792 4111
rect 219752 4004 219804 4010
rect 219752 3946 219804 3952
rect 220028 3664 220080 3670
rect 220028 3606 220080 3612
rect 220040 2650 220068 3606
rect 220028 2644 220080 2650
rect 220028 2586 220080 2592
rect 219672 1278 219884 1306
rect 219856 480 219884 1278
rect 221236 610 221264 329190
rect 224732 209778 224760 459750
rect 227480 458992 227532 458998
rect 227480 458934 227532 458940
rect 226192 458856 226244 458862
rect 226192 458798 226244 458804
rect 226100 458788 226152 458794
rect 226100 458730 226152 458736
rect 225364 336320 225416 336326
rect 225364 336262 225416 336268
rect 225376 309126 225404 336262
rect 226112 310486 226140 458730
rect 226204 411194 226232 458798
rect 226192 411188 226244 411194
rect 226192 411130 226244 411136
rect 226926 337648 226982 337657
rect 226926 337583 226982 337592
rect 226940 337482 226968 337583
rect 226928 337476 226980 337482
rect 226928 337418 226980 337424
rect 226100 310480 226152 310486
rect 226100 310422 226152 310428
rect 225364 309120 225416 309126
rect 225364 309062 225416 309068
rect 225364 299532 225416 299538
rect 225364 299474 225416 299480
rect 225376 270502 225404 299474
rect 225364 270496 225416 270502
rect 225364 270438 225416 270444
rect 225364 260908 225416 260914
rect 225364 260850 225416 260856
rect 225376 251190 225404 260850
rect 225364 251184 225416 251190
rect 225364 251126 225416 251132
rect 225364 241664 225416 241670
rect 225364 241606 225416 241612
rect 225376 212537 225404 241606
rect 225362 212528 225418 212537
rect 225362 212463 225418 212472
rect 225546 212528 225602 212537
rect 225546 212463 225602 212472
rect 224720 209772 224772 209778
rect 224720 209714 224772 209720
rect 225560 203046 225588 212463
rect 225364 203040 225416 203046
rect 225364 202982 225416 202988
rect 225548 203040 225600 203046
rect 225548 202982 225600 202988
rect 225376 173913 225404 202982
rect 225362 173904 225418 173913
rect 225362 173839 225418 173848
rect 225362 164248 225418 164257
rect 225362 164183 225418 164192
rect 225376 144906 225404 164183
rect 225364 144900 225416 144906
rect 225364 144842 225416 144848
rect 227492 143546 227520 458934
rect 227584 394670 227612 460022
rect 227572 394664 227624 394670
rect 227572 394606 227624 394612
rect 228872 244186 228900 460294
rect 228964 343602 228992 461518
rect 240268 461440 240320 461446
rect 240268 461382 240320 461388
rect 235024 461236 235076 461242
rect 235024 461178 235076 461184
rect 235036 459884 235064 461178
rect 240280 459884 240308 461382
rect 243488 460148 243540 460154
rect 243488 460090 243540 460096
rect 243500 459884 243528 460090
rect 252780 459944 252832 459950
rect 247746 459882 248128 459898
rect 252832 459892 252990 459898
rect 252780 459886 252990 459892
rect 247746 459876 248140 459882
rect 247746 459870 248088 459876
rect 252792 459870 252990 459886
rect 253988 459884 254016 463286
rect 255080 462868 255132 462874
rect 255080 462810 255132 462816
rect 255092 459884 255120 462810
rect 257116 459884 257144 463558
rect 258208 463412 258260 463418
rect 258208 463354 258260 463360
rect 258220 459884 258248 463354
rect 261336 463140 261388 463146
rect 261336 463082 261388 463088
rect 259220 461168 259272 461174
rect 259220 461110 259272 461116
rect 259232 459884 259260 461110
rect 260324 460964 260376 460970
rect 260324 460906 260376 460912
rect 260336 459884 260364 460906
rect 261348 459884 261376 463082
rect 262636 459898 262664 476070
rect 264016 460034 264044 507826
rect 265384 492720 265436 492726
rect 265384 492662 265436 492668
rect 265396 463078 265424 492662
rect 266684 463078 266712 522990
rect 264556 463072 264608 463078
rect 264556 463014 264608 463020
rect 265384 463072 265436 463078
rect 265384 463014 265436 463020
rect 265568 463072 265620 463078
rect 265568 463014 265620 463020
rect 266672 463072 266724 463078
rect 266672 463014 266724 463020
rect 263740 460006 264044 460034
rect 263740 459898 263768 460006
rect 262466 459870 262664 459898
rect 263478 459870 263768 459898
rect 264568 459884 264596 463014
rect 265580 459884 265608 463014
rect 266776 459898 266804 554746
rect 268144 539776 268196 539782
rect 268144 539718 268196 539724
rect 268156 460034 268184 539718
rect 269536 463078 269564 569910
rect 268696 463072 268748 463078
rect 268696 463014 268748 463020
rect 269524 463072 269576 463078
rect 269524 463014 269576 463020
rect 269800 463072 269852 463078
rect 269800 463014 269852 463020
rect 268064 460006 268184 460034
rect 268064 459898 268092 460006
rect 266606 459870 266804 459898
rect 267710 459870 268092 459898
rect 268708 459884 268736 463014
rect 269812 459884 269840 463014
rect 270824 459884 270852 586502
rect 270916 463078 270944 601734
rect 270904 463072 270956 463078
rect 270904 463014 270956 463020
rect 272296 459898 272324 616966
rect 273676 463078 273704 648586
rect 274952 633480 275004 633486
rect 274952 633422 275004 633428
rect 274964 463078 274992 633422
rect 272928 463072 272980 463078
rect 272928 463014 272980 463020
rect 273664 463072 273716 463078
rect 273664 463014 273716 463020
rect 273940 463072 273992 463078
rect 273940 463014 273992 463020
rect 274952 463072 275004 463078
rect 274952 463014 275004 463020
rect 271942 459870 272324 459898
rect 272940 459884 272968 463014
rect 273952 459884 273980 463014
rect 275056 459884 275084 663750
rect 276436 459898 276464 695506
rect 277804 680400 277856 680406
rect 277804 680342 277856 680348
rect 277816 460034 277844 680342
rect 278172 463140 278224 463146
rect 278172 463082 278224 463088
rect 277540 460006 277844 460034
rect 277540 459898 277568 460006
rect 276082 459870 276464 459898
rect 277186 459870 277568 459898
rect 278184 459884 278212 463082
rect 279276 463072 279328 463078
rect 279276 463014 279328 463020
rect 279288 459884 279316 463014
rect 280484 459898 280512 700334
rect 280576 463078 280604 700402
rect 283324 699916 283376 699922
rect 283324 699858 283376 699864
rect 283336 463146 283364 699858
rect 283600 463276 283652 463282
rect 283600 463218 283652 463224
rect 283612 463185 283640 463218
rect 283598 463176 283654 463185
rect 282312 463140 282364 463146
rect 282312 463082 282364 463088
rect 282404 463140 282456 463146
rect 282404 463082 282456 463088
rect 283324 463140 283376 463146
rect 283324 463082 283376 463088
rect 283416 463140 283468 463146
rect 283598 463111 283654 463120
rect 283416 463082 283468 463088
rect 280564 463072 280616 463078
rect 280564 463014 280616 463020
rect 281392 463072 281444 463078
rect 282324 463049 282352 463082
rect 281392 463014 281444 463020
rect 282310 463040 282366 463049
rect 280314 459870 280512 459898
rect 281404 459884 281432 463014
rect 282310 462975 282366 462984
rect 282416 459884 282444 463082
rect 283428 463049 283456 463082
rect 284716 463078 284744 700878
rect 286084 700868 286136 700874
rect 286084 700810 286136 700816
rect 288844 700868 288896 700874
rect 288844 700810 288896 700816
rect 283784 463072 283836 463078
rect 283414 463040 283470 463049
rect 283784 463014 283836 463020
rect 284704 463072 284756 463078
rect 284704 463014 284756 463020
rect 283414 462975 283470 462984
rect 283796 459898 283824 463014
rect 284704 462256 284756 462262
rect 284704 462198 284756 462204
rect 284716 459898 284744 462198
rect 283442 459870 283824 459898
rect 284546 459870 284744 459898
rect 248088 459818 248140 459824
rect 286096 459762 286124 700810
rect 287464 699984 287516 699990
rect 287464 699926 287516 699932
rect 287476 463078 287504 699926
rect 288198 463176 288254 463185
rect 288382 463176 288438 463185
rect 288198 463111 288200 463120
rect 288252 463111 288254 463120
rect 288304 463134 288382 463162
rect 288200 463082 288252 463088
rect 286636 463072 286688 463078
rect 286636 463014 286688 463020
rect 287464 463072 287516 463078
rect 287464 463014 287516 463020
rect 286648 459884 286676 463014
rect 288304 460034 288332 463134
rect 288382 463111 288438 463120
rect 288120 460006 288332 460034
rect 288120 459898 288148 460006
rect 288856 459898 288884 700810
rect 290224 699848 290276 699854
rect 290224 699790 290276 699796
rect 287674 459870 288148 459898
rect 288778 459870 288884 459898
rect 290236 459762 290264 699790
rect 291788 699780 291840 699786
rect 291788 699722 291840 699728
rect 291696 699712 291748 699718
rect 291696 699654 291748 699660
rect 291708 463146 291736 699654
rect 291696 463140 291748 463146
rect 291696 463082 291748 463088
rect 291144 462324 291196 462330
rect 291144 462266 291196 462272
rect 291156 459898 291184 462266
rect 290894 459870 291184 459898
rect 291800 459898 291828 699722
rect 292444 699718 292472 703520
rect 314064 703474 314092 703520
rect 313972 703446 314092 703474
rect 299976 701004 300028 701010
rect 299976 700946 300028 700952
rect 298596 700256 298648 700262
rect 298596 700198 298648 700204
rect 294456 699916 294508 699922
rect 294456 699858 294508 699864
rect 292524 699848 292576 699854
rect 292524 699790 292576 699796
rect 292536 699718 292564 699790
rect 292432 699712 292484 699718
rect 292432 699654 292484 699660
rect 292524 699712 292576 699718
rect 292524 699654 292576 699660
rect 293076 463276 293128 463282
rect 293076 463218 293128 463224
rect 293168 463276 293220 463282
rect 293168 463218 293220 463224
rect 292524 463140 292576 463146
rect 292524 463082 292576 463088
rect 292536 459898 292564 463082
rect 293088 459898 293116 463218
rect 293180 463185 293208 463218
rect 293166 463176 293222 463185
rect 293166 463111 293222 463120
rect 291800 459870 291906 459898
rect 292536 459870 292918 459898
rect 293088 459870 294022 459898
rect 285558 459734 286124 459762
rect 289790 459734 290264 459762
rect 294468 459762 294496 699858
rect 295928 699780 295980 699786
rect 295928 699722 295980 699728
rect 297216 699780 297268 699786
rect 297216 699722 297268 699728
rect 295940 459898 295968 699722
rect 296756 462188 296808 462194
rect 296756 462130 296808 462136
rect 296768 459898 296796 462130
rect 297228 460034 297256 699722
rect 297228 460006 297716 460034
rect 295940 459870 296138 459898
rect 296768 459870 297150 459898
rect 297688 459762 297716 460006
rect 298608 459762 298636 700198
rect 299988 459898 300016 700946
rect 301356 700800 301408 700806
rect 301356 700742 301408 700748
rect 301368 463146 301396 700742
rect 301448 700596 301500 700602
rect 301448 700538 301500 700544
rect 301356 463140 301408 463146
rect 301356 463082 301408 463088
rect 301460 459898 301488 700538
rect 302736 700528 302788 700534
rect 302736 700470 302788 700476
rect 302092 463140 302144 463146
rect 302092 463082 302144 463088
rect 299988 459870 300278 459898
rect 301382 459870 301488 459898
rect 302104 459898 302132 463082
rect 302748 460034 302776 700470
rect 304114 700360 304170 700369
rect 304114 700295 304170 700304
rect 305496 700324 305548 700330
rect 302748 460006 302960 460034
rect 302104 459870 302394 459898
rect 302932 459762 302960 460006
rect 304128 459898 304156 700295
rect 305496 700266 305548 700272
rect 305508 459898 305536 700266
rect 305588 694272 305640 694278
rect 305588 694214 305640 694220
rect 305600 460306 305628 694214
rect 313972 688650 314000 703446
rect 335684 699854 335712 703520
rect 335672 699848 335724 699854
rect 335672 699790 335724 699796
rect 357304 699718 357332 703520
rect 378924 702386 378952 703520
rect 378740 702358 378952 702386
rect 357292 699712 357344 699718
rect 357292 699654 357344 699660
rect 378740 695502 378768 702358
rect 400636 699922 400664 703520
rect 422256 699990 422284 703520
rect 443876 703474 443904 703520
rect 443692 703446 443904 703474
rect 422244 699984 422296 699990
rect 422244 699926 422296 699932
rect 400624 699916 400676 699922
rect 400624 699858 400676 699864
rect 378728 695496 378780 695502
rect 378728 695438 378780 695444
rect 443692 688650 443720 703446
rect 465496 700942 465524 703520
rect 465484 700936 465536 700942
rect 465484 700878 465536 700884
rect 487116 700874 487144 703520
rect 508736 702386 508764 703520
rect 508460 702358 508764 702386
rect 487104 700868 487156 700874
rect 487104 700810 487156 700816
rect 508460 695502 508488 702358
rect 530356 700466 530384 703520
rect 530344 700460 530396 700466
rect 530344 700402 530396 700408
rect 551976 700398 552004 703520
rect 573596 703474 573624 703520
rect 573412 703446 573624 703474
rect 551964 700392 552016 700398
rect 551964 700334 552016 700340
rect 508448 695496 508500 695502
rect 508448 695438 508500 695444
rect 573412 688650 573440 703446
rect 580114 696008 580170 696017
rect 580114 695943 580170 695952
rect 580128 695570 580156 695943
rect 580116 695564 580168 695570
rect 580116 695506 580168 695512
rect 313972 688634 314092 688650
rect 443692 688634 443812 688650
rect 573412 688634 573532 688650
rect 313972 688628 314104 688634
rect 313972 688622 314052 688628
rect 314052 688570 314104 688576
rect 314236 688628 314288 688634
rect 443692 688628 443824 688634
rect 443692 688622 443772 688628
rect 314236 688570 314288 688576
rect 443772 688570 443824 688576
rect 443956 688628 444008 688634
rect 573412 688628 573544 688634
rect 573412 688622 573492 688628
rect 443956 688570 444008 688576
rect 573492 688570 573544 688576
rect 573676 688628 573728 688634
rect 573676 688570 573728 688576
rect 314064 688539 314092 688570
rect 314248 681034 314276 688570
rect 443784 688539 443812 688570
rect 378820 685908 378872 685914
rect 378820 685850 378872 685856
rect 314156 681006 314276 681034
rect 308256 677612 308308 677618
rect 308256 677554 308308 677560
rect 306876 661088 306928 661094
rect 306876 661030 306928 661036
rect 305600 460278 306364 460306
rect 306336 459898 306364 460278
rect 306888 459898 306916 661030
rect 308268 459898 308296 677554
rect 314156 676122 314184 681006
rect 378832 679130 378860 685850
rect 443968 681034 443996 688570
rect 573504 688539 573532 688570
rect 508540 685908 508592 685914
rect 508540 685850 508592 685856
rect 378740 679102 378860 679130
rect 443876 681006 443996 681034
rect 378740 678858 378768 679102
rect 378648 678830 378768 678858
rect 378648 676122 378676 678830
rect 443876 676122 443904 681006
rect 508552 679130 508580 685850
rect 573688 681034 573716 688570
rect 508460 679102 508580 679130
rect 573596 681006 573716 681034
rect 508460 678858 508488 679102
rect 508368 678830 508488 678858
rect 508368 676122 508396 678830
rect 573596 676122 573624 681006
rect 580116 680400 580168 680406
rect 580114 680368 580116 680377
rect 580168 680368 580170 680377
rect 580114 680303 580170 680312
rect 314144 676116 314196 676122
rect 314144 676058 314196 676064
rect 378636 676116 378688 676122
rect 378636 676058 378688 676064
rect 443864 676116 443916 676122
rect 443864 676058 443916 676064
rect 508356 676116 508408 676122
rect 508356 676058 508408 676064
rect 573584 676116 573636 676122
rect 573584 676058 573636 676064
rect 314236 666596 314288 666602
rect 314236 666538 314288 666544
rect 378728 666596 378780 666602
rect 378728 666538 378780 666544
rect 443956 666596 444008 666602
rect 443956 666538 444008 666544
rect 508448 666596 508500 666602
rect 508448 666538 508500 666544
rect 573676 666596 573728 666602
rect 573676 666538 573728 666544
rect 314248 659682 314276 666538
rect 378740 659734 378768 666538
rect 314064 659654 314276 659682
rect 378728 659728 378780 659734
rect 378728 659670 378780 659676
rect 378820 659728 378872 659734
rect 443968 659682 443996 666538
rect 508460 659734 508488 666538
rect 378820 659670 378872 659676
rect 314064 647290 314092 659654
rect 378832 654158 378860 659670
rect 443784 659654 443996 659682
rect 508448 659728 508500 659734
rect 508448 659670 508500 659676
rect 508540 659728 508592 659734
rect 573688 659682 573716 666538
rect 580114 664728 580170 664737
rect 580114 664663 580170 664672
rect 580128 663814 580156 664663
rect 580116 663808 580168 663814
rect 580116 663750 580168 663756
rect 508540 659670 508592 659676
rect 378636 654152 378688 654158
rect 378636 654094 378688 654100
rect 378820 654152 378872 654158
rect 378820 654094 378872 654100
rect 313960 647284 314012 647290
rect 313960 647226 314012 647232
rect 314052 647284 314104 647290
rect 314052 647226 314104 647232
rect 309636 644496 309688 644502
rect 309636 644438 309688 644444
rect 309648 459898 309676 644438
rect 313972 640370 314000 647226
rect 378648 644450 378676 654094
rect 443784 647290 443812 659654
rect 508552 654158 508580 659670
rect 573504 659654 573716 659682
rect 508356 654152 508408 654158
rect 508356 654094 508408 654100
rect 508540 654152 508592 654158
rect 508540 654094 508592 654100
rect 443680 647284 443732 647290
rect 443680 647226 443732 647232
rect 443772 647284 443824 647290
rect 443772 647226 443824 647232
rect 378648 644422 378860 644450
rect 313972 640342 314184 640370
rect 314156 637498 314184 640342
rect 314144 637492 314196 637498
rect 314144 637434 314196 637440
rect 311016 627972 311068 627978
rect 311016 627914 311068 627920
rect 314236 627972 314288 627978
rect 314236 627914 314288 627920
rect 309728 611380 309780 611386
rect 309728 611322 309780 611328
rect 309740 460442 309768 611322
rect 309740 460414 310596 460442
rect 310568 459898 310596 460414
rect 304128 459870 304510 459898
rect 305508 459870 305614 459898
rect 306336 459870 306626 459898
rect 306888 459870 307730 459898
rect 308268 459870 308742 459898
rect 309648 459870 309754 459898
rect 310568 459870 310858 459898
rect 311028 459762 311056 627914
rect 314248 618322 314276 627914
rect 314052 618316 314104 618322
rect 314052 618258 314104 618264
rect 314236 618316 314288 618322
rect 314236 618258 314288 618264
rect 314064 618225 314092 618258
rect 313774 618216 313830 618225
rect 313774 618151 313830 618160
rect 314050 618216 314106 618225
rect 314050 618151 314106 618160
rect 313788 608666 313816 618151
rect 378832 615534 378860 644422
rect 443692 640370 443720 647226
rect 508368 644450 508396 654094
rect 573504 647290 573532 659654
rect 580114 649088 580170 649097
rect 580114 649023 580170 649032
rect 580128 648650 580156 649023
rect 580116 648644 580168 648650
rect 580116 648586 580168 648592
rect 573400 647284 573452 647290
rect 573400 647226 573452 647232
rect 573492 647284 573544 647290
rect 573492 647226 573544 647232
rect 508368 644422 508580 644450
rect 443692 640342 443904 640370
rect 443876 637498 443904 640342
rect 443864 637492 443916 637498
rect 443864 637434 443916 637440
rect 443956 627972 444008 627978
rect 443956 627914 444008 627920
rect 443968 618322 443996 627914
rect 443772 618316 443824 618322
rect 443772 618258 443824 618264
rect 443956 618316 444008 618322
rect 443956 618258 444008 618264
rect 443784 618225 443812 618258
rect 443770 618216 443826 618225
rect 443770 618151 443826 618160
rect 508552 615534 508580 644422
rect 573412 640370 573440 647226
rect 573412 640342 573624 640370
rect 573596 637498 573624 640342
rect 573584 637492 573636 637498
rect 573584 637434 573636 637440
rect 580116 633480 580168 633486
rect 580114 633448 580116 633457
rect 580168 633448 580170 633457
rect 580114 633383 580170 633392
rect 573676 627972 573728 627978
rect 573676 627914 573728 627920
rect 573688 618322 573716 627914
rect 573492 618316 573544 618322
rect 573492 618258 573544 618264
rect 573676 618316 573728 618322
rect 573676 618258 573728 618264
rect 573504 618186 573532 618258
rect 573492 618180 573544 618186
rect 573492 618122 573544 618128
rect 573768 618180 573820 618186
rect 573768 618122 573820 618128
rect 378636 615528 378688 615534
rect 378636 615470 378688 615476
rect 378820 615528 378872 615534
rect 378820 615470 378872 615476
rect 508356 615528 508408 615534
rect 508356 615470 508408 615476
rect 508540 615528 508592 615534
rect 508540 615470 508592 615476
rect 313776 608660 313828 608666
rect 313776 608602 313828 608608
rect 313960 608660 314012 608666
rect 313960 608602 314012 608608
rect 313972 601746 314000 608602
rect 378648 605826 378676 615470
rect 443678 608696 443734 608705
rect 443678 608631 443734 608640
rect 443692 608598 443720 608631
rect 443680 608592 443732 608598
rect 443680 608534 443732 608540
rect 508368 605826 508396 615470
rect 573780 608705 573808 618122
rect 580114 617808 580170 617817
rect 580114 617743 580170 617752
rect 580128 617030 580156 617743
rect 580116 617024 580168 617030
rect 580116 616966 580168 616972
rect 573398 608696 573454 608705
rect 573398 608631 573454 608640
rect 573766 608696 573822 608705
rect 573766 608631 573822 608640
rect 573412 608598 573440 608631
rect 573400 608592 573452 608598
rect 573400 608534 573452 608540
rect 378648 605798 378860 605826
rect 508368 605798 508580 605826
rect 313880 601718 314000 601746
rect 313880 598874 313908 601718
rect 313868 598868 313920 598874
rect 313868 598810 313920 598816
rect 312396 594856 312448 594862
rect 312396 594798 312448 594804
rect 312408 460034 312436 594798
rect 378832 591954 378860 605798
rect 443864 601588 443916 601594
rect 443864 601530 443916 601536
rect 443876 598874 443904 601530
rect 443864 598868 443916 598874
rect 443864 598810 443916 598816
rect 508552 591954 508580 605798
rect 580114 602168 580170 602177
rect 580114 602103 580170 602112
rect 580128 601798 580156 602103
rect 580116 601792 580168 601798
rect 580116 601734 580168 601740
rect 573584 601588 573636 601594
rect 573584 601530 573636 601536
rect 573596 598874 573624 601530
rect 573584 598868 573636 598874
rect 573584 598810 573636 598816
rect 378740 591926 378860 591954
rect 508460 591926 508580 591954
rect 314052 589348 314104 589354
rect 314052 589290 314104 589296
rect 314064 582418 314092 589290
rect 378740 589286 378768 591926
rect 443956 589348 444008 589354
rect 443956 589290 444008 589296
rect 378728 589280 378780 589286
rect 378728 589222 378780 589228
rect 443968 582486 443996 589290
rect 508460 589286 508488 591926
rect 573676 589348 573728 589354
rect 573676 589290 573728 589296
rect 508448 589280 508500 589286
rect 508448 589222 508500 589228
rect 573688 582486 573716 589290
rect 580116 586560 580168 586566
rect 580114 586528 580116 586537
rect 580168 586528 580170 586537
rect 580114 586463 580170 586472
rect 443956 582480 444008 582486
rect 443956 582422 444008 582428
rect 573676 582480 573728 582486
rect 573676 582422 573728 582428
rect 314052 582412 314104 582418
rect 314052 582354 314104 582360
rect 314144 582344 314196 582350
rect 314144 582286 314196 582292
rect 443864 582344 443916 582350
rect 443864 582286 443916 582292
rect 573584 582344 573636 582350
rect 573584 582286 573636 582292
rect 314156 579630 314184 582286
rect 378636 579692 378688 579698
rect 378636 579634 378688 579640
rect 314144 579624 314196 579630
rect 314144 579566 314196 579572
rect 313868 576904 313920 576910
rect 313868 576846 313920 576852
rect 313774 557560 313830 557569
rect 313774 557495 313830 557504
rect 313788 552634 313816 557495
rect 313776 552628 313828 552634
rect 313776 552570 313828 552576
rect 313776 538280 313828 538286
rect 313776 538222 313828 538228
rect 313788 528562 313816 538222
rect 313776 528556 313828 528562
rect 313776 528498 313828 528504
rect 313774 518936 313830 518945
rect 313774 518871 313830 518880
rect 313788 514010 313816 518871
rect 313776 514004 313828 514010
rect 313776 513946 313828 513952
rect 313776 499588 313828 499594
rect 313776 499530 313828 499536
rect 313788 489870 313816 499530
rect 313776 489864 313828 489870
rect 313776 489806 313828 489812
rect 313776 480276 313828 480282
rect 313776 480218 313828 480224
rect 313788 475386 313816 480218
rect 313776 475380 313828 475386
rect 313776 475322 313828 475328
rect 313880 462330 313908 576846
rect 378648 572642 378676 579634
rect 443876 572642 443904 582286
rect 508356 579692 508408 579698
rect 508356 579634 508408 579640
rect 378648 572614 378768 572642
rect 313960 570036 314012 570042
rect 313960 569978 314012 569984
rect 313972 565162 314000 569978
rect 378740 569906 378768 572614
rect 443692 572614 443904 572642
rect 508368 572642 508396 579634
rect 573596 572642 573624 582286
rect 508368 572614 508488 572642
rect 378728 569900 378780 569906
rect 378728 569842 378780 569848
rect 313972 565134 314184 565162
rect 314156 562986 314184 565134
rect 443692 563122 443720 572614
rect 508460 569906 508488 572614
rect 573412 572614 573624 572642
rect 508448 569900 508500 569906
rect 508448 569842 508500 569848
rect 573412 563122 573440 572614
rect 580114 570888 580170 570897
rect 580114 570823 580170 570832
rect 580128 569974 580156 570823
rect 580116 569968 580168 569974
rect 580116 569910 580168 569916
rect 314064 562958 314184 562986
rect 443600 563094 443720 563122
rect 573320 563094 573440 563122
rect 378912 562964 378964 562970
rect 313960 560448 314012 560454
rect 313960 560390 314012 560396
rect 313868 462324 313920 462330
rect 313868 462266 313920 462272
rect 312408 460006 312620 460034
rect 312592 459898 312620 460006
rect 312592 459870 312974 459898
rect 313972 459884 314000 560390
rect 314064 557569 314092 562958
rect 378912 562906 378964 562912
rect 378924 560289 378952 562906
rect 378726 560280 378782 560289
rect 378726 560215 378782 560224
rect 378910 560280 378966 560289
rect 443600 560266 443628 563094
rect 508632 562964 508684 562970
rect 508632 562906 508684 562912
rect 508644 560289 508672 562906
rect 378910 560215 378966 560224
rect 443508 560238 443628 560266
rect 508446 560280 508502 560289
rect 314050 557560 314106 557569
rect 314050 557495 314106 557504
rect 314052 552628 314104 552634
rect 314052 552570 314104 552576
rect 314064 538286 314092 552570
rect 378740 550662 378768 560215
rect 443508 553450 443536 560238
rect 508446 560215 508502 560224
rect 508630 560280 508686 560289
rect 573320 560266 573348 563094
rect 508630 560215 508686 560224
rect 573228 560238 573348 560266
rect 443496 553444 443548 553450
rect 443496 553386 443548 553392
rect 508460 550662 508488 560215
rect 573228 553450 573256 560238
rect 580114 555248 580170 555257
rect 580114 555183 580170 555192
rect 580128 554810 580156 555183
rect 580116 554804 580168 554810
rect 580116 554746 580168 554752
rect 573216 553444 573268 553450
rect 573216 553386 573268 553392
rect 378728 550656 378780 550662
rect 378728 550598 378780 550604
rect 379004 550656 379056 550662
rect 379004 550598 379056 550604
rect 443496 550656 443548 550662
rect 443496 550598 443548 550604
rect 508448 550656 508500 550662
rect 508448 550598 508500 550604
rect 508724 550656 508776 550662
rect 508724 550598 508776 550604
rect 573216 550656 573268 550662
rect 573216 550598 573268 550604
rect 379016 543862 379044 550598
rect 379004 543856 379056 543862
rect 379004 543798 379056 543804
rect 443508 543794 443536 550598
rect 508736 543862 508764 550598
rect 508724 543856 508776 543862
rect 508724 543798 508776 543804
rect 573228 543794 573256 550598
rect 315156 543788 315208 543794
rect 315156 543730 315208 543736
rect 443496 543788 443548 543794
rect 443496 543730 443548 543736
rect 573216 543788 573268 543794
rect 573216 543730 573268 543736
rect 314052 538280 314104 538286
rect 314052 538222 314104 538228
rect 314052 528556 314104 528562
rect 314052 528498 314104 528504
rect 314064 518945 314092 528498
rect 314050 518936 314106 518945
rect 314050 518871 314106 518880
rect 314052 514004 314104 514010
rect 314052 513946 314104 513952
rect 314064 499594 314092 513946
rect 314052 499588 314104 499594
rect 314052 499530 314104 499536
rect 314052 489864 314104 489870
rect 314052 489806 314104 489812
rect 314064 480282 314092 489806
rect 314052 480276 314104 480282
rect 314052 480218 314104 480224
rect 314052 475380 314104 475386
rect 314052 475322 314104 475328
rect 314064 463758 314092 475322
rect 314052 463752 314104 463758
rect 314052 463694 314104 463700
rect 314788 462324 314840 462330
rect 314788 462266 314840 462272
rect 314800 459898 314828 462266
rect 315168 460034 315196 543730
rect 378912 543720 378964 543726
rect 378912 543662 378964 543668
rect 508632 543720 508684 543726
rect 508632 543662 508684 543668
rect 378924 534138 378952 543662
rect 443588 543652 443640 543658
rect 443588 543594 443640 543600
rect 443600 540954 443628 543594
rect 443508 540926 443628 540954
rect 443508 534138 443536 540926
rect 508644 534138 508672 543662
rect 573308 543652 573360 543658
rect 573308 543594 573360 543600
rect 573320 540954 573348 543594
rect 573228 540926 573348 540954
rect 573228 534138 573256 540926
rect 580116 539776 580168 539782
rect 580116 539718 580168 539724
rect 580128 539617 580156 539718
rect 580114 539608 580170 539617
rect 580114 539543 580170 539552
rect 378912 534132 378964 534138
rect 378912 534074 378964 534080
rect 443496 534132 443548 534138
rect 443496 534074 443548 534080
rect 508632 534132 508684 534138
rect 508632 534074 508684 534080
rect 573216 534132 573268 534138
rect 573216 534074 573268 534080
rect 379004 533996 379056 534002
rect 379004 533938 379056 533944
rect 508724 533996 508776 534002
rect 508724 533938 508776 533944
rect 379016 529825 379044 533938
rect 443508 531350 443536 531381
rect 443496 531344 443548 531350
rect 443548 531292 443628 531298
rect 443496 531286 443628 531292
rect 443508 531282 443628 531286
rect 443508 531276 443640 531282
rect 443508 531270 443588 531276
rect 443588 531218 443640 531224
rect 508736 529825 508764 533938
rect 573228 531350 573256 531381
rect 573216 531344 573268 531350
rect 573268 531292 573348 531298
rect 573216 531286 573348 531292
rect 573228 531282 573348 531286
rect 573228 531276 573360 531282
rect 573228 531270 573308 531276
rect 573308 531218 573360 531224
rect 379002 529816 379058 529825
rect 379002 529751 379058 529760
rect 508722 529816 508778 529825
rect 508722 529751 508778 529760
rect 317916 527264 317968 527270
rect 317916 527206 317968 527212
rect 316536 510672 316588 510678
rect 316536 510614 316588 510620
rect 316548 460034 316576 510614
rect 315168 460006 315748 460034
rect 316548 460006 316852 460034
rect 315720 459898 315748 460006
rect 316824 459898 316852 460006
rect 317928 459898 317956 527206
rect 443588 524340 443640 524346
rect 443588 524282 443640 524288
rect 573308 524340 573360 524346
rect 573308 524282 573360 524288
rect 379186 520296 379242 520305
rect 379186 520231 379242 520240
rect 379200 514554 379228 520231
rect 443600 514706 443628 524282
rect 508906 520296 508962 520305
rect 508906 520231 508962 520240
rect 443600 514678 443720 514706
rect 379004 514548 379056 514554
rect 379004 514490 379056 514496
rect 379188 514548 379240 514554
rect 379188 514490 379240 514496
rect 379016 502382 379044 514490
rect 443692 512009 443720 514678
rect 508920 514554 508948 520231
rect 573320 514706 573348 524282
rect 580114 523968 580170 523977
rect 580114 523903 580170 523912
rect 580128 523054 580156 523903
rect 580116 523048 580168 523054
rect 580116 522990 580168 522996
rect 573320 514678 573440 514706
rect 508724 514548 508776 514554
rect 508724 514490 508776 514496
rect 508908 514548 508960 514554
rect 508908 514490 508960 514496
rect 443494 512000 443550 512009
rect 443494 511935 443550 511944
rect 443678 512000 443734 512009
rect 443678 511935 443734 511944
rect 443508 502382 443536 511935
rect 508736 502382 508764 514490
rect 573412 512009 573440 514678
rect 573214 512000 573270 512009
rect 573214 511935 573270 511944
rect 573398 512000 573454 512009
rect 573398 511935 573454 511944
rect 573228 502382 573256 511935
rect 580114 508328 580170 508337
rect 580114 508263 580170 508272
rect 580128 507890 580156 508263
rect 580116 507884 580168 507890
rect 580116 507826 580168 507832
rect 378820 502376 378872 502382
rect 378542 502344 378598 502353
rect 378542 502279 378598 502288
rect 378818 502344 378820 502353
rect 379004 502376 379056 502382
rect 378872 502344 378874 502353
rect 379004 502318 379056 502324
rect 443496 502376 443548 502382
rect 443496 502318 443548 502324
rect 443772 502376 443824 502382
rect 508540 502376 508592 502382
rect 443772 502318 443824 502324
rect 508262 502344 508318 502353
rect 378818 502279 378874 502288
rect 318008 494080 318060 494086
rect 318008 494022 318060 494028
rect 318020 460442 318048 494022
rect 378556 492697 378584 502279
rect 378542 492688 378598 492697
rect 378542 492623 378598 492632
rect 378726 492688 378782 492697
rect 378726 492623 378782 492632
rect 378740 489954 378768 492623
rect 378740 489926 378860 489954
rect 378832 480282 378860 489926
rect 443784 485926 443812 502318
rect 508262 502279 508318 502288
rect 508538 502344 508540 502353
rect 508724 502376 508776 502382
rect 508592 502344 508594 502353
rect 508724 502318 508776 502324
rect 573216 502376 573268 502382
rect 573216 502318 573268 502324
rect 573492 502376 573544 502382
rect 573492 502318 573544 502324
rect 508538 502279 508594 502288
rect 508276 492697 508304 502279
rect 508262 492688 508318 492697
rect 508262 492623 508318 492632
rect 508446 492688 508502 492697
rect 508446 492623 508502 492632
rect 508460 489954 508488 492623
rect 508460 489926 508580 489954
rect 443772 485920 443824 485926
rect 443772 485862 443824 485868
rect 443496 485716 443548 485722
rect 443496 485658 443548 485664
rect 378636 480276 378688 480282
rect 378636 480218 378688 480224
rect 378820 480276 378872 480282
rect 378820 480218 378872 480224
rect 378648 480162 378676 480218
rect 378648 480134 378768 480162
rect 320676 477556 320728 477562
rect 320676 477498 320728 477504
rect 318020 460414 318876 460442
rect 318848 459898 318876 460414
rect 320688 460034 320716 477498
rect 378740 470642 378768 480134
rect 443508 475946 443536 485658
rect 508552 480282 508580 489926
rect 573504 485926 573532 502318
rect 580116 492720 580168 492726
rect 580114 492688 580116 492697
rect 580168 492688 580170 492697
rect 580114 492623 580170 492632
rect 573492 485920 573544 485926
rect 573492 485862 573544 485868
rect 573216 485716 573268 485722
rect 573216 485658 573268 485664
rect 508356 480276 508408 480282
rect 508356 480218 508408 480224
rect 508540 480276 508592 480282
rect 508540 480218 508592 480224
rect 508368 480162 508396 480218
rect 508368 480134 508488 480162
rect 443508 475918 443628 475946
rect 443600 471986 443628 475918
rect 443588 471980 443640 471986
rect 443588 471922 443640 471928
rect 508460 470642 508488 480134
rect 573228 475946 573256 485658
rect 580114 477048 580170 477057
rect 580114 476983 580170 476992
rect 580128 476134 580156 476983
rect 580116 476128 580168 476134
rect 580116 476070 580168 476076
rect 573228 475918 573348 475946
rect 573320 471986 573348 475918
rect 573308 471980 573360 471986
rect 573308 471922 573360 471928
rect 378740 470614 378860 470642
rect 508460 470614 508580 470642
rect 359960 463684 360012 463690
rect 359960 463626 360012 463632
rect 355912 463616 355964 463622
rect 355912 463558 355964 463564
rect 354532 463344 354584 463350
rect 354532 463286 354584 463292
rect 330796 462800 330848 462806
rect 330796 462742 330848 462748
rect 328680 461576 328732 461582
rect 328680 461518 328732 461524
rect 324540 461508 324592 461514
rect 324540 461450 324592 461456
rect 322424 461032 322476 461038
rect 322424 460974 322476 460980
rect 320688 460006 321084 460034
rect 321056 459898 321084 460006
rect 314800 459870 315090 459898
rect 315720 459870 316102 459898
rect 316824 459870 317114 459898
rect 317928 459870 318218 459898
rect 318848 459870 319230 459898
rect 321056 459870 321346 459898
rect 322436 459884 322464 460974
rect 324552 459884 324580 461450
rect 325276 460080 325328 460086
rect 325276 460022 325328 460028
rect 325288 459898 325316 460022
rect 326380 460012 326432 460018
rect 326380 459954 326432 459960
rect 326392 459898 326420 459954
rect 325288 459870 325578 459898
rect 326392 459870 326590 459898
rect 328692 459884 328720 461518
rect 330808 459884 330836 462742
rect 333924 462732 333976 462738
rect 333924 462674 333976 462680
rect 332912 461100 332964 461106
rect 332912 461042 332964 461048
rect 332924 459884 332952 461042
rect 333936 459884 333964 462674
rect 337144 462664 337196 462670
rect 337144 462606 337196 462612
rect 335028 460352 335080 460358
rect 335028 460294 335080 460300
rect 335040 459884 335068 460294
rect 337156 459884 337184 462606
rect 339260 462596 339312 462602
rect 339260 462538 339312 462544
rect 339272 459884 339300 462538
rect 340272 462528 340324 462534
rect 340272 462470 340324 462476
rect 342386 462496 342442 462505
rect 340284 459884 340312 462470
rect 342386 462431 342442 462440
rect 342400 459884 342428 462431
rect 351680 461440 351732 461446
rect 351680 461382 351732 461388
rect 335856 459808 335908 459814
rect 294468 459734 295034 459762
rect 297688 459734 298254 459762
rect 298608 459734 299266 459762
rect 302932 459734 303498 459762
rect 311028 459734 311870 459762
rect 319952 459746 320334 459762
rect 335908 459756 336066 459762
rect 335856 459750 336066 459756
rect 319940 459740 320334 459746
rect 319992 459734 320334 459740
rect 335868 459734 336066 459750
rect 319940 459682 319992 459688
rect 234288 459672 234340 459678
rect 232170 459640 232226 459649
rect 229608 459598 230910 459626
rect 231922 459598 232170 459626
rect 228952 343596 229004 343602
rect 228952 343538 229004 343544
rect 229504 325100 229556 325106
rect 229504 325042 229556 325048
rect 228860 244180 228912 244186
rect 228860 244122 228912 244128
rect 227480 143540 227532 143546
rect 227480 143482 227532 143488
rect 225364 135380 225416 135386
rect 225364 135322 225416 135328
rect 225376 57934 225404 135322
rect 225180 57928 225232 57934
rect 225180 57870 225232 57876
rect 225364 57928 225416 57934
rect 225364 57870 225416 57876
rect 225192 48385 225220 57870
rect 225178 48376 225234 48385
rect 225178 48311 225234 48320
rect 225362 48376 225418 48385
rect 225362 48311 225418 48320
rect 225376 46918 225404 48311
rect 225364 46912 225416 46918
rect 225364 46854 225416 46860
rect 225456 37324 225508 37330
rect 225456 37266 225508 37272
rect 225468 29050 225496 37266
rect 225376 29022 225496 29050
rect 225376 27606 225404 29022
rect 225364 27600 225416 27606
rect 225364 27542 225416 27548
rect 225088 18080 225140 18086
rect 225088 18022 225140 18028
rect 225100 9761 225128 18022
rect 225454 10704 225510 10713
rect 225454 10639 225510 10648
rect 225468 10198 225496 10639
rect 225638 10432 225694 10441
rect 225638 10367 225694 10376
rect 225652 10266 225680 10367
rect 225640 10260 225692 10266
rect 225640 10202 225692 10208
rect 225456 10192 225508 10198
rect 225456 10134 225508 10140
rect 225640 10124 225692 10130
rect 225640 10066 225692 10072
rect 225652 10033 225680 10066
rect 225638 10024 225694 10033
rect 225638 9959 225694 9968
rect 225086 9752 225142 9761
rect 225086 9687 225142 9696
rect 225270 9752 225326 9761
rect 225270 9687 225326 9696
rect 222512 8424 222564 8430
rect 222512 8366 222564 8372
rect 222524 626 222552 8366
rect 225284 7993 225312 9687
rect 229410 8936 229466 8945
rect 229410 8871 229466 8880
rect 225822 8800 225878 8809
rect 225822 8735 225878 8744
rect 224626 7984 224682 7993
rect 224626 7919 224682 7928
rect 225270 7984 225326 7993
rect 225270 7919 225326 7928
rect 225454 7984 225510 7993
rect 225454 7919 225510 7928
rect 224536 3664 224588 3670
rect 224536 3606 224588 3612
rect 224548 3233 224576 3606
rect 224534 3224 224590 3233
rect 224534 3159 224590 3168
rect 223432 2644 223484 2650
rect 223432 2586 223484 2592
rect 221040 604 221092 610
rect 221040 546 221092 552
rect 221224 604 221276 610
rect 221224 546 221276 552
rect 222248 598 222552 626
rect 221052 480 221080 546
rect 222248 480 222276 598
rect 223444 480 223472 2586
rect 224640 480 224668 7919
rect 225468 7886 225496 7919
rect 225272 7880 225324 7886
rect 225272 7822 225324 7828
rect 225364 7880 225416 7886
rect 225364 7822 225416 7828
rect 225456 7880 225508 7886
rect 225456 7822 225508 7828
rect 225548 7880 225600 7886
rect 225548 7822 225600 7828
rect 225284 7721 225312 7822
rect 225270 7712 225326 7721
rect 225270 7647 225326 7656
rect 225376 7585 225404 7822
rect 225560 7721 225588 7822
rect 225546 7712 225602 7721
rect 225546 7647 225602 7656
rect 225362 7576 225418 7585
rect 225362 7511 225418 7520
rect 225454 6488 225510 6497
rect 225454 6423 225510 6432
rect 225178 6352 225234 6361
rect 225178 6287 225234 6296
rect 225192 6254 225220 6287
rect 225180 6248 225232 6254
rect 225180 6190 225232 6196
rect 225272 6248 225324 6254
rect 225272 6190 225324 6196
rect 225284 5817 225312 6190
rect 225468 5953 225496 6423
rect 225454 5944 225510 5953
rect 225454 5879 225510 5888
rect 225270 5808 225326 5817
rect 225270 5743 225326 5752
rect 225270 5264 225326 5273
rect 225270 5199 225326 5208
rect 225284 4826 225312 5199
rect 225272 4820 225324 4826
rect 225272 4762 225324 4768
rect 225364 4820 225416 4826
rect 225364 4762 225416 4768
rect 225270 4720 225326 4729
rect 225376 4706 225404 4762
rect 225326 4678 225404 4706
rect 225270 4655 225326 4664
rect 225454 4312 225510 4321
rect 225454 4247 225510 4256
rect 225468 3670 225496 4247
rect 225180 3664 225232 3670
rect 225180 3606 225232 3612
rect 225456 3664 225508 3670
rect 225456 3606 225508 3612
rect 225192 3097 225220 3606
rect 225640 3596 225692 3602
rect 225640 3538 225692 3544
rect 225652 3233 225680 3538
rect 225638 3224 225694 3233
rect 225638 3159 225694 3168
rect 225178 3088 225234 3097
rect 225178 3023 225234 3032
rect 225836 480 225864 8735
rect 226926 5264 226982 5273
rect 226926 5199 226982 5208
rect 226940 5166 226968 5199
rect 226928 5160 226980 5166
rect 226928 5102 226980 5108
rect 227020 5160 227072 5166
rect 227020 5102 227072 5108
rect 227032 480 227060 5102
rect 228124 4072 228176 4078
rect 228124 4014 228176 4020
rect 228216 4072 228268 4078
rect 228216 4014 228268 4020
rect 228136 3641 228164 4014
rect 228122 3632 228178 3641
rect 228122 3567 228178 3576
rect 228228 480 228256 4014
rect 229424 480 229452 8871
rect 229516 4078 229544 325042
rect 229608 7177 229636 459598
rect 233182 459640 233238 459649
rect 232934 459598 233182 459626
rect 232170 459575 232226 459584
rect 234038 459620 234288 459626
rect 250112 459672 250164 459678
rect 236218 459640 236274 459649
rect 234038 459614 234340 459620
rect 234038 459598 234328 459614
rect 236154 459598 236218 459626
rect 233182 459575 233238 459584
rect 237414 459640 237470 459649
rect 237166 459598 237414 459626
rect 236218 459575 236274 459584
rect 238518 459640 238574 459649
rect 238270 459598 238518 459626
rect 237414 459575 237470 459584
rect 239622 459640 239678 459649
rect 239282 459598 239622 459626
rect 238518 459575 238574 459584
rect 241646 459640 241702 459649
rect 241398 459598 241646 459626
rect 239622 459575 239678 459584
rect 242750 459640 242806 459649
rect 242410 459598 242750 459626
rect 241646 459575 241702 459584
rect 244590 459640 244646 459649
rect 244526 459598 244590 459626
rect 242750 459575 242806 459584
rect 245878 459640 245934 459649
rect 245630 459598 245878 459626
rect 244590 459575 244646 459584
rect 246982 459640 247038 459649
rect 246642 459598 246982 459626
rect 245878 459575 245934 459584
rect 248822 459640 248878 459649
rect 248758 459598 248822 459626
rect 246982 459575 247038 459584
rect 249770 459620 250112 459626
rect 256368 459672 256420 459678
rect 251214 459640 251270 459649
rect 249770 459614 250164 459620
rect 249770 459598 250152 459614
rect 250874 459598 251214 459626
rect 248822 459575 248878 459584
rect 252134 459640 252190 459649
rect 251886 459598 252134 459626
rect 251214 459575 251270 459584
rect 256118 459620 256368 459626
rect 323528 459672 323580 459678
rect 256118 459614 256420 459620
rect 323462 459620 323528 459626
rect 323462 459614 323580 459620
rect 327484 459672 327536 459678
rect 329508 459672 329560 459678
rect 327536 459620 327694 459626
rect 327484 459614 327694 459620
rect 331716 459672 331768 459678
rect 329560 459620 329810 459626
rect 329508 459614 329810 459620
rect 337788 459672 337840 459678
rect 331768 459620 331926 459626
rect 331716 459614 331926 459620
rect 341192 459672 341244 459678
rect 337840 459620 338182 459626
rect 337788 459614 338182 459620
rect 345608 459672 345660 459678
rect 343122 459640 343178 459649
rect 341244 459620 341402 459626
rect 341192 459614 341402 459620
rect 256118 459598 256408 459614
rect 323462 459598 323568 459614
rect 327496 459598 327694 459614
rect 329520 459598 329810 459614
rect 331728 459598 331926 459614
rect 337800 459598 338182 459614
rect 341204 459598 341402 459614
rect 252134 459575 252190 459584
rect 344226 459640 344282 459649
rect 343178 459598 343426 459626
rect 343122 459575 343178 459584
rect 344282 459598 344530 459626
rect 345542 459620 345608 459626
rect 345542 459614 345660 459620
rect 346250 459640 346306 459649
rect 345542 459598 345648 459614
rect 344226 459575 344282 459584
rect 347354 459640 347410 459649
rect 346306 459598 346646 459626
rect 346250 459575 346306 459584
rect 348458 459640 348514 459649
rect 347410 459598 347658 459626
rect 347354 459575 347410 459584
rect 348514 459598 348762 459626
rect 349774 459598 350064 459626
rect 348458 459575 348514 459584
rect 273400 340190 273598 340218
rect 319676 340190 319874 340218
rect 229700 340054 230542 340082
rect 229594 7168 229650 7177
rect 229594 7103 229650 7112
rect 229700 5030 229728 340054
rect 230056 337680 230108 337686
rect 230056 337622 230108 337628
rect 230068 337482 230096 337622
rect 230056 337476 230108 337482
rect 230056 337418 230108 337424
rect 230712 335578 230740 340068
rect 231002 340054 231108 340082
rect 231186 340054 231292 340082
rect 231080 335782 231108 340054
rect 231068 335776 231120 335782
rect 231068 335718 231120 335724
rect 229964 335572 230016 335578
rect 229964 335514 230016 335520
rect 230700 335572 230752 335578
rect 230700 335514 230752 335520
rect 229976 328438 230004 335514
rect 231068 335504 231120 335510
rect 231068 335446 231120 335452
rect 229964 328432 230016 328438
rect 229964 328374 230016 328380
rect 229872 321428 229924 321434
rect 229872 321370 229924 321376
rect 229884 311930 229912 321370
rect 229884 311902 230004 311930
rect 229976 307766 230004 311902
rect 229872 307760 229924 307766
rect 229872 307702 229924 307708
rect 229964 307760 230016 307766
rect 229964 307702 230016 307708
rect 229884 298042 229912 307702
rect 229872 298036 229924 298042
rect 229872 297978 229924 297984
rect 230240 298036 230292 298042
rect 230240 297978 230292 297984
rect 230252 296698 230280 297978
rect 230160 296670 230280 296698
rect 230160 287094 230188 296670
rect 229964 287088 230016 287094
rect 229964 287030 230016 287036
rect 230148 287088 230200 287094
rect 230148 287030 230200 287036
rect 229976 278798 230004 287030
rect 229964 278792 230016 278798
rect 229964 278734 230016 278740
rect 230056 278792 230108 278798
rect 230056 278734 230108 278740
rect 230068 273306 230096 278734
rect 229884 273278 230096 273306
rect 229884 269142 229912 273278
rect 229780 269136 229832 269142
rect 229780 269078 229832 269084
rect 229872 269136 229924 269142
rect 229872 269078 229924 269084
rect 229792 265690 229820 269078
rect 229792 265662 229912 265690
rect 229884 253994 229912 265662
rect 229884 253966 230004 253994
rect 229976 251190 230004 253966
rect 229964 251184 230016 251190
rect 229964 251126 230016 251132
rect 229964 244180 230016 244186
rect 229964 244122 230016 244128
rect 229976 225010 230004 244122
rect 229780 225004 229832 225010
rect 229780 224946 229832 224952
rect 229964 225004 230016 225010
rect 229964 224946 230016 224952
rect 229792 224890 229820 224946
rect 229792 224862 229912 224890
rect 229884 215370 229912 224862
rect 229884 215342 230004 215370
rect 229976 212514 230004 215342
rect 229976 212486 230096 212514
rect 230068 205834 230096 212486
rect 230056 205828 230108 205834
rect 230056 205770 230108 205776
rect 229964 205556 230016 205562
rect 229964 205498 230016 205504
rect 229976 186386 230004 205498
rect 229780 186380 229832 186386
rect 229780 186322 229832 186328
rect 229964 186380 230016 186386
rect 229964 186322 230016 186328
rect 229792 186266 229820 186322
rect 229792 186238 229912 186266
rect 229884 182170 229912 186238
rect 229872 182164 229924 182170
rect 229872 182106 229924 182112
rect 229872 176588 229924 176594
rect 229872 176530 229924 176536
rect 229884 166954 229912 176530
rect 229884 166926 230004 166954
rect 229976 164234 230004 166926
rect 229976 164206 230096 164234
rect 230068 162858 230096 164206
rect 230056 162852 230108 162858
rect 230056 162794 230108 162800
rect 230056 157140 230108 157146
rect 230056 157082 230108 157088
rect 230068 144922 230096 157082
rect 229884 144894 230096 144922
rect 229884 138038 229912 144894
rect 229872 138032 229924 138038
rect 229872 137974 229924 137980
rect 229780 137964 229832 137970
rect 229780 137906 229832 137912
rect 229792 135289 229820 137906
rect 229778 135280 229834 135289
rect 229778 135215 229834 135224
rect 229962 135280 230018 135289
rect 229962 135215 230018 135224
rect 229976 128330 230004 135215
rect 229884 128302 230004 128330
rect 229884 118794 229912 128302
rect 229872 118788 229924 118794
rect 229872 118730 229924 118736
rect 229780 114708 229832 114714
rect 229780 114650 229832 114656
rect 229792 109070 229820 114650
rect 229780 109064 229832 109070
rect 229780 109006 229832 109012
rect 229872 108996 229924 109002
rect 229872 108938 229924 108944
rect 229884 103494 229912 108938
rect 229872 103488 229924 103494
rect 229872 103430 229924 103436
rect 230056 85604 230108 85610
rect 230056 85546 230108 85552
rect 230068 80170 230096 85546
rect 230056 80164 230108 80170
rect 230056 80106 230108 80112
rect 229964 79892 230016 79898
rect 229964 79834 230016 79840
rect 229976 66298 230004 79834
rect 229872 66292 229924 66298
rect 229872 66234 229924 66240
rect 229964 66292 230016 66298
rect 229964 66234 230016 66240
rect 229884 60858 229912 66234
rect 229872 60852 229924 60858
rect 229872 60794 229924 60800
rect 229780 60716 229832 60722
rect 229780 60658 229832 60664
rect 229792 53122 229820 60658
rect 229792 53094 229912 53122
rect 229884 41426 229912 53094
rect 229884 41398 230004 41426
rect 229976 31822 230004 41398
rect 229964 31816 230016 31822
rect 229964 31758 230016 31764
rect 229964 31680 230016 31686
rect 229964 31622 230016 31628
rect 229976 24206 230004 31622
rect 229964 24200 230016 24206
rect 229964 24142 230016 24148
rect 230148 24200 230200 24206
rect 230148 24142 230200 24148
rect 230160 5030 230188 24142
rect 231080 5273 231108 335446
rect 231264 7886 231292 340054
rect 231448 337385 231476 340068
rect 231540 340054 231738 340082
rect 231816 340054 231922 340082
rect 232000 340054 232198 340082
rect 232368 340054 232474 340082
rect 231434 337376 231490 337385
rect 231434 337311 231490 337320
rect 231344 335572 231396 335578
rect 231344 335514 231396 335520
rect 231356 8974 231384 335514
rect 231344 8968 231396 8974
rect 231344 8910 231396 8916
rect 231252 7880 231304 7886
rect 231344 7880 231396 7886
rect 231252 7822 231304 7828
rect 231342 7848 231344 7857
rect 231396 7848 231398 7857
rect 231342 7783 231398 7792
rect 231540 6089 231568 340054
rect 231620 335776 231672 335782
rect 231620 335718 231672 335724
rect 231526 6080 231582 6089
rect 231526 6015 231582 6024
rect 231632 5409 231660 335718
rect 231816 335510 231844 340054
rect 232000 335578 232028 340054
rect 232368 338162 232396 340054
rect 232356 338156 232408 338162
rect 232356 338098 232408 338104
rect 232644 337754 232672 340068
rect 232736 340054 232934 340082
rect 233104 340054 233210 340082
rect 233288 340054 233394 340082
rect 233472 340054 233670 340082
rect 233946 340054 234052 340082
rect 232632 337748 232684 337754
rect 232632 337690 232684 337696
rect 232736 335594 232764 340054
rect 232814 337784 232870 337793
rect 232814 337719 232816 337728
rect 232868 337719 232870 337728
rect 232816 337690 232868 337696
rect 231988 335572 232040 335578
rect 231988 335514 232040 335520
rect 232552 335566 232764 335594
rect 233000 335572 233052 335578
rect 231804 335504 231856 335510
rect 231804 335446 231856 335452
rect 232172 17264 232224 17270
rect 232172 17206 232224 17212
rect 232184 9761 232212 17206
rect 232448 10260 232500 10266
rect 232448 10202 232500 10208
rect 232460 10033 232488 10202
rect 232446 10024 232502 10033
rect 232446 9959 232502 9968
rect 231894 9752 231950 9761
rect 231894 9687 231950 9696
rect 232170 9752 232226 9761
rect 232170 9687 232226 9696
rect 231618 5400 231674 5409
rect 231618 5335 231674 5344
rect 231066 5264 231122 5273
rect 231066 5199 231122 5208
rect 229688 5024 229740 5030
rect 229688 4966 229740 4972
rect 230148 5024 230200 5030
rect 230148 4966 230200 4972
rect 230608 5024 230660 5030
rect 230608 4966 230660 4972
rect 231908 4978 231936 9687
rect 232552 7886 232580 335566
rect 233000 335514 233052 335520
rect 232724 335504 232776 335510
rect 232724 335446 232776 335452
rect 232540 7880 232592 7886
rect 232540 7822 232592 7828
rect 232446 7440 232502 7449
rect 232446 7375 232502 7384
rect 232354 7168 232410 7177
rect 232354 7103 232410 7112
rect 232368 7018 232396 7103
rect 232460 7018 232488 7375
rect 232368 6990 232488 7018
rect 230146 4176 230202 4185
rect 230146 4111 230202 4120
rect 230160 4078 230188 4111
rect 229504 4072 229556 4078
rect 229504 4014 229556 4020
rect 230148 4072 230200 4078
rect 230148 4014 230200 4020
rect 230424 3732 230476 3738
rect 230424 3674 230476 3680
rect 230436 3641 230464 3674
rect 230422 3632 230478 3641
rect 230422 3567 230478 3576
rect 230620 480 230648 4966
rect 231908 4950 232028 4978
rect 232000 610 232028 4950
rect 232736 3369 232764 335446
rect 233012 9058 233040 335514
rect 233104 312594 233132 340054
rect 233288 335510 233316 340054
rect 233472 335578 233500 340054
rect 233460 335572 233512 335578
rect 233460 335514 233512 335520
rect 233828 335572 233880 335578
rect 233828 335514 233880 335520
rect 233276 335504 233328 335510
rect 233276 335446 233328 335452
rect 233092 312588 233144 312594
rect 233092 312530 233144 312536
rect 232920 9030 233040 9058
rect 233840 9042 233868 335514
rect 233828 9036 233880 9042
rect 232920 3505 232948 9030
rect 233828 8978 233880 8984
rect 233000 8968 233052 8974
rect 233000 8910 233052 8916
rect 232906 3496 232962 3505
rect 232906 3431 232962 3440
rect 232722 3360 232778 3369
rect 232722 3295 232778 3304
rect 231804 604 231856 610
rect 231804 546 231856 552
rect 231988 604 232040 610
rect 231988 546 232040 552
rect 231816 480 231844 546
rect 233012 480 233040 8910
rect 234024 7993 234052 340054
rect 234116 273970 234144 340068
rect 234208 340054 234406 340082
rect 234208 338230 234236 340054
rect 234196 338224 234248 338230
rect 234196 338166 234248 338172
rect 234668 337754 234696 340068
rect 234760 340054 234866 340082
rect 234656 337748 234708 337754
rect 234656 337690 234708 337696
rect 234760 335578 234788 340054
rect 234748 335572 234800 335578
rect 234748 335514 234800 335520
rect 235128 330546 235156 340068
rect 235208 335776 235260 335782
rect 235208 335718 235260 335724
rect 235116 330540 235168 330546
rect 235116 330482 235168 330488
rect 234104 273964 234156 273970
rect 234104 273906 234156 273912
rect 234932 11076 234984 11082
rect 234932 11018 234984 11024
rect 234944 10962 234972 11018
rect 234852 10934 234972 10962
rect 234656 10804 234708 10810
rect 234656 10746 234708 10752
rect 234668 10577 234696 10746
rect 234852 10742 234880 10934
rect 235024 10804 235076 10810
rect 235220 10792 235248 335718
rect 235300 335572 235352 335578
rect 235300 335514 235352 335520
rect 235312 11286 235340 335514
rect 235404 335458 235432 340068
rect 235496 340054 235602 340082
rect 235680 340054 235878 340082
rect 236048 340054 236154 340082
rect 235496 335782 235524 340054
rect 235484 335776 235536 335782
rect 235484 335718 235536 335724
rect 235680 335578 235708 340054
rect 236048 335594 236076 340054
rect 236324 338026 236352 340068
rect 236312 338020 236364 338026
rect 236312 337962 236364 337968
rect 235668 335572 235720 335578
rect 235668 335514 235720 335520
rect 235772 335566 236076 335594
rect 235404 335430 235616 335458
rect 235588 328438 235616 335430
rect 235576 328432 235628 328438
rect 235576 328374 235628 328380
rect 235772 321978 235800 335566
rect 235760 321972 235812 321978
rect 235760 321914 235812 321920
rect 235484 318912 235536 318918
rect 235484 318854 235536 318860
rect 235668 318912 235720 318918
rect 235668 318854 235720 318860
rect 235496 318714 235524 318854
rect 235680 318714 235708 318854
rect 235484 318708 235536 318714
rect 235484 318650 235536 318656
rect 235668 318708 235720 318714
rect 235668 318650 235720 318656
rect 235944 318708 235996 318714
rect 235944 318650 235996 318656
rect 235576 311840 235628 311846
rect 235576 311782 235628 311788
rect 235588 289882 235616 311782
rect 235956 309210 235984 318650
rect 235772 309182 235984 309210
rect 235772 302326 235800 309182
rect 235760 302320 235812 302326
rect 235760 302262 235812 302268
rect 235668 302184 235720 302190
rect 235668 302126 235720 302132
rect 235680 299470 235708 302126
rect 235668 299464 235720 299470
rect 235668 299406 235720 299412
rect 235484 289876 235536 289882
rect 235484 289818 235536 289824
rect 235576 289876 235628 289882
rect 235576 289818 235628 289824
rect 235496 285326 235524 289818
rect 235484 285320 235536 285326
rect 235484 285262 235536 285268
rect 235576 282804 235628 282810
rect 235576 282746 235628 282752
rect 235588 278769 235616 282746
rect 235390 278760 235446 278769
rect 235390 278695 235446 278704
rect 235574 278760 235630 278769
rect 235574 278695 235630 278704
rect 235404 269142 235432 278695
rect 235392 269136 235444 269142
rect 235392 269078 235444 269084
rect 235576 269136 235628 269142
rect 235576 269078 235628 269084
rect 235588 263702 235616 269078
rect 235576 263696 235628 263702
rect 235576 263638 235628 263644
rect 235576 263492 235628 263498
rect 235576 263434 235628 263440
rect 235588 260846 235616 263434
rect 235576 260840 235628 260846
rect 235576 260782 235628 260788
rect 235576 253836 235628 253842
rect 235576 253778 235628 253784
rect 235588 244361 235616 253778
rect 235574 244352 235630 244361
rect 235574 244287 235630 244296
rect 235482 241632 235538 241641
rect 235482 241567 235538 241576
rect 235496 240106 235524 241567
rect 235484 240100 235536 240106
rect 235484 240042 235536 240048
rect 235668 230512 235720 230518
rect 235668 230454 235720 230460
rect 235680 221105 235708 230454
rect 235666 221096 235722 221105
rect 235666 221031 235722 221040
rect 235574 220960 235630 220969
rect 235574 220895 235630 220904
rect 235588 220833 235616 220895
rect 235390 220824 235446 220833
rect 235390 220759 235446 220768
rect 235574 220824 235630 220833
rect 235574 220759 235630 220768
rect 235404 211206 235432 220759
rect 235392 211200 235444 211206
rect 235392 211142 235444 211148
rect 235484 211200 235536 211206
rect 235484 211142 235536 211148
rect 235496 205766 235524 211142
rect 235484 205760 235536 205766
rect 235484 205702 235536 205708
rect 235484 203040 235536 203046
rect 235484 202982 235536 202988
rect 235496 202858 235524 202982
rect 235496 202842 235616 202858
rect 235496 202836 235628 202842
rect 235496 202830 235576 202836
rect 235576 202778 235628 202784
rect 235576 195764 235628 195770
rect 235576 195706 235628 195712
rect 235588 191826 235616 195706
rect 235576 191820 235628 191826
rect 235576 191762 235628 191768
rect 235760 191820 235812 191826
rect 235760 191762 235812 191768
rect 235772 182209 235800 191762
rect 235574 182200 235630 182209
rect 235496 182158 235574 182186
rect 235496 176730 235524 182158
rect 235574 182135 235630 182144
rect 235758 182200 235814 182209
rect 235758 182135 235814 182144
rect 235484 176724 235536 176730
rect 235484 176666 235536 176672
rect 235576 176588 235628 176594
rect 235576 176530 235628 176536
rect 235588 167210 235616 176530
rect 235576 167204 235628 167210
rect 235576 167146 235628 167152
rect 235484 166932 235536 166938
rect 235484 166874 235536 166880
rect 235496 159322 235524 166874
rect 235484 159316 235536 159322
rect 235484 159258 235536 159264
rect 235576 157140 235628 157146
rect 235576 157082 235628 157088
rect 235588 154465 235616 157082
rect 235574 154456 235630 154465
rect 235574 154391 235630 154400
rect 235850 154456 235906 154465
rect 235850 154391 235906 154400
rect 235864 144945 235892 154391
rect 235482 144936 235538 144945
rect 235482 144871 235538 144880
rect 235850 144936 235906 144945
rect 235850 144871 235906 144880
rect 235496 138038 235524 144871
rect 235484 138032 235536 138038
rect 235484 137974 235536 137980
rect 235576 137964 235628 137970
rect 235576 137906 235628 137912
rect 235588 135250 235616 137906
rect 235576 135244 235628 135250
rect 235576 135186 235628 135192
rect 235760 135244 235812 135250
rect 235760 135186 235812 135192
rect 235772 125633 235800 135186
rect 235574 125624 235630 125633
rect 235496 125582 235574 125610
rect 235496 118538 235524 125582
rect 235574 125559 235630 125568
rect 235758 125624 235814 125633
rect 235758 125559 235814 125568
rect 235496 118510 235616 118538
rect 235588 115802 235616 118510
rect 235576 115796 235628 115802
rect 235576 115738 235628 115744
rect 235576 108996 235628 109002
rect 235576 108938 235628 108944
rect 235588 106298 235616 108938
rect 235496 106282 235616 106298
rect 235484 106276 235616 106282
rect 235536 106270 235616 106276
rect 235484 106218 235536 106224
rect 235484 96688 235536 96694
rect 235536 96636 235616 96642
rect 235484 96630 235616 96636
rect 235496 96626 235616 96630
rect 235496 96620 235628 96626
rect 235496 96614 235576 96620
rect 235576 96562 235628 96568
rect 235588 96531 235616 96562
rect 235576 89684 235628 89690
rect 235576 89626 235628 89632
rect 235588 86986 235616 89626
rect 235496 86958 235616 86986
rect 235496 79914 235524 86958
rect 235496 79886 235616 79914
rect 235588 77178 235616 79886
rect 235576 77172 235628 77178
rect 235576 77114 235628 77120
rect 235484 67652 235536 67658
rect 235484 67594 235536 67600
rect 235496 60790 235524 67594
rect 235484 60784 235536 60790
rect 235484 60726 235536 60732
rect 235576 60648 235628 60654
rect 235576 60590 235628 60596
rect 235588 57934 235616 60590
rect 235576 57928 235628 57934
rect 235576 57870 235628 57876
rect 235392 48340 235444 48346
rect 235392 48282 235444 48288
rect 235404 48249 235432 48282
rect 235390 48240 235446 48249
rect 235390 48175 235446 48184
rect 235666 48104 235722 48113
rect 235666 48039 235722 48048
rect 235680 38706 235708 48039
rect 235588 38678 235708 38706
rect 235588 38570 235616 38678
rect 235496 38542 235616 38570
rect 235496 31822 235524 38542
rect 235484 31816 235536 31822
rect 235484 31758 235536 31764
rect 235484 29028 235536 29034
rect 235484 28970 235536 28976
rect 235496 22166 235524 28970
rect 235484 22160 235536 22166
rect 235484 22102 235536 22108
rect 235576 22024 235628 22030
rect 235576 21966 235628 21972
rect 235300 11280 235352 11286
rect 235300 11222 235352 11228
rect 235220 10764 235340 10792
rect 235024 10746 235076 10752
rect 234840 10736 234892 10742
rect 235036 10713 235064 10746
rect 234840 10678 234892 10684
rect 235022 10704 235078 10713
rect 235022 10639 235078 10648
rect 234654 10568 234710 10577
rect 234654 10503 234710 10512
rect 235022 10160 235078 10169
rect 235022 10095 235024 10104
rect 235076 10095 235078 10104
rect 235024 10066 235076 10072
rect 234932 9036 234984 9042
rect 234932 8978 234984 8984
rect 234944 8945 234972 8978
rect 235024 8968 235076 8974
rect 234930 8936 234986 8945
rect 235024 8910 235076 8916
rect 234930 8871 234986 8880
rect 235036 8809 235064 8910
rect 235022 8800 235078 8809
rect 235022 8735 235078 8744
rect 234010 7984 234066 7993
rect 234010 7919 234066 7928
rect 235114 6624 235170 6633
rect 235114 6559 235170 6568
rect 235128 6322 235156 6559
rect 235116 6316 235168 6322
rect 235116 6258 235168 6264
rect 235312 4298 235340 10764
rect 235392 10668 235444 10674
rect 235392 10610 235444 10616
rect 235404 10577 235432 10610
rect 235390 10568 235446 10577
rect 235390 10503 235446 10512
rect 235220 4270 235340 4298
rect 234930 4176 234986 4185
rect 234930 4111 234986 4120
rect 235114 4176 235170 4185
rect 235114 4111 235116 4120
rect 234944 3670 234972 4111
rect 235168 4111 235170 4120
rect 235116 4082 235168 4088
rect 235220 3913 235248 4270
rect 235300 4140 235352 4146
rect 235300 4082 235352 4088
rect 235206 3904 235262 3913
rect 235206 3839 235262 3848
rect 235208 3732 235260 3738
rect 235208 3674 235260 3680
rect 234840 3664 234892 3670
rect 234840 3606 234892 3612
rect 234932 3664 234984 3670
rect 235220 3641 235248 3674
rect 234932 3606 234984 3612
rect 235206 3632 235262 3641
rect 234748 3596 234800 3602
rect 234748 3538 234800 3544
rect 234760 3233 234788 3538
rect 234852 3369 234880 3606
rect 235206 3567 235262 3576
rect 235114 3496 235170 3505
rect 235114 3431 235170 3440
rect 235128 3398 235156 3431
rect 235116 3392 235168 3398
rect 234838 3360 234894 3369
rect 235116 3334 235168 3340
rect 235208 3392 235260 3398
rect 235208 3334 235260 3340
rect 234838 3295 234894 3304
rect 235220 3233 235248 3334
rect 234746 3224 234802 3233
rect 234746 3159 234802 3168
rect 235206 3224 235262 3233
rect 235206 3159 235262 3168
rect 234196 604 234248 610
rect 234196 546 234248 552
rect 234208 480 234236 546
rect 235312 480 235340 4082
rect 235588 3777 235616 21966
rect 236404 18624 236456 18630
rect 236404 18566 236456 18572
rect 235666 4312 235722 4321
rect 235666 4247 235722 4256
rect 235680 4078 235708 4247
rect 236416 4146 236444 18566
rect 236600 10305 236628 340068
rect 236890 340054 236996 340082
rect 236772 335572 236824 335578
rect 236772 335514 236824 335520
rect 236680 333600 236732 333606
rect 236680 333542 236732 333548
rect 236586 10296 236642 10305
rect 236586 10231 236642 10240
rect 236404 4140 236456 4146
rect 236404 4082 236456 4088
rect 236496 4140 236548 4146
rect 236496 4082 236548 4088
rect 235668 4072 235720 4078
rect 235668 4014 235720 4020
rect 235574 3768 235630 3777
rect 235574 3703 235630 3712
rect 235392 3596 235444 3602
rect 235392 3538 235444 3544
rect 235404 3369 235432 3538
rect 235390 3360 235446 3369
rect 235390 3295 235446 3304
rect 236508 480 236536 4082
rect 236692 3534 236720 333542
rect 236784 11014 236812 335514
rect 236772 11008 236824 11014
rect 236772 10950 236824 10956
rect 236968 4049 236996 340054
rect 236954 4040 237010 4049
rect 236954 3975 237010 3984
rect 236770 3632 236826 3641
rect 236770 3567 236826 3576
rect 236784 3534 236812 3567
rect 236680 3528 236732 3534
rect 236680 3470 236732 3476
rect 236772 3528 236824 3534
rect 236772 3470 236824 3476
rect 237060 3398 237088 340068
rect 237152 340054 237350 340082
rect 237428 340054 237626 340082
rect 237152 335578 237180 340054
rect 237140 335572 237192 335578
rect 237140 335514 237192 335520
rect 237428 333606 237456 340054
rect 237796 337958 237824 340068
rect 238086 340054 238284 340082
rect 237784 337952 237836 337958
rect 237784 337894 237836 337900
rect 237968 335776 238020 335782
rect 237968 335718 238020 335724
rect 237876 335504 237928 335510
rect 237876 335446 237928 335452
rect 237416 333600 237468 333606
rect 237416 333542 237468 333548
rect 237782 9208 237838 9217
rect 237782 9143 237838 9152
rect 237690 5264 237746 5273
rect 237690 5199 237746 5208
rect 237138 3496 237194 3505
rect 237138 3431 237194 3440
rect 237152 3398 237180 3431
rect 237048 3392 237100 3398
rect 237048 3334 237100 3340
rect 237140 3392 237192 3398
rect 237140 3334 237192 3340
rect 237704 480 237732 5199
rect 237796 4146 237824 9143
rect 237888 7886 237916 335446
rect 237876 7880 237928 7886
rect 237876 7822 237928 7828
rect 237784 4140 237836 4146
rect 237784 4082 237836 4088
rect 237980 4078 238008 335718
rect 238152 335572 238204 335578
rect 238152 335514 238204 335520
rect 238164 10810 238192 335514
rect 238152 10804 238204 10810
rect 238152 10746 238204 10752
rect 238256 10674 238284 340054
rect 238348 10792 238376 340068
rect 238440 340054 238546 340082
rect 238624 340054 238822 340082
rect 238900 340054 239098 340082
rect 238440 335782 238468 340054
rect 238428 335776 238480 335782
rect 238428 335718 238480 335724
rect 238624 335578 238652 340054
rect 238612 335572 238664 335578
rect 238612 335514 238664 335520
rect 238900 335510 238928 340054
rect 239268 337618 239296 340068
rect 239256 337612 239308 337618
rect 239256 337554 239308 337560
rect 239348 335776 239400 335782
rect 239348 335718 239400 335724
rect 238888 335504 238940 335510
rect 238888 335446 238940 335452
rect 239256 321632 239308 321638
rect 239256 321574 239308 321580
rect 239268 302326 239296 321574
rect 239360 302326 239388 335718
rect 239440 335504 239492 335510
rect 239440 335446 239492 335452
rect 239452 321638 239480 335446
rect 239440 321632 239492 321638
rect 239440 321574 239492 321580
rect 239256 302320 239308 302326
rect 239256 302262 239308 302268
rect 239348 302320 239400 302326
rect 239348 302262 239400 302268
rect 239256 302184 239308 302190
rect 239256 302126 239308 302132
rect 239348 302184 239400 302190
rect 239348 302126 239400 302132
rect 239268 299470 239296 302126
rect 239256 299464 239308 299470
rect 239256 299406 239308 299412
rect 239256 273284 239308 273290
rect 239256 273226 239308 273232
rect 239268 263634 239296 273226
rect 239256 263628 239308 263634
rect 239256 263570 239308 263576
rect 239256 244384 239308 244390
rect 239256 244326 239308 244332
rect 239268 244186 239296 244326
rect 239256 244180 239308 244186
rect 239256 244122 239308 244128
rect 239256 225684 239308 225690
rect 239256 225626 239308 225632
rect 239268 205562 239296 225626
rect 239360 222290 239388 302126
rect 239440 299464 239492 299470
rect 239440 299406 239492 299412
rect 239452 273290 239480 299406
rect 239440 273284 239492 273290
rect 239440 273226 239492 273232
rect 239440 263628 239492 263634
rect 239440 263570 239492 263576
rect 239452 244390 239480 263570
rect 239440 244384 239492 244390
rect 239440 244326 239492 244332
rect 239440 244180 239492 244186
rect 239440 244122 239492 244128
rect 239452 225690 239480 244122
rect 239440 225684 239492 225690
rect 239440 225626 239492 225632
rect 239348 222284 239400 222290
rect 239348 222226 239400 222232
rect 239348 222148 239400 222154
rect 239348 222090 239400 222096
rect 239256 205556 239308 205562
rect 239256 205498 239308 205504
rect 239256 167136 239308 167142
rect 239256 167078 239308 167084
rect 239268 166938 239296 167078
rect 239256 166932 239308 166938
rect 239256 166874 239308 166880
rect 239256 128512 239308 128518
rect 239256 128454 239308 128460
rect 239268 128314 239296 128454
rect 239256 128308 239308 128314
rect 239256 128250 239308 128256
rect 239256 106276 239308 106282
rect 239256 106218 239308 106224
rect 239268 96665 239296 106218
rect 239254 96656 239310 96665
rect 239254 96591 239310 96600
rect 239254 51096 239310 51105
rect 239254 51031 239256 51040
rect 239308 51031 239310 51040
rect 239256 51002 239308 51008
rect 239256 17332 239308 17338
rect 239256 17274 239308 17280
rect 238520 10804 238572 10810
rect 238348 10764 238468 10792
rect 238244 10668 238296 10674
rect 238244 10610 238296 10616
rect 238058 4176 238114 4185
rect 238058 4111 238060 4120
rect 238112 4111 238114 4120
rect 238060 4082 238112 4088
rect 237968 4072 238020 4078
rect 237968 4014 238020 4020
rect 238440 3602 238468 10764
rect 238520 10746 238572 10752
rect 238532 10169 238560 10746
rect 239268 10742 239296 17274
rect 239256 10736 239308 10742
rect 239256 10678 239308 10684
rect 238518 10160 238574 10169
rect 238518 10095 238574 10104
rect 238888 7880 238940 7886
rect 238888 7822 238940 7828
rect 238428 3596 238480 3602
rect 238428 3538 238480 3544
rect 238900 480 238928 7822
rect 239360 4010 239388 222090
rect 239440 205556 239492 205562
rect 239440 205498 239492 205504
rect 239452 167142 239480 205498
rect 239440 167136 239492 167142
rect 239440 167078 239492 167084
rect 239440 166932 239492 166938
rect 239440 166874 239492 166880
rect 239452 128518 239480 166874
rect 239440 128512 239492 128518
rect 239440 128454 239492 128460
rect 239440 128308 239492 128314
rect 239440 128250 239492 128256
rect 239452 106282 239480 128250
rect 239440 106276 239492 106282
rect 239440 106218 239492 106224
rect 239438 96656 239494 96665
rect 239438 96591 239494 96600
rect 239452 51105 239480 96591
rect 239438 51096 239494 51105
rect 239438 51031 239440 51040
rect 239492 51031 239494 51040
rect 239440 51002 239492 51008
rect 239452 6225 239480 51002
rect 239544 17338 239572 340068
rect 239728 340054 239834 340082
rect 239912 340054 240018 340082
rect 240096 340054 240294 340082
rect 240372 340054 240570 340082
rect 240754 340054 240860 340082
rect 239624 335572 239676 335578
rect 239624 335514 239676 335520
rect 239532 17332 239584 17338
rect 239532 17274 239584 17280
rect 239636 10266 239664 335514
rect 239624 10260 239676 10266
rect 239624 10202 239676 10208
rect 239438 6216 239494 6225
rect 239438 6151 239494 6160
rect 239348 4004 239400 4010
rect 239348 3946 239400 3952
rect 239728 3738 239756 340054
rect 239912 335782 239940 340054
rect 239900 335776 239952 335782
rect 239900 335718 239952 335724
rect 240096 335510 240124 340054
rect 240372 335578 240400 340054
rect 240832 335578 240860 340054
rect 240912 339108 240964 339114
rect 240912 339050 240964 339056
rect 240360 335572 240412 335578
rect 240360 335514 240412 335520
rect 240820 335572 240872 335578
rect 240820 335514 240872 335520
rect 240084 335504 240136 335510
rect 240084 335446 240136 335452
rect 240820 335436 240872 335442
rect 240820 335378 240872 335384
rect 240082 9344 240138 9353
rect 240082 9279 240138 9288
rect 239716 3732 239768 3738
rect 239716 3674 239768 3680
rect 240096 480 240124 9279
rect 240832 6361 240860 335378
rect 240924 10198 240952 339050
rect 240912 10192 240964 10198
rect 240912 10134 240964 10140
rect 241016 6633 241044 340068
rect 241292 339114 241320 340068
rect 241280 339108 241332 339114
rect 241280 339050 241332 339056
rect 241476 337754 241504 340068
rect 241568 340054 241766 340082
rect 241464 337748 241516 337754
rect 241464 337690 241516 337696
rect 241096 335572 241148 335578
rect 241096 335514 241148 335520
rect 241002 6624 241058 6633
rect 241002 6559 241058 6568
rect 240818 6352 240874 6361
rect 240818 6287 240874 6296
rect 241108 3534 241136 335514
rect 241568 335442 241596 340054
rect 242028 335510 242056 340068
rect 242226 340054 242424 340082
rect 242108 339108 242160 339114
rect 242108 339050 242160 339056
rect 242016 335504 242068 335510
rect 242016 335446 242068 335452
rect 241556 335436 241608 335442
rect 241556 335378 241608 335384
rect 242120 331242 242148 339050
rect 242396 335730 242424 340054
rect 242488 339114 242516 340068
rect 242580 340054 242778 340082
rect 242476 339108 242528 339114
rect 242476 339050 242528 339056
rect 242396 335702 242516 335730
rect 242384 335572 242436 335578
rect 242384 335514 242436 335520
rect 242292 335504 242344 335510
rect 242292 335446 242344 335452
rect 242120 331214 242240 331242
rect 242212 319025 242240 331214
rect 242198 319016 242254 319025
rect 242198 318951 242254 318960
rect 242198 318880 242254 318889
rect 242198 318815 242254 318824
rect 242212 285682 242240 318815
rect 242120 285654 242240 285682
rect 242120 278866 242148 285654
rect 242108 278860 242160 278866
rect 242108 278802 242160 278808
rect 242108 277364 242160 277370
rect 242108 277306 242160 277312
rect 242120 254946 242148 277306
rect 242120 254918 242240 254946
rect 242212 246378 242240 254918
rect 242120 246350 242240 246378
rect 242120 231878 242148 246350
rect 242108 231872 242160 231878
rect 242108 231814 242160 231820
rect 242200 231872 242252 231878
rect 242200 231814 242252 231820
rect 242212 222290 242240 231814
rect 242200 222284 242252 222290
rect 242200 222226 242252 222232
rect 242108 222148 242160 222154
rect 242108 222090 242160 222096
rect 242120 213194 242148 222090
rect 242120 213166 242240 213194
rect 242212 203402 242240 213166
rect 242120 203374 242240 203402
rect 242120 193882 242148 203374
rect 242120 193854 242240 193882
rect 242212 182170 242240 193854
rect 242108 182164 242160 182170
rect 242108 182106 242160 182112
rect 242200 182164 242252 182170
rect 242200 182106 242252 182112
rect 242120 164218 242148 182106
rect 242108 164212 242160 164218
rect 242108 164154 242160 164160
rect 242200 164144 242252 164150
rect 242200 164086 242252 164092
rect 242212 162858 242240 164086
rect 242016 162852 242068 162858
rect 242016 162794 242068 162800
rect 242200 162852 242252 162858
rect 242200 162794 242252 162800
rect 242028 153241 242056 162794
rect 242014 153232 242070 153241
rect 242014 153167 242070 153176
rect 242198 153232 242254 153241
rect 242198 153167 242254 153176
rect 242212 149682 242240 153167
rect 242120 149654 242240 149682
rect 242120 144906 242148 149654
rect 242108 144900 242160 144906
rect 242108 144842 242160 144848
rect 242200 144900 242252 144906
rect 242200 144842 242252 144848
rect 242212 143546 242240 144842
rect 242016 143540 242068 143546
rect 242016 143482 242068 143488
rect 242200 143540 242252 143546
rect 242200 143482 242252 143488
rect 241830 134056 241886 134065
rect 241830 133991 241886 134000
rect 241844 132841 241872 133991
rect 242028 133929 242056 143482
rect 242014 133920 242070 133929
rect 242014 133855 242070 133864
rect 242198 133920 242254 133929
rect 242198 133855 242254 133864
rect 241830 132832 241886 132841
rect 241830 132767 241886 132776
rect 242212 125769 242240 133855
rect 242198 125760 242254 125769
rect 242198 125695 242254 125704
rect 242106 125624 242162 125633
rect 242106 125559 242162 125568
rect 242120 115818 242148 125559
rect 242120 115790 242240 115818
rect 242212 106457 242240 115790
rect 242198 106448 242254 106457
rect 242198 106383 242254 106392
rect 242106 106312 242162 106321
rect 242106 106247 242162 106256
rect 242120 101454 242148 106247
rect 242108 101448 242160 101454
rect 242108 101390 242160 101396
rect 242016 93900 242068 93906
rect 242016 93842 242068 93848
rect 242028 86850 242056 93842
rect 242028 86822 242240 86850
rect 242212 80730 242240 86822
rect 242028 80702 242240 80730
rect 242028 67658 242056 80702
rect 242016 67652 242068 67658
rect 242016 67594 242068 67600
rect 242108 67652 242160 67658
rect 242108 67594 242160 67600
rect 242120 46918 242148 67594
rect 242016 46912 242068 46918
rect 242016 46854 242068 46860
rect 242108 46912 242160 46918
rect 242108 46854 242160 46860
rect 242028 37262 242056 46854
rect 242016 37256 242068 37262
rect 242016 37198 242068 37204
rect 242108 37256 242160 37262
rect 242108 37198 242160 37204
rect 242120 22794 242148 37198
rect 242120 22766 242240 22794
rect 241924 10124 241976 10130
rect 241924 10066 241976 10072
rect 241936 10033 241964 10066
rect 241922 10024 241978 10033
rect 241922 9959 241978 9968
rect 242212 6497 242240 22766
rect 242304 11014 242332 335446
rect 242292 11008 242344 11014
rect 242292 10950 242344 10956
rect 242396 10130 242424 335514
rect 242488 321450 242516 335702
rect 242580 335578 242608 340054
rect 242948 338094 242976 340068
rect 243132 340054 243238 340082
rect 243514 340054 243620 340082
rect 243698 340054 243896 340082
rect 242936 338088 242988 338094
rect 242936 338030 242988 338036
rect 243132 335594 243160 340054
rect 242568 335572 242620 335578
rect 242568 335514 242620 335520
rect 242764 335566 243160 335594
rect 243592 335594 243620 340054
rect 243592 335566 243804 335594
rect 242764 321722 242792 335566
rect 243580 335504 243632 335510
rect 243580 335446 243632 335452
rect 242672 321694 242792 321722
rect 242488 321422 242608 321450
rect 242580 309194 242608 321422
rect 242672 314022 242700 321694
rect 242660 314016 242712 314022
rect 242660 313958 242712 313964
rect 242844 314016 242896 314022
rect 242844 313958 242896 313964
rect 242476 309188 242528 309194
rect 242476 309130 242528 309136
rect 242568 309188 242620 309194
rect 242568 309130 242620 309136
rect 242488 299538 242516 309130
rect 242856 304314 242884 313958
rect 242764 304286 242884 304314
rect 242476 299532 242528 299538
rect 242476 299474 242528 299480
rect 242568 299532 242620 299538
rect 242568 299474 242620 299480
rect 242580 267850 242608 299474
rect 242764 285682 242792 304286
rect 242672 285654 242792 285682
rect 242672 276185 242700 285654
rect 242658 276176 242714 276185
rect 242658 276111 242714 276120
rect 242750 276040 242806 276049
rect 242750 275975 242806 275984
rect 242764 269754 242792 275975
rect 242752 269748 242804 269754
rect 242752 269690 242804 269696
rect 242568 267844 242620 267850
rect 242568 267786 242620 267792
rect 242476 267776 242528 267782
rect 242476 267718 242528 267724
rect 242488 264738 242516 267718
rect 242936 267572 242988 267578
rect 242936 267514 242988 267520
rect 242948 264858 242976 267514
rect 242936 264852 242988 264858
rect 242936 264794 242988 264800
rect 242488 264710 242608 264738
rect 242580 255270 242608 264710
rect 242844 255332 242896 255338
rect 242844 255274 242896 255280
rect 242568 255264 242620 255270
rect 242856 255218 242884 255274
rect 242568 255206 242620 255212
rect 242764 255190 242884 255218
rect 242764 246838 242792 255190
rect 242752 246832 242804 246838
rect 242752 246774 242804 246780
rect 242660 245676 242712 245682
rect 242660 245618 242712 245624
rect 242672 242026 242700 245618
rect 242488 241998 242700 242026
rect 242752 242004 242804 242010
rect 242488 237386 242516 241998
rect 242752 241946 242804 241952
rect 242476 237380 242528 237386
rect 242476 237322 242528 237328
rect 242764 229106 242792 241946
rect 242672 229078 242792 229106
rect 242672 228834 242700 229078
rect 242672 228806 242792 228834
rect 242474 218104 242530 218113
rect 242474 218039 242530 218048
rect 242488 216646 242516 218039
rect 242476 216640 242528 216646
rect 242476 216582 242528 216588
rect 242476 207052 242528 207058
rect 242476 206994 242528 207000
rect 242488 201550 242516 206994
rect 242476 201544 242528 201550
rect 242476 201486 242528 201492
rect 242568 201408 242620 201414
rect 242568 201350 242620 201356
rect 242580 198694 242608 201350
rect 242568 198688 242620 198694
rect 242568 198630 242620 198636
rect 242764 191842 242792 228806
rect 242844 227792 242896 227798
rect 242844 227734 242896 227740
rect 242856 218249 242884 227734
rect 242842 218240 242898 218249
rect 242842 218175 242898 218184
rect 242764 191814 242884 191842
rect 242476 189100 242528 189106
rect 242476 189042 242528 189048
rect 242488 182209 242516 189042
rect 242856 189038 242884 191814
rect 242844 189032 242896 189038
rect 242844 188974 242896 188980
rect 242474 182200 242530 182209
rect 242474 182135 242530 182144
rect 242844 182028 242896 182034
rect 242844 181970 242896 181976
rect 242856 164257 242884 181970
rect 242658 164248 242714 164257
rect 242658 164183 242660 164192
rect 242712 164183 242714 164192
rect 242842 164248 242898 164257
rect 242842 164183 242898 164192
rect 242660 164154 242712 164160
rect 242566 163024 242622 163033
rect 242566 162959 242622 162968
rect 242580 162926 242608 162959
rect 242568 162920 242620 162926
rect 242568 162862 242620 162868
rect 242476 157956 242528 157962
rect 242476 157898 242528 157904
rect 242488 157865 242516 157898
rect 242474 157856 242530 157865
rect 242474 157791 242530 157800
rect 242660 157140 242712 157146
rect 242660 157082 242712 157088
rect 242474 144936 242530 144945
rect 242474 144871 242530 144880
rect 242488 143546 242516 144871
rect 242672 144838 242700 157082
rect 242660 144832 242712 144838
rect 242660 144774 242712 144780
rect 242752 144832 242804 144838
rect 242752 144774 242804 144780
rect 242476 143540 242528 143546
rect 242476 143482 242528 143488
rect 242568 143540 242620 143546
rect 242568 143482 242620 143488
rect 242580 119406 242608 143482
rect 242764 130370 242792 144774
rect 242764 130342 242884 130370
rect 242856 125594 242884 130342
rect 242844 125588 242896 125594
rect 242844 125530 242896 125536
rect 242568 119400 242620 119406
rect 242568 119342 242620 119348
rect 242936 119400 242988 119406
rect 242936 119342 242988 119348
rect 242844 116748 242896 116754
rect 242844 116690 242896 116696
rect 242856 114510 242884 116690
rect 242844 114504 242896 114510
rect 242844 114446 242896 114452
rect 242948 111178 242976 119342
rect 242936 111172 242988 111178
rect 242936 111114 242988 111120
rect 242936 110560 242988 110566
rect 242936 110502 242988 110508
rect 242660 104916 242712 104922
rect 242660 104858 242712 104864
rect 242672 96665 242700 104858
rect 242948 101402 242976 110502
rect 242856 101374 242976 101402
rect 242474 96656 242530 96665
rect 242474 96591 242530 96600
rect 242658 96656 242714 96665
rect 242658 96591 242714 96600
rect 242488 87242 242516 96591
rect 242476 87236 242528 87242
rect 242476 87178 242528 87184
rect 242856 86970 242884 101374
rect 242844 86964 242896 86970
rect 242844 86906 242896 86912
rect 242936 86964 242988 86970
rect 242936 86906 242988 86912
rect 242476 86896 242528 86902
rect 242476 86838 242528 86844
rect 242488 85542 242516 86838
rect 242476 85536 242528 85542
rect 242476 85478 242528 85484
rect 242568 85332 242620 85338
rect 242568 85274 242620 85280
rect 242580 65006 242608 85274
rect 242948 77353 242976 86906
rect 242750 77344 242806 77353
rect 242750 77279 242806 77288
rect 242934 77344 242990 77353
rect 242934 77279 242990 77288
rect 242764 72434 242792 77279
rect 242672 72406 242792 72434
rect 242568 65000 242620 65006
rect 242568 64942 242620 64948
rect 242476 64932 242528 64938
rect 242476 64874 242528 64880
rect 242488 63510 242516 64874
rect 242476 63504 242528 63510
rect 242476 63446 242528 63452
rect 242672 57882 242700 72406
rect 242672 57854 242792 57882
rect 242764 48346 242792 57854
rect 242752 48340 242804 48346
rect 242752 48282 242804 48288
rect 242844 48340 242896 48346
rect 242844 48282 242896 48288
rect 242568 45620 242620 45626
rect 242568 45562 242620 45568
rect 242580 41834 242608 45562
rect 242580 41806 242700 41834
rect 242672 29102 242700 41806
rect 242660 29096 242712 29102
rect 242660 29038 242712 29044
rect 242856 29034 242884 48282
rect 242752 29028 242804 29034
rect 242752 28970 242804 28976
rect 242844 29028 242896 29034
rect 242844 28970 242896 28976
rect 242568 28960 242620 28966
rect 242568 28902 242620 28908
rect 242580 27606 242608 28902
rect 242568 27600 242620 27606
rect 242568 27542 242620 27548
rect 242568 22704 242620 22710
rect 242568 22646 242620 22652
rect 242580 18057 242608 22646
rect 242764 18154 242792 28970
rect 242752 18148 242804 18154
rect 242752 18090 242804 18096
rect 242660 18080 242712 18086
rect 242566 18048 242622 18057
rect 242660 18022 242712 18028
rect 242750 18048 242806 18057
rect 242566 17983 242622 17992
rect 242672 17338 242700 18022
rect 242750 17983 242806 17992
rect 242476 17332 242528 17338
rect 242476 17274 242528 17280
rect 242660 17332 242712 17338
rect 242660 17274 242712 17280
rect 242384 10124 242436 10130
rect 242384 10066 242436 10072
rect 242488 8106 242516 17274
rect 242396 8078 242516 8106
rect 242396 7954 242424 8078
rect 242384 7948 242436 7954
rect 242384 7890 242436 7896
rect 242476 7948 242528 7954
rect 242476 7890 242528 7896
rect 242198 6488 242254 6497
rect 242198 6423 242254 6432
rect 241280 4072 241332 4078
rect 241280 4014 241332 4020
rect 241096 3528 241148 3534
rect 241096 3470 241148 3476
rect 241292 480 241320 4014
rect 242488 480 242516 7890
rect 242764 4146 242792 17983
rect 243592 8022 243620 335446
rect 243776 10674 243804 335566
rect 243764 10668 243816 10674
rect 243764 10610 243816 10616
rect 243580 8016 243632 8022
rect 243580 7958 243632 7964
rect 242752 4140 242804 4146
rect 242752 4082 242804 4088
rect 243672 3664 243724 3670
rect 243672 3606 243724 3612
rect 243684 480 243712 3606
rect 243868 3398 243896 340054
rect 243960 335510 243988 340068
rect 244144 340054 244250 340082
rect 244040 335572 244092 335578
rect 244040 335514 244092 335520
rect 243948 335504 244000 335510
rect 243948 335446 244000 335452
rect 244052 8090 244080 335514
rect 244144 10810 244172 340054
rect 244420 337210 244448 340068
rect 244512 340054 244710 340082
rect 244408 337204 244460 337210
rect 244408 337146 244460 337152
rect 244512 335578 244540 340054
rect 244500 335572 244552 335578
rect 244500 335514 244552 335520
rect 244868 335572 244920 335578
rect 244868 335514 244920 335520
rect 244880 11830 244908 335514
rect 244868 11824 244920 11830
rect 244868 11766 244920 11772
rect 244972 11762 245000 340068
rect 245052 335776 245104 335782
rect 245052 335718 245104 335724
rect 245064 324970 245092 335718
rect 245052 324964 245104 324970
rect 245052 324906 245104 324912
rect 244960 11756 245012 11762
rect 244960 11698 245012 11704
rect 244132 10804 244184 10810
rect 244132 10746 244184 10752
rect 244776 10124 244828 10130
rect 244776 10066 244828 10072
rect 244788 9178 244816 10066
rect 244868 9376 244920 9382
rect 244866 9344 244868 9353
rect 244920 9344 244922 9353
rect 244866 9279 244922 9288
rect 244866 9208 244922 9217
rect 244776 9172 244828 9178
rect 244866 9143 244868 9152
rect 244776 9114 244828 9120
rect 244920 9143 244922 9152
rect 244868 9114 244920 9120
rect 244040 8084 244092 8090
rect 244040 8026 244092 8032
rect 244774 5536 244830 5545
rect 244774 5471 244830 5480
rect 244788 5302 244816 5471
rect 244866 5400 244922 5409
rect 244866 5335 244922 5344
rect 244776 5296 244828 5302
rect 244776 5238 244828 5244
rect 244880 5234 244908 5335
rect 244958 5264 245014 5273
rect 244868 5228 244920 5234
rect 244958 5199 244960 5208
rect 244868 5170 244920 5176
rect 245012 5199 245014 5208
rect 244960 5170 245012 5176
rect 244868 4140 244920 4146
rect 244868 4082 244920 4088
rect 243856 3392 243908 3398
rect 243856 3334 243908 3340
rect 244880 480 244908 4082
rect 245156 3194 245184 340068
rect 245248 340054 245446 340082
rect 245524 340054 245630 340082
rect 245248 335782 245276 340054
rect 245420 336864 245472 336870
rect 245420 336806 245472 336812
rect 245236 335776 245288 335782
rect 245236 335718 245288 335724
rect 245432 291854 245460 336806
rect 245524 335578 245552 340054
rect 245892 337142 245920 340068
rect 245880 337136 245932 337142
rect 245880 337078 245932 337084
rect 245512 335572 245564 335578
rect 245512 335514 245564 335520
rect 246168 327758 246196 340068
rect 246260 340054 246366 340082
rect 246156 327752 246208 327758
rect 246156 327694 246208 327700
rect 245420 291848 245472 291854
rect 245420 291790 245472 291796
rect 246064 14544 246116 14550
rect 246064 14486 246116 14492
rect 245972 8016 246024 8022
rect 245972 7958 246024 7964
rect 245984 4026 246012 7958
rect 246076 4146 246104 14486
rect 246260 11898 246288 340054
rect 246628 338314 246656 340068
rect 246536 338286 246656 338314
rect 246720 340054 246918 340082
rect 246996 340054 247102 340082
rect 246536 338178 246564 338286
rect 246536 338150 246656 338178
rect 246432 331084 246484 331090
rect 246432 331026 246484 331032
rect 246444 294642 246472 331026
rect 246628 328522 246656 338150
rect 246720 331090 246748 340054
rect 246996 333282 247024 340054
rect 247364 337074 247392 340068
rect 247352 337068 247404 337074
rect 247352 337010 247404 337016
rect 247640 336870 247668 340068
rect 247838 340054 248036 340082
rect 247628 336864 247680 336870
rect 247628 336806 247680 336812
rect 247904 335776 247956 335782
rect 247904 335718 247956 335724
rect 247720 335572 247772 335578
rect 247720 335514 247772 335520
rect 246812 333254 247024 333282
rect 246708 331084 246760 331090
rect 246708 331026 246760 331032
rect 246628 328494 246748 328522
rect 246720 327146 246748 328494
rect 246524 327140 246576 327146
rect 246524 327082 246576 327088
rect 246708 327140 246760 327146
rect 246708 327082 246760 327088
rect 246432 294636 246484 294642
rect 246432 294578 246484 294584
rect 246536 285841 246564 327082
rect 246522 285832 246578 285841
rect 246522 285767 246578 285776
rect 246614 285696 246670 285705
rect 246614 285631 246670 285640
rect 246628 278866 246656 285631
rect 246616 278860 246668 278866
rect 246616 278802 246668 278808
rect 246616 277364 246668 277370
rect 246616 277306 246668 277312
rect 246628 254182 246656 277306
rect 246812 273358 246840 333254
rect 247732 276690 247760 335514
rect 247720 276684 247772 276690
rect 247720 276626 247772 276632
rect 246800 273352 246852 273358
rect 246800 273294 246852 273300
rect 246708 273216 246760 273222
rect 246708 273158 246760 273164
rect 246720 263514 246748 273158
rect 246720 263486 246840 263514
rect 246616 254176 246668 254182
rect 246616 254118 246668 254124
rect 246524 249824 246576 249830
rect 246444 249772 246524 249778
rect 246444 249766 246576 249772
rect 246444 249750 246564 249766
rect 246444 241466 246472 249750
rect 246432 241460 246484 241466
rect 246432 241402 246484 241408
rect 246708 241460 246760 241466
rect 246708 241402 246760 241408
rect 246720 231878 246748 241402
rect 246616 231872 246668 231878
rect 246616 231814 246668 231820
rect 246708 231872 246760 231878
rect 246708 231814 246760 231820
rect 246628 222290 246656 231814
rect 246616 222284 246668 222290
rect 246616 222226 246668 222232
rect 246812 222222 246840 263486
rect 246800 222216 246852 222222
rect 246800 222158 246852 222164
rect 246524 222148 246576 222154
rect 246524 222090 246576 222096
rect 246536 213058 246564 222090
rect 246800 222080 246852 222086
rect 246800 222022 246852 222028
rect 246444 213030 246564 213058
rect 246444 203538 246472 213030
rect 246812 208434 246840 222022
rect 246352 203510 246472 203538
rect 246720 208406 246840 208434
rect 246352 198801 246380 203510
rect 246338 198792 246394 198801
rect 246338 198727 246394 198736
rect 246430 198520 246486 198529
rect 246430 198455 246486 198464
rect 246444 189106 246472 198455
rect 246720 193934 246748 208406
rect 246708 193928 246760 193934
rect 246708 193870 246760 193876
rect 246984 193928 247036 193934
rect 246984 193870 247036 193876
rect 246432 189100 246484 189106
rect 246432 189042 246484 189048
rect 246616 189100 246668 189106
rect 246616 189042 246668 189048
rect 246628 182170 246656 189042
rect 246524 182164 246576 182170
rect 246524 182106 246576 182112
rect 246616 182164 246668 182170
rect 246616 182106 246668 182112
rect 246536 164218 246564 182106
rect 246996 169318 247024 193870
rect 246984 169312 247036 169318
rect 246984 169254 247036 169260
rect 246524 164212 246576 164218
rect 246524 164154 246576 164160
rect 246616 164144 246668 164150
rect 246616 164086 246668 164092
rect 246628 162858 246656 164086
rect 246616 162852 246668 162858
rect 246616 162794 246668 162800
rect 246892 161492 246944 161498
rect 246892 161434 246944 161440
rect 246904 159526 246932 161434
rect 246892 159520 246944 159526
rect 246892 159462 246944 159468
rect 246800 157140 246852 157146
rect 246800 157082 246852 157088
rect 246616 153264 246668 153270
rect 246616 153206 246668 153212
rect 246628 147762 246656 153206
rect 246812 147778 246840 157082
rect 246616 147756 246668 147762
rect 246616 147698 246668 147704
rect 246720 147750 246840 147778
rect 246720 147642 246748 147750
rect 246524 147620 246576 147626
rect 246720 147614 246932 147642
rect 246524 147562 246576 147568
rect 246536 135318 246564 147562
rect 246904 138106 246932 147614
rect 246892 138100 246944 138106
rect 246892 138042 246944 138048
rect 246800 137964 246852 137970
rect 246800 137906 246852 137912
rect 246524 135312 246576 135318
rect 246524 135254 246576 135260
rect 246524 135176 246576 135182
rect 246524 135118 246576 135124
rect 246536 125594 246564 135118
rect 246812 128466 246840 137906
rect 246720 128438 246840 128466
rect 246720 128330 246748 128438
rect 246720 128302 246840 128330
rect 246812 128194 246840 128302
rect 246812 128166 246932 128194
rect 246524 125588 246576 125594
rect 246524 125530 246576 125536
rect 246616 125520 246668 125526
rect 246616 125462 246668 125468
rect 246628 109154 246656 125462
rect 246628 109126 246748 109154
rect 246720 109018 246748 109126
rect 246628 108990 246748 109018
rect 246628 99482 246656 108990
rect 246616 99476 246668 99482
rect 246616 99418 246668 99424
rect 246616 99340 246668 99346
rect 246616 99282 246668 99288
rect 246628 90098 246656 99282
rect 246904 96801 246932 128166
rect 246890 96792 246946 96801
rect 246890 96727 246946 96736
rect 246798 96656 246854 96665
rect 246798 96591 246854 96600
rect 246616 90092 246668 90098
rect 246616 90034 246668 90040
rect 246524 88460 246576 88466
rect 246524 88402 246576 88408
rect 246536 82498 246564 88402
rect 246536 82470 246748 82498
rect 246720 70514 246748 82470
rect 246708 70508 246760 70514
rect 246708 70450 246760 70456
rect 246812 70394 246840 96591
rect 246720 70366 246840 70394
rect 246720 70258 246748 70366
rect 246720 70230 246840 70258
rect 246708 66292 246760 66298
rect 246708 66234 246760 66240
rect 246720 57746 246748 66234
rect 246812 60330 246840 70230
rect 246812 60302 247024 60330
rect 246996 60058 247024 60302
rect 246536 57718 246748 57746
rect 246904 60030 247024 60058
rect 246536 46866 246564 57718
rect 246904 55214 246932 60030
rect 246892 55208 246944 55214
rect 246892 55150 246944 55156
rect 246536 46838 246656 46866
rect 246628 29034 246656 46838
rect 246892 45620 246944 45626
rect 246892 45562 246944 45568
rect 246904 29102 246932 45562
rect 246892 29096 246944 29102
rect 246892 29038 246944 29044
rect 246524 29028 246576 29034
rect 246524 28970 246576 28976
rect 246616 29028 246668 29034
rect 246616 28970 246668 28976
rect 246708 29028 246760 29034
rect 246708 28970 246760 28976
rect 246536 27606 246564 28970
rect 246524 27600 246576 27606
rect 246524 27542 246576 27548
rect 246616 27600 246668 27606
rect 246616 27542 246668 27548
rect 246248 11892 246300 11898
rect 246248 11834 246300 11840
rect 246064 4140 246116 4146
rect 246064 4082 246116 4088
rect 245984 3998 246104 4026
rect 245144 3188 245196 3194
rect 245144 3130 245196 3136
rect 246076 480 246104 3998
rect 246628 3126 246656 27542
rect 246720 21842 246748 28970
rect 246720 21814 246840 21842
rect 246812 12458 246840 21814
rect 246720 12430 246840 12458
rect 246720 12102 246748 12430
rect 246708 12096 246760 12102
rect 246708 12038 246760 12044
rect 247260 3664 247312 3670
rect 247260 3606 247312 3612
rect 246616 3120 246668 3126
rect 246616 3062 246668 3068
rect 247272 480 247300 3606
rect 247916 3058 247944 335718
rect 248008 335594 248036 340054
rect 248100 337006 248128 340068
rect 248284 340054 248390 340082
rect 248468 340054 248574 340082
rect 248652 340054 248850 340082
rect 249126 340054 249232 340082
rect 248088 337000 248140 337006
rect 248088 336942 248140 336948
rect 248008 335566 248220 335594
rect 248192 12170 248220 335566
rect 248284 289134 248312 340054
rect 248468 335578 248496 340054
rect 248652 335782 248680 340054
rect 248640 335776 248692 335782
rect 248640 335718 248692 335724
rect 248456 335572 248508 335578
rect 248456 335514 248508 335520
rect 249008 335572 249060 335578
rect 249008 335514 249060 335520
rect 248272 289128 248324 289134
rect 248272 289070 248324 289076
rect 249020 89010 249048 335514
rect 249204 286346 249232 340054
rect 249192 286340 249244 286346
rect 249192 286282 249244 286288
rect 249008 89004 249060 89010
rect 249008 88946 249060 88952
rect 249296 12238 249324 340068
rect 249572 336938 249600 340068
rect 249664 340054 249862 340082
rect 249940 340054 250046 340082
rect 250322 340054 250428 340082
rect 249560 336932 249612 336938
rect 249560 336874 249612 336880
rect 249664 335594 249692 340054
rect 249744 336864 249796 336870
rect 249744 336806 249796 336812
rect 249480 335566 249692 335594
rect 249480 311846 249508 335566
rect 249756 335458 249784 336806
rect 249940 335578 249968 340054
rect 249928 335572 249980 335578
rect 249928 335514 249980 335520
rect 249572 335430 249784 335458
rect 250400 335458 250428 340054
rect 250584 336870 250612 340068
rect 250572 336864 250624 336870
rect 250572 336806 250624 336812
rect 250400 335430 250704 335458
rect 249468 311840 249520 311846
rect 249468 311782 249520 311788
rect 249376 295316 249428 295322
rect 249376 295258 249428 295264
rect 249388 283626 249416 295258
rect 249376 283620 249428 283626
rect 249376 283562 249428 283568
rect 249572 279478 249600 335430
rect 250388 335368 250440 335374
rect 250388 335310 250440 335316
rect 249652 311840 249704 311846
rect 249652 311782 249704 311788
rect 249664 295322 249692 311782
rect 249652 295316 249704 295322
rect 249652 295258 249704 295264
rect 249560 279472 249612 279478
rect 249560 279414 249612 279420
rect 249284 12232 249336 12238
rect 249284 12174 249336 12180
rect 248180 12164 248232 12170
rect 248180 12106 248232 12112
rect 248824 11756 248876 11762
rect 248824 11698 248876 11704
rect 247904 3052 247956 3058
rect 247904 2994 247956 3000
rect 248836 610 248864 11698
rect 250400 10062 250428 335310
rect 250480 335300 250532 335306
rect 250480 335242 250532 335248
rect 250492 12306 250520 335242
rect 250480 12300 250532 12306
rect 250480 12242 250532 12248
rect 250388 10056 250440 10062
rect 250388 9998 250440 10004
rect 249652 8084 249704 8090
rect 249652 8026 249704 8032
rect 248456 604 248508 610
rect 248456 546 248508 552
rect 248824 604 248876 610
rect 248824 546 248876 552
rect 248468 480 248496 546
rect 249664 480 249692 8026
rect 250676 2990 250704 335430
rect 250768 335306 250796 340068
rect 251044 337210 251072 340068
rect 251136 340054 251334 340082
rect 251412 340054 251518 340082
rect 251794 340054 251992 340082
rect 252070 340054 252176 340082
rect 252254 340054 252452 340082
rect 251032 337204 251084 337210
rect 251032 337146 251084 337152
rect 251136 335374 251164 340054
rect 251124 335368 251176 335374
rect 251124 335310 251176 335316
rect 250756 335300 250808 335306
rect 250756 335242 250808 335248
rect 251412 335186 251440 340054
rect 251584 337612 251636 337618
rect 251584 337554 251636 337560
rect 250952 335158 251440 335186
rect 250952 307086 250980 335158
rect 250940 307080 250992 307086
rect 250940 307022 250992 307028
rect 251596 3058 251624 337554
rect 251964 335458 251992 340054
rect 252148 335594 252176 340054
rect 252148 335566 252360 335594
rect 251964 335430 252176 335458
rect 251860 335368 251912 335374
rect 251860 335310 251912 335316
rect 251676 241800 251728 241806
rect 251674 241768 251676 241777
rect 251728 241768 251730 241777
rect 251674 241703 251730 241712
rect 251674 179616 251730 179625
rect 251674 179551 251730 179560
rect 251688 179450 251716 179551
rect 251676 179444 251728 179450
rect 251676 179386 251728 179392
rect 251766 132968 251822 132977
rect 251766 132903 251822 132912
rect 251780 132705 251808 132903
rect 251766 132696 251822 132705
rect 251766 132631 251822 132640
rect 251676 100904 251728 100910
rect 251674 100872 251676 100881
rect 251728 100872 251730 100881
rect 251674 100807 251730 100816
rect 251872 9926 251900 335310
rect 251952 335300 252004 335306
rect 251952 335242 252004 335248
rect 251964 12374 251992 335242
rect 251952 12368 252004 12374
rect 251952 12310 252004 12316
rect 251860 9920 251912 9926
rect 251860 9862 251912 9868
rect 251952 4140 252004 4146
rect 251952 4082 252004 4088
rect 250848 3052 250900 3058
rect 250848 2994 250900 3000
rect 251584 3052 251636 3058
rect 251584 2994 251636 3000
rect 250664 2984 250716 2990
rect 250664 2926 250716 2932
rect 250860 480 250888 2994
rect 251964 480 251992 4082
rect 252148 2922 252176 335430
rect 252332 9994 252360 335566
rect 252424 335306 252452 340054
rect 252516 337414 252544 340068
rect 252608 340054 252806 340082
rect 252884 340054 252990 340082
rect 253266 340054 253464 340082
rect 252504 337408 252556 337414
rect 252504 337350 252556 337356
rect 252608 335374 252636 340054
rect 252596 335368 252648 335374
rect 252596 335310 252648 335316
rect 252412 335300 252464 335306
rect 252412 335242 252464 335248
rect 252884 328506 252912 340054
rect 253148 335776 253200 335782
rect 253148 335718 253200 335724
rect 252504 328500 252556 328506
rect 252504 328442 252556 328448
rect 252872 328500 252924 328506
rect 252872 328442 252924 328448
rect 252516 320890 252544 328442
rect 252504 320884 252556 320890
rect 252504 320826 252556 320832
rect 252964 14476 253016 14482
rect 252964 14418 253016 14424
rect 252320 9988 252372 9994
rect 252320 9930 252372 9936
rect 252976 4146 253004 14418
rect 253160 10470 253188 335718
rect 253332 335572 253384 335578
rect 253332 335514 253384 335520
rect 253344 12442 253372 335514
rect 253332 12436 253384 12442
rect 253332 12378 253384 12384
rect 253148 10464 253200 10470
rect 253148 10406 253200 10412
rect 252964 4140 253016 4146
rect 252964 4082 253016 4088
rect 253148 3188 253200 3194
rect 253148 3130 253200 3136
rect 252136 2916 252188 2922
rect 252136 2858 252188 2864
rect 253160 480 253188 3130
rect 253436 2854 253464 340054
rect 253528 10198 253556 340068
rect 253620 340054 253726 340082
rect 253620 335578 253648 340054
rect 253988 337550 254016 340068
rect 254080 340054 254278 340082
rect 253976 337544 254028 337550
rect 253976 337486 254028 337492
rect 254080 335782 254108 340054
rect 254344 337544 254396 337550
rect 254344 337486 254396 337492
rect 254252 337408 254304 337414
rect 254252 337350 254304 337356
rect 254068 335776 254120 335782
rect 254068 335718 254120 335724
rect 253608 335572 253660 335578
rect 253608 335514 253660 335520
rect 254160 320544 254212 320550
rect 254158 320512 254160 320521
rect 254212 320512 254214 320521
rect 254158 320447 254214 320456
rect 253516 10192 253568 10198
rect 253516 10134 253568 10140
rect 254264 9330 254292 337350
rect 254172 9302 254292 9330
rect 254172 3194 254200 9302
rect 254250 9208 254306 9217
rect 254250 9143 254252 9152
rect 254304 9143 254306 9152
rect 254252 9114 254304 9120
rect 254160 3188 254212 3194
rect 254160 3130 254212 3136
rect 253424 2848 253476 2854
rect 253424 2790 253476 2796
rect 254356 480 254384 337486
rect 254448 331974 254476 340068
rect 254540 340054 254738 340082
rect 254436 331968 254488 331974
rect 254436 331910 254488 331916
rect 254540 9330 254568 340054
rect 254804 338564 254856 338570
rect 254804 338506 254856 338512
rect 254620 335776 254672 335782
rect 254620 335718 254672 335724
rect 254632 10538 254660 335718
rect 254712 335572 254764 335578
rect 254712 335514 254764 335520
rect 254724 331226 254752 335514
rect 254712 331220 254764 331226
rect 254712 331162 254764 331168
rect 254816 316742 254844 338506
rect 254896 331220 254948 331226
rect 254896 331162 254948 331168
rect 254804 316736 254856 316742
rect 254804 316678 254856 316684
rect 254908 273306 254936 331162
rect 254816 273278 254936 273306
rect 254816 195922 254844 273278
rect 254816 195894 254936 195922
rect 254908 167090 254936 195894
rect 254816 167062 254936 167090
rect 254816 157162 254844 167062
rect 254816 157134 254936 157162
rect 254908 128466 254936 157134
rect 254816 128438 254936 128466
rect 254816 109018 254844 128438
rect 254816 108990 254936 109018
rect 254908 89842 254936 108990
rect 254816 89814 254936 89842
rect 254816 79914 254844 89814
rect 254816 79886 254936 79914
rect 254908 60738 254936 79886
rect 254816 60710 254936 60738
rect 254816 60602 254844 60710
rect 254816 60574 254936 60602
rect 254908 28966 254936 60574
rect 254896 28960 254948 28966
rect 254896 28902 254948 28908
rect 254804 21412 254856 21418
rect 254804 21354 254856 21360
rect 254620 10532 254672 10538
rect 254620 10474 254672 10480
rect 254540 9302 254752 9330
rect 254526 9208 254582 9217
rect 254436 9172 254488 9178
rect 254526 9143 254528 9152
rect 254436 9114 254488 9120
rect 254580 9143 254582 9152
rect 254528 9114 254580 9120
rect 254448 8945 254476 9114
rect 254434 8936 254490 8945
rect 254434 8871 254490 8880
rect 254724 3466 254752 9302
rect 254816 3738 254844 21354
rect 255000 10606 255028 340068
rect 255184 338570 255212 340068
rect 255276 340054 255474 340082
rect 255552 340054 255750 340082
rect 255172 338564 255224 338570
rect 255172 338506 255224 338512
rect 255276 335578 255304 340054
rect 255552 335782 255580 340054
rect 255540 335776 255592 335782
rect 255540 335718 255592 335724
rect 255264 335572 255316 335578
rect 255264 335514 255316 335520
rect 255920 271182 255948 340068
rect 256196 337482 256224 340068
rect 256184 337476 256236 337482
rect 256184 337418 256236 337424
rect 256472 336054 256500 340068
rect 256564 340054 256670 340082
rect 256748 340054 256946 340082
rect 257222 340054 257328 340082
rect 256460 336048 256512 336054
rect 256460 335990 256512 335996
rect 256564 335730 256592 340054
rect 256012 335702 256592 335730
rect 256012 304298 256040 335702
rect 256748 335594 256776 340054
rect 257104 337476 257156 337482
rect 257104 337418 257156 337424
rect 256828 336864 256880 336870
rect 256828 336806 256880 336812
rect 256104 335566 256776 335594
rect 256000 304292 256052 304298
rect 256000 304234 256052 304240
rect 255908 271176 255960 271182
rect 255908 271118 255960 271124
rect 254988 10600 255040 10606
rect 254988 10542 255040 10548
rect 255724 10464 255776 10470
rect 255724 10406 255776 10412
rect 254894 8936 254950 8945
rect 254894 8871 254950 8880
rect 254908 8838 254936 8871
rect 254896 8832 254948 8838
rect 254896 8774 254948 8780
rect 255078 7576 255134 7585
rect 255078 7511 255134 7520
rect 255092 7177 255120 7511
rect 255078 7168 255134 7177
rect 255078 7103 255134 7112
rect 254804 3732 254856 3738
rect 254804 3674 254856 3680
rect 254712 3460 254764 3466
rect 254712 3402 254764 3408
rect 255736 626 255764 10406
rect 256104 8294 256132 335566
rect 256840 335458 256868 336806
rect 256472 335430 256868 335458
rect 256472 318102 256500 335430
rect 256460 318096 256512 318102
rect 256460 318038 256512 318044
rect 256092 8288 256144 8294
rect 256092 8230 256144 8236
rect 255552 598 255764 626
rect 257116 610 257144 337418
rect 257300 5409 257328 340054
rect 257392 6390 257420 340068
rect 257576 340054 257682 340082
rect 257760 340054 257958 340082
rect 257472 335572 257524 335578
rect 257472 335514 257524 335520
rect 257484 9654 257512 335514
rect 257576 319462 257604 340054
rect 257564 319456 257616 319462
rect 257564 319398 257616 319404
rect 257472 9648 257524 9654
rect 257472 9590 257524 9596
rect 257380 6384 257432 6390
rect 257380 6326 257432 6332
rect 257760 5545 257788 340054
rect 258128 332058 258156 340068
rect 258220 340054 258418 340082
rect 258220 335578 258248 340054
rect 258680 336870 258708 340068
rect 258668 336864 258720 336870
rect 258668 336806 258720 336812
rect 258208 335572 258260 335578
rect 258208 335514 258260 335520
rect 258760 335572 258812 335578
rect 258760 335514 258812 335520
rect 257944 332030 258156 332058
rect 257944 322250 257972 332030
rect 257932 322244 257984 322250
rect 257932 322186 257984 322192
rect 258772 300150 258800 335514
rect 258864 301510 258892 340068
rect 259140 331430 259168 340068
rect 259232 340054 259430 340082
rect 259508 340054 259614 340082
rect 259784 340054 259890 340082
rect 259232 338094 259260 340054
rect 259220 338088 259272 338094
rect 259220 338030 259272 338036
rect 259508 335578 259536 340054
rect 259496 335572 259548 335578
rect 259496 335514 259548 335520
rect 259128 331424 259180 331430
rect 259128 331366 259180 331372
rect 259036 331220 259088 331226
rect 259036 331162 259088 331168
rect 258944 321632 258996 321638
rect 258944 321574 258996 321580
rect 258956 315314 258984 321574
rect 258944 315308 258996 315314
rect 258944 315250 258996 315256
rect 258852 301504 258904 301510
rect 258852 301446 258904 301452
rect 258760 300144 258812 300150
rect 258760 300086 258812 300092
rect 259048 9518 259076 331162
rect 259128 331152 259180 331158
rect 259128 331094 259180 331100
rect 259140 321638 259168 331094
rect 259784 328506 259812 340054
rect 260048 335776 260100 335782
rect 260048 335718 260100 335724
rect 259312 328500 259364 328506
rect 259312 328442 259364 328448
rect 259772 328500 259824 328506
rect 259772 328442 259824 328448
rect 259128 321632 259180 321638
rect 259128 321574 259180 321580
rect 259324 309126 259352 328442
rect 259312 309120 259364 309126
rect 259312 309062 259364 309068
rect 259404 299532 259456 299538
rect 259404 299474 259456 299480
rect 259416 289814 259444 299474
rect 259404 289808 259456 289814
rect 259404 289750 259456 289756
rect 259404 280288 259456 280294
rect 259404 280230 259456 280236
rect 259416 273358 259444 280230
rect 259404 273352 259456 273358
rect 259404 273294 259456 273300
rect 259312 270564 259364 270570
rect 259312 270506 259364 270512
rect 259324 263650 259352 270506
rect 259232 263622 259352 263650
rect 259232 263514 259260 263622
rect 259232 263486 259352 263514
rect 259324 244338 259352 263486
rect 259232 244310 259352 244338
rect 259232 244202 259260 244310
rect 259232 244174 259352 244202
rect 259324 225026 259352 244174
rect 259232 224998 259352 225026
rect 259232 224890 259260 224998
rect 259232 224862 259352 224890
rect 259324 205714 259352 224862
rect 259232 205686 259352 205714
rect 259232 205578 259260 205686
rect 259232 205550 259352 205578
rect 259324 186402 259352 205550
rect 259232 186374 259352 186402
rect 259232 186266 259260 186374
rect 259232 186238 259352 186266
rect 259324 167090 259352 186238
rect 259864 179444 259916 179450
rect 259864 179386 259916 179392
rect 259876 179353 259904 179386
rect 259862 179344 259918 179353
rect 259862 179279 259918 179288
rect 259232 167062 259352 167090
rect 259232 166954 259260 167062
rect 259232 166926 259352 166954
rect 259324 164218 259352 166926
rect 259312 164212 259364 164218
rect 259312 164154 259364 164160
rect 259312 157344 259364 157350
rect 259312 157286 259364 157292
rect 259324 154578 259352 157286
rect 259324 154550 259444 154578
rect 259416 147642 259444 154550
rect 259324 147614 259444 147642
rect 259324 138038 259352 147614
rect 259312 138032 259364 138038
rect 259312 137974 259364 137980
rect 259404 137828 259456 137834
rect 259404 137770 259456 137776
rect 259416 135250 259444 137770
rect 259404 135244 259456 135250
rect 259404 135186 259456 135192
rect 259404 128308 259456 128314
rect 259404 128250 259456 128256
rect 259416 125610 259444 128250
rect 259416 125582 259536 125610
rect 259508 116006 259536 125582
rect 259312 116000 259364 116006
rect 259312 115942 259364 115948
rect 259496 116000 259548 116006
rect 259496 115942 259548 115948
rect 259324 89842 259352 115942
rect 259232 89814 259352 89842
rect 259232 89706 259260 89814
rect 259232 89678 259352 89706
rect 259324 70394 259352 89678
rect 259232 70366 259352 70394
rect 259232 70258 259260 70366
rect 259232 70230 259352 70258
rect 259324 51082 259352 70230
rect 259232 51066 259352 51082
rect 259220 51060 259352 51066
rect 259272 51054 259352 51060
rect 259404 51060 259456 51066
rect 259220 51002 259272 51008
rect 259404 51002 259456 51008
rect 259232 50971 259260 51002
rect 259416 48278 259444 51002
rect 259404 48272 259456 48278
rect 259404 48214 259456 48220
rect 259312 38752 259364 38758
rect 259312 38694 259364 38700
rect 259324 31770 259352 38694
rect 259232 31742 259352 31770
rect 259232 31634 259260 31742
rect 259232 31606 259352 31634
rect 259324 12458 259352 31606
rect 259232 12430 259352 12458
rect 259036 9512 259088 9518
rect 259036 9454 259088 9460
rect 259232 9450 259260 12430
rect 259220 9444 259272 9450
rect 259220 9386 259272 9392
rect 260060 7478 260088 335718
rect 260152 333266 260180 340068
rect 260232 335572 260284 335578
rect 260232 335514 260284 335520
rect 260140 333260 260192 333266
rect 260140 333202 260192 333208
rect 260244 312662 260272 335514
rect 260232 312656 260284 312662
rect 260232 312598 260284 312604
rect 260336 7546 260364 340068
rect 260428 340054 260626 340082
rect 260704 340054 260810 340082
rect 260888 340054 261086 340082
rect 260428 8838 260456 340054
rect 260704 335578 260732 340054
rect 260888 335782 260916 340054
rect 261244 337068 261296 337074
rect 261244 337010 261296 337016
rect 260876 335776 260928 335782
rect 260876 335718 260928 335724
rect 260692 335572 260744 335578
rect 260692 335514 260744 335520
rect 261256 320686 261284 337010
rect 261348 334506 261376 340068
rect 261532 334694 261560 340068
rect 261704 335572 261756 335578
rect 261704 335514 261756 335520
rect 261520 334688 261572 334694
rect 261520 334630 261572 334636
rect 261348 334478 261652 334506
rect 261244 320680 261296 320686
rect 261244 320622 261296 320628
rect 261152 320544 261204 320550
rect 261152 320486 261204 320492
rect 261164 320362 261192 320486
rect 261242 320376 261298 320385
rect 261164 320334 261242 320362
rect 261242 320311 261298 320320
rect 261244 320272 261296 320278
rect 261244 320214 261296 320220
rect 261150 242040 261206 242049
rect 261150 241975 261206 241984
rect 261164 241806 261192 241975
rect 261152 241800 261204 241806
rect 261152 241742 261204 241748
rect 261150 179752 261206 179761
rect 261150 179687 261206 179696
rect 261164 179353 261192 179687
rect 261150 179344 261206 179353
rect 261150 179279 261206 179288
rect 261150 101144 261206 101153
rect 261150 101079 261206 101088
rect 261164 100910 261192 101079
rect 261152 100904 261204 100910
rect 261152 100846 261204 100852
rect 261060 38752 261112 38758
rect 261058 38720 261060 38729
rect 261112 38720 261114 38729
rect 261058 38655 261114 38664
rect 260416 8832 260468 8838
rect 260416 8774 260468 8780
rect 260324 7540 260376 7546
rect 260324 7482 260376 7488
rect 260048 7472 260100 7478
rect 260048 7414 260100 7420
rect 259954 7168 260010 7177
rect 259954 7103 260010 7112
rect 259968 6769 259996 7103
rect 259954 6760 260010 6769
rect 259954 6695 260010 6704
rect 257746 5536 257802 5545
rect 257746 5471 257802 5480
rect 257286 5400 257342 5409
rect 257286 5335 257342 5344
rect 259128 4752 259180 4758
rect 259128 4694 259180 4700
rect 257932 3392 257984 3398
rect 257932 3334 257984 3340
rect 256736 604 256788 610
rect 255552 480 255580 598
rect 256736 546 256788 552
rect 257104 604 257156 610
rect 257104 546 257156 552
rect 256748 480 256776 546
rect 257944 480 257972 3334
rect 259140 480 259168 4694
rect 261256 4146 261284 320214
rect 261624 9586 261652 334478
rect 261612 9580 261664 9586
rect 261612 9522 261664 9528
rect 261716 7342 261744 335514
rect 261808 7410 261836 340068
rect 261900 340054 262098 340082
rect 261900 8906 261928 340054
rect 262268 335594 262296 340068
rect 262084 335566 262296 335594
rect 262360 340054 262558 340082
rect 262360 335578 262388 340054
rect 262348 335572 262400 335578
rect 262084 330614 262112 335566
rect 262348 335514 262400 335520
rect 262624 333260 262676 333266
rect 262624 333202 262676 333208
rect 262072 330608 262124 330614
rect 262072 330550 262124 330556
rect 261888 8900 261940 8906
rect 261888 8842 261940 8848
rect 261796 7404 261848 7410
rect 261796 7346 261848 7352
rect 261704 7336 261756 7342
rect 261704 7278 261756 7284
rect 260324 4140 260376 4146
rect 260324 4082 260376 4088
rect 261244 4140 261296 4146
rect 261244 4082 261296 4088
rect 260336 480 260364 4082
rect 262636 3466 262664 333202
rect 262820 9654 262848 340068
rect 263018 340054 263124 340082
rect 262900 335572 262952 335578
rect 262900 335514 262952 335520
rect 262808 9648 262860 9654
rect 262808 9590 262860 9596
rect 262912 9518 262940 335514
rect 263096 307154 263124 340054
rect 263176 334960 263228 334966
rect 263176 334902 263228 334908
rect 263084 307148 263136 307154
rect 263084 307090 263136 307096
rect 262900 9512 262952 9518
rect 262900 9454 262952 9460
rect 263188 6458 263216 334902
rect 263280 7274 263308 340068
rect 263372 340054 263570 340082
rect 263372 335578 263400 340054
rect 263360 335572 263412 335578
rect 263360 335514 263412 335520
rect 263740 333334 263768 340068
rect 263832 340054 264030 340082
rect 263832 334966 263860 340054
rect 264188 335776 264240 335782
rect 264188 335718 264240 335724
rect 264096 335572 264148 335578
rect 264096 335514 264148 335520
rect 263820 334960 263872 334966
rect 263820 334902 263872 334908
rect 263728 333328 263780 333334
rect 263728 333270 263780 333276
rect 264108 330682 264136 335514
rect 264096 330676 264148 330682
rect 264096 330618 264148 330624
rect 263268 7268 263320 7274
rect 263268 7210 263320 7216
rect 264200 7002 264228 335718
rect 264292 7206 264320 340068
rect 264384 340054 264490 340082
rect 264568 340054 264766 340082
rect 264844 340054 265042 340082
rect 265120 340054 265226 340082
rect 265502 340054 265608 340082
rect 264384 335578 264412 340054
rect 264372 335572 264424 335578
rect 264372 335514 264424 335520
rect 264372 335436 264424 335442
rect 264372 335378 264424 335384
rect 264384 327826 264412 335378
rect 264372 327820 264424 327826
rect 264372 327762 264424 327768
rect 264280 7200 264332 7206
rect 264280 7142 264332 7148
rect 264188 6996 264240 7002
rect 264188 6938 264240 6944
rect 264568 6662 264596 340054
rect 264740 337748 264792 337754
rect 264740 337690 264792 337696
rect 264752 14550 264780 337690
rect 264844 335782 264872 340054
rect 264832 335776 264884 335782
rect 264832 335718 264884 335724
rect 265120 335442 265148 340054
rect 265108 335436 265160 335442
rect 265108 335378 265160 335384
rect 264740 14544 264792 14550
rect 264740 14486 264792 14492
rect 265580 6730 265608 340054
rect 265660 335776 265712 335782
rect 265660 335718 265712 335724
rect 265672 7750 265700 335718
rect 265660 7744 265712 7750
rect 265660 7686 265712 7692
rect 265764 6934 265792 340068
rect 265844 335572 265896 335578
rect 265844 335514 265896 335520
rect 265856 322318 265884 335514
rect 265948 325038 265976 340068
rect 266040 340054 266238 340082
rect 266316 340054 266514 340082
rect 266592 340054 266698 340082
rect 265936 325032 265988 325038
rect 265936 324974 265988 324980
rect 265844 322312 265896 322318
rect 265844 322254 265896 322260
rect 265752 6928 265804 6934
rect 265752 6870 265804 6876
rect 266040 6798 266068 340054
rect 266316 335782 266344 340054
rect 266304 335776 266356 335782
rect 266304 335718 266356 335724
rect 266592 335578 266620 340054
rect 266580 335572 266632 335578
rect 266580 335514 266632 335520
rect 266960 6866 266988 340068
rect 267052 340054 267250 340082
rect 267052 7818 267080 340054
rect 267420 336122 267448 340068
rect 267604 340054 267710 340082
rect 267788 340054 267986 340082
rect 267408 336116 267460 336122
rect 267408 336058 267460 336064
rect 267604 335594 267632 340054
rect 267132 335572 267184 335578
rect 267132 335514 267184 335520
rect 267328 335566 267632 335594
rect 267788 335578 267816 340054
rect 267776 335572 267828 335578
rect 267144 297498 267172 335514
rect 267132 297492 267184 297498
rect 267132 297434 267184 297440
rect 267040 7812 267092 7818
rect 267040 7754 267092 7760
rect 266948 6860 267000 6866
rect 266948 6802 267000 6808
rect 266028 6792 266080 6798
rect 266028 6734 266080 6740
rect 265568 6724 265620 6730
rect 265568 6666 265620 6672
rect 264556 6656 264608 6662
rect 264556 6598 264608 6604
rect 263176 6452 263228 6458
rect 263176 6394 263228 6400
rect 264004 6316 264056 6322
rect 264004 6258 264056 6264
rect 264016 5302 264044 6258
rect 267328 6118 267356 335566
rect 267776 335514 267828 335520
rect 268156 335458 268184 340068
rect 268236 339108 268288 339114
rect 268236 339050 268288 339056
rect 267604 335430 268184 335458
rect 267604 319530 267632 335430
rect 268248 326534 268276 339050
rect 268432 336002 268460 340068
rect 268708 339114 268736 340068
rect 268696 339108 268748 339114
rect 268696 339050 268748 339056
rect 268432 335974 268644 336002
rect 268328 335776 268380 335782
rect 268616 335730 268644 335974
rect 268328 335718 268380 335724
rect 268236 326528 268288 326534
rect 268236 326470 268288 326476
rect 267592 319524 267644 319530
rect 267592 319466 267644 319472
rect 268144 38752 268196 38758
rect 268142 38720 268144 38729
rect 268196 38720 268198 38729
rect 268142 38655 268198 38664
rect 267316 6112 267368 6118
rect 267316 6054 267368 6060
rect 268340 5846 268368 335718
rect 268432 335702 268644 335730
rect 268432 5914 268460 335702
rect 268512 335572 268564 335578
rect 268512 335514 268564 335520
rect 268524 309806 268552 335514
rect 268892 333282 268920 340068
rect 268984 340054 269182 340082
rect 269260 340054 269458 340082
rect 269642 340054 269748 340082
rect 268984 335782 269012 340054
rect 268972 335776 269024 335782
rect 268972 335718 269024 335724
rect 269260 335578 269288 340054
rect 269248 335572 269300 335578
rect 269248 335514 269300 335520
rect 268616 333254 268920 333282
rect 268616 328438 268644 333254
rect 268604 328432 268656 328438
rect 268604 328374 268656 328380
rect 268696 321428 268748 321434
rect 268696 321370 268748 321376
rect 268708 311982 268736 321370
rect 268696 311976 268748 311982
rect 268696 311918 268748 311924
rect 268696 311636 268748 311642
rect 268696 311578 268748 311584
rect 268512 309800 268564 309806
rect 268512 309742 268564 309748
rect 268708 292534 268736 311578
rect 268696 292528 268748 292534
rect 268696 292470 268748 292476
rect 268696 292392 268748 292398
rect 268696 292334 268748 292340
rect 268708 284986 268736 292334
rect 268696 284980 268748 284986
rect 268696 284922 268748 284928
rect 268788 282804 268840 282810
rect 268788 282746 268840 282752
rect 268800 278746 268828 282746
rect 268708 278718 268828 278746
rect 268708 269142 268736 278718
rect 268604 269136 268656 269142
rect 268604 269078 268656 269084
rect 268696 269136 268748 269142
rect 268696 269078 268748 269084
rect 268616 263514 268644 269078
rect 268616 263486 268828 263514
rect 268800 253722 268828 263486
rect 268708 253694 268828 253722
rect 268708 227050 268736 253694
rect 268696 227044 268748 227050
rect 268696 226986 268748 226992
rect 268788 222216 268840 222222
rect 268788 222158 268840 222164
rect 268800 212650 268828 222158
rect 268708 212622 268828 212650
rect 268708 207738 268736 212622
rect 268696 207732 268748 207738
rect 268696 207674 268748 207680
rect 268788 205556 268840 205562
rect 268788 205498 268840 205504
rect 268800 201482 268828 205498
rect 268512 201476 268564 201482
rect 268512 201418 268564 201424
rect 268788 201476 268840 201482
rect 268788 201418 268840 201424
rect 268524 191865 268552 201418
rect 268510 191856 268566 191865
rect 268510 191791 268566 191800
rect 268694 191856 268750 191865
rect 268694 191791 268750 191800
rect 268708 183569 268736 191791
rect 268510 183560 268566 183569
rect 268510 183495 268566 183504
rect 268694 183560 268750 183569
rect 268694 183495 268750 183504
rect 268524 173942 268552 183495
rect 268512 173936 268564 173942
rect 268512 173878 268564 173884
rect 268696 173936 268748 173942
rect 268696 173878 268748 173884
rect 268708 166954 268736 173878
rect 268524 166926 268736 166954
rect 268524 161294 268552 166926
rect 268512 161288 268564 161294
rect 268512 161230 268564 161236
rect 268696 157140 268748 157146
rect 268696 157082 268748 157088
rect 268708 154426 268736 157082
rect 268696 154420 268748 154426
rect 268696 154362 268748 154368
rect 268696 147620 268748 147626
rect 268696 147562 268748 147568
rect 268708 144922 268736 147562
rect 268708 144894 268828 144922
rect 268800 138038 268828 144894
rect 268788 138032 268840 138038
rect 268788 137974 268840 137980
rect 268696 137964 268748 137970
rect 268696 137906 268748 137912
rect 268708 135250 268736 137906
rect 268696 135244 268748 135250
rect 268696 135186 268748 135192
rect 268696 128308 268748 128314
rect 268696 128250 268748 128256
rect 268708 125610 268736 128250
rect 268708 125582 268828 125610
rect 268800 115954 268828 125582
rect 268708 115926 268828 115954
rect 268708 99414 268736 115926
rect 268696 99408 268748 99414
rect 268696 99350 268748 99356
rect 268696 99272 268748 99278
rect 268696 99214 268748 99220
rect 268708 96626 268736 99214
rect 268696 96620 268748 96626
rect 268696 96562 268748 96568
rect 268696 89684 268748 89690
rect 268696 89626 268748 89632
rect 268708 86986 268736 89626
rect 268708 86958 268828 86986
rect 268800 79914 268828 86958
rect 268708 79886 268828 79914
rect 268708 52562 268736 79886
rect 268604 52556 268656 52562
rect 268604 52498 268656 52504
rect 268696 52556 268748 52562
rect 268696 52498 268748 52504
rect 268616 42786 268644 52498
rect 268616 42758 268828 42786
rect 268800 41290 268828 42758
rect 268708 41262 268828 41290
rect 268420 5908 268472 5914
rect 268420 5850 268472 5856
rect 268328 5840 268380 5846
rect 268328 5782 268380 5788
rect 264004 5296 264056 5302
rect 264004 5238 264056 5244
rect 268708 4865 268736 41262
rect 269522 7032 269578 7041
rect 269522 6967 269578 6976
rect 269536 6769 269564 6967
rect 269522 6760 269578 6769
rect 269522 6695 269578 6704
rect 268694 4856 268750 4865
rect 268694 4791 268750 4800
rect 264280 4616 264332 4622
rect 264280 4558 264332 4564
rect 264370 4584 264426 4593
rect 264292 4486 264320 4558
rect 269720 4554 269748 340054
rect 269800 335776 269852 335782
rect 269800 335718 269852 335724
rect 269812 5710 269840 335718
rect 269904 5778 269932 340068
rect 269984 335572 270036 335578
rect 269984 335514 270036 335520
rect 269996 318170 270024 335514
rect 270076 335504 270128 335510
rect 270076 335446 270128 335452
rect 269984 318164 270036 318170
rect 269984 318106 270036 318112
rect 270088 6390 270116 335446
rect 270180 323610 270208 340068
rect 270272 340054 270378 340082
rect 270456 340054 270654 340082
rect 270732 340054 270930 340082
rect 271008 340054 271114 340082
rect 271284 340054 271390 340082
rect 270272 335510 270300 340054
rect 270456 335782 270484 340054
rect 270444 335776 270496 335782
rect 270444 335718 270496 335724
rect 270732 335578 270760 340054
rect 270720 335572 270772 335578
rect 270720 335514 270772 335520
rect 270260 335504 270312 335510
rect 270260 335446 270312 335452
rect 270168 323604 270220 323610
rect 270168 323546 270220 323552
rect 270902 226672 270958 226681
rect 270902 226607 270958 226616
rect 270916 226273 270944 226607
rect 270902 226264 270958 226273
rect 270902 226199 270958 226208
rect 270076 6384 270128 6390
rect 270076 6326 270128 6332
rect 269892 5772 269944 5778
rect 269892 5714 269944 5720
rect 269800 5704 269852 5710
rect 269800 5646 269852 5652
rect 269798 4584 269854 4593
rect 264370 4519 264372 4528
rect 264424 4519 264426 4528
rect 269708 4548 269760 4554
rect 264372 4490 264424 4496
rect 269798 4519 269800 4528
rect 269708 4490 269760 4496
rect 269852 4519 269854 4528
rect 269800 4490 269852 4496
rect 271008 4486 271036 340054
rect 271180 335776 271232 335782
rect 271180 335718 271232 335724
rect 271192 5574 271220 335718
rect 271284 5642 271312 340054
rect 271364 331084 271416 331090
rect 271364 331026 271416 331032
rect 271376 316010 271404 331026
rect 271376 315982 271496 316010
rect 271468 304994 271496 315982
rect 271652 315382 271680 340068
rect 271744 340054 271850 340082
rect 271928 340054 272126 340082
rect 271744 331090 271772 340054
rect 271928 335782 271956 340054
rect 271916 335776 271968 335782
rect 271916 335718 271968 335724
rect 272388 333402 272416 340068
rect 272480 340054 272586 340082
rect 272862 340054 272968 340082
rect 272376 333396 272428 333402
rect 272376 333338 272428 333344
rect 271732 331084 271784 331090
rect 271732 331026 271784 331032
rect 271640 315376 271692 315382
rect 271640 315318 271692 315324
rect 271376 304966 271496 304994
rect 271376 299538 271404 304966
rect 271364 299532 271416 299538
rect 271364 299474 271416 299480
rect 271456 299396 271508 299402
rect 271456 299338 271508 299344
rect 271468 283082 271496 299338
rect 271456 283076 271508 283082
rect 271456 283018 271508 283024
rect 271456 282804 271508 282810
rect 271456 282746 271508 282752
rect 271468 270450 271496 282746
rect 271468 270422 271588 270450
rect 271560 256034 271588 270422
rect 271468 256006 271588 256034
rect 271468 244338 271496 256006
rect 271376 244310 271496 244338
rect 271376 244202 271404 244310
rect 271376 244174 271496 244202
rect 271468 225026 271496 244174
rect 271376 224998 271496 225026
rect 271376 224942 271404 224998
rect 271364 224936 271416 224942
rect 271364 224878 271416 224884
rect 271548 224936 271600 224942
rect 271548 224878 271600 224884
rect 271560 217410 271588 224878
rect 271468 217382 271588 217410
rect 271468 205766 271496 217382
rect 271456 205760 271508 205766
rect 271456 205702 271508 205708
rect 271456 205556 271508 205562
rect 271456 205498 271508 205504
rect 271468 167090 271496 205498
rect 271376 167062 271496 167090
rect 271376 166954 271404 167062
rect 271376 166926 271588 166954
rect 271560 149190 271588 166926
rect 271456 149184 271508 149190
rect 271456 149126 271508 149132
rect 271548 149184 271600 149190
rect 271548 149126 271600 149132
rect 271468 149002 271496 149126
rect 271468 148974 271588 149002
rect 271560 139466 271588 148974
rect 271456 139460 271508 139466
rect 271456 139402 271508 139408
rect 271548 139460 271600 139466
rect 271548 139402 271600 139408
rect 271468 137970 271496 139402
rect 271456 137964 271508 137970
rect 271456 137906 271508 137912
rect 271456 128512 271508 128518
rect 271456 128454 271508 128460
rect 271468 125746 271496 128454
rect 271468 125718 271588 125746
rect 271560 124930 271588 125718
rect 271376 124902 271588 124930
rect 271376 109041 271404 124902
rect 271362 109032 271418 109041
rect 271362 108967 271418 108976
rect 271638 109032 271694 109041
rect 271638 108967 271694 108976
rect 271652 99414 271680 108967
rect 271456 99408 271508 99414
rect 271456 99350 271508 99356
rect 271640 99408 271692 99414
rect 271640 99350 271692 99356
rect 271468 81530 271496 99350
rect 271456 81524 271508 81530
rect 271456 81466 271508 81472
rect 271364 80096 271416 80102
rect 271364 80038 271416 80044
rect 271376 76634 271404 80038
rect 271364 76628 271416 76634
rect 271364 76570 271416 76576
rect 271456 63572 271508 63578
rect 271456 63514 271508 63520
rect 271468 51082 271496 63514
rect 271376 51066 271496 51082
rect 271364 51060 271496 51066
rect 271416 51054 271496 51060
rect 271548 51060 271600 51066
rect 271364 51002 271416 51008
rect 271548 51002 271600 51008
rect 271376 50971 271404 51002
rect 271560 37330 271588 51002
rect 271456 37324 271508 37330
rect 271456 37266 271508 37272
rect 271548 37324 271600 37330
rect 271548 37266 271600 37272
rect 271468 18034 271496 37266
rect 271376 18006 271496 18034
rect 271376 9738 271404 18006
rect 271376 9710 271588 9738
rect 271560 9602 271588 9710
rect 271376 9574 271588 9602
rect 271272 5636 271324 5642
rect 271272 5578 271324 5584
rect 271180 5568 271232 5574
rect 271180 5510 271232 5516
rect 264188 4480 264240 4486
rect 264186 4448 264188 4457
rect 264280 4480 264332 4486
rect 264240 4448 264242 4457
rect 264280 4422 264332 4428
rect 270996 4480 271048 4486
rect 270996 4422 271048 4428
rect 264186 4383 264242 4392
rect 271376 4214 271404 9574
rect 272480 4554 272508 340054
rect 272652 338496 272704 338502
rect 272652 338438 272704 338444
rect 272664 335594 272692 338438
rect 272940 336818 272968 340054
rect 273124 338502 273152 340068
rect 273112 338496 273164 338502
rect 273112 338438 273164 338444
rect 273308 336977 273336 340068
rect 273294 336968 273350 336977
rect 273294 336903 273350 336912
rect 272572 335566 272692 335594
rect 272848 336790 272968 336818
rect 273294 336832 273350 336841
rect 272572 321638 272600 335566
rect 272652 335504 272704 335510
rect 272652 335446 272704 335452
rect 272560 321632 272612 321638
rect 272560 321574 272612 321580
rect 272560 304972 272612 304978
rect 272560 304914 272612 304920
rect 272572 298790 272600 304914
rect 272560 298784 272612 298790
rect 272560 298726 272612 298732
rect 272664 295594 272692 335446
rect 272744 321632 272796 321638
rect 272744 321574 272796 321580
rect 272652 295588 272704 295594
rect 272652 295530 272704 295536
rect 272756 295526 272784 321574
rect 272848 316010 272876 336790
rect 273294 336767 273350 336776
rect 273308 333985 273336 336767
rect 273400 335510 273428 340190
rect 273874 340054 273980 340082
rect 274058 340054 274256 340082
rect 273756 335776 273808 335782
rect 273756 335718 273808 335724
rect 273388 335504 273440 335510
rect 273388 335446 273440 335452
rect 272926 333976 272982 333985
rect 272926 333911 272982 333920
rect 273294 333976 273350 333985
rect 273294 333911 273350 333920
rect 272940 324358 272968 333911
rect 273768 327894 273796 335718
rect 273756 327888 273808 327894
rect 273756 327830 273808 327836
rect 272928 324352 272980 324358
rect 272928 324294 272980 324300
rect 273020 324352 273072 324358
rect 273020 324294 273072 324300
rect 273032 316010 273060 324294
rect 272848 315982 272968 316010
rect 273032 315982 273152 316010
rect 272940 304994 272968 315982
rect 273124 304994 273152 315982
rect 272848 304978 272968 304994
rect 273032 304978 273152 304994
rect 272836 304972 272968 304978
rect 272888 304966 272968 304972
rect 273020 304972 273152 304978
rect 272836 304914 272888 304920
rect 273072 304966 273152 304972
rect 273204 304972 273256 304978
rect 273020 304914 273072 304920
rect 273204 304914 273256 304920
rect 272848 304883 272876 304914
rect 273032 304883 273060 304914
rect 272928 298784 272980 298790
rect 272928 298726 272980 298732
rect 272744 295520 272796 295526
rect 272744 295462 272796 295468
rect 272744 295316 272796 295322
rect 272744 295258 272796 295264
rect 272652 295248 272704 295254
rect 272652 295190 272704 295196
rect 272664 6254 272692 295190
rect 272756 8634 272784 295258
rect 272940 295202 272968 298726
rect 273216 295361 273244 304914
rect 273018 295352 273074 295361
rect 273018 295287 273074 295296
rect 273202 295352 273258 295361
rect 273202 295287 273258 295296
rect 272848 295174 272968 295202
rect 272848 284306 272876 295174
rect 272836 284300 272888 284306
rect 272836 284242 272888 284248
rect 272928 284300 272980 284306
rect 272928 284242 272980 284248
rect 272940 274825 272968 284242
rect 273032 276010 273060 295287
rect 273020 276004 273072 276010
rect 273020 275946 273072 275952
rect 273112 276004 273164 276010
rect 273112 275946 273164 275952
rect 272926 274816 272982 274825
rect 272926 274751 272982 274760
rect 272834 274680 272890 274689
rect 272834 274615 272836 274624
rect 272888 274615 272890 274624
rect 273020 274644 273072 274650
rect 272836 274586 272888 274592
rect 273020 274586 273072 274592
rect 273032 265033 273060 274586
rect 272834 265024 272890 265033
rect 272834 264959 272890 264968
rect 273018 265024 273074 265033
rect 273018 264959 273074 264968
rect 272848 235958 272876 264959
rect 273124 264874 273152 275946
rect 273032 264846 273152 264874
rect 273032 256902 273060 264846
rect 273020 256896 273072 256902
rect 273020 256838 273072 256844
rect 273020 255332 273072 255338
rect 273020 255274 273072 255280
rect 273032 253910 273060 255274
rect 273020 253904 273072 253910
rect 273020 253846 273072 253852
rect 273020 236020 273072 236026
rect 273020 235962 273072 235968
rect 272836 235952 272888 235958
rect 272836 235894 272888 235900
rect 272928 231600 272980 231606
rect 272928 231542 272980 231548
rect 272940 224942 272968 231542
rect 273032 227066 273060 235962
rect 273032 227038 273244 227066
rect 272928 224936 272980 224942
rect 273216 224890 273244 227038
rect 272928 224878 272980 224884
rect 273124 224862 273244 224890
rect 272928 218000 272980 218006
rect 272928 217942 272980 217948
rect 272940 215370 272968 217942
rect 272848 215342 272968 215370
rect 272848 215286 272876 215342
rect 272836 215280 272888 215286
rect 272836 215222 272888 215228
rect 273124 211154 273152 224862
rect 273032 211126 273152 211154
rect 272836 210452 272888 210458
rect 272836 210394 272888 210400
rect 272848 197282 272876 210394
rect 273032 206990 273060 211126
rect 273020 206984 273072 206990
rect 273020 206926 273072 206932
rect 273112 206916 273164 206922
rect 273112 206858 273164 206864
rect 272848 197254 272968 197282
rect 272940 189106 272968 197254
rect 272928 189100 272980 189106
rect 272928 189042 272980 189048
rect 272928 188964 272980 188970
rect 272928 188906 272980 188912
rect 272940 179330 272968 188906
rect 273124 187762 273152 206858
rect 273032 187734 273152 187762
rect 273032 180810 273060 187734
rect 273020 180804 273072 180810
rect 273020 180746 273072 180752
rect 273112 180804 273164 180810
rect 273112 180746 273164 180752
rect 272848 179302 272968 179330
rect 272848 171034 272876 179302
rect 272848 171006 273060 171034
rect 273032 167770 273060 171006
rect 273124 168366 273152 180746
rect 273112 168360 273164 168366
rect 273112 168302 273164 168308
rect 272940 167742 273060 167770
rect 272940 166326 272968 167742
rect 272928 166320 272980 166326
rect 272928 166262 272980 166268
rect 272836 166252 272888 166258
rect 272836 166194 272888 166200
rect 272848 121446 272876 166194
rect 273020 163532 273072 163538
rect 273020 163474 273072 163480
rect 273032 158710 273060 163474
rect 273020 158704 273072 158710
rect 273020 158646 273072 158652
rect 273112 158704 273164 158710
rect 273112 158646 273164 158652
rect 273124 157350 273152 158646
rect 273112 157344 273164 157350
rect 273112 157286 273164 157292
rect 273020 147688 273072 147694
rect 273020 147630 273072 147636
rect 273032 143750 273060 147630
rect 273020 143744 273072 143750
rect 273020 143686 273072 143692
rect 273020 139460 273072 139466
rect 273020 139402 273072 139408
rect 273032 134586 273060 139402
rect 273032 134558 273152 134586
rect 273124 121446 273152 134558
rect 272836 121440 272888 121446
rect 272836 121382 272888 121388
rect 273020 121440 273072 121446
rect 273020 121382 273072 121388
rect 273112 121440 273164 121446
rect 273112 121382 273164 121388
rect 272836 111852 272888 111858
rect 272836 111794 272888 111800
rect 272848 57934 272876 111794
rect 273032 98682 273060 121382
rect 273032 98654 273152 98682
rect 273124 62150 273152 98654
rect 273020 62144 273072 62150
rect 273020 62086 273072 62092
rect 273112 62144 273164 62150
rect 273112 62086 273164 62092
rect 272836 57928 272888 57934
rect 272836 57870 272888 57876
rect 273032 57338 273060 62086
rect 272940 57310 273060 57338
rect 272940 52465 272968 57310
rect 272926 52456 272982 52465
rect 272926 52391 272982 52400
rect 273294 52456 273350 52465
rect 273294 52391 273350 52400
rect 272836 48340 272888 48346
rect 272836 48282 272888 48288
rect 272848 46918 272876 48282
rect 272836 46912 272888 46918
rect 272836 46854 272888 46860
rect 273308 42838 273336 52391
rect 273112 42832 273164 42838
rect 273112 42774 273164 42780
rect 273296 42832 273348 42838
rect 273296 42774 273348 42780
rect 273124 42702 273152 42774
rect 273112 42696 273164 42702
rect 273112 42638 273164 42644
rect 273020 42628 273072 42634
rect 273020 42570 273072 42576
rect 272836 37324 272888 37330
rect 272836 37266 272888 37272
rect 272848 27606 272876 37266
rect 273032 33289 273060 42570
rect 273018 33280 273074 33289
rect 273018 33215 273074 33224
rect 273202 33280 273258 33289
rect 273202 33215 273258 33224
rect 272836 27600 272888 27606
rect 272836 27542 272888 27548
rect 273216 18834 273244 33215
rect 273020 18828 273072 18834
rect 273020 18770 273072 18776
rect 273204 18828 273256 18834
rect 273204 18770 273256 18776
rect 272836 18080 272888 18086
rect 272836 18022 272888 18028
rect 272744 8628 272796 8634
rect 272744 8570 272796 8576
rect 272848 8294 272876 18022
rect 273032 11370 273060 18770
rect 272940 11342 273060 11370
rect 272836 8288 272888 8294
rect 272836 8230 272888 8236
rect 272652 6248 272704 6254
rect 272652 6190 272704 6196
rect 272468 4548 272520 4554
rect 272468 4490 272520 4496
rect 272940 4457 272968 11342
rect 273952 8566 273980 340054
rect 274124 335572 274176 335578
rect 274124 335514 274176 335520
rect 273940 8560 273992 8566
rect 273940 8502 273992 8508
rect 274136 4622 274164 335514
rect 274124 4616 274176 4622
rect 274124 4558 274176 4564
rect 272926 4448 272982 4457
rect 272926 4383 272982 4392
rect 274228 4282 274256 340054
rect 274320 332042 274348 340068
rect 274412 340054 274610 340082
rect 274688 340054 274794 340082
rect 274872 340054 275070 340082
rect 274308 332036 274360 332042
rect 274308 331978 274360 331984
rect 274412 8498 274440 340054
rect 274688 335578 274716 340054
rect 274872 335782 274900 340054
rect 275228 335912 275280 335918
rect 275228 335854 275280 335860
rect 275136 335844 275188 335850
rect 275136 335786 275188 335792
rect 274860 335776 274912 335782
rect 274860 335718 274912 335724
rect 274676 335572 274728 335578
rect 274676 335514 274728 335520
rect 275148 329254 275176 335786
rect 275136 329248 275188 329254
rect 275136 329190 275188 329196
rect 274400 8492 274452 8498
rect 274400 8434 274452 8440
rect 275240 4826 275268 335854
rect 275332 8430 275360 340068
rect 275424 340054 275530 340082
rect 275608 340054 275806 340082
rect 275884 340054 275990 340082
rect 276068 340054 276266 340082
rect 275424 335918 275452 340054
rect 275412 335912 275464 335918
rect 275412 335854 275464 335860
rect 275608 335850 275636 340054
rect 275596 335844 275648 335850
rect 275596 335786 275648 335792
rect 275884 335730 275912 340054
rect 275424 335702 275912 335730
rect 275320 8424 275372 8430
rect 275320 8366 275372 8372
rect 275424 8362 275452 335702
rect 276068 333962 276096 340054
rect 276148 336864 276200 336870
rect 276148 336806 276200 336812
rect 275976 333934 276096 333962
rect 275780 324420 275832 324426
rect 275780 324362 275832 324368
rect 275688 324352 275740 324358
rect 275502 324320 275558 324329
rect 275502 324255 275558 324264
rect 275686 324320 275688 324329
rect 275740 324320 275742 324329
rect 275686 324255 275742 324264
rect 275516 314702 275544 324255
rect 275504 314696 275556 314702
rect 275504 314638 275556 314644
rect 275688 314696 275740 314702
rect 275688 314638 275740 314644
rect 275700 305130 275728 314638
rect 275608 305102 275728 305130
rect 275608 304994 275636 305102
rect 275608 304966 275728 304994
rect 275700 299538 275728 304966
rect 275688 299532 275740 299538
rect 275688 299474 275740 299480
rect 275504 296948 275556 296954
rect 275504 296890 275556 296896
rect 275516 285274 275544 296890
rect 275516 285246 275636 285274
rect 275608 275346 275636 285246
rect 275608 275318 275728 275346
rect 275700 265690 275728 275318
rect 275608 265662 275728 265690
rect 275608 256034 275636 265662
rect 275608 256006 275728 256034
rect 275700 255270 275728 256006
rect 275688 255264 275740 255270
rect 275688 255206 275740 255212
rect 275596 245676 275648 245682
rect 275596 245618 275648 245624
rect 275608 236042 275636 245618
rect 275608 236014 275728 236042
rect 275700 234598 275728 236014
rect 275688 234592 275740 234598
rect 275688 234534 275740 234540
rect 275688 225004 275740 225010
rect 275688 224946 275740 224952
rect 275700 224874 275728 224946
rect 275688 224868 275740 224874
rect 275688 224810 275740 224816
rect 275596 215348 275648 215354
rect 275596 215290 275648 215296
rect 275608 211274 275636 215290
rect 275596 211268 275648 211274
rect 275596 211210 275648 211216
rect 275596 210452 275648 210458
rect 275596 210394 275648 210400
rect 275608 197606 275636 210394
rect 275596 197600 275648 197606
rect 275596 197542 275648 197548
rect 275688 197396 275740 197402
rect 275688 197338 275740 197344
rect 275700 197282 275728 197338
rect 275608 197254 275728 197282
rect 275608 187921 275636 197254
rect 275594 187912 275650 187921
rect 275594 187847 275650 187856
rect 275686 187776 275742 187785
rect 275686 187711 275742 187720
rect 275700 177970 275728 187711
rect 275608 177942 275728 177970
rect 275608 173262 275636 177942
rect 275596 173256 275648 173262
rect 275596 173198 275648 173204
rect 275596 163532 275648 163538
rect 275596 163474 275648 163480
rect 275608 157350 275636 163474
rect 275596 157344 275648 157350
rect 275596 157286 275648 157292
rect 275688 147688 275740 147694
rect 275688 147630 275740 147636
rect 275700 139602 275728 147630
rect 275504 139596 275556 139602
rect 275504 139538 275556 139544
rect 275688 139596 275740 139602
rect 275688 139538 275740 139544
rect 275516 129878 275544 139538
rect 275504 129872 275556 129878
rect 275504 129814 275556 129820
rect 275688 129872 275740 129878
rect 275688 129814 275740 129820
rect 275700 129742 275728 129814
rect 275596 129736 275648 129742
rect 275596 129678 275648 129684
rect 275688 129736 275740 129742
rect 275688 129678 275740 129684
rect 275608 120170 275636 129678
rect 275608 120142 275728 120170
rect 275700 118697 275728 120142
rect 275502 118688 275558 118697
rect 275502 118623 275558 118632
rect 275686 118688 275742 118697
rect 275686 118623 275742 118632
rect 275516 109070 275544 118623
rect 275504 109064 275556 109070
rect 275504 109006 275556 109012
rect 275596 109064 275648 109070
rect 275596 109006 275648 109012
rect 275608 106350 275636 109006
rect 275596 106344 275648 106350
rect 275596 106286 275648 106292
rect 275504 100768 275556 100774
rect 275504 100710 275556 100716
rect 275516 91118 275544 100710
rect 275504 91112 275556 91118
rect 275504 91054 275556 91060
rect 275688 91112 275740 91118
rect 275688 91054 275740 91060
rect 275700 73166 275728 91054
rect 275688 73160 275740 73166
rect 275688 73102 275740 73108
rect 275596 63572 275648 63578
rect 275596 63514 275648 63520
rect 275608 62778 275636 63514
rect 275516 62750 275636 62778
rect 275516 62506 275544 62750
rect 275516 62478 275728 62506
rect 275700 62098 275728 62478
rect 275608 62070 275728 62098
rect 275608 58002 275636 62070
rect 275596 57996 275648 58002
rect 275596 57938 275648 57944
rect 275596 52488 275648 52494
rect 275596 52430 275648 52436
rect 275608 46986 275636 52430
rect 275596 46980 275648 46986
rect 275596 46922 275648 46928
rect 275608 42838 275636 42869
rect 275596 42832 275648 42838
rect 275516 42780 275596 42786
rect 275516 42774 275648 42780
rect 275516 42758 275636 42774
rect 275516 38010 275544 42758
rect 275504 38004 275556 38010
rect 275504 37946 275556 37952
rect 275688 24880 275740 24886
rect 275688 24822 275740 24828
rect 275412 8356 275464 8362
rect 275412 8298 275464 8304
rect 275700 5098 275728 24822
rect 275792 18630 275820 324362
rect 275976 324358 276004 333934
rect 276160 324426 276188 336806
rect 276528 336326 276556 340068
rect 276620 340054 276726 340082
rect 276804 340054 277002 340082
rect 277080 340054 277278 340082
rect 277356 340054 277462 340082
rect 277540 340054 277738 340082
rect 277908 340054 278014 340082
rect 276516 336320 276568 336326
rect 276516 336262 276568 336268
rect 276516 335776 276568 335782
rect 276516 335718 276568 335724
rect 276528 333946 276556 335718
rect 276516 333940 276568 333946
rect 276516 333882 276568 333888
rect 276620 329474 276648 340054
rect 276804 335782 276832 340054
rect 276792 335776 276844 335782
rect 276792 335718 276844 335724
rect 277080 335594 277108 340054
rect 276792 335572 276844 335578
rect 276792 335514 276844 335520
rect 276896 335566 277108 335594
rect 277356 335578 277384 340054
rect 277344 335572 277396 335578
rect 276620 329446 276740 329474
rect 276148 324420 276200 324426
rect 276148 324362 276200 324368
rect 276608 324420 276660 324426
rect 276608 324362 276660 324368
rect 275964 324352 276016 324358
rect 275964 324294 276016 324300
rect 276620 304978 276648 324362
rect 276712 304978 276740 329446
rect 276608 304972 276660 304978
rect 276608 304914 276660 304920
rect 276700 304972 276752 304978
rect 276700 304914 276752 304920
rect 276514 295352 276570 295361
rect 276698 295352 276754 295361
rect 276570 295310 276648 295338
rect 276514 295287 276570 295296
rect 276620 295254 276648 295310
rect 276698 295287 276700 295296
rect 276752 295287 276754 295296
rect 276700 295258 276752 295264
rect 276608 295248 276660 295254
rect 276608 295190 276660 295196
rect 276608 285728 276660 285734
rect 276608 285670 276660 285676
rect 276620 232626 276648 285670
rect 276804 280498 276832 335514
rect 276896 325106 276924 335566
rect 277344 335514 277396 335520
rect 277540 335306 277568 340054
rect 277908 336818 277936 340054
rect 277632 336790 277936 336818
rect 277068 335300 277120 335306
rect 277068 335242 277120 335248
rect 277528 335300 277580 335306
rect 277528 335242 277580 335248
rect 276884 325100 276936 325106
rect 276884 325042 276936 325048
rect 277080 318918 277108 335242
rect 277632 335186 277660 336790
rect 278080 335572 278132 335578
rect 278080 335514 278132 335520
rect 277172 335158 277660 335186
rect 277068 318912 277120 318918
rect 277068 318854 277120 318860
rect 276976 318708 277028 318714
rect 276976 318650 277028 318656
rect 276988 311250 277016 318650
rect 276988 311222 277108 311250
rect 276976 304972 277028 304978
rect 276976 304914 277028 304920
rect 276988 295361 277016 304914
rect 276974 295352 277030 295361
rect 276974 295287 277030 295296
rect 276976 285728 277028 285734
rect 276976 285670 277028 285676
rect 276988 285190 277016 285670
rect 276976 285184 277028 285190
rect 276976 285126 277028 285132
rect 277080 285002 277108 311222
rect 276988 284974 277108 285002
rect 276792 280492 276844 280498
rect 276792 280434 276844 280440
rect 276792 280084 276844 280090
rect 276792 280026 276844 280032
rect 276700 280016 276752 280022
rect 276700 279958 276752 279964
rect 276712 237386 276740 279958
rect 276700 237380 276752 237386
rect 276700 237322 276752 237328
rect 276608 232620 276660 232626
rect 276608 232562 276660 232568
rect 276804 227905 276832 280026
rect 276988 275346 277016 284974
rect 276988 275318 277108 275346
rect 277080 265690 277108 275318
rect 276988 265662 277108 265690
rect 276988 256034 277016 265662
rect 276988 256006 277108 256034
rect 277080 246378 277108 256006
rect 276988 246350 277108 246378
rect 276988 241482 277016 246350
rect 276988 241454 277108 241482
rect 276884 237380 276936 237386
rect 276884 237322 276936 237328
rect 276790 227896 276846 227905
rect 276790 227831 276846 227840
rect 276516 227792 276568 227798
rect 276516 227734 276568 227740
rect 276790 227760 276846 227769
rect 276528 221513 276556 227734
rect 276790 227695 276846 227704
rect 276700 222216 276752 222222
rect 276700 222158 276752 222164
rect 276514 221504 276570 221513
rect 276514 221439 276570 221448
rect 276712 220794 276740 222158
rect 276700 220788 276752 220794
rect 276700 220730 276752 220736
rect 276700 211200 276752 211206
rect 276700 211142 276752 211148
rect 276514 208448 276570 208457
rect 276514 208383 276570 208392
rect 276528 208298 276556 208383
rect 276528 208270 276648 208298
rect 276620 198098 276648 208270
rect 276528 198070 276648 198098
rect 276528 193202 276556 198070
rect 276528 193174 276648 193202
rect 276620 178786 276648 193174
rect 276528 178758 276648 178786
rect 276528 173890 276556 178758
rect 276436 173862 276556 173890
rect 276436 164234 276464 173862
rect 276712 169538 276740 211142
rect 276620 169510 276740 169538
rect 276620 164370 276648 169510
rect 276804 169402 276832 227695
rect 276896 222222 276924 237322
rect 277080 232558 277108 241454
rect 277068 232552 277120 232558
rect 277068 232494 277120 232500
rect 276974 227760 277030 227769
rect 276974 227695 277030 227704
rect 276884 222216 276936 222222
rect 276884 222158 276936 222164
rect 276988 217410 277016 227695
rect 276988 217382 277108 217410
rect 277080 207754 277108 217382
rect 276988 207726 277108 207754
rect 276988 198150 277016 207726
rect 276976 198144 277028 198150
rect 276976 198086 277028 198092
rect 276976 189100 277028 189106
rect 276976 189042 277028 189048
rect 276988 183546 277016 189042
rect 276988 183518 277108 183546
rect 276712 169374 276832 169402
rect 276712 164529 276740 169374
rect 276698 164520 276754 164529
rect 276698 164455 276754 164464
rect 276790 164384 276846 164393
rect 276620 164342 276740 164370
rect 276436 164206 276648 164234
rect 276620 157434 276648 164206
rect 276528 157406 276648 157434
rect 276528 149682 276556 157406
rect 276528 149654 276648 149682
rect 276620 138122 276648 149654
rect 276712 143546 276740 164342
rect 276790 164319 276846 164328
rect 276700 143540 276752 143546
rect 276700 143482 276752 143488
rect 276528 138094 276648 138122
rect 276528 130370 276556 138094
rect 276698 133920 276754 133929
rect 276698 133855 276754 133864
rect 276528 130342 276648 130370
rect 276620 114730 276648 130342
rect 276528 114702 276648 114730
rect 276528 102218 276556 114702
rect 276528 102190 276648 102218
rect 276620 100722 276648 102190
rect 276528 100694 276648 100722
rect 276528 93906 276556 100694
rect 276516 93900 276568 93906
rect 276516 93842 276568 93848
rect 276608 93832 276660 93838
rect 276608 93774 276660 93780
rect 276620 82822 276648 93774
rect 276608 82816 276660 82822
rect 276608 82758 276660 82764
rect 276608 73228 276660 73234
rect 276608 73170 276660 73176
rect 276620 62121 276648 73170
rect 276422 62112 276478 62121
rect 276422 62047 276478 62056
rect 276606 62112 276662 62121
rect 276606 62047 276662 62056
rect 276436 57322 276464 62047
rect 276424 57316 276476 57322
rect 276424 57258 276476 57264
rect 276608 44192 276660 44198
rect 276608 44134 276660 44140
rect 276620 38010 276648 44134
rect 276240 38004 276292 38010
rect 276240 37946 276292 37952
rect 276608 38004 276660 38010
rect 276608 37946 276660 37952
rect 276252 27674 276280 37946
rect 276240 27668 276292 27674
rect 276240 27610 276292 27616
rect 276516 27668 276568 27674
rect 276516 27610 276568 27616
rect 275780 18624 275832 18630
rect 275780 18566 275832 18572
rect 276528 5166 276556 27610
rect 276712 8974 276740 133855
rect 276804 9042 276832 164319
rect 276884 143540 276936 143546
rect 276884 143482 276936 143488
rect 276896 133929 276924 143482
rect 276882 133920 276938 133929
rect 276882 133855 276938 133864
rect 277080 93820 277108 183518
rect 276988 93792 277108 93820
rect 276988 82958 277016 93792
rect 276976 82952 277028 82958
rect 276976 82894 277028 82900
rect 277068 82884 277120 82890
rect 277068 82826 277120 82832
rect 277080 71754 277108 82826
rect 276988 71726 277108 71754
rect 276988 67658 277016 71726
rect 276976 67652 277028 67658
rect 276976 67594 277028 67600
rect 277068 62756 277120 62762
rect 277068 62698 277120 62704
rect 277080 51048 277108 62698
rect 276988 51020 277108 51048
rect 276988 37330 277016 51020
rect 276976 37324 277028 37330
rect 276976 37266 277028 37272
rect 277068 37324 277120 37330
rect 277068 37266 277120 37272
rect 277080 22166 277108 37266
rect 277068 22160 277120 22166
rect 277068 22102 277120 22108
rect 276976 22092 277028 22098
rect 276976 22034 277028 22040
rect 276792 9036 276844 9042
rect 276792 8978 276844 8984
rect 276700 8968 276752 8974
rect 276700 8910 276752 8916
rect 276516 5160 276568 5166
rect 276516 5102 276568 5108
rect 275688 5092 275740 5098
rect 275688 5034 275740 5040
rect 276988 5030 277016 22034
rect 277172 17270 277200 335158
rect 277252 304904 277304 304910
rect 277252 304846 277304 304852
rect 277264 295497 277292 304846
rect 277250 295488 277306 295497
rect 277250 295423 277306 295432
rect 277252 232552 277304 232558
rect 277252 232494 277304 232500
rect 277264 227769 277292 232494
rect 277250 227760 277306 227769
rect 277250 227695 277306 227704
rect 277160 17264 277212 17270
rect 277160 17206 277212 17212
rect 278092 9178 278120 335514
rect 278080 9172 278132 9178
rect 278080 9114 278132 9120
rect 278184 9110 278212 340068
rect 278276 340054 278474 340082
rect 278172 9104 278224 9110
rect 278172 9046 278224 9052
rect 278276 5302 278304 340054
rect 278540 337136 278592 337142
rect 278540 337078 278592 337084
rect 278448 295316 278500 295322
rect 278448 295258 278500 295264
rect 278460 277545 278488 295258
rect 278446 277536 278502 277545
rect 278446 277471 278502 277480
rect 278446 277400 278502 277409
rect 278446 277335 278502 277344
rect 278460 270298 278488 277335
rect 278448 270292 278500 270298
rect 278448 270234 278500 270240
rect 278446 16552 278502 16561
rect 278446 16487 278502 16496
rect 278460 6934 278488 16487
rect 278448 6928 278500 6934
rect 278448 6870 278500 6876
rect 278264 5296 278316 5302
rect 278264 5238 278316 5244
rect 276976 5024 277028 5030
rect 276976 4966 277028 4972
rect 275228 4820 275280 4826
rect 275228 4762 275280 4768
rect 274216 4276 274268 4282
rect 274216 4218 274268 4224
rect 271364 4208 271416 4214
rect 271364 4150 271416 4156
rect 269800 4140 269852 4146
rect 269800 4082 269852 4088
rect 268604 4072 268656 4078
rect 268604 4014 268656 4020
rect 267500 4004 267552 4010
rect 267500 3946 267552 3952
rect 266304 3936 266356 3942
rect 266304 3878 266356 3884
rect 263912 3732 263964 3738
rect 263912 3674 263964 3680
rect 261520 3460 261572 3466
rect 261520 3402 261572 3408
rect 262624 3460 262676 3466
rect 262624 3402 262676 3408
rect 262728 3454 262940 3482
rect 261532 480 261560 3402
rect 262728 480 262756 3454
rect 262912 3398 262940 3454
rect 262900 3392 262952 3398
rect 262900 3334 262952 3340
rect 263924 480 263952 3674
rect 265108 3528 265160 3534
rect 265108 3470 265160 3476
rect 265120 480 265148 3470
rect 266316 480 266344 3878
rect 267512 480 267540 3946
rect 268616 480 268644 4014
rect 269812 480 269840 4082
rect 273388 3596 273440 3602
rect 273388 3538 273440 3544
rect 278448 3596 278500 3602
rect 278552 3584 278580 337078
rect 278736 336870 278764 340068
rect 278828 340054 278934 340082
rect 278724 336864 278776 336870
rect 278724 336806 278776 336812
rect 278828 335578 278856 340054
rect 279196 338502 279224 340068
rect 279486 340054 279592 340082
rect 278908 338496 278960 338502
rect 278908 338438 278960 338444
rect 279184 338496 279236 338502
rect 279184 338438 279236 338444
rect 278816 335572 278868 335578
rect 278816 335514 278868 335520
rect 278920 335322 278948 338438
rect 279276 335572 279328 335578
rect 279276 335514 279328 335520
rect 278828 335294 278948 335322
rect 278828 331974 278856 335294
rect 278816 331968 278868 331974
rect 278816 331910 278868 331916
rect 278724 326868 278776 326874
rect 278724 326810 278776 326816
rect 278736 316282 278764 326810
rect 278736 316254 278856 316282
rect 278828 316146 278856 316254
rect 278736 316118 278856 316146
rect 278736 306377 278764 316118
rect 278722 306368 278778 306377
rect 278722 306303 278778 306312
rect 278906 306368 278962 306377
rect 278906 306303 278962 306312
rect 278920 296750 278948 306303
rect 278724 296744 278776 296750
rect 278724 296686 278776 296692
rect 278908 296744 278960 296750
rect 278908 296686 278960 296692
rect 278736 295322 278764 296686
rect 278724 295316 278776 295322
rect 278724 295258 278776 295264
rect 278630 277536 278686 277545
rect 278630 277471 278686 277480
rect 278644 277409 278672 277471
rect 278630 277400 278686 277409
rect 278630 277335 278686 277344
rect 278816 270292 278868 270298
rect 278816 270234 278868 270240
rect 278828 267753 278856 270234
rect 278814 267744 278870 267753
rect 278814 267679 278870 267688
rect 278998 267744 279054 267753
rect 278998 267679 279054 267688
rect 279012 260794 279040 267679
rect 278828 260766 279040 260794
rect 278828 251258 278856 260766
rect 278816 251252 278868 251258
rect 278816 251194 278868 251200
rect 278816 251116 278868 251122
rect 278816 251058 278868 251064
rect 278828 236722 278856 251058
rect 278736 236694 278856 236722
rect 278736 231826 278764 236694
rect 278736 231798 278856 231826
rect 278828 211018 278856 231798
rect 278828 210990 278948 211018
rect 278920 206122 278948 210990
rect 278828 206094 278948 206122
rect 278828 180810 278856 206094
rect 278816 180804 278868 180810
rect 278816 180746 278868 180752
rect 278816 171148 278868 171154
rect 278816 171090 278868 171096
rect 278828 163033 278856 171090
rect 278814 163024 278870 163033
rect 278814 162959 278870 162968
rect 278722 162888 278778 162897
rect 278722 162823 278778 162832
rect 278736 149870 278764 162823
rect 278724 149864 278776 149870
rect 278724 149806 278776 149812
rect 278816 142180 278868 142186
rect 278816 142122 278868 142128
rect 278828 93974 278856 142122
rect 278816 93968 278868 93974
rect 278816 93910 278868 93916
rect 278724 93900 278776 93906
rect 278724 93842 278776 93848
rect 278736 67726 278764 93842
rect 278724 67720 278776 67726
rect 278724 67662 278776 67668
rect 278632 67584 278684 67590
rect 278632 67526 278684 67532
rect 278644 64870 278672 67526
rect 278632 64864 278684 64870
rect 278632 64806 278684 64812
rect 278724 55276 278776 55282
rect 278724 55218 278776 55224
rect 278736 55162 278764 55218
rect 278736 55134 278856 55162
rect 278828 48346 278856 55134
rect 278816 48340 278868 48346
rect 278816 48282 278868 48288
rect 278724 45620 278776 45626
rect 278724 45562 278776 45568
rect 278736 37262 278764 45562
rect 278724 37256 278776 37262
rect 278724 37198 278776 37204
rect 278908 37256 278960 37262
rect 278908 37198 278960 37204
rect 278920 35850 278948 37198
rect 278828 35822 278948 35850
rect 278828 27674 278856 35822
rect 278816 27668 278868 27674
rect 278816 27610 278868 27616
rect 278816 26308 278868 26314
rect 278816 26250 278868 26256
rect 278828 16658 278856 26250
rect 278632 16652 278684 16658
rect 278632 16594 278684 16600
rect 278816 16652 278868 16658
rect 278816 16594 278868 16600
rect 278644 16561 278672 16594
rect 278630 16552 278686 16561
rect 278630 16487 278686 16496
rect 278724 6928 278776 6934
rect 278724 6870 278776 6876
rect 278736 5234 278764 6870
rect 278724 5228 278776 5234
rect 278724 5170 278776 5176
rect 278500 3556 278580 3584
rect 278448 3538 278500 3544
rect 272192 3392 272244 3398
rect 272192 3334 272244 3340
rect 270996 3188 271048 3194
rect 270996 3130 271048 3136
rect 271008 480 271036 3130
rect 272204 480 272232 3334
rect 273400 480 273428 3538
rect 275780 3460 275832 3466
rect 275780 3402 275832 3408
rect 274584 2984 274636 2990
rect 274584 2926 274636 2932
rect 274596 480 274624 2926
rect 275792 480 275820 3402
rect 278172 3188 278224 3194
rect 278172 3130 278224 3136
rect 276976 2916 277028 2922
rect 276976 2858 277028 2864
rect 276988 480 277016 2858
rect 278184 480 278212 3130
rect 279288 2854 279316 335514
rect 279368 332852 279420 332858
rect 279368 332794 279420 332800
rect 279380 4758 279408 332794
rect 279458 249792 279514 249801
rect 279458 249727 279514 249736
rect 279472 240174 279500 249727
rect 279460 240168 279512 240174
rect 279460 240110 279512 240116
rect 279564 7886 279592 340054
rect 279656 9382 279684 340068
rect 279748 340054 279946 340082
rect 280024 340054 280222 340082
rect 280300 340054 280406 340082
rect 279748 332858 279776 340054
rect 280024 334354 280052 340054
rect 280104 337204 280156 337210
rect 280104 337146 280156 337152
rect 280012 334348 280064 334354
rect 280012 334290 280064 334296
rect 280116 334234 280144 337146
rect 280300 335578 280328 340054
rect 280668 337754 280696 340068
rect 280852 340054 280958 340082
rect 281036 340054 281142 340082
rect 281312 340054 281418 340082
rect 281496 340054 281694 340082
rect 280656 337748 280708 337754
rect 280656 337690 280708 337696
rect 280288 335572 280340 335578
rect 280288 335514 280340 335520
rect 280748 335572 280800 335578
rect 280748 335514 280800 335520
rect 279932 334206 280144 334234
rect 279736 332852 279788 332858
rect 279736 332794 279788 332800
rect 279828 327140 279880 327146
rect 279828 327082 279880 327088
rect 279840 285002 279868 327082
rect 279748 284974 279868 285002
rect 279748 278769 279776 284974
rect 279734 278760 279790 278769
rect 279734 278695 279790 278704
rect 279828 269136 279880 269142
rect 279828 269078 279880 269084
rect 279840 260914 279868 269078
rect 279736 260908 279788 260914
rect 279736 260850 279788 260856
rect 279828 260908 279880 260914
rect 279828 260850 279880 260856
rect 279748 256086 279776 260850
rect 279736 256080 279788 256086
rect 279736 256022 279788 256028
rect 279828 256012 279880 256018
rect 279828 255954 279880 255960
rect 279840 249801 279868 255954
rect 279826 249792 279882 249801
rect 279826 249727 279882 249736
rect 279736 240168 279788 240174
rect 279736 240110 279788 240116
rect 279748 236722 279776 240110
rect 279748 236694 279868 236722
rect 279840 219502 279868 236694
rect 279736 219496 279788 219502
rect 279736 219438 279788 219444
rect 279828 219496 279880 219502
rect 279828 219438 279880 219444
rect 279748 212498 279776 219438
rect 279736 212492 279788 212498
rect 279736 212434 279788 212440
rect 279828 212492 279880 212498
rect 279828 212434 279880 212440
rect 279840 200122 279868 212434
rect 279828 200116 279880 200122
rect 279828 200058 279880 200064
rect 279828 190528 279880 190534
rect 279828 190470 279880 190476
rect 279840 183666 279868 190470
rect 279828 183660 279880 183666
rect 279828 183602 279880 183608
rect 279736 183524 279788 183530
rect 279736 183466 279788 183472
rect 279748 164234 279776 183466
rect 279748 164206 279868 164234
rect 279840 139482 279868 164206
rect 279748 139454 279868 139482
rect 279748 139398 279776 139454
rect 279736 139392 279788 139398
rect 279736 139334 279788 139340
rect 279828 129804 279880 129810
rect 279828 129746 279880 129752
rect 279840 121446 279868 129746
rect 279736 121440 279788 121446
rect 279736 121382 279788 121388
rect 279828 121440 279880 121446
rect 279828 121382 279880 121388
rect 279748 100774 279776 121382
rect 279736 100768 279788 100774
rect 279736 100710 279788 100716
rect 279826 100736 279882 100745
rect 279826 100671 279882 100680
rect 279840 91118 279868 100671
rect 279828 91112 279880 91118
rect 279828 91054 279880 91060
rect 279828 86828 279880 86834
rect 279828 86770 279880 86776
rect 279840 82822 279868 86770
rect 279932 84266 279960 334206
rect 280010 278760 280066 278769
rect 280010 278695 280066 278704
rect 280024 269142 280052 278695
rect 280012 269136 280064 269142
rect 280012 269078 280064 269084
rect 280012 100768 280064 100774
rect 280010 100736 280012 100745
rect 280064 100736 280066 100745
rect 280010 100671 280066 100680
rect 280012 91112 280064 91118
rect 280012 91054 280064 91060
rect 280024 86834 280052 91054
rect 280012 86828 280064 86834
rect 280012 86770 280064 86776
rect 279932 84250 280052 84266
rect 279932 84244 280064 84250
rect 279932 84238 280012 84244
rect 280012 84186 280064 84192
rect 279920 84176 279972 84182
rect 279920 84118 279972 84124
rect 279828 82816 279880 82822
rect 279828 82758 279880 82764
rect 279932 74662 279960 84118
rect 280104 82816 280156 82822
rect 280104 82758 280156 82764
rect 279920 74656 279972 74662
rect 279920 74598 279972 74604
rect 280116 74474 280144 82758
rect 279920 74452 279972 74458
rect 279920 74394 279972 74400
rect 280024 74446 280144 74474
rect 279734 64968 279790 64977
rect 279734 64903 279790 64912
rect 279748 64870 279776 64903
rect 279736 64864 279788 64870
rect 279736 64806 279788 64812
rect 279736 55276 279788 55282
rect 279736 55218 279788 55224
rect 279748 51814 279776 55218
rect 279736 51808 279788 51814
rect 279736 51750 279788 51756
rect 279828 37256 279880 37262
rect 279828 37198 279880 37204
rect 279644 9376 279696 9382
rect 279644 9318 279696 9324
rect 279840 7954 279868 37198
rect 279828 7948 279880 7954
rect 279828 7890 279880 7896
rect 279552 7880 279604 7886
rect 279552 7822 279604 7828
rect 279368 4752 279420 4758
rect 279368 4694 279420 4700
rect 279932 2922 279960 74394
rect 280024 64977 280052 74446
rect 280010 64968 280066 64977
rect 280010 64903 280066 64912
rect 280012 51808 280064 51814
rect 280012 51750 280064 51756
rect 280024 37330 280052 51750
rect 280012 37324 280064 37330
rect 280012 37266 280064 37272
rect 280760 8090 280788 335514
rect 280748 8084 280800 8090
rect 280748 8026 280800 8032
rect 280852 8022 280880 340054
rect 280840 8016 280892 8022
rect 280840 7958 280892 7964
rect 281036 3602 281064 340054
rect 281312 11762 281340 340054
rect 281496 335578 281524 340054
rect 281864 337618 281892 340068
rect 282154 340054 282260 340082
rect 281852 337612 281904 337618
rect 281852 337554 281904 337560
rect 281484 335572 281536 335578
rect 281484 335514 281536 335520
rect 282232 14482 282260 340054
rect 282416 337414 282444 340068
rect 282600 337550 282628 340068
rect 282692 340054 282890 340082
rect 282588 337544 282640 337550
rect 282588 337486 282640 337492
rect 282404 337408 282456 337414
rect 282404 337350 282456 337356
rect 282692 335594 282720 340054
rect 283152 337482 283180 340068
rect 283244 340054 283350 340082
rect 283140 337476 283192 337482
rect 283140 337418 283192 337424
rect 282508 335566 282720 335594
rect 282312 331628 282364 331634
rect 282312 331570 282364 331576
rect 282220 14476 282272 14482
rect 282220 14418 282272 14424
rect 281300 11756 281352 11762
rect 281300 11698 281352 11704
rect 281024 3596 281076 3602
rect 281024 3538 281076 3544
rect 282324 3534 282352 331570
rect 282508 10470 282536 335566
rect 283244 331634 283272 340054
rect 283508 337068 283560 337074
rect 283508 337010 283560 337016
rect 283232 331628 283284 331634
rect 283232 331570 283284 331576
rect 282496 10464 282548 10470
rect 282496 10406 282548 10412
rect 283520 4690 283548 337010
rect 283612 5370 283640 340068
rect 283888 338094 283916 340068
rect 283876 338088 283928 338094
rect 283876 338030 283928 338036
rect 284072 337754 284100 340068
rect 284164 340054 284362 340082
rect 284440 340054 284638 340082
rect 284822 340054 285020 340082
rect 284060 337748 284112 337754
rect 284060 337690 284112 337696
rect 284164 337074 284192 340054
rect 284152 337068 284204 337074
rect 284152 337010 284204 337016
rect 284440 336954 284468 340054
rect 283704 336926 284468 336954
rect 283600 5364 283652 5370
rect 283600 5306 283652 5312
rect 283508 4684 283560 4690
rect 283508 4626 283560 4632
rect 283704 3738 283732 336926
rect 284060 336864 284112 336870
rect 284060 336806 284112 336812
rect 284152 336864 284204 336870
rect 284152 336806 284204 336812
rect 284072 4434 284100 336806
rect 283980 4406 284100 4434
rect 283692 3732 283744 3738
rect 283692 3674 283744 3680
rect 282956 3596 283008 3602
rect 282956 3538 283008 3544
rect 282312 3528 282364 3534
rect 282312 3470 282364 3476
rect 280104 3460 280156 3466
rect 280104 3402 280156 3408
rect 279920 2916 279972 2922
rect 279920 2858 279972 2864
rect 279276 2848 279328 2854
rect 279276 2790 279328 2796
rect 280116 1850 280144 3402
rect 280564 2916 280616 2922
rect 280564 2858 280616 2864
rect 279380 1822 280144 1850
rect 279380 480 279408 1822
rect 280576 480 280604 2858
rect 281760 2848 281812 2854
rect 281760 2790 281812 2796
rect 281772 480 281800 2790
rect 282968 480 282996 3538
rect 283980 2922 284008 4406
rect 284164 4298 284192 336806
rect 284992 336462 285020 340054
rect 285084 336870 285112 340068
rect 285176 340054 285374 340082
rect 285452 340054 285558 340082
rect 285636 340054 285834 340082
rect 286004 340054 286110 340082
rect 286294 340054 286400 340082
rect 285072 336864 285124 336870
rect 285072 336806 285124 336812
rect 284980 336456 285032 336462
rect 284980 336398 285032 336404
rect 284980 335504 285032 335510
rect 284980 335446 285032 335452
rect 284888 333328 284940 333334
rect 284888 333270 284940 333276
rect 284796 164416 284848 164422
rect 284796 164358 284848 164364
rect 284808 164257 284836 164358
rect 284794 164248 284850 164257
rect 284794 164183 284850 164192
rect 284072 4270 284192 4298
rect 284072 3942 284100 4270
rect 284152 4140 284204 4146
rect 284152 4082 284204 4088
rect 284060 3936 284112 3942
rect 284060 3878 284112 3884
rect 283968 2916 284020 2922
rect 283968 2858 284020 2864
rect 284164 480 284192 4082
rect 284900 4010 284928 333270
rect 284992 4078 285020 335446
rect 285176 333334 285204 340054
rect 285164 333328 285216 333334
rect 285164 333270 285216 333276
rect 285452 331498 285480 340054
rect 285636 335510 285664 340054
rect 285624 335504 285676 335510
rect 285624 335446 285676 335452
rect 285440 331492 285492 331498
rect 285440 331434 285492 331440
rect 285164 331152 285216 331158
rect 285164 331094 285216 331100
rect 285440 331152 285492 331158
rect 285440 331094 285492 331100
rect 285176 318594 285204 331094
rect 285348 328500 285400 328506
rect 285348 328442 285400 328448
rect 285360 321586 285388 328442
rect 285268 321558 285388 321586
rect 285268 318714 285296 321558
rect 285256 318708 285308 318714
rect 285256 318650 285308 318656
rect 285084 318566 285204 318594
rect 285084 313698 285112 318566
rect 285084 313670 285204 313698
rect 285176 279886 285204 313670
rect 285452 309330 285480 331094
rect 286004 328506 286032 340054
rect 285716 328500 285768 328506
rect 285716 328442 285768 328448
rect 285992 328500 286044 328506
rect 285992 328442 286044 328448
rect 285728 323626 285756 328442
rect 285636 323598 285756 323626
rect 285636 318714 285664 323598
rect 285624 318708 285676 318714
rect 285624 318650 285676 318656
rect 285440 309324 285492 309330
rect 285440 309266 285492 309272
rect 285348 309188 285400 309194
rect 285348 309130 285400 309136
rect 285440 309188 285492 309194
rect 285440 309130 285492 309136
rect 285716 309188 285768 309194
rect 285716 309130 285768 309136
rect 285360 302326 285388 309130
rect 285348 302320 285400 302326
rect 285348 302262 285400 302268
rect 285256 302184 285308 302190
rect 285256 302126 285308 302132
rect 285268 279886 285296 302126
rect 285164 279880 285216 279886
rect 285164 279822 285216 279828
rect 285256 279880 285308 279886
rect 285256 279822 285308 279828
rect 285348 270564 285400 270570
rect 285348 270506 285400 270512
rect 285164 269136 285216 269142
rect 285164 269078 285216 269084
rect 285072 198756 285124 198762
rect 285072 198698 285124 198704
rect 285084 186318 285112 198698
rect 285072 186312 285124 186318
rect 285072 186254 285124 186260
rect 285176 182170 285204 269078
rect 285360 263702 285388 270506
rect 285348 263696 285400 263702
rect 285348 263638 285400 263644
rect 285256 263560 285308 263566
rect 285256 263502 285308 263508
rect 285268 260778 285296 263502
rect 285256 260772 285308 260778
rect 285256 260714 285308 260720
rect 285348 251252 285400 251258
rect 285348 251194 285400 251200
rect 285360 244390 285388 251194
rect 285348 244384 285400 244390
rect 285348 244326 285400 244332
rect 285348 244180 285400 244186
rect 285348 244122 285400 244128
rect 285360 236774 285388 244122
rect 285348 236768 285400 236774
rect 285348 236710 285400 236716
rect 285348 231940 285400 231946
rect 285348 231882 285400 231888
rect 285360 225010 285388 231882
rect 285348 225004 285400 225010
rect 285348 224946 285400 224952
rect 285256 219496 285308 219502
rect 285256 219438 285308 219444
rect 285268 208622 285296 219438
rect 285256 208616 285308 208622
rect 285256 208558 285308 208564
rect 285256 208480 285308 208486
rect 285256 208422 285308 208428
rect 285268 208282 285296 208422
rect 285256 208276 285308 208282
rect 285256 208218 285308 208224
rect 285256 186312 285308 186318
rect 285256 186254 285308 186260
rect 285164 182164 285216 182170
rect 285164 182106 285216 182112
rect 285268 177313 285296 186254
rect 285254 177304 285310 177313
rect 285254 177239 285310 177248
rect 285164 172576 285216 172582
rect 285164 172518 285216 172524
rect 285176 164529 285204 172518
rect 285162 164520 285218 164529
rect 285162 164455 285218 164464
rect 285162 164384 285218 164393
rect 285162 164319 285218 164328
rect 285176 156806 285204 164319
rect 285346 164112 285402 164121
rect 285346 164047 285402 164056
rect 285360 161498 285388 164047
rect 285256 161492 285308 161498
rect 285256 161434 285308 161440
rect 285348 161492 285400 161498
rect 285348 161434 285400 161440
rect 285268 161378 285296 161434
rect 285268 161350 285388 161378
rect 285360 157418 285388 161350
rect 285348 157412 285400 157418
rect 285348 157354 285400 157360
rect 285164 156800 285216 156806
rect 285164 156742 285216 156748
rect 285348 138100 285400 138106
rect 285348 138042 285400 138048
rect 285164 137896 285216 137902
rect 285164 137838 285216 137844
rect 285072 46912 285124 46918
rect 285072 46854 285124 46860
rect 285084 29034 285112 46854
rect 285072 29028 285124 29034
rect 285072 28970 285124 28976
rect 285176 28966 285204 137838
rect 285360 128466 285388 138042
rect 285452 135590 285480 309130
rect 285728 302326 285756 309130
rect 285716 302320 285768 302326
rect 285716 302262 285768 302268
rect 285808 302116 285860 302122
rect 285808 302058 285860 302064
rect 285820 278730 285848 302058
rect 285716 278724 285768 278730
rect 285716 278666 285768 278672
rect 285808 278724 285860 278730
rect 285808 278666 285860 278672
rect 285728 260930 285756 278666
rect 285636 260902 285756 260930
rect 285636 260846 285664 260902
rect 285624 260840 285676 260846
rect 285624 260782 285676 260788
rect 285716 251252 285768 251258
rect 285716 251194 285768 251200
rect 285728 246378 285756 251194
rect 285728 246350 285940 246378
rect 285912 244202 285940 246350
rect 285820 244174 285940 244202
rect 285820 231878 285848 244174
rect 285716 231872 285768 231878
rect 285716 231814 285768 231820
rect 285808 231872 285860 231878
rect 285808 231814 285860 231820
rect 285728 225010 285756 231814
rect 285532 225004 285584 225010
rect 285532 224946 285584 224952
rect 285716 225004 285768 225010
rect 285716 224946 285768 224952
rect 285544 224890 285572 224946
rect 285544 224862 285664 224890
rect 285636 215370 285664 224862
rect 285636 215342 285756 215370
rect 285728 201550 285756 215342
rect 285624 201544 285676 201550
rect 285624 201486 285676 201492
rect 285716 201544 285768 201550
rect 285716 201486 285768 201492
rect 285636 196058 285664 201486
rect 285544 196030 285664 196058
rect 285544 186386 285572 196030
rect 285532 186380 285584 186386
rect 285532 186322 285584 186328
rect 285624 186244 285676 186250
rect 285624 186186 285676 186192
rect 285636 182170 285664 186186
rect 285624 182164 285676 182170
rect 285624 182106 285676 182112
rect 285716 182164 285768 182170
rect 285716 182106 285768 182112
rect 285728 166870 285756 182106
rect 285716 166864 285768 166870
rect 285716 166806 285768 166812
rect 285716 166728 285768 166734
rect 285716 166670 285768 166676
rect 285624 164416 285676 164422
rect 285624 164358 285676 164364
rect 285636 164257 285664 164358
rect 285622 164248 285678 164257
rect 285622 164183 285678 164192
rect 285728 147694 285756 166670
rect 285532 147688 285584 147694
rect 285716 147688 285768 147694
rect 285584 147636 285664 147642
rect 285532 147630 285664 147636
rect 285716 147630 285768 147636
rect 285544 147614 285664 147630
rect 285636 144906 285664 147614
rect 285624 144900 285676 144906
rect 285624 144842 285676 144848
rect 285624 137964 285676 137970
rect 285624 137906 285676 137912
rect 285440 135584 285492 135590
rect 285440 135526 285492 135532
rect 285532 135312 285584 135318
rect 285268 128438 285388 128466
rect 285452 135260 285532 135266
rect 285452 135254 285584 135260
rect 285636 135266 285664 137906
rect 285452 135238 285572 135254
rect 285636 135238 285756 135266
rect 285268 111858 285296 128438
rect 285256 111852 285308 111858
rect 285256 111794 285308 111800
rect 285348 111852 285400 111858
rect 285348 111794 285400 111800
rect 285360 102406 285388 111794
rect 285348 102400 285400 102406
rect 285348 102342 285400 102348
rect 285256 102196 285308 102202
rect 285256 102138 285308 102144
rect 285268 93906 285296 102138
rect 285256 93900 285308 93906
rect 285256 93842 285308 93848
rect 285348 93900 285400 93906
rect 285348 93842 285400 93848
rect 285360 84266 285388 93842
rect 285268 84238 285388 84266
rect 285268 82822 285296 84238
rect 285256 82816 285308 82822
rect 285256 82758 285308 82764
rect 285256 77988 285308 77994
rect 285256 77930 285308 77936
rect 285268 64870 285296 77930
rect 285256 64864 285308 64870
rect 285256 64806 285308 64812
rect 285256 56500 285308 56506
rect 285256 56442 285308 56448
rect 285268 46918 285296 56442
rect 285256 46912 285308 46918
rect 285256 46854 285308 46860
rect 285256 29028 285308 29034
rect 285256 28970 285308 28976
rect 285164 28960 285216 28966
rect 285070 28928 285126 28937
rect 285268 28937 285296 28970
rect 285164 28902 285216 28908
rect 285254 28928 285310 28937
rect 285070 28863 285126 28872
rect 285254 28863 285310 28872
rect 285084 19446 285112 28863
rect 285072 19440 285124 19446
rect 285072 19382 285124 19388
rect 285164 19372 285216 19378
rect 285164 19314 285216 19320
rect 285348 19372 285400 19378
rect 285348 19314 285400 19320
rect 285070 19272 285126 19281
rect 285070 19207 285126 19216
rect 285084 9722 285112 19207
rect 285072 9716 285124 9722
rect 285072 9658 285124 9664
rect 284980 4072 285032 4078
rect 284980 4014 285032 4020
rect 284888 4004 284940 4010
rect 284888 3946 284940 3952
rect 285176 3670 285204 19314
rect 285360 19281 285388 19314
rect 285346 19272 285402 19281
rect 285346 19207 285402 19216
rect 285256 9716 285308 9722
rect 285256 9658 285308 9664
rect 285268 3942 285296 9658
rect 285452 4146 285480 135238
rect 285728 124114 285756 135238
rect 285636 124086 285756 124114
rect 285636 120086 285664 124086
rect 285624 120080 285676 120086
rect 285624 120022 285676 120028
rect 285624 111308 285676 111314
rect 285624 111250 285676 111256
rect 285636 106978 285664 111250
rect 285636 106950 285756 106978
rect 285728 66450 285756 106950
rect 285728 66422 285848 66450
rect 285820 66298 285848 66422
rect 285624 66292 285676 66298
rect 285624 66234 285676 66240
rect 285808 66292 285860 66298
rect 285808 66234 285860 66240
rect 285636 60874 285664 66234
rect 285636 60846 285756 60874
rect 285728 60058 285756 60846
rect 285636 60030 285756 60058
rect 285636 42090 285664 60030
rect 285624 42084 285676 42090
rect 285624 42026 285676 42032
rect 285808 29028 285860 29034
rect 285808 28970 285860 28976
rect 285820 24206 285848 28970
rect 285808 24200 285860 24206
rect 285808 24142 285860 24148
rect 285716 19372 285768 19378
rect 285716 19314 285768 19320
rect 285728 12458 285756 19314
rect 285544 12430 285756 12458
rect 285440 4140 285492 4146
rect 285440 4082 285492 4088
rect 285256 3936 285308 3942
rect 285256 3878 285308 3884
rect 285164 3664 285216 3670
rect 285164 3606 285216 3612
rect 285256 3664 285308 3670
rect 285256 3606 285308 3612
rect 285268 480 285296 3606
rect 285544 3126 285572 12430
rect 285532 3120 285584 3126
rect 285532 3062 285584 3068
rect 286372 3058 286400 340054
rect 286556 337142 286584 340068
rect 286648 340054 286846 340082
rect 286924 340054 287030 340082
rect 286544 337136 286596 337142
rect 286544 337078 286596 337084
rect 286452 4004 286504 4010
rect 286452 3946 286504 3952
rect 286360 3052 286412 3058
rect 286360 2994 286412 3000
rect 286464 480 286492 3946
rect 286648 2990 286676 340054
rect 286924 333010 286952 340054
rect 287292 337210 287320 340068
rect 287280 337204 287332 337210
rect 287280 337146 287332 337152
rect 287568 336870 287596 340068
rect 287766 340054 287964 340082
rect 287096 336864 287148 336870
rect 287096 336806 287148 336812
rect 287556 336864 287608 336870
rect 287556 336806 287608 336812
rect 286740 332982 286952 333010
rect 286740 3398 286768 332982
rect 287108 332874 287136 336806
rect 287936 335594 287964 340054
rect 288028 337006 288056 340068
rect 288212 340054 288318 340082
rect 288396 340054 288502 340082
rect 288016 337000 288068 337006
rect 288016 336942 288068 336948
rect 287936 335566 288148 335594
rect 286832 332846 287136 332874
rect 286728 3392 286780 3398
rect 286728 3334 286780 3340
rect 286832 3194 286860 332846
rect 287924 332036 287976 332042
rect 287924 331978 287976 331984
rect 287648 4140 287700 4146
rect 287648 4082 287700 4088
rect 286820 3188 286872 3194
rect 286820 3130 286872 3136
rect 286636 2984 286688 2990
rect 286636 2926 286688 2932
rect 287660 480 287688 4082
rect 287936 3602 287964 331978
rect 287924 3596 287976 3602
rect 287924 3538 287976 3544
rect 288120 3466 288148 335566
rect 288108 3460 288160 3466
rect 288108 3402 288160 3408
rect 288212 2854 288240 340054
rect 288396 332042 288424 340054
rect 288384 332036 288436 332042
rect 288384 331978 288436 331984
rect 288764 331158 288792 340068
rect 288844 336864 288896 336870
rect 288844 336806 288896 336812
rect 288752 331152 288804 331158
rect 288752 331094 288804 331100
rect 288856 4282 288884 336806
rect 289040 335510 289068 340068
rect 289132 340054 289238 340082
rect 289028 335504 289080 335510
rect 289028 335446 289080 335452
rect 288844 4276 288896 4282
rect 288844 4218 288896 4224
rect 288844 4140 288896 4146
rect 288844 4082 288896 4088
rect 288200 2848 288252 2854
rect 288200 2790 288252 2796
rect 288856 480 288884 4082
rect 289132 4010 289160 340054
rect 289500 336870 289528 340068
rect 289592 340054 289790 340082
rect 289868 340054 289974 340082
rect 289488 336864 289540 336870
rect 289488 336806 289540 336812
rect 289592 335730 289620 340054
rect 289408 335702 289620 335730
rect 289408 4146 289436 335702
rect 289868 335594 289896 340054
rect 290236 336818 290264 340068
rect 290512 337006 290540 340068
rect 290500 337000 290552 337006
rect 290500 336942 290552 336948
rect 290696 336870 290724 340068
rect 290972 336938 291000 340068
rect 291156 337074 291184 340068
rect 291432 337142 291460 340068
rect 291420 337136 291472 337142
rect 291420 337078 291472 337084
rect 291144 337068 291196 337074
rect 291144 337010 291196 337016
rect 291512 337000 291564 337006
rect 291512 336942 291564 336948
rect 290960 336932 291012 336938
rect 290960 336874 291012 336880
rect 290684 336864 290736 336870
rect 290236 336790 290632 336818
rect 290684 336806 290736 336812
rect 291420 336864 291472 336870
rect 291420 336806 291472 336812
rect 289592 335566 289896 335594
rect 289592 4146 289620 335566
rect 289672 335504 289724 335510
rect 289672 335446 289724 335452
rect 289396 4140 289448 4146
rect 289396 4082 289448 4088
rect 289580 4140 289632 4146
rect 289580 4082 289632 4088
rect 289120 4004 289172 4010
rect 289120 3946 289172 3952
rect 289684 3670 289712 335446
rect 290316 320272 290368 320278
rect 290314 320240 290316 320249
rect 290368 320240 290370 320249
rect 290314 320175 290370 320184
rect 289946 241768 290002 241777
rect 290002 241726 290080 241754
rect 289946 241703 290002 241712
rect 290052 241641 290080 241726
rect 290316 241664 290368 241670
rect 290038 241632 290094 241641
rect 290038 241567 290094 241576
rect 290314 241632 290316 241641
rect 290368 241632 290370 241641
rect 290314 241567 290370 241576
rect 290316 132864 290368 132870
rect 290314 132832 290316 132841
rect 290368 132832 290370 132841
rect 290314 132767 290370 132776
rect 290222 101144 290278 101153
rect 290406 101144 290462 101153
rect 290278 101102 290406 101130
rect 290222 101079 290278 101088
rect 290406 101079 290462 101088
rect 290040 4140 290092 4146
rect 290040 4082 290092 4088
rect 289672 3664 289724 3670
rect 289672 3606 289724 3612
rect 290052 480 290080 4082
rect 290604 610 290632 336790
rect 291432 3466 291460 336806
rect 291524 4146 291552 336942
rect 291708 336938 291736 340068
rect 291892 337006 291920 340068
rect 292182 340054 292380 340082
rect 292248 337068 292300 337074
rect 292248 337010 292300 337016
rect 291880 337000 291932 337006
rect 291880 336942 291932 336948
rect 291604 336932 291656 336938
rect 291604 336874 291656 336880
rect 291696 336932 291748 336938
rect 291696 336874 291748 336880
rect 291512 4140 291564 4146
rect 291512 4082 291564 4088
rect 291420 3460 291472 3466
rect 291420 3402 291472 3408
rect 291616 2990 291644 336874
rect 292260 335458 292288 337010
rect 292352 335594 292380 340054
rect 292444 336870 292472 340068
rect 292628 338026 292656 340068
rect 292616 338020 292668 338026
rect 292616 337962 292668 337968
rect 292904 337686 292932 340068
rect 292892 337680 292944 337686
rect 292892 337622 292944 337628
rect 293180 337210 293208 340068
rect 293364 337754 293392 340068
rect 293352 337748 293404 337754
rect 293352 337690 293404 337696
rect 293640 337618 293668 340068
rect 293812 338020 293864 338026
rect 293812 337962 293864 337968
rect 293720 337680 293772 337686
rect 293720 337622 293772 337628
rect 293628 337612 293680 337618
rect 293628 337554 293680 337560
rect 293168 337204 293220 337210
rect 293168 337146 293220 337152
rect 292892 337000 292944 337006
rect 292892 336942 292944 336948
rect 292800 336932 292852 336938
rect 292800 336874 292852 336880
rect 292432 336864 292484 336870
rect 292432 336806 292484 336812
rect 292352 335566 292748 335594
rect 292260 335430 292380 335458
rect 292352 3126 292380 335430
rect 292432 4140 292484 4146
rect 292432 4082 292484 4088
rect 292340 3120 292392 3126
rect 292340 3062 292392 3068
rect 291604 2984 291656 2990
rect 291604 2926 291656 2932
rect 290592 604 290644 610
rect 290592 546 290644 552
rect 291236 604 291288 610
rect 291236 546 291288 552
rect 291248 480 291276 546
rect 292444 480 292472 4082
rect 292720 3534 292748 335566
rect 292812 3942 292840 336874
rect 292800 3936 292852 3942
rect 292800 3878 292852 3884
rect 292904 3738 292932 336942
rect 292984 336864 293036 336870
rect 292984 336806 293036 336812
rect 292892 3732 292944 3738
rect 292892 3674 292944 3680
rect 292708 3528 292760 3534
rect 292708 3470 292760 3476
rect 292996 2922 293024 336806
rect 293626 180024 293682 180033
rect 293626 179959 293682 179968
rect 293640 179761 293668 179959
rect 293626 179752 293682 179761
rect 293626 179687 293682 179696
rect 293260 132864 293312 132870
rect 293260 132806 293312 132812
rect 293272 132705 293300 132806
rect 293258 132696 293314 132705
rect 293258 132631 293314 132640
rect 293628 3460 293680 3466
rect 293628 3402 293680 3408
rect 292984 2916 293036 2922
rect 292984 2858 293036 2864
rect 293640 480 293668 3402
rect 293732 3398 293760 337622
rect 293720 3392 293772 3398
rect 293720 3334 293772 3340
rect 293824 2854 293852 337962
rect 293916 337686 293944 340068
rect 293904 337680 293956 337686
rect 293904 337622 293956 337628
rect 293904 337136 293956 337142
rect 293904 337078 293956 337084
rect 293916 4146 293944 337078
rect 293904 4140 293956 4146
rect 293904 4082 293956 4088
rect 294100 3194 294128 340068
rect 294284 340054 294390 340082
rect 294180 337748 294232 337754
rect 294180 337690 294232 337696
rect 294088 3188 294140 3194
rect 294088 3130 294140 3136
rect 294192 3058 294220 337690
rect 294284 4078 294312 340054
rect 294364 337612 294416 337618
rect 294364 337554 294416 337560
rect 294272 4072 294324 4078
rect 294272 4014 294324 4020
rect 294376 3466 294404 337554
rect 294652 337482 294680 340068
rect 294836 337754 294864 340068
rect 294824 337748 294876 337754
rect 294824 337690 294876 337696
rect 294640 337476 294692 337482
rect 294640 337418 294692 337424
rect 295112 337414 295140 340068
rect 295388 337686 295416 340068
rect 295586 340054 295692 340082
rect 295192 337680 295244 337686
rect 295192 337622 295244 337628
rect 295376 337680 295428 337686
rect 295376 337622 295428 337628
rect 295560 337680 295612 337686
rect 295560 337622 295612 337628
rect 295100 337408 295152 337414
rect 295100 337350 295152 337356
rect 295100 337204 295152 337210
rect 295100 337146 295152 337152
rect 294638 320512 294694 320521
rect 294638 320447 294694 320456
rect 294652 320278 294680 320447
rect 294640 320272 294692 320278
rect 294640 320214 294692 320220
rect 294822 241904 294878 241913
rect 294822 241839 294878 241848
rect 294836 241670 294864 241839
rect 294824 241664 294876 241670
rect 294824 241606 294876 241612
rect 295112 4010 295140 337146
rect 295204 181490 295232 337622
rect 295192 181484 295244 181490
rect 295192 181426 295244 181432
rect 295572 11830 295600 337622
rect 295560 11824 295612 11830
rect 295560 11766 295612 11772
rect 295664 5098 295692 340054
rect 295744 337748 295796 337754
rect 295744 337690 295796 337696
rect 295652 5092 295704 5098
rect 295652 5034 295704 5040
rect 295100 4004 295152 4010
rect 295100 3946 295152 3952
rect 295756 3670 295784 337690
rect 295848 337550 295876 340068
rect 296124 337618 296152 340068
rect 296308 337754 296336 340068
rect 296296 337748 296348 337754
rect 296296 337690 296348 337696
rect 296584 337686 296612 340068
rect 296874 340054 296980 340082
rect 296756 337748 296808 337754
rect 296756 337690 296808 337696
rect 296848 337748 296900 337754
rect 296848 337690 296900 337696
rect 296572 337680 296624 337686
rect 296572 337622 296624 337628
rect 296112 337612 296164 337618
rect 296112 337554 296164 337560
rect 295836 337544 295888 337550
rect 295836 337486 295888 337492
rect 296768 5234 296796 337690
rect 296756 5228 296808 5234
rect 296756 5170 296808 5176
rect 296860 5166 296888 337690
rect 296848 5160 296900 5166
rect 296848 5102 296900 5108
rect 296952 4826 296980 340054
rect 297044 337754 297072 340068
rect 297320 338026 297348 340068
rect 297308 338020 297360 338026
rect 297308 337962 297360 337968
rect 297596 337754 297624 340068
rect 297032 337748 297084 337754
rect 297032 337690 297084 337696
rect 297584 337748 297636 337754
rect 297584 337690 297636 337696
rect 297780 337618 297808 340068
rect 297032 337612 297084 337618
rect 297032 337554 297084 337560
rect 297768 337612 297820 337618
rect 297768 337554 297820 337560
rect 296940 4820 296992 4826
rect 296940 4762 296992 4768
rect 297044 4758 297072 337554
rect 297124 337544 297176 337550
rect 297124 337486 297176 337492
rect 297032 4752 297084 4758
rect 297032 4694 297084 4700
rect 295744 3664 295796 3670
rect 295744 3606 295796 3612
rect 297136 3602 297164 337486
rect 298056 337006 298084 340068
rect 298346 340054 298452 340082
rect 298228 337952 298280 337958
rect 298228 337894 298280 337900
rect 298044 337000 298096 337006
rect 298044 336942 298096 336948
rect 298240 4282 298268 337894
rect 298320 337748 298372 337754
rect 298424 337736 298452 340054
rect 298516 337958 298544 340068
rect 298504 337952 298556 337958
rect 298504 337894 298556 337900
rect 298792 337754 298820 340068
rect 298780 337748 298832 337754
rect 298424 337708 298544 337736
rect 298320 337690 298372 337696
rect 298228 4276 298280 4282
rect 298228 4218 298280 4224
rect 298332 4214 298360 337690
rect 298412 337612 298464 337618
rect 298412 337554 298464 337560
rect 298424 4554 298452 337554
rect 298412 4548 298464 4554
rect 298412 4490 298464 4496
rect 298516 4486 298544 337708
rect 298780 337690 298832 337696
rect 299068 337618 299096 340068
rect 299252 337686 299280 340068
rect 299542 340054 299648 340082
rect 299516 337748 299568 337754
rect 299516 337690 299568 337696
rect 299240 337680 299292 337686
rect 299240 337622 299292 337628
rect 299056 337612 299108 337618
rect 299056 337554 299108 337560
rect 299528 322250 299556 337690
rect 299516 322244 299568 322250
rect 299516 322186 299568 322192
rect 298594 38856 298650 38865
rect 298594 38791 298596 38800
rect 298648 38791 298650 38800
rect 298596 38762 298648 38768
rect 299620 18630 299648 340054
rect 299712 340054 299818 340082
rect 299608 18624 299660 18630
rect 299608 18566 299660 18572
rect 299712 4622 299740 340054
rect 299988 337686 300016 340068
rect 300264 337958 300292 340068
rect 300252 337952 300304 337958
rect 300252 337894 300304 337900
rect 299884 337680 299936 337686
rect 299884 337622 299936 337628
rect 299976 337680 300028 337686
rect 299976 337622 300028 337628
rect 299792 337612 299844 337618
rect 299792 337554 299844 337560
rect 299804 5302 299832 337554
rect 299792 5296 299844 5302
rect 299792 5238 299844 5244
rect 299896 4690 299924 337622
rect 300540 337074 300568 340068
rect 300724 337754 300752 340068
rect 300908 340054 301014 340082
rect 301092 340054 301290 340082
rect 300712 337748 300764 337754
rect 300712 337690 300764 337696
rect 300528 337068 300580 337074
rect 300528 337010 300580 337016
rect 300908 265674 300936 340054
rect 300988 337068 301040 337074
rect 300988 337010 301040 337016
rect 300896 265668 300948 265674
rect 300896 265610 300948 265616
rect 300434 226672 300490 226681
rect 300434 226607 300436 226616
rect 300488 226607 300490 226616
rect 300436 226578 300488 226584
rect 301000 5030 301028 337010
rect 301092 5370 301120 340054
rect 301172 337748 301224 337754
rect 301172 337690 301224 337696
rect 301080 5364 301132 5370
rect 301080 5306 301132 5312
rect 300988 5024 301040 5030
rect 300988 4966 301040 4972
rect 301184 4826 301212 337690
rect 301264 337680 301316 337686
rect 301264 337622 301316 337628
rect 301276 5166 301304 337622
rect 301460 337618 301488 340068
rect 301448 337612 301500 337618
rect 301448 337554 301500 337560
rect 301736 337210 301764 340068
rect 302012 337686 302040 340068
rect 302196 337754 302224 340068
rect 302380 340054 302486 340082
rect 302184 337748 302236 337754
rect 302184 337690 302236 337696
rect 302000 337680 302052 337686
rect 302000 337622 302052 337628
rect 301724 337204 301776 337210
rect 301724 337146 301776 337152
rect 302380 253230 302408 340054
rect 302460 337748 302512 337754
rect 302460 337690 302512 337696
rect 302368 253224 302420 253230
rect 302368 253166 302420 253172
rect 302472 6254 302500 337690
rect 302552 337680 302604 337686
rect 302552 337622 302604 337628
rect 302460 6248 302512 6254
rect 302460 6190 302512 6196
rect 301264 5160 301316 5166
rect 301264 5102 301316 5108
rect 302564 4865 302592 337622
rect 302644 337612 302696 337618
rect 302644 337554 302696 337560
rect 302656 5098 302684 337554
rect 302748 336326 302776 340068
rect 302932 337754 302960 340068
rect 303116 340054 303222 340082
rect 303498 340054 303604 340082
rect 303682 340054 303788 340082
rect 302920 337748 302972 337754
rect 302920 337690 302972 337696
rect 302736 336320 302788 336326
rect 302736 336262 302788 336268
rect 303116 333402 303144 340054
rect 303472 337952 303524 337958
rect 303472 337894 303524 337900
rect 303380 337544 303432 337550
rect 303380 337486 303432 337492
rect 303104 333396 303156 333402
rect 303104 333338 303156 333344
rect 303392 14482 303420 337486
rect 303484 294642 303512 337894
rect 303576 330682 303604 340054
rect 303564 330676 303616 330682
rect 303564 330618 303616 330624
rect 303472 294636 303524 294642
rect 303472 294578 303524 294584
rect 303380 14476 303432 14482
rect 303380 14418 303432 14424
rect 303760 9042 303788 340054
rect 303944 338094 303972 340068
rect 303932 338088 303984 338094
rect 303932 338030 303984 338036
rect 303932 337748 303984 337754
rect 303932 337690 303984 337696
rect 303748 9036 303800 9042
rect 303748 8978 303800 8984
rect 303944 8974 303972 337690
rect 304220 336122 304248 340068
rect 304404 337686 304432 340068
rect 304680 337754 304708 340068
rect 304970 340054 305076 340082
rect 304760 338020 304812 338026
rect 304760 337962 304812 337968
rect 304668 337748 304720 337754
rect 304668 337690 304720 337696
rect 304392 337680 304444 337686
rect 304392 337622 304444 337628
rect 304208 336116 304260 336122
rect 304208 336058 304260 336064
rect 304772 11762 304800 337962
rect 304944 337952 304996 337958
rect 304944 337894 304996 337900
rect 304956 335322 304984 337894
rect 305048 337736 305076 340054
rect 305140 337958 305168 340068
rect 305416 338026 305444 340068
rect 305404 338020 305456 338026
rect 305404 337962 305456 337968
rect 305128 337952 305180 337958
rect 305128 337894 305180 337900
rect 305220 337748 305272 337754
rect 305048 337708 305168 337736
rect 304956 335294 305076 335322
rect 305048 321586 305076 335294
rect 305140 327894 305168 337708
rect 305220 337690 305272 337696
rect 305128 327888 305180 327894
rect 305128 327830 305180 327836
rect 305048 321558 305168 321586
rect 305140 302274 305168 321558
rect 305232 314022 305260 337690
rect 305312 337680 305364 337686
rect 305312 337622 305364 337628
rect 305220 314016 305272 314022
rect 305220 313958 305272 313964
rect 305048 302246 305168 302274
rect 305048 302138 305076 302246
rect 305048 302110 305168 302138
rect 305140 282962 305168 302110
rect 305048 282934 305168 282962
rect 305048 282826 305076 282934
rect 305048 282798 305168 282826
rect 305140 263650 305168 282798
rect 305048 263622 305168 263650
rect 305048 259418 305076 263622
rect 305036 259412 305088 259418
rect 305036 259354 305088 259360
rect 305128 249824 305180 249830
rect 305128 249766 305180 249772
rect 305140 230489 305168 249766
rect 304942 230480 304998 230489
rect 304942 230415 304998 230424
rect 305126 230480 305182 230489
rect 305126 230415 305182 230424
rect 304956 225010 304984 230415
rect 304944 225004 304996 225010
rect 304944 224946 304996 224952
rect 304944 224868 304996 224874
rect 304944 224810 304996 224816
rect 304956 207754 304984 224810
rect 304956 207726 305168 207754
rect 305140 205578 305168 207726
rect 305048 205550 305168 205578
rect 305048 196058 305076 205550
rect 305048 196030 305260 196058
rect 305232 186386 305260 196030
rect 305036 186380 305088 186386
rect 305036 186322 305088 186328
rect 305220 186380 305272 186386
rect 305220 186322 305272 186328
rect 305048 186266 305076 186322
rect 305048 186238 305168 186266
rect 305140 178770 305168 186238
rect 304852 178764 304904 178770
rect 304852 178706 304904 178712
rect 305128 178764 305180 178770
rect 305128 178706 305180 178712
rect 304864 173913 304892 178706
rect 304850 173904 304906 173913
rect 304850 173839 304906 173848
rect 305126 173904 305182 173913
rect 305126 173839 305182 173848
rect 305140 164218 305168 173839
rect 305128 164212 305180 164218
rect 305128 164154 305180 164160
rect 305128 157344 305180 157350
rect 305128 157286 305180 157292
rect 305140 154578 305168 157286
rect 305140 154550 305260 154578
rect 305232 147694 305260 154550
rect 305036 147688 305088 147694
rect 305036 147630 305088 147636
rect 305220 147688 305272 147694
rect 305220 147630 305272 147636
rect 305048 138038 305076 147630
rect 305036 138032 305088 138038
rect 305036 137974 305088 137980
rect 305128 137964 305180 137970
rect 305128 137906 305180 137912
rect 305140 125594 305168 137906
rect 305128 125588 305180 125594
rect 305128 125530 305180 125536
rect 305128 118516 305180 118522
rect 305128 118458 305180 118464
rect 305140 115954 305168 118458
rect 305140 115926 305260 115954
rect 305232 109070 305260 115926
rect 305036 109064 305088 109070
rect 305036 109006 305088 109012
rect 305220 109064 305272 109070
rect 305220 109006 305272 109012
rect 305048 104854 305076 109006
rect 305036 104848 305088 104854
rect 305036 104790 305088 104796
rect 305128 99340 305180 99346
rect 305128 99282 305180 99288
rect 305140 86970 305168 99282
rect 305128 86964 305180 86970
rect 305128 86906 305180 86912
rect 305128 79892 305180 79898
rect 305128 79834 305180 79840
rect 305140 77330 305168 79834
rect 305140 77302 305260 77330
rect 305232 53122 305260 77302
rect 305140 53094 305260 53122
rect 305140 41426 305168 53094
rect 305140 41398 305260 41426
rect 305232 29050 305260 41398
rect 305140 29022 305260 29050
rect 305140 27606 305168 29022
rect 305128 27600 305180 27606
rect 305128 27542 305180 27548
rect 305128 18080 305180 18086
rect 305128 18022 305180 18028
rect 304760 11756 304812 11762
rect 304760 11698 304812 11704
rect 305140 9722 305168 18022
rect 305036 9716 305088 9722
rect 305036 9658 305088 9664
rect 305128 9716 305180 9722
rect 305128 9658 305180 9664
rect 303932 8968 303984 8974
rect 303932 8910 303984 8916
rect 305048 8430 305076 9658
rect 305036 8424 305088 8430
rect 305036 8366 305088 8372
rect 305324 8362 305352 337622
rect 305600 334762 305628 340068
rect 305876 337686 305904 340068
rect 305864 337680 305916 337686
rect 305864 337622 305916 337628
rect 306152 337618 306180 340068
rect 306350 340054 306548 340082
rect 306416 337748 306468 337754
rect 306416 337690 306468 337696
rect 306140 337612 306192 337618
rect 306140 337554 306192 337560
rect 306140 337000 306192 337006
rect 306140 336942 306192 336948
rect 305588 334756 305640 334762
rect 305588 334698 305640 334704
rect 306152 17270 306180 336942
rect 306140 17264 306192 17270
rect 306140 17206 306192 17212
rect 306428 8566 306456 337690
rect 306520 325106 306548 340054
rect 306612 337754 306640 340068
rect 306600 337748 306652 337754
rect 306600 337690 306652 337696
rect 306692 337680 306744 337686
rect 306692 337622 306744 337628
rect 306600 337612 306652 337618
rect 306600 337554 306652 337560
rect 306508 325100 306560 325106
rect 306508 325042 306560 325048
rect 306612 311302 306640 337554
rect 306600 311296 306652 311302
rect 306600 311238 306652 311244
rect 306416 8560 306468 8566
rect 306416 8502 306468 8508
rect 306704 8498 306732 337622
rect 306888 337550 306916 340068
rect 306876 337544 306928 337550
rect 306876 337486 306928 337492
rect 307072 332042 307100 340068
rect 307348 337754 307376 340068
rect 307336 337748 307388 337754
rect 307336 337690 307388 337696
rect 307624 336938 307652 340068
rect 307612 336932 307664 336938
rect 307612 336874 307664 336880
rect 307060 332036 307112 332042
rect 307060 331978 307112 331984
rect 306692 8492 306744 8498
rect 306692 8434 306744 8440
rect 305312 8356 305364 8362
rect 305312 8298 305364 8304
rect 307808 6186 307836 340068
rect 307980 337748 308032 337754
rect 307980 337690 308032 337696
rect 307888 336932 307940 336938
rect 307888 336874 307940 336880
rect 307900 297498 307928 336874
rect 307888 297492 307940 297498
rect 307888 297434 307940 297440
rect 307888 96620 307940 96626
rect 307888 96562 307940 96568
rect 307900 87009 307928 96562
rect 307886 87000 307942 87009
rect 307886 86935 307942 86944
rect 307992 8634 308020 337690
rect 308084 8838 308112 340068
rect 308360 337006 308388 340068
rect 308544 337414 308572 340068
rect 308834 340054 309032 340082
rect 308900 338156 308952 338162
rect 308900 338098 308952 338104
rect 308532 337408 308584 337414
rect 308532 337350 308584 337356
rect 308348 337000 308400 337006
rect 308348 336942 308400 336948
rect 308912 335322 308940 338098
rect 309004 337770 309032 340054
rect 309096 337958 309124 340068
rect 309294 340054 309492 340082
rect 309084 337952 309136 337958
rect 309084 337894 309136 337900
rect 309004 337742 309308 337770
rect 308912 335294 309032 335322
rect 309004 335186 309032 335294
rect 309004 335158 309216 335186
rect 309188 311846 309216 335158
rect 309176 311840 309228 311846
rect 309176 311782 309228 311788
rect 309176 309188 309228 309194
rect 309176 309130 309228 309136
rect 309188 299470 309216 309130
rect 309176 299464 309228 299470
rect 309176 299406 309228 299412
rect 309176 289876 309228 289882
rect 309176 289818 309228 289824
rect 309188 280090 309216 289818
rect 309176 280084 309228 280090
rect 309176 280026 309228 280032
rect 309176 270564 309228 270570
rect 309176 270506 309228 270512
rect 309188 259434 309216 270506
rect 309004 259406 309216 259434
rect 309004 253978 309032 259406
rect 308992 253972 309044 253978
rect 308992 253914 309044 253920
rect 309084 253904 309136 253910
rect 309084 253846 309136 253852
rect 309096 241482 309124 253846
rect 309096 241466 309216 241482
rect 309096 241460 309228 241466
rect 309096 241454 309176 241460
rect 309176 241402 309228 241408
rect 309176 234388 309228 234394
rect 309176 234330 309228 234336
rect 308164 226636 308216 226642
rect 308164 226578 308216 226584
rect 308176 226545 308204 226578
rect 308162 226536 308218 226545
rect 308162 226471 308218 226480
rect 309188 224890 309216 234330
rect 309096 224862 309216 224890
rect 309096 205766 309124 224862
rect 309084 205760 309136 205766
rect 309084 205702 309136 205708
rect 309084 205556 309136 205562
rect 309084 205498 309136 205504
rect 309096 196058 309124 205498
rect 309096 196030 309216 196058
rect 309188 193202 309216 196030
rect 309096 193174 309216 193202
rect 309096 186386 309124 193174
rect 309084 186380 309136 186386
rect 309084 186322 309136 186328
rect 308992 183592 309044 183598
rect 308992 183534 309044 183540
rect 308256 181484 308308 181490
rect 308256 181426 308308 181432
rect 308268 96626 308296 181426
rect 309004 173942 309032 183534
rect 308992 173936 309044 173942
rect 308992 173878 309044 173884
rect 309084 173936 309136 173942
rect 309084 173878 309136 173884
rect 309096 169130 309124 173878
rect 308912 169102 309124 169130
rect 308912 166954 308940 169102
rect 308912 166926 309032 166954
rect 309004 164218 309032 166926
rect 308992 164212 309044 164218
rect 308992 164154 309044 164160
rect 309084 164212 309136 164218
rect 309084 164154 309136 164160
rect 309096 157162 309124 164154
rect 309096 157134 309216 157162
rect 309188 151745 309216 157134
rect 309174 151736 309230 151745
rect 309174 151671 309230 151680
rect 309174 142216 309230 142225
rect 309096 142174 309174 142202
rect 309096 140758 309124 142174
rect 309174 142151 309230 142160
rect 309084 140752 309136 140758
rect 309084 140694 309136 140700
rect 309084 134700 309136 134706
rect 309084 134642 309136 134648
rect 309096 128466 309124 134642
rect 309004 128438 309124 128466
rect 309004 125594 309032 128438
rect 308992 125588 309044 125594
rect 308992 125530 309044 125536
rect 309176 119400 309228 119406
rect 309176 119342 309228 119348
rect 309188 106350 309216 119342
rect 309176 106344 309228 106350
rect 309176 106286 309228 106292
rect 309084 106276 309136 106282
rect 309084 106218 309136 106224
rect 309096 103494 309124 106218
rect 309084 103488 309136 103494
rect 309084 103430 309136 103436
rect 308256 96620 308308 96626
rect 308256 96562 308308 96568
rect 308900 93900 308952 93906
rect 308900 93842 308952 93848
rect 308912 87009 308940 93842
rect 308162 87000 308218 87009
rect 308898 87000 308954 87009
rect 308218 86958 308296 86986
rect 308162 86935 308218 86944
rect 308164 38820 308216 38826
rect 308164 38762 308216 38768
rect 308176 38729 308204 38762
rect 308162 38720 308218 38729
rect 308162 38655 308218 38664
rect 308268 19310 308296 86958
rect 308898 86935 308954 86944
rect 309082 87000 309138 87009
rect 309082 86935 309138 86944
rect 309096 80050 309124 86935
rect 309004 80022 309124 80050
rect 309004 70258 309032 80022
rect 309004 70230 309124 70258
rect 309096 66230 309124 70230
rect 309084 66224 309136 66230
rect 309084 66166 309136 66172
rect 308900 56704 308952 56710
rect 308900 56646 308952 56652
rect 308912 48362 308940 56646
rect 308912 48334 309032 48362
rect 309004 46918 309032 48334
rect 308992 46912 309044 46918
rect 308992 46854 309044 46860
rect 309176 46912 309228 46918
rect 309176 46854 309228 46860
rect 309188 29034 309216 46854
rect 308992 29028 309044 29034
rect 308992 28970 309044 28976
rect 309176 29028 309228 29034
rect 309176 28970 309228 28976
rect 309004 22114 309032 28970
rect 309004 22086 309216 22114
rect 308256 19304 308308 19310
rect 308256 19246 308308 19252
rect 308256 9716 308308 9722
rect 308256 9658 308308 9664
rect 308072 8832 308124 8838
rect 308072 8774 308124 8780
rect 307980 8628 308032 8634
rect 307980 8570 308032 8576
rect 307796 6180 307848 6186
rect 307796 6122 307848 6128
rect 302736 5160 302788 5166
rect 302736 5102 302788 5108
rect 307520 5160 307572 5166
rect 307520 5102 307572 5108
rect 302644 5092 302696 5098
rect 302644 5034 302696 5040
rect 302550 4856 302606 4865
rect 301172 4820 301224 4826
rect 302550 4791 302606 4800
rect 301172 4762 301224 4768
rect 299884 4684 299936 4690
rect 299884 4626 299936 4632
rect 299700 4616 299752 4622
rect 299700 4558 299752 4564
rect 302550 4584 302606 4593
rect 302550 4519 302552 4528
rect 302604 4519 302606 4528
rect 302552 4490 302604 4496
rect 298504 4480 298556 4486
rect 298504 4422 298556 4428
rect 302458 4448 302514 4457
rect 302458 4383 302514 4392
rect 302472 4214 302500 4383
rect 302644 4276 302696 4282
rect 302644 4218 302696 4224
rect 298320 4208 298372 4214
rect 298320 4150 298372 4156
rect 302460 4208 302512 4214
rect 302460 4150 302512 4156
rect 297216 4140 297268 4146
rect 297216 4082 297268 4088
rect 297124 3596 297176 3602
rect 297124 3538 297176 3544
rect 294364 3460 294416 3466
rect 294364 3402 294416 3408
rect 296020 3120 296072 3126
rect 296020 3062 296072 3068
rect 294180 3052 294232 3058
rect 294180 2994 294232 3000
rect 294824 2984 294876 2990
rect 294824 2926 294876 2932
rect 293812 2848 293864 2854
rect 293812 2790 293864 2796
rect 294836 480 294864 2926
rect 296032 480 296060 3062
rect 297228 480 297256 4082
rect 302552 4072 302604 4078
rect 302656 4060 302684 4218
rect 302748 4078 302776 5102
rect 307532 5030 307560 5102
rect 307520 5024 307572 5030
rect 302826 4992 302882 5001
rect 307520 4966 307572 4972
rect 302826 4927 302882 4936
rect 302840 4554 302868 4927
rect 303102 4584 303158 4593
rect 302828 4548 302880 4554
rect 303102 4519 303104 4528
rect 302828 4490 302880 4496
rect 303156 4519 303158 4528
rect 303104 4490 303156 4496
rect 303012 4480 303064 4486
rect 303010 4448 303012 4457
rect 303064 4448 303066 4457
rect 303010 4383 303066 4392
rect 305496 4140 305548 4146
rect 305496 4082 305548 4088
rect 302604 4032 302684 4060
rect 302736 4072 302788 4078
rect 302552 4014 302604 4020
rect 302736 4014 302788 4020
rect 304300 4004 304352 4010
rect 304300 3946 304352 3952
rect 298412 3936 298464 3942
rect 298412 3878 298464 3884
rect 298424 480 298452 3878
rect 299608 3732 299660 3738
rect 299608 3674 299660 3680
rect 299620 480 299648 3674
rect 300804 3528 300856 3534
rect 300804 3470 300856 3476
rect 300816 480 300844 3470
rect 303104 3392 303156 3398
rect 303104 3334 303156 3340
rect 301908 2916 301960 2922
rect 301908 2858 301960 2864
rect 301920 480 301948 2858
rect 303116 480 303144 3334
rect 304312 480 304340 3946
rect 305508 480 305536 4082
rect 307888 3596 307940 3602
rect 307888 3538 307940 3544
rect 306692 2916 306744 2922
rect 306692 2858 306744 2864
rect 306704 480 306732 2858
rect 307900 480 307928 3538
rect 308268 2854 308296 9658
rect 309188 9654 309216 22086
rect 309176 9648 309228 9654
rect 309176 9590 309228 9596
rect 309280 8906 309308 337742
rect 309360 337408 309412 337414
rect 309360 337350 309412 337356
rect 309268 8900 309320 8906
rect 309268 8842 309320 8848
rect 309372 6118 309400 337350
rect 309360 6112 309412 6118
rect 309360 6054 309412 6060
rect 309464 5574 309492 340054
rect 309556 338162 309584 340068
rect 309544 338156 309596 338162
rect 309544 338098 309596 338104
rect 309544 337952 309596 337958
rect 309544 337894 309596 337900
rect 309452 5568 309504 5574
rect 309452 5510 309504 5516
rect 309556 3602 309584 337894
rect 309832 337074 309860 340068
rect 310016 337754 310044 340068
rect 310004 337748 310056 337754
rect 310004 337690 310056 337696
rect 310292 337686 310320 340068
rect 310280 337680 310332 337686
rect 310280 337622 310332 337628
rect 310568 337550 310596 340068
rect 310648 337680 310700 337686
rect 310648 337622 310700 337628
rect 310556 337544 310608 337550
rect 310556 337486 310608 337492
rect 310280 337476 310332 337482
rect 310280 337418 310332 337424
rect 309820 337068 309872 337074
rect 309820 337010 309872 337016
rect 309634 242448 309690 242457
rect 309634 242383 309690 242392
rect 309648 241777 309676 242383
rect 309634 241768 309690 241777
rect 309634 241703 309690 241712
rect 309634 227216 309690 227225
rect 309634 227151 309690 227160
rect 309648 226545 309676 227151
rect 309634 226536 309690 226545
rect 309634 226471 309690 226480
rect 310292 8294 310320 337418
rect 310660 9586 310688 337622
rect 310648 9580 310700 9586
rect 310648 9522 310700 9528
rect 310280 8288 310332 8294
rect 310280 8230 310332 8236
rect 310752 6390 310780 340068
rect 310832 337748 310884 337754
rect 310832 337690 310884 337696
rect 310740 6384 310792 6390
rect 310740 6326 310792 6332
rect 310844 6322 310872 337690
rect 311028 337618 311056 340068
rect 311016 337612 311068 337618
rect 311016 337554 311068 337560
rect 311304 337550 311332 340068
rect 311488 337686 311516 340068
rect 311672 340054 311778 340082
rect 311476 337680 311528 337686
rect 311476 337622 311528 337628
rect 310924 337544 310976 337550
rect 310924 337486 310976 337492
rect 311292 337544 311344 337550
rect 311292 337486 311344 337492
rect 310832 6316 310884 6322
rect 310832 6258 310884 6264
rect 309544 3596 309596 3602
rect 309544 3538 309596 3544
rect 310936 3466 310964 337486
rect 311672 335322 311700 340054
rect 312040 337754 312068 340068
rect 312028 337748 312080 337754
rect 312028 337690 312080 337696
rect 312120 337680 312172 337686
rect 312120 337622 312172 337628
rect 312028 337612 312080 337618
rect 312028 337554 312080 337560
rect 311672 335294 311792 335322
rect 311764 335186 311792 335294
rect 311764 335158 311976 335186
rect 311948 319598 311976 335158
rect 311936 319592 311988 319598
rect 311936 319534 311988 319540
rect 312040 9518 312068 337554
rect 312028 9512 312080 9518
rect 312028 9454 312080 9460
rect 312132 5914 312160 337622
rect 312224 5914 312252 340068
rect 312304 337748 312356 337754
rect 312304 337690 312356 337696
rect 312120 5908 312172 5914
rect 312120 5850 312172 5856
rect 312212 5908 312264 5914
rect 312212 5850 312264 5856
rect 312316 5794 312344 337690
rect 312500 336870 312528 340068
rect 312776 337414 312804 340068
rect 312974 340054 313172 340082
rect 313250 340054 313448 340082
rect 312764 337408 312816 337414
rect 312764 337350 312816 337356
rect 313040 337204 313092 337210
rect 313040 337146 313092 337152
rect 312488 336864 312540 336870
rect 312488 336806 312540 336812
rect 313052 21418 313080 337146
rect 313144 335510 313172 340054
rect 313316 336864 313368 336870
rect 313316 336806 313368 336812
rect 313132 335504 313184 335510
rect 313132 335446 313184 335452
rect 313328 323610 313356 336806
rect 313316 323604 313368 323610
rect 313316 323546 313368 323552
rect 313420 312662 313448 340054
rect 313512 336870 313540 340068
rect 313604 340054 313710 340082
rect 313500 336864 313552 336870
rect 313500 336806 313552 336812
rect 313604 335594 313632 340054
rect 313684 337408 313736 337414
rect 313684 337350 313736 337356
rect 313696 337210 313724 337350
rect 313684 337204 313736 337210
rect 313684 337146 313736 337152
rect 313972 336938 314000 340068
rect 314248 337550 314276 340068
rect 314236 337544 314288 337550
rect 314236 337486 314288 337492
rect 314144 337136 314196 337142
rect 314144 337078 314196 337084
rect 313960 336932 314012 336938
rect 313960 336874 314012 336880
rect 313684 336864 313736 336870
rect 313684 336806 313736 336812
rect 313512 335566 313632 335594
rect 313408 312656 313460 312662
rect 313408 312598 313460 312604
rect 313040 21412 313092 21418
rect 313040 21354 313092 21360
rect 312672 8288 312724 8294
rect 312672 8230 312724 8236
rect 311948 5766 312344 5794
rect 311476 3732 311528 3738
rect 311476 3674 311528 3680
rect 310280 3460 310332 3466
rect 310280 3402 310332 3408
rect 310924 3460 310976 3466
rect 310924 3402 310976 3408
rect 308256 2848 308308 2854
rect 308256 2790 308308 2796
rect 309084 604 309136 610
rect 309084 546 309136 552
rect 309096 480 309124 546
rect 310292 480 310320 3402
rect 311488 480 311516 3674
rect 311948 2854 311976 5766
rect 312028 5636 312080 5642
rect 312028 5578 312080 5584
rect 312040 5386 312068 5578
rect 312040 5358 312344 5386
rect 312212 5092 312264 5098
rect 312212 5034 312264 5040
rect 312224 5001 312252 5034
rect 312210 4992 312266 5001
rect 312210 4927 312266 4936
rect 312316 4690 312344 5358
rect 312580 5296 312632 5302
rect 312578 5264 312580 5273
rect 312632 5264 312634 5273
rect 312578 5199 312634 5208
rect 312304 4684 312356 4690
rect 312304 4626 312356 4632
rect 311936 2848 311988 2854
rect 311936 2790 311988 2796
rect 312684 480 312712 8230
rect 313512 6866 313540 335566
rect 313592 335504 313644 335510
rect 313592 335446 313644 335452
rect 313500 6860 313552 6866
rect 313500 6802 313552 6808
rect 313604 6458 313632 335446
rect 313592 6452 313644 6458
rect 313592 6394 313644 6400
rect 313696 2922 313724 336806
rect 313868 3664 313920 3670
rect 313868 3606 313920 3612
rect 313684 2916 313736 2922
rect 313684 2858 313736 2864
rect 313880 480 313908 3606
rect 314156 2836 314184 337078
rect 314432 336870 314460 340068
rect 314722 340054 314920 340082
rect 314998 340054 315104 340082
rect 314788 336932 314840 336938
rect 314788 336874 314840 336880
rect 314420 336864 314472 336870
rect 314420 336806 314472 336812
rect 314800 318170 314828 336874
rect 314788 318164 314840 318170
rect 314788 318106 314840 318112
rect 314892 286414 314920 340054
rect 314972 336864 315024 336870
rect 314972 336806 315024 336812
rect 314880 286408 314932 286414
rect 314880 286350 314932 286356
rect 314984 6798 315012 336806
rect 314972 6792 315024 6798
rect 314972 6734 315024 6740
rect 315076 2990 315104 340054
rect 315168 337006 315196 340068
rect 315156 337000 315208 337006
rect 315156 336942 315208 336948
rect 315444 336870 315472 340068
rect 315720 337414 315748 340068
rect 315708 337408 315760 337414
rect 315708 337350 315760 337356
rect 315904 336938 315932 340068
rect 315892 336932 315944 336938
rect 315892 336874 315944 336880
rect 315432 336864 315484 336870
rect 315432 336806 315484 336812
rect 316076 336864 316128 336870
rect 316076 336806 316128 336812
rect 316088 315382 316116 336806
rect 316076 315376 316128 315382
rect 316076 315318 316128 315324
rect 316180 283694 316208 340068
rect 316352 337000 316404 337006
rect 316352 336942 316404 336948
rect 316260 336932 316312 336938
rect 316260 336874 316312 336880
rect 316168 283688 316220 283694
rect 316168 283630 316220 283636
rect 316168 11824 316220 11830
rect 316168 11766 316220 11772
rect 316180 6474 316208 11766
rect 316272 6662 316300 336874
rect 316364 6730 316392 336942
rect 316352 6724 316404 6730
rect 316352 6666 316404 6672
rect 316260 6656 316312 6662
rect 316260 6598 316312 6604
rect 316180 6446 316300 6474
rect 315064 2984 315116 2990
rect 315064 2926 315116 2932
rect 314156 2808 315104 2836
rect 315076 480 315104 2808
rect 316272 480 316300 6446
rect 316456 3058 316484 340068
rect 316640 337006 316668 340068
rect 316628 337000 316680 337006
rect 316628 336942 316680 336948
rect 316916 336870 316944 340068
rect 317192 336938 317220 340068
rect 317180 336932 317232 336938
rect 317180 336874 317232 336880
rect 317376 336870 317404 340068
rect 317560 340054 317666 340082
rect 317942 340054 318048 340082
rect 316904 336864 316956 336870
rect 316904 336806 316956 336812
rect 317272 336864 317324 336870
rect 317272 336806 317324 336812
rect 317364 336864 317416 336870
rect 317364 336806 317416 336812
rect 317284 335594 317312 336806
rect 317284 335566 317496 335594
rect 317468 316742 317496 335566
rect 317456 316736 317508 316742
rect 317456 316678 317508 316684
rect 317560 10538 317588 340054
rect 317640 337000 317692 337006
rect 317640 336942 317692 336948
rect 317548 10532 317600 10538
rect 317548 10474 317600 10480
rect 317652 7274 317680 336942
rect 317824 336932 317876 336938
rect 317824 336874 317876 336880
rect 317732 336864 317784 336870
rect 317732 336806 317784 336812
rect 317640 7268 317692 7274
rect 317640 7210 317692 7216
rect 317744 6458 317772 336806
rect 317732 6452 317784 6458
rect 317732 6394 317784 6400
rect 317454 5264 317510 5273
rect 317454 5199 317510 5208
rect 316444 3052 316496 3058
rect 316444 2994 316496 3000
rect 317468 480 317496 5199
rect 317836 3126 317864 336874
rect 318020 335510 318048 340054
rect 318112 336870 318140 340068
rect 318388 337074 318416 340068
rect 318376 337068 318428 337074
rect 318376 337010 318428 337016
rect 318664 337006 318692 340068
rect 318862 340054 319060 340082
rect 318836 337068 318888 337074
rect 318836 337010 318888 337016
rect 318652 337000 318704 337006
rect 318652 336942 318704 336948
rect 318100 336864 318152 336870
rect 318100 336806 318152 336812
rect 318650 335744 318706 335753
rect 318650 335679 318706 335688
rect 318008 335504 318060 335510
rect 318008 335446 318060 335452
rect 318664 328438 318692 335679
rect 318652 328432 318704 328438
rect 318652 328374 318704 328380
rect 318652 321428 318704 321434
rect 318652 321370 318704 321376
rect 318664 318866 318692 321370
rect 318664 318838 318784 318866
rect 318756 311982 318784 318838
rect 318744 311976 318796 311982
rect 318744 311918 318796 311924
rect 318744 311840 318796 311846
rect 318744 311782 318796 311788
rect 318756 282962 318784 311782
rect 318664 282934 318784 282962
rect 318664 282826 318692 282934
rect 318664 282798 318784 282826
rect 318756 263650 318784 282798
rect 318664 263622 318784 263650
rect 318664 263514 318692 263622
rect 318664 263486 318784 263514
rect 318756 244338 318784 263486
rect 318664 244310 318784 244338
rect 318664 244202 318692 244310
rect 318664 244174 318784 244202
rect 318756 225026 318784 244174
rect 318664 224998 318784 225026
rect 318664 224890 318692 224998
rect 318664 224862 318784 224890
rect 318756 205714 318784 224862
rect 318664 205686 318784 205714
rect 318664 205578 318692 205686
rect 318664 205550 318784 205578
rect 318756 186402 318784 205550
rect 318664 186374 318784 186402
rect 318664 186266 318692 186374
rect 318664 186238 318784 186266
rect 318756 167090 318784 186238
rect 318664 167062 318784 167090
rect 318664 166954 318692 167062
rect 318664 166926 318784 166954
rect 318756 147778 318784 166926
rect 318664 147750 318784 147778
rect 318664 147642 318692 147750
rect 318664 147614 318784 147642
rect 318756 128466 318784 147614
rect 318664 128438 318784 128466
rect 318664 128330 318692 128438
rect 318664 128302 318784 128330
rect 318756 109154 318784 128302
rect 318664 109126 318784 109154
rect 318664 109018 318692 109126
rect 318664 108990 318784 109018
rect 318756 89842 318784 108990
rect 318664 89814 318784 89842
rect 318664 89706 318692 89814
rect 318664 89678 318784 89706
rect 318756 70394 318784 89678
rect 318664 70366 318784 70394
rect 318664 70258 318692 70366
rect 318664 70230 318784 70258
rect 318756 51082 318784 70230
rect 318664 51054 318784 51082
rect 318664 50946 318692 51054
rect 318664 50918 318784 50946
rect 318756 31770 318784 50918
rect 318664 31742 318784 31770
rect 318664 31634 318692 31742
rect 318664 31606 318784 31634
rect 318756 12458 318784 31606
rect 318664 12430 318784 12458
rect 318664 10470 318692 12430
rect 318848 10606 318876 337010
rect 318928 336864 318980 336870
rect 318928 336806 318980 336812
rect 318940 318714 318968 336806
rect 319032 318753 319060 340054
rect 319124 335753 319152 340068
rect 319414 340054 319520 340082
rect 319204 337000 319256 337006
rect 319204 336942 319256 336948
rect 319110 335744 319166 335753
rect 319110 335679 319166 335688
rect 319216 335594 319244 336942
rect 319124 335566 319244 335594
rect 319018 318744 319074 318753
rect 318928 318708 318980 318714
rect 319124 318714 319152 335566
rect 319492 335510 319520 340054
rect 319584 336938 319612 340068
rect 319572 336932 319624 336938
rect 319572 336874 319624 336880
rect 319676 336870 319704 340190
rect 320136 337006 320164 340068
rect 320334 340054 320440 340082
rect 320124 337000 320176 337006
rect 320124 336942 320176 336948
rect 320308 336932 320360 336938
rect 320308 336874 320360 336880
rect 319664 336864 319716 336870
rect 320032 336864 320084 336870
rect 319664 336806 319716 336812
rect 319952 336824 320032 336852
rect 319204 335504 319256 335510
rect 319204 335446 319256 335452
rect 319480 335504 319532 335510
rect 319480 335446 319532 335452
rect 319018 318679 319074 318688
rect 319112 318708 319164 318714
rect 318928 318650 318980 318656
rect 319112 318650 319164 318656
rect 319216 318646 319244 335446
rect 319952 335306 319980 336824
rect 320032 336806 320084 336812
rect 320216 336864 320268 336870
rect 320216 336806 320268 336812
rect 319940 335300 319992 335306
rect 319940 335242 319992 335248
rect 319204 318640 319256 318646
rect 319204 318582 319256 318588
rect 319204 318504 319256 318510
rect 318926 318472 318982 318481
rect 319204 318446 319256 318452
rect 318926 318407 318982 318416
rect 318940 314242 318968 318407
rect 318940 314214 319060 314242
rect 318928 314084 318980 314090
rect 318928 314026 318980 314032
rect 318836 10600 318888 10606
rect 318836 10542 318888 10548
rect 318652 10464 318704 10470
rect 318652 10406 318704 10412
rect 318940 6497 318968 314026
rect 318926 6488 318982 6497
rect 318926 6423 318982 6432
rect 318836 6384 318888 6390
rect 318834 6352 318836 6361
rect 318888 6352 318890 6361
rect 319032 6322 319060 314214
rect 319112 309868 319164 309874
rect 319112 309810 319164 309816
rect 318834 6287 318890 6296
rect 319020 6316 319072 6322
rect 319020 6258 319072 6264
rect 318560 3528 318612 3534
rect 318560 3470 318612 3476
rect 317824 3120 317876 3126
rect 317824 3062 317876 3068
rect 318572 480 318600 3470
rect 319124 3398 319152 309810
rect 319112 3392 319164 3398
rect 319112 3334 319164 3340
rect 319216 3194 319244 318446
rect 320124 317484 320176 317490
rect 320124 317426 320176 317432
rect 320136 307834 320164 317426
rect 319940 307828 319992 307834
rect 319940 307770 319992 307776
rect 320124 307828 320176 307834
rect 320124 307770 320176 307776
rect 319952 298042 319980 307770
rect 319940 298036 319992 298042
rect 319940 297978 319992 297984
rect 320124 292460 320176 292466
rect 320124 292402 320176 292408
rect 320136 282985 320164 292402
rect 320122 282976 320178 282985
rect 320122 282911 320178 282920
rect 320030 278896 320086 278905
rect 320030 278831 320086 278840
rect 320044 273306 320072 278831
rect 319952 273278 320072 273306
rect 319952 272762 319980 273278
rect 319952 272734 320164 272762
rect 320136 267730 320164 272734
rect 320044 267702 320164 267730
rect 320044 263634 320072 267702
rect 320032 263628 320084 263634
rect 320032 263570 320084 263576
rect 320032 258120 320084 258126
rect 320032 258062 320084 258068
rect 320044 251161 320072 258062
rect 320030 251152 320086 251161
rect 320030 251087 320086 251096
rect 320030 241632 320086 241641
rect 320030 241567 320086 241576
rect 320044 235362 320072 241567
rect 319952 235334 320072 235362
rect 319952 234394 319980 235334
rect 319940 234388 319992 234394
rect 319940 234330 319992 234336
rect 320124 234388 320176 234394
rect 320124 234330 320176 234336
rect 320136 230466 320164 234330
rect 320044 230438 320164 230466
rect 320044 225010 320072 230438
rect 320032 225004 320084 225010
rect 320032 224946 320084 224952
rect 320032 220992 320084 220998
rect 320032 220934 320084 220940
rect 320044 216073 320072 220934
rect 320030 216064 320086 216073
rect 320030 215999 320086 216008
rect 320030 206272 320086 206281
rect 320030 206207 320086 206216
rect 320044 200122 320072 206207
rect 320032 200116 320084 200122
rect 320032 200058 320084 200064
rect 320032 195968 320084 195974
rect 320032 195910 320084 195916
rect 320044 190482 320072 195910
rect 320044 190454 320164 190482
rect 320136 186946 320164 190454
rect 319952 186918 320164 186946
rect 319952 186266 319980 186918
rect 319952 186238 320072 186266
rect 320044 177274 320072 186238
rect 319756 177268 319808 177274
rect 319756 177210 319808 177216
rect 320032 177268 320084 177274
rect 320032 177210 320084 177216
rect 319768 172553 319796 177210
rect 319754 172544 319810 172553
rect 319754 172479 319810 172488
rect 319938 172544 319994 172553
rect 319938 172479 319994 172488
rect 319952 168994 319980 172479
rect 319952 168966 320072 168994
rect 320044 164150 320072 168966
rect 320032 164144 320084 164150
rect 320032 164086 320084 164092
rect 320124 164144 320176 164150
rect 320124 164086 320176 164092
rect 320136 158030 320164 164086
rect 319848 158024 319900 158030
rect 319848 157966 319900 157972
rect 320124 158024 320176 158030
rect 320124 157966 320176 157972
rect 319860 153241 319888 157966
rect 319846 153232 319902 153241
rect 319846 153167 319902 153176
rect 320030 153232 320086 153241
rect 320030 153167 320086 153176
rect 320044 145042 320072 153167
rect 320032 145036 320084 145042
rect 320032 144978 320084 144984
rect 320124 145036 320176 145042
rect 320124 144978 320176 144984
rect 320136 143546 320164 144978
rect 320124 143540 320176 143546
rect 320124 143482 320176 143488
rect 319940 133952 319992 133958
rect 319940 133894 319992 133900
rect 319952 114578 319980 133894
rect 319940 114572 319992 114578
rect 319940 114514 319992 114520
rect 320124 114572 320176 114578
rect 320124 114514 320176 114520
rect 320136 109070 320164 114514
rect 320124 109064 320176 109070
rect 320124 109006 320176 109012
rect 320124 104916 320176 104922
rect 320124 104858 320176 104864
rect 320136 103494 320164 104858
rect 320124 103488 320176 103494
rect 320124 103430 320176 103436
rect 319940 93900 319992 93906
rect 319940 93842 319992 93848
rect 319952 85542 319980 93842
rect 319940 85536 319992 85542
rect 319940 85478 319992 85484
rect 320124 75948 320176 75954
rect 320124 75890 320176 75896
rect 320136 66230 320164 75890
rect 320124 66224 320176 66230
rect 320124 66166 320176 66172
rect 320124 56704 320176 56710
rect 320124 56646 320176 56652
rect 320136 56545 320164 56646
rect 319846 56536 319902 56545
rect 319846 56471 319902 56480
rect 320122 56536 320178 56545
rect 320122 56471 320178 56480
rect 319860 47054 319888 56471
rect 319848 47048 319900 47054
rect 319848 46990 319900 46996
rect 320032 47048 320084 47054
rect 320032 46990 320084 46996
rect 320044 46918 320072 46990
rect 320032 46912 320084 46918
rect 320032 46854 320084 46860
rect 319940 37324 319992 37330
rect 319940 37266 319992 37272
rect 319952 24206 319980 37266
rect 319940 24200 319992 24206
rect 319940 24142 319992 24148
rect 320124 24200 320176 24206
rect 320124 24142 320176 24148
rect 320136 9722 320164 24142
rect 320228 9926 320256 336806
rect 320320 38554 320348 336874
rect 320308 38548 320360 38554
rect 320308 38490 320360 38496
rect 320308 31884 320360 31890
rect 320308 31826 320360 31832
rect 320216 9920 320268 9926
rect 320216 9862 320268 9868
rect 320124 9716 320176 9722
rect 320124 9658 320176 9664
rect 320320 7206 320348 31826
rect 320308 7200 320360 7206
rect 320308 7142 320360 7148
rect 320412 6225 320440 340054
rect 320492 337000 320544 337006
rect 320492 336942 320544 336948
rect 320504 335594 320532 336942
rect 320596 336870 320624 340068
rect 320780 337006 320808 340068
rect 321056 337074 321084 340068
rect 321044 337068 321096 337074
rect 321044 337010 321096 337016
rect 320768 337000 320820 337006
rect 320768 336942 320820 336948
rect 321332 336938 321360 340068
rect 321320 336932 321372 336938
rect 321320 336874 321372 336880
rect 321516 336870 321544 340068
rect 321700 340054 321806 340082
rect 322082 340054 322188 340082
rect 321596 337068 321648 337074
rect 321596 337010 321648 337016
rect 320584 336864 320636 336870
rect 320584 336806 320636 336812
rect 321504 336864 321556 336870
rect 321504 336806 321556 336812
rect 320504 335566 320624 335594
rect 320492 335504 320544 335510
rect 320492 335446 320544 335452
rect 320398 6216 320454 6225
rect 320398 6151 320454 6160
rect 319756 4140 319808 4146
rect 319756 4082 319808 4088
rect 319204 3188 319256 3194
rect 319204 3130 319256 3136
rect 319768 480 319796 4082
rect 320504 3942 320532 335446
rect 320596 4146 320624 335566
rect 321608 309874 321636 337010
rect 321596 309868 321648 309874
rect 321596 309810 321648 309816
rect 321700 307154 321728 340054
rect 321964 337000 322016 337006
rect 321964 336942 322016 336948
rect 321780 336932 321832 336938
rect 321780 336874 321832 336880
rect 321688 307148 321740 307154
rect 321688 307090 321740 307096
rect 321792 9994 321820 336874
rect 321872 336864 321924 336870
rect 321872 336806 321924 336812
rect 321780 9988 321832 9994
rect 321780 9930 321832 9936
rect 321884 8378 321912 336806
rect 321792 8350 321912 8378
rect 320584 4140 320636 4146
rect 320584 4082 320636 4088
rect 320952 4072 321004 4078
rect 320952 4014 321004 4020
rect 320492 3936 320544 3942
rect 320492 3878 320544 3884
rect 320964 480 320992 4014
rect 321792 3534 321820 8350
rect 321976 8242 322004 336942
rect 322160 335510 322188 340054
rect 322252 336870 322280 340068
rect 322240 336864 322292 336870
rect 322240 336806 322292 336812
rect 322148 335504 322200 335510
rect 322148 335446 322200 335452
rect 322528 329254 322556 340068
rect 322804 336938 322832 340068
rect 322792 336932 322844 336938
rect 322792 336874 322844 336880
rect 322988 336870 323016 340068
rect 323080 340054 323278 340082
rect 322884 336864 322936 336870
rect 322884 336806 322936 336812
rect 322976 336864 323028 336870
rect 322976 336806 323028 336812
rect 322516 329248 322568 329254
rect 322516 329190 322568 329196
rect 322056 14476 322108 14482
rect 322056 14418 322108 14424
rect 321884 8214 322004 8242
rect 321884 4010 321912 8214
rect 321962 6352 322018 6361
rect 321962 6287 322018 6296
rect 321976 6118 322004 6287
rect 321964 6112 322016 6118
rect 321964 6054 322016 6060
rect 321964 4820 322016 4826
rect 321964 4762 322016 4768
rect 321976 4729 322004 4762
rect 321962 4720 322018 4729
rect 321962 4655 322018 4664
rect 321872 4004 321924 4010
rect 321872 3946 321924 3952
rect 321780 3528 321832 3534
rect 321780 3470 321832 3476
rect 322068 626 322096 14418
rect 322896 8106 322924 336806
rect 323080 335594 323108 340054
rect 323540 336938 323568 340068
rect 323160 336932 323212 336938
rect 323160 336874 323212 336880
rect 323528 336932 323580 336938
rect 323528 336874 323580 336880
rect 322988 335566 323108 335594
rect 322988 304366 323016 335566
rect 323068 335504 323120 335510
rect 323068 335446 323120 335452
rect 322976 304360 323028 304366
rect 322976 304302 323028 304308
rect 323080 10742 323108 335446
rect 323172 11014 323200 336874
rect 323724 336870 323752 340068
rect 323252 336864 323304 336870
rect 323252 336806 323304 336812
rect 323712 336864 323764 336870
rect 323712 336806 323764 336812
rect 323160 11008 323212 11014
rect 323160 10950 323212 10956
rect 323068 10736 323120 10742
rect 323068 10678 323120 10684
rect 322896 8078 323016 8106
rect 322240 6928 322292 6934
rect 322240 6870 322292 6876
rect 322252 6361 322280 6870
rect 322238 6352 322294 6361
rect 322238 6287 322294 6296
rect 322148 4820 322200 4826
rect 322148 4762 322200 4768
rect 322160 4729 322188 4762
rect 322146 4720 322202 4729
rect 322146 4655 322202 4664
rect 322988 3942 323016 8078
rect 322976 3936 323028 3942
rect 322976 3878 323028 3884
rect 323264 3670 323292 336806
rect 324000 336054 324028 340068
rect 324290 340054 324396 340082
rect 324474 340054 324672 340082
rect 324368 337056 324396 340054
rect 324368 337028 324580 337056
rect 324448 336932 324500 336938
rect 324448 336874 324500 336880
rect 324172 336864 324224 336870
rect 324172 336806 324224 336812
rect 324264 336864 324316 336870
rect 324264 336806 324316 336812
rect 323988 336048 324040 336054
rect 323988 335990 324040 335996
rect 324184 331242 324212 336806
rect 324276 333010 324304 336806
rect 324276 332982 324396 333010
rect 324184 331214 324304 331242
rect 323344 4208 323396 4214
rect 323344 4150 323396 4156
rect 323252 3664 323304 3670
rect 323252 3606 323304 3612
rect 322068 598 322188 626
rect 322160 480 322188 598
rect 323356 480 323384 4150
rect 324276 3942 324304 331214
rect 324368 301578 324396 332982
rect 324356 301572 324408 301578
rect 324356 301514 324408 301520
rect 324460 10674 324488 336874
rect 324448 10668 324500 10674
rect 324448 10610 324500 10616
rect 324552 10062 324580 337028
rect 324540 10056 324592 10062
rect 324540 9998 324592 10004
rect 324540 4276 324592 4282
rect 324540 4218 324592 4224
rect 324264 3936 324316 3942
rect 324264 3878 324316 3884
rect 324552 480 324580 4218
rect 324644 3738 324672 340054
rect 324736 336870 324764 340068
rect 325012 336870 325040 340068
rect 325196 336938 325224 340068
rect 325184 336932 325236 336938
rect 325184 336874 325236 336880
rect 324724 336864 324776 336870
rect 324724 336806 324776 336812
rect 325000 336864 325052 336870
rect 325000 336806 325052 336812
rect 325472 335322 325500 340068
rect 325762 340054 325868 340082
rect 325946 340054 326052 340082
rect 325736 336864 325788 336870
rect 325736 336806 325788 336812
rect 325748 335458 325776 336806
rect 325840 335594 325868 340054
rect 325840 335566 325960 335594
rect 325748 335430 325868 335458
rect 325472 335294 325776 335322
rect 325748 300218 325776 335294
rect 325736 300212 325788 300218
rect 325736 300154 325788 300160
rect 324816 11756 324868 11762
rect 324816 11698 324868 11704
rect 324632 3732 324684 3738
rect 324632 3674 324684 3680
rect 324828 610 324856 11698
rect 325840 10198 325868 335430
rect 325828 10192 325880 10198
rect 325828 10134 325880 10140
rect 325932 10130 325960 335566
rect 325920 10124 325972 10130
rect 325920 10066 325972 10072
rect 326024 4049 326052 340054
rect 326104 336932 326156 336938
rect 326104 336874 326156 336880
rect 326010 4040 326066 4049
rect 326010 3975 326066 3984
rect 326116 3534 326144 336874
rect 326208 336870 326236 340068
rect 326484 337006 326512 340068
rect 326668 337074 326696 340068
rect 326656 337068 326708 337074
rect 326656 337010 326708 337016
rect 326472 337000 326524 337006
rect 326472 336942 326524 336948
rect 326944 336938 326972 340068
rect 327128 340054 327234 340082
rect 327418 340054 327524 340082
rect 327694 340054 327892 340082
rect 326932 336932 326984 336938
rect 326932 336874 326984 336880
rect 326196 336864 326248 336870
rect 326196 336806 326248 336812
rect 327024 336864 327076 336870
rect 327024 336806 327076 336812
rect 327036 326534 327064 336806
rect 327024 326528 327076 326534
rect 327024 326470 327076 326476
rect 327128 10266 327156 340054
rect 327392 337068 327444 337074
rect 327392 337010 327444 337016
rect 327208 337000 327260 337006
rect 327208 336942 327260 336948
rect 327220 10810 327248 336942
rect 327300 336932 327352 336938
rect 327300 336874 327352 336880
rect 327208 10804 327260 10810
rect 327208 10746 327260 10752
rect 327116 10260 327168 10266
rect 327116 10202 327168 10208
rect 327312 7818 327340 336874
rect 327300 7812 327352 7818
rect 327300 7754 327352 7760
rect 326932 4480 326984 4486
rect 326932 4422 326984 4428
rect 326104 3528 326156 3534
rect 326104 3470 326156 3476
rect 324816 604 324868 610
rect 324816 546 324868 552
rect 325736 604 325788 610
rect 325736 546 325788 552
rect 325748 480 325776 546
rect 326944 480 326972 4422
rect 327404 3913 327432 337010
rect 327390 3904 327446 3913
rect 327390 3839 327446 3848
rect 327496 3777 327524 340054
rect 327864 335578 327892 340054
rect 327956 336870 327984 340068
rect 328140 337006 328168 340068
rect 328430 340054 328628 340082
rect 328128 337000 328180 337006
rect 328128 336942 328180 336948
rect 327944 336864 327996 336870
rect 327944 336806 327996 336812
rect 328496 336864 328548 336870
rect 328496 336806 328548 336812
rect 328220 335776 328272 335782
rect 328220 335718 328272 335724
rect 327852 335572 327904 335578
rect 327852 335514 327904 335520
rect 328232 328438 328260 335718
rect 328128 328432 328180 328438
rect 328128 328374 328180 328380
rect 328220 328432 328272 328438
rect 328220 328374 328272 328380
rect 328140 327078 328168 328374
rect 328128 327072 328180 327078
rect 328128 327014 328180 327020
rect 328404 317484 328456 317490
rect 328404 317426 328456 317432
rect 328416 317370 328444 317426
rect 328232 317342 328444 317370
rect 328232 288561 328260 317342
rect 328218 288552 328274 288561
rect 328218 288487 328274 288496
rect 328402 288552 328458 288561
rect 328402 288487 328458 288496
rect 328416 288402 328444 288487
rect 328324 288374 328444 288402
rect 328324 277386 328352 288374
rect 328324 277358 328444 277386
rect 328416 276010 328444 277358
rect 328220 276004 328272 276010
rect 328220 275946 328272 275952
rect 328404 276004 328456 276010
rect 328404 275946 328456 275952
rect 328232 266393 328260 275946
rect 328218 266384 328274 266393
rect 328218 266319 328274 266328
rect 328402 266384 328458 266393
rect 328402 266319 328458 266328
rect 328416 263702 328444 266319
rect 328404 263696 328456 263702
rect 328404 263638 328456 263644
rect 328312 263560 328364 263566
rect 328312 263502 328364 263508
rect 328324 256698 328352 263502
rect 328312 256692 328364 256698
rect 328312 256634 328364 256640
rect 328312 253904 328364 253910
rect 328312 253846 328364 253852
rect 328324 247058 328352 253846
rect 328324 247030 328444 247058
rect 328416 243506 328444 247030
rect 328312 243500 328364 243506
rect 328312 243442 328364 243448
rect 328404 243500 328456 243506
rect 328404 243442 328456 243448
rect 328324 235958 328352 243442
rect 328312 235952 328364 235958
rect 328312 235894 328364 235900
rect 328312 211200 328364 211206
rect 328364 211148 328444 211154
rect 328312 211142 328444 211148
rect 328324 211126 328444 211142
rect 328416 209778 328444 211126
rect 328404 209772 328456 209778
rect 328404 209714 328456 209720
rect 328404 204944 328456 204950
rect 328404 204886 328456 204892
rect 328416 200054 328444 204886
rect 328404 200048 328456 200054
rect 328404 199990 328456 199996
rect 328404 195764 328456 195770
rect 328404 195706 328456 195712
rect 328416 186946 328444 195706
rect 328232 186918 328444 186946
rect 328232 186266 328260 186918
rect 328232 186238 328352 186266
rect 328324 182170 328352 186238
rect 328312 182164 328364 182170
rect 328312 182106 328364 182112
rect 328404 176588 328456 176594
rect 328404 176530 328456 176536
rect 328416 164234 328444 176530
rect 328324 164206 328444 164234
rect 328324 164098 328352 164206
rect 328324 164070 328444 164098
rect 328416 147744 328444 164070
rect 328324 147716 328444 147744
rect 328324 145042 328352 147716
rect 328312 145036 328364 145042
rect 328312 144978 328364 144984
rect 328404 145036 328456 145042
rect 328404 144978 328456 144984
rect 328416 143546 328444 144978
rect 328404 143540 328456 143546
rect 328404 143482 328456 143488
rect 328404 133952 328456 133958
rect 328404 133894 328456 133900
rect 328416 130234 328444 133894
rect 328232 130206 328444 130234
rect 328232 115977 328260 130206
rect 328218 115968 328274 115977
rect 328218 115903 328274 115912
rect 328402 115968 328458 115977
rect 328402 115903 328458 115912
rect 328416 109070 328444 115903
rect 328404 109064 328456 109070
rect 328404 109006 328456 109012
rect 328404 104916 328456 104922
rect 328404 104858 328456 104864
rect 328416 87122 328444 104858
rect 328508 95169 328536 336806
rect 328494 95160 328550 95169
rect 328600 95130 328628 340054
rect 328692 335782 328720 340068
rect 328772 337000 328824 337006
rect 328772 336942 328824 336948
rect 328680 335776 328732 335782
rect 328680 335718 328732 335724
rect 328680 335572 328732 335578
rect 328680 335514 328732 335520
rect 328494 95095 328550 95104
rect 328588 95124 328640 95130
rect 328588 95066 328640 95072
rect 328494 95024 328550 95033
rect 328494 94959 328550 94968
rect 328588 94988 328640 94994
rect 328232 87094 328444 87122
rect 328232 77353 328260 87094
rect 328218 77344 328274 77353
rect 328218 77279 328274 77288
rect 328402 77344 328458 77353
rect 328402 77279 328458 77288
rect 328416 58177 328444 77279
rect 328402 58168 328458 58177
rect 328402 58103 328458 58112
rect 328402 58032 328458 58041
rect 328402 57967 328458 57976
rect 328416 46918 328444 57967
rect 328404 46912 328456 46918
rect 328404 46854 328456 46860
rect 328220 37324 328272 37330
rect 328220 37266 328272 37272
rect 328232 19258 328260 37266
rect 328232 19230 328444 19258
rect 328416 11014 328444 19230
rect 328404 11008 328456 11014
rect 328404 10950 328456 10956
rect 328508 10742 328536 94959
rect 328588 94930 328640 94936
rect 328404 10736 328456 10742
rect 328404 10678 328456 10684
rect 328496 10736 328548 10742
rect 328496 10678 328548 10684
rect 328416 10033 328444 10678
rect 328402 10024 328458 10033
rect 328402 9959 328458 9968
rect 328600 6934 328628 94930
rect 328692 7750 328720 335514
rect 328680 7744 328732 7750
rect 328680 7686 328732 7692
rect 328588 6928 328640 6934
rect 328588 6870 328640 6876
rect 328678 6488 328734 6497
rect 328678 6423 328734 6432
rect 328692 6322 328720 6423
rect 328680 6316 328732 6322
rect 328680 6258 328732 6264
rect 328128 4548 328180 4554
rect 328128 4490 328180 4496
rect 327482 3768 327538 3777
rect 327482 3703 327538 3712
rect 328140 480 328168 4490
rect 328784 3641 328812 336942
rect 328770 3632 328826 3641
rect 328770 3567 328826 3576
rect 328876 3505 328904 340068
rect 329152 336938 329180 340068
rect 329140 336932 329192 336938
rect 329140 336874 329192 336880
rect 329428 336870 329456 340068
rect 329626 340054 329732 340082
rect 329416 336864 329468 336870
rect 329416 336806 329468 336812
rect 329704 331242 329732 340054
rect 329888 333334 329916 340068
rect 330060 336932 330112 336938
rect 330060 336874 330112 336880
rect 329968 336864 330020 336870
rect 329968 336806 330020 336812
rect 329876 333328 329928 333334
rect 329876 333270 329928 333276
rect 329704 331214 329916 331242
rect 328956 17264 329008 17270
rect 328956 17206 329008 17212
rect 328862 3496 328918 3505
rect 328862 3431 328918 3440
rect 328968 2802 328996 17206
rect 329888 10826 329916 331214
rect 329796 10798 329916 10826
rect 329796 2961 329824 10798
rect 329980 10674 330008 336806
rect 329876 10668 329928 10674
rect 329876 10610 329928 10616
rect 329968 10668 330020 10674
rect 329968 10610 330020 10616
rect 329888 10577 329916 10610
rect 329874 10568 329930 10577
rect 329874 10503 329930 10512
rect 330072 7886 330100 336874
rect 330060 7880 330112 7886
rect 330060 7822 330112 7828
rect 330164 7206 330192 340068
rect 330348 336938 330376 340068
rect 330532 340054 330638 340082
rect 330336 336932 330388 336938
rect 330336 336874 330388 336880
rect 330532 330614 330560 340054
rect 330900 337006 330928 340068
rect 330888 337000 330940 337006
rect 330888 336942 330940 336948
rect 331084 336870 331112 340068
rect 331268 340054 331374 340082
rect 331544 340054 331650 340082
rect 331164 337000 331216 337006
rect 331164 336942 331216 336948
rect 331072 336864 331124 336870
rect 331072 336806 331124 336812
rect 330520 330608 330572 330614
rect 330520 330550 330572 330556
rect 331176 326346 331204 336942
rect 331268 327826 331296 340054
rect 331440 336932 331492 336938
rect 331440 336874 331492 336880
rect 331348 336864 331400 336870
rect 331348 336806 331400 336812
rect 331256 327820 331308 327826
rect 331256 327762 331308 327768
rect 331176 326318 331296 326346
rect 331268 318730 331296 326318
rect 331176 318702 331296 318730
rect 331176 311982 331204 318702
rect 331164 311976 331216 311982
rect 331164 311918 331216 311924
rect 331256 309256 331308 309262
rect 331176 309204 331256 309210
rect 331176 309198 331308 309204
rect 331176 309182 331296 309198
rect 331176 302258 331204 309182
rect 331164 302252 331216 302258
rect 331164 302194 331216 302200
rect 331256 302184 331308 302190
rect 331256 302126 331308 302132
rect 331268 298058 331296 302126
rect 331176 298030 331296 298058
rect 331176 292602 331204 298030
rect 331164 292596 331216 292602
rect 331164 292538 331216 292544
rect 331256 292528 331308 292534
rect 331256 292470 331308 292476
rect 331268 280090 331296 292470
rect 331256 280084 331308 280090
rect 331256 280026 331308 280032
rect 331256 270564 331308 270570
rect 331256 270506 331308 270512
rect 331268 260846 331296 270506
rect 331256 260840 331308 260846
rect 331256 260782 331308 260788
rect 331256 251252 331308 251258
rect 331256 251194 331308 251200
rect 331268 241505 331296 251194
rect 331070 241496 331126 241505
rect 331070 241431 331126 241440
rect 331254 241496 331310 241505
rect 331254 241431 331310 241440
rect 331084 231878 331112 241431
rect 331072 231872 331124 231878
rect 331072 231814 331124 231820
rect 331256 231872 331308 231878
rect 331256 231814 331308 231820
rect 331268 222193 331296 231814
rect 331070 222184 331126 222193
rect 331070 222119 331126 222128
rect 331254 222184 331310 222193
rect 331254 222119 331310 222128
rect 331084 212566 331112 222119
rect 331072 212560 331124 212566
rect 331072 212502 331124 212508
rect 331256 212560 331308 212566
rect 331256 212502 331308 212508
rect 331268 202881 331296 212502
rect 331070 202872 331126 202881
rect 331070 202807 331126 202816
rect 331254 202872 331310 202881
rect 331254 202807 331310 202816
rect 331084 193254 331112 202807
rect 331072 193248 331124 193254
rect 331072 193190 331124 193196
rect 331256 193248 331308 193254
rect 331256 193190 331308 193196
rect 331268 183569 331296 193190
rect 331070 183560 331126 183569
rect 331070 183495 331126 183504
rect 331254 183560 331310 183569
rect 331254 183495 331310 183504
rect 331084 173942 331112 183495
rect 331072 173936 331124 173942
rect 331072 173878 331124 173884
rect 331256 173936 331308 173942
rect 331256 173878 331308 173884
rect 331268 164218 331296 173878
rect 331072 164212 331124 164218
rect 331072 164154 331124 164160
rect 331256 164212 331308 164218
rect 331256 164154 331308 164160
rect 331084 154601 331112 164154
rect 331070 154592 331126 154601
rect 331070 154527 331126 154536
rect 331254 154592 331310 154601
rect 331254 154527 331310 154536
rect 331268 144906 331296 154527
rect 331072 144900 331124 144906
rect 331072 144842 331124 144848
rect 331256 144900 331308 144906
rect 331256 144842 331308 144848
rect 331084 135289 331112 144842
rect 331070 135280 331126 135289
rect 331070 135215 331126 135224
rect 331254 135280 331310 135289
rect 331254 135215 331310 135224
rect 331268 125594 331296 135215
rect 331072 125588 331124 125594
rect 331072 125530 331124 125536
rect 331256 125588 331308 125594
rect 331256 125530 331308 125536
rect 331084 115977 331112 125530
rect 331070 115968 331126 115977
rect 331070 115903 331126 115912
rect 331254 115968 331310 115977
rect 331254 115903 331310 115912
rect 331268 106282 331296 115903
rect 331072 106276 331124 106282
rect 331072 106218 331124 106224
rect 331256 106276 331308 106282
rect 331256 106218 331308 106224
rect 330978 100872 331034 100881
rect 330978 100807 331034 100816
rect 330992 100609 331020 100807
rect 330978 100600 331034 100609
rect 330978 100535 331034 100544
rect 331084 96665 331112 106218
rect 331070 96656 331126 96665
rect 331070 96591 331126 96600
rect 331254 96656 331310 96665
rect 331254 96591 331310 96600
rect 331268 86970 331296 96591
rect 331072 86964 331124 86970
rect 331072 86906 331124 86912
rect 331256 86964 331308 86970
rect 331256 86906 331308 86912
rect 331084 77353 331112 86906
rect 331070 77344 331126 77353
rect 331070 77279 331126 77288
rect 331254 77344 331310 77353
rect 331254 77279 331310 77288
rect 331268 67590 331296 77279
rect 331256 67584 331308 67590
rect 331256 67526 331308 67532
rect 331256 62824 331308 62830
rect 331256 62766 331308 62772
rect 331268 41426 331296 62766
rect 331176 41398 331296 41426
rect 331176 41290 331204 41398
rect 331176 41262 331296 41290
rect 331268 12458 331296 41262
rect 331176 12430 331296 12458
rect 331176 7274 331204 12430
rect 331360 11694 331388 336806
rect 331348 11688 331400 11694
rect 331348 11630 331400 11636
rect 331452 11370 331480 336874
rect 331268 11342 331480 11370
rect 331268 10305 331296 11342
rect 331348 11076 331400 11082
rect 331348 11018 331400 11024
rect 331254 10296 331310 10305
rect 331254 10231 331310 10240
rect 331360 10130 331388 11018
rect 331544 10826 331572 340054
rect 331820 337006 331848 340068
rect 332096 337074 332124 340068
rect 332084 337068 332136 337074
rect 332084 337010 332136 337016
rect 331808 337000 331860 337006
rect 331808 336942 331860 336948
rect 332372 336938 332400 340068
rect 332360 336932 332412 336938
rect 332360 336874 332412 336880
rect 332556 336870 332584 340068
rect 332740 340054 332846 340082
rect 333122 340054 333228 340082
rect 332636 337068 332688 337074
rect 332636 337010 332688 337016
rect 332544 336864 332596 336870
rect 332544 336806 332596 336812
rect 332648 325038 332676 337010
rect 332636 325032 332688 325038
rect 332636 324974 332688 324980
rect 332740 322318 332768 340054
rect 332912 337000 332964 337006
rect 332912 336942 332964 336948
rect 332820 336864 332872 336870
rect 332820 336806 332872 336812
rect 332728 322312 332780 322318
rect 332728 322254 332780 322260
rect 331716 322244 331768 322250
rect 331716 322186 331768 322192
rect 331452 10798 331572 10826
rect 331348 10124 331400 10130
rect 331348 10066 331400 10072
rect 331452 7342 331480 10798
rect 331622 10568 331678 10577
rect 331622 10503 331678 10512
rect 331636 10198 331664 10503
rect 331624 10192 331676 10198
rect 331624 10134 331676 10140
rect 331624 10056 331676 10062
rect 331622 10024 331624 10033
rect 331676 10024 331678 10033
rect 331622 9959 331678 9968
rect 331728 7546 331756 322186
rect 332832 12374 332860 336806
rect 332924 12442 332952 336942
rect 333004 336932 333056 336938
rect 333004 336874 333056 336880
rect 332912 12436 332964 12442
rect 332912 12378 332964 12384
rect 332820 12368 332872 12374
rect 332820 12310 332872 12316
rect 333016 8022 333044 336874
rect 333200 335578 333228 340054
rect 333292 336938 333320 340068
rect 333568 338065 333596 340068
rect 333370 338056 333426 338065
rect 333370 337991 333426 338000
rect 333554 338056 333610 338065
rect 333554 337991 333610 338000
rect 333280 336932 333332 336938
rect 333280 336874 333332 336880
rect 333188 335572 333240 335578
rect 333188 335514 333240 335520
rect 333384 328506 333412 337991
rect 333844 337006 333872 340068
rect 334042 340054 334148 340082
rect 333832 337000 333884 337006
rect 333832 336942 333884 336948
rect 334016 336864 334068 336870
rect 334016 336806 334068 336812
rect 333372 328500 333424 328506
rect 333372 328442 333424 328448
rect 333924 328500 333976 328506
rect 333924 328442 333976 328448
rect 333738 320648 333794 320657
rect 333738 320583 333794 320592
rect 333752 320249 333780 320583
rect 333738 320240 333794 320249
rect 333738 320175 333794 320184
rect 333936 319530 333964 328442
rect 333924 319524 333976 319530
rect 333924 319466 333976 319472
rect 334028 318102 334056 336806
rect 334016 318096 334068 318102
rect 334016 318038 334068 318044
rect 334120 12238 334148 340054
rect 334200 336932 334252 336938
rect 334200 336874 334252 336880
rect 334212 12306 334240 336874
rect 334304 336870 334332 340068
rect 334580 337006 334608 340068
rect 334384 337000 334436 337006
rect 334384 336942 334436 336948
rect 334568 337000 334620 337006
rect 334568 336942 334620 336948
rect 334292 336864 334344 336870
rect 334292 336806 334344 336812
rect 334292 335572 334344 335578
rect 334292 335514 334344 335520
rect 334200 12300 334252 12306
rect 334200 12242 334252 12248
rect 334108 12232 334160 12238
rect 334108 12174 334160 12180
rect 333004 8016 333056 8022
rect 333004 7958 333056 7964
rect 334304 7954 334332 335514
rect 334292 7948 334344 7954
rect 334292 7890 334344 7896
rect 331716 7540 331768 7546
rect 331716 7482 331768 7488
rect 332912 7540 332964 7546
rect 332912 7482 332964 7488
rect 331440 7336 331492 7342
rect 331440 7278 331492 7284
rect 331164 7268 331216 7274
rect 331164 7210 331216 7216
rect 330152 7200 330204 7206
rect 330152 7142 330204 7148
rect 331716 6996 331768 7002
rect 331716 6938 331768 6944
rect 331728 6089 331756 6938
rect 331714 6080 331770 6089
rect 331714 6015 331770 6024
rect 331716 5092 331768 5098
rect 331716 5034 331768 5040
rect 330520 4616 330572 4622
rect 330520 4558 330572 4564
rect 329782 2952 329838 2961
rect 329782 2887 329838 2896
rect 328968 2774 329272 2802
rect 329244 2666 329272 2774
rect 329244 2638 329364 2666
rect 329336 480 329364 2638
rect 330532 480 330560 4558
rect 331728 480 331756 5034
rect 332924 480 332952 7482
rect 334396 7410 334424 336942
rect 334764 336870 334792 340068
rect 334752 336864 334804 336870
rect 334752 336806 334804 336812
rect 335040 335594 335068 340068
rect 335316 336938 335344 340068
rect 335304 336932 335356 336938
rect 335304 336874 335356 336880
rect 335396 336864 335448 336870
rect 335396 336806 335448 336812
rect 335040 335566 335344 335594
rect 335316 315314 335344 335566
rect 335304 315308 335356 315314
rect 335304 315250 335356 315256
rect 335408 279478 335436 336806
rect 335396 279472 335448 279478
rect 335396 279414 335448 279420
rect 335500 12170 335528 340068
rect 335672 337000 335724 337006
rect 335672 336942 335724 336948
rect 335580 336932 335632 336938
rect 335580 336874 335632 336880
rect 335488 12164 335540 12170
rect 335488 12106 335540 12112
rect 335592 7478 335620 336874
rect 335684 7546 335712 336942
rect 335672 7540 335724 7546
rect 335672 7482 335724 7488
rect 335580 7472 335632 7478
rect 335580 7414 335632 7420
rect 334384 7404 334436 7410
rect 334384 7346 334436 7352
rect 335776 5030 335804 340068
rect 335960 337006 335988 340068
rect 336236 337074 336264 340068
rect 336224 337068 336276 337074
rect 336224 337010 336276 337016
rect 335948 337000 336000 337006
rect 335948 336942 336000 336948
rect 336512 336938 336540 340068
rect 336500 336932 336552 336938
rect 336500 336874 336552 336880
rect 336696 336870 336724 340068
rect 336880 340054 336986 340082
rect 336776 337068 336828 337074
rect 336776 337010 336828 337016
rect 336684 336864 336736 336870
rect 336684 336806 336736 336812
rect 336788 276690 336816 337010
rect 336776 276684 336828 276690
rect 336776 276626 336828 276632
rect 336132 18624 336184 18630
rect 336132 18566 336184 18572
rect 335212 5024 335264 5030
rect 335212 4966 335264 4972
rect 335764 5024 335816 5030
rect 335764 4966 335816 4972
rect 334108 4684 334160 4690
rect 334108 4626 334160 4632
rect 334120 480 334148 4626
rect 335224 480 335252 4966
rect 336144 4842 336172 18566
rect 336880 12102 336908 340054
rect 336960 337000 337012 337006
rect 336960 336942 337012 336948
rect 336868 12096 336920 12102
rect 336868 12038 336920 12044
rect 336972 8090 337000 336942
rect 337144 336932 337196 336938
rect 337144 336874 337196 336880
rect 337052 336864 337104 336870
rect 337052 336806 337104 336812
rect 337064 8294 337092 336806
rect 337052 8288 337104 8294
rect 337052 8230 337104 8236
rect 336960 8084 337012 8090
rect 336960 8026 337012 8032
rect 336144 4814 336448 4842
rect 336420 480 336448 4814
rect 337156 4690 337184 336874
rect 337248 336870 337276 340068
rect 337432 336938 337460 340068
rect 337420 336932 337472 336938
rect 337420 336874 337472 336880
rect 337236 336864 337288 336870
rect 337236 336806 337288 336812
rect 337708 331974 337736 340068
rect 337984 335578 338012 340068
rect 338182 340054 338380 340082
rect 338248 336932 338300 336938
rect 338248 336874 338300 336880
rect 338064 336864 338116 336870
rect 338064 336806 338116 336812
rect 338156 336864 338208 336870
rect 338156 336806 338208 336812
rect 337972 335572 338024 335578
rect 337972 335514 338024 335520
rect 337696 331968 337748 331974
rect 337696 331910 337748 331916
rect 337234 39264 337290 39273
rect 337234 39199 337290 39208
rect 337248 39001 337276 39199
rect 337234 38992 337290 39001
rect 337234 38927 337290 38936
rect 337234 6488 337290 6497
rect 337234 6423 337290 6432
rect 337248 6322 337276 6423
rect 337236 6316 337288 6322
rect 337236 6258 337288 6264
rect 338076 5302 338104 336806
rect 338168 11898 338196 336806
rect 338156 11892 338208 11898
rect 338156 11834 338208 11840
rect 338156 8016 338208 8022
rect 338156 7958 338208 7964
rect 338168 7449 338196 7958
rect 338260 7886 338288 336874
rect 338352 8022 338380 340054
rect 338444 336870 338472 340068
rect 338734 340054 338840 340082
rect 338432 336864 338484 336870
rect 338432 336806 338484 336812
rect 338432 335572 338484 335578
rect 338432 335514 338484 335520
rect 338340 8016 338392 8022
rect 338340 7958 338392 7964
rect 338248 7880 338300 7886
rect 338248 7822 338300 7828
rect 338154 7440 338210 7449
rect 338154 7375 338210 7384
rect 338064 5296 338116 5302
rect 338064 5238 338116 5244
rect 337604 4820 337656 4826
rect 337604 4762 337656 4768
rect 337144 4684 337196 4690
rect 337144 4626 337196 4632
rect 336684 4276 336736 4282
rect 336684 4218 336736 4224
rect 336696 3505 336724 4218
rect 336682 3496 336738 3505
rect 336682 3431 336738 3440
rect 337616 480 337644 4762
rect 338444 4214 338472 335514
rect 338812 335374 338840 340054
rect 338904 337006 338932 340068
rect 338892 337000 338944 337006
rect 338892 336942 338944 336948
rect 339180 336870 339208 340068
rect 339352 336932 339404 336938
rect 339352 336874 339404 336880
rect 339168 336864 339220 336870
rect 339168 336806 339220 336812
rect 338800 335368 338852 335374
rect 338800 335310 338852 335316
rect 339364 330478 339392 336874
rect 339352 330472 339404 330478
rect 339352 330414 339404 330420
rect 338798 6488 338854 6497
rect 338798 6423 338854 6432
rect 338812 6322 338840 6423
rect 338800 6316 338852 6322
rect 338800 6258 338852 6264
rect 338800 4752 338852 4758
rect 338800 4694 338852 4700
rect 338432 4208 338484 4214
rect 338432 4150 338484 4156
rect 338522 3360 338578 3369
rect 338352 3318 338522 3346
rect 338352 3233 338380 3318
rect 338522 3295 338578 3304
rect 338338 3224 338394 3233
rect 338338 3159 338394 3168
rect 338812 480 338840 4694
rect 339456 4282 339484 340068
rect 339640 336938 339668 340068
rect 339732 340054 339930 340082
rect 339628 336932 339680 336938
rect 339628 336874 339680 336880
rect 339536 336864 339588 336870
rect 339536 336806 339588 336812
rect 339548 307086 339576 336806
rect 339732 335594 339760 340054
rect 340192 337006 340220 340068
rect 340390 340054 340588 340082
rect 339812 337000 339864 337006
rect 339812 336942 339864 336948
rect 340180 337000 340232 337006
rect 340180 336942 340232 336948
rect 339640 335566 339760 335594
rect 339536 307080 339588 307086
rect 339536 307022 339588 307028
rect 339640 11830 339668 335566
rect 339824 335458 339852 336942
rect 340560 335594 340588 340054
rect 340652 336938 340680 340068
rect 340640 336932 340692 336938
rect 340640 336874 340692 336880
rect 340928 336870 340956 340068
rect 341020 340054 341126 340082
rect 340916 336864 340968 336870
rect 340916 336806 340968 336812
rect 340560 335566 340956 335594
rect 339732 335430 339852 335458
rect 339628 11824 339680 11830
rect 339628 11766 339680 11772
rect 339732 7954 339760 335430
rect 339812 335368 339864 335374
rect 339812 335310 339864 335316
rect 339720 7948 339772 7954
rect 339720 7890 339772 7896
rect 339824 4826 339852 335310
rect 340824 331220 340876 331226
rect 340824 331162 340876 331168
rect 340836 321638 340864 331162
rect 340824 321632 340876 321638
rect 340824 321574 340876 321580
rect 340824 321428 340876 321434
rect 340824 321370 340876 321376
rect 340836 309194 340864 321370
rect 340824 309188 340876 309194
rect 340824 309130 340876 309136
rect 340824 302184 340876 302190
rect 340824 302126 340876 302132
rect 340836 294982 340864 302126
rect 340928 297430 340956 335566
rect 340916 297424 340968 297430
rect 340916 297366 340968 297372
rect 340824 294976 340876 294982
rect 340824 294918 340876 294924
rect 341020 294642 341048 340054
rect 341388 337142 341416 340068
rect 341376 337136 341428 337142
rect 341376 337078 341428 337084
rect 341664 337074 341692 340068
rect 341652 337068 341704 337074
rect 341652 337010 341704 337016
rect 341284 337000 341336 337006
rect 341284 336942 341336 336948
rect 341100 336932 341152 336938
rect 341100 336874 341152 336880
rect 339996 294636 340048 294642
rect 339996 294578 340048 294584
rect 341008 294636 341060 294642
rect 341008 294578 341060 294584
rect 339812 4820 339864 4826
rect 339812 4762 339864 4768
rect 339444 4276 339496 4282
rect 339444 4218 339496 4224
rect 340008 480 340036 294578
rect 341112 290193 341140 336874
rect 341192 336864 341244 336870
rect 341192 336806 341244 336812
rect 341204 331226 341232 336806
rect 341192 331220 341244 331226
rect 341192 331162 341244 331168
rect 341192 321632 341244 321638
rect 341192 321574 341244 321580
rect 341204 321434 341232 321574
rect 341192 321428 341244 321434
rect 341192 321370 341244 321376
rect 341192 309188 341244 309194
rect 341192 309130 341244 309136
rect 341204 302190 341232 309130
rect 341192 302184 341244 302190
rect 341192 302126 341244 302132
rect 341192 294976 341244 294982
rect 341192 294918 341244 294924
rect 341098 290184 341154 290193
rect 341098 290119 341154 290128
rect 341098 289912 341154 289921
rect 341098 289847 341154 289856
rect 341112 283014 341140 289847
rect 341204 289814 341232 294918
rect 341192 289808 341244 289814
rect 341192 289750 341244 289756
rect 341100 283008 341152 283014
rect 341100 282950 341152 282956
rect 341100 282804 341152 282810
rect 341100 282746 341152 282752
rect 340916 280288 340968 280294
rect 340916 280230 340968 280236
rect 340928 270881 340956 280230
rect 341112 271182 341140 282746
rect 341100 271176 341152 271182
rect 341100 271118 341152 271124
rect 340914 270872 340970 270881
rect 340914 270807 340970 270816
rect 341190 270600 341246 270609
rect 341190 270535 341246 270544
rect 341204 263702 341232 270535
rect 341192 263696 341244 263702
rect 341192 263638 341244 263644
rect 341100 263560 341152 263566
rect 341100 263502 341152 263508
rect 341112 260846 341140 263502
rect 341100 260840 341152 260846
rect 341100 260782 341152 260788
rect 341192 251252 341244 251258
rect 341192 251194 341244 251200
rect 341204 241482 341232 251194
rect 341112 241454 341232 241482
rect 341112 234818 341140 241454
rect 341020 234790 341140 234818
rect 341020 231878 341048 234790
rect 341008 231872 341060 231878
rect 341008 231814 341060 231820
rect 341100 231872 341152 231878
rect 341100 231814 341152 231820
rect 341112 225078 341140 231814
rect 341100 225072 341152 225078
rect 341100 225014 341152 225020
rect 341008 224936 341060 224942
rect 341008 224878 341060 224884
rect 341020 220794 341048 224878
rect 341008 220788 341060 220794
rect 341008 220730 341060 220736
rect 341100 215280 341152 215286
rect 341100 215222 341152 215228
rect 341112 211154 341140 215222
rect 341112 211126 341232 211154
rect 341204 205834 341232 211126
rect 341192 205828 341244 205834
rect 341192 205770 341244 205776
rect 341100 205556 341152 205562
rect 341100 205498 341152 205504
rect 341112 202842 341140 205498
rect 341100 202836 341152 202842
rect 341100 202778 341152 202784
rect 341192 193384 341244 193390
rect 341192 193326 341244 193332
rect 341204 193202 341232 193326
rect 341112 193174 341232 193202
rect 341112 186386 341140 193174
rect 341100 186380 341152 186386
rect 341100 186322 341152 186328
rect 341100 183660 341152 183666
rect 341100 183602 341152 183608
rect 341112 183530 341140 183602
rect 341100 183524 341152 183530
rect 341100 183466 341152 183472
rect 341190 174040 341246 174049
rect 341190 173975 341246 173984
rect 341204 173913 341232 173975
rect 341190 173904 341246 173913
rect 341190 173839 341246 173848
rect 341098 164384 341154 164393
rect 341098 164319 341154 164328
rect 341112 164218 341140 164319
rect 341008 164212 341060 164218
rect 341008 164154 341060 164160
rect 341100 164212 341152 164218
rect 341100 164154 341152 164160
rect 341020 157298 341048 164154
rect 341020 157270 341140 157298
rect 341112 154578 341140 157270
rect 341112 154550 341232 154578
rect 341204 147762 341232 154550
rect 341192 147756 341244 147762
rect 341192 147698 341244 147704
rect 341100 147620 341152 147626
rect 341100 147562 341152 147568
rect 341112 144906 341140 147562
rect 341008 144900 341060 144906
rect 341008 144842 341060 144848
rect 341100 144900 341152 144906
rect 341100 144842 341152 144848
rect 341020 137986 341048 144842
rect 341020 137958 341140 137986
rect 341112 135266 341140 137958
rect 341112 135250 341232 135266
rect 341112 135244 341244 135250
rect 341112 135238 341192 135244
rect 341192 135186 341244 135192
rect 341204 135155 341232 135186
rect 341190 125624 341246 125633
rect 341112 125594 341190 125610
rect 341100 125588 341190 125594
rect 341152 125582 341190 125588
rect 341190 125559 341246 125568
rect 341100 125530 341152 125536
rect 341192 116068 341244 116074
rect 341192 116010 341244 116016
rect 341204 115841 341232 116010
rect 341190 115832 341246 115841
rect 341190 115767 341246 115776
rect 341190 106312 341246 106321
rect 341112 106282 341190 106298
rect 341008 106276 341060 106282
rect 341008 106218 341060 106224
rect 341100 106276 341190 106282
rect 341152 106270 341190 106276
rect 341190 106247 341246 106256
rect 341100 106218 341152 106224
rect 341020 99362 341048 106218
rect 341020 99334 341140 99362
rect 341112 96642 341140 99334
rect 341112 96626 341232 96642
rect 341112 96620 341244 96626
rect 341112 96614 341192 96620
rect 341192 96562 341244 96568
rect 341204 96531 341232 96562
rect 341190 87000 341246 87009
rect 341112 86970 341190 86986
rect 341100 86964 341190 86970
rect 341152 86958 341190 86964
rect 341190 86935 341246 86944
rect 341100 86906 341152 86912
rect 341192 77444 341244 77450
rect 341192 77386 341244 77392
rect 341204 77178 341232 77386
rect 341192 77172 341244 77178
rect 341192 77114 341244 77120
rect 341100 67652 341152 67658
rect 341100 67594 341152 67600
rect 341112 67538 341140 67594
rect 341112 67510 341232 67538
rect 341204 60790 341232 67510
rect 341192 60784 341244 60790
rect 341192 60726 341244 60732
rect 341100 60716 341152 60722
rect 341100 60658 341152 60664
rect 341112 58018 341140 60658
rect 341112 57990 341232 58018
rect 341204 57934 341232 57990
rect 340916 57928 340968 57934
rect 340916 57870 340968 57876
rect 341192 57928 341244 57934
rect 341192 57870 341244 57876
rect 340928 48385 340956 57870
rect 340914 48376 340970 48385
rect 340914 48311 340970 48320
rect 341098 48376 341154 48385
rect 341098 48311 341154 48320
rect 341112 48278 341140 48311
rect 341008 48272 341060 48278
rect 341008 48214 341060 48220
rect 341100 48272 341152 48278
rect 341100 48214 341152 48220
rect 341020 38706 341048 48214
rect 341020 38678 341232 38706
rect 341204 38570 341232 38678
rect 341112 38542 341232 38570
rect 341112 31890 341140 38542
rect 341100 31884 341152 31890
rect 341100 31826 341152 31832
rect 341008 29028 341060 29034
rect 341008 28970 341060 28976
rect 341020 22250 341048 28970
rect 340928 22222 341048 22250
rect 340928 19394 340956 22222
rect 340928 19366 341048 19394
rect 341020 19310 341048 19366
rect 340732 19304 340784 19310
rect 340732 19246 340784 19252
rect 341008 19304 341060 19310
rect 341008 19246 341060 19252
rect 340744 9761 340772 19246
rect 340730 9752 340786 9761
rect 340730 9687 340786 9696
rect 340914 9752 340970 9761
rect 340914 9687 340970 9696
rect 340822 8256 340878 8265
rect 340822 8191 340878 8200
rect 340730 8120 340786 8129
rect 340730 8055 340786 8064
rect 340744 7478 340772 8055
rect 340836 7546 340864 8191
rect 340824 7540 340876 7546
rect 340824 7482 340876 7488
rect 340732 7472 340784 7478
rect 340732 7414 340784 7420
rect 340928 4758 340956 9687
rect 341296 9382 341324 336942
rect 341848 327758 341876 340068
rect 342032 340054 342138 340082
rect 342414 340054 342520 340082
rect 342598 340054 342704 340082
rect 342032 330546 342060 340054
rect 342492 337770 342520 340054
rect 342492 337742 342612 337770
rect 342388 337204 342440 337210
rect 342388 337146 342440 337152
rect 342400 330698 342428 337146
rect 342480 337136 342532 337142
rect 342480 337078 342532 337084
rect 342308 330670 342428 330698
rect 342020 330540 342072 330546
rect 342020 330482 342072 330488
rect 341836 327752 341888 327758
rect 341836 327694 341888 327700
rect 342204 316804 342256 316810
rect 342204 316746 342256 316752
rect 342216 306406 342244 316746
rect 342204 306400 342256 306406
rect 342204 306342 342256 306348
rect 342204 296744 342256 296750
rect 342204 296686 342256 296692
rect 342216 282962 342244 296686
rect 342308 291854 342336 330670
rect 342388 330540 342440 330546
rect 342388 330482 342440 330488
rect 342400 316810 342428 330482
rect 342388 316804 342440 316810
rect 342388 316746 342440 316752
rect 342388 306400 342440 306406
rect 342388 306342 342440 306348
rect 342400 296750 342428 306342
rect 342388 296744 342440 296750
rect 342388 296686 342440 296692
rect 342296 291848 342348 291854
rect 342296 291790 342348 291796
rect 342216 282934 342428 282962
rect 342400 268394 342428 282934
rect 342388 268388 342440 268394
rect 342388 268330 342440 268336
rect 341468 183524 341520 183530
rect 341468 183466 341520 183472
rect 341480 174049 341508 183466
rect 341466 174040 341522 174049
rect 341466 173975 341522 173984
rect 341374 173904 341430 173913
rect 341374 173839 341430 173848
rect 341388 164393 341416 173839
rect 341374 164384 341430 164393
rect 341374 164319 341430 164328
rect 341376 135244 341428 135250
rect 341376 135186 341428 135192
rect 341388 125633 341416 135186
rect 341374 125624 341430 125633
rect 341374 125559 341430 125568
rect 341466 115832 341522 115841
rect 341466 115767 341522 115776
rect 341480 106321 341508 115767
rect 341466 106312 341522 106321
rect 341466 106247 341522 106256
rect 341376 96620 341428 96626
rect 341376 96562 341428 96568
rect 341388 87009 341416 96562
rect 341374 87000 341430 87009
rect 341374 86935 341430 86944
rect 342492 11762 342520 337078
rect 342480 11756 342532 11762
rect 342480 11698 342532 11704
rect 341468 11212 341520 11218
rect 341468 11154 341520 11160
rect 341480 10441 341508 11154
rect 341466 10432 341522 10441
rect 341466 10367 341522 10376
rect 341284 9376 341336 9382
rect 341284 9318 341336 9324
rect 341284 8288 341336 8294
rect 341282 8256 341284 8265
rect 341336 8256 341338 8265
rect 341282 8191 341338 8200
rect 341374 8120 341430 8129
rect 341374 8055 341376 8064
rect 341428 8055 341430 8064
rect 341376 8026 341428 8032
rect 341192 5364 341244 5370
rect 341192 5306 341244 5312
rect 340916 4752 340968 4758
rect 340916 4694 340968 4700
rect 341204 480 341232 5306
rect 342388 5160 342440 5166
rect 342388 5102 342440 5108
rect 341468 3528 341520 3534
rect 341466 3496 341468 3505
rect 341520 3496 341522 3505
rect 341466 3431 341522 3440
rect 342400 480 342428 5102
rect 342584 5098 342612 337742
rect 342676 337210 342704 340054
rect 342860 337210 342888 340068
rect 342664 337204 342716 337210
rect 342664 337146 342716 337152
rect 342848 337204 342900 337210
rect 342848 337146 342900 337152
rect 343136 337074 343164 340068
rect 342664 337068 342716 337074
rect 342664 337010 342716 337016
rect 343124 337068 343176 337074
rect 343124 337010 343176 337016
rect 342572 5092 342624 5098
rect 342572 5034 342624 5040
rect 342676 4457 342704 337010
rect 343320 336938 343348 340068
rect 343610 340054 343808 340082
rect 343886 340054 343992 340082
rect 343780 337770 343808 340054
rect 343780 337742 343900 337770
rect 343768 337204 343820 337210
rect 343768 337146 343820 337152
rect 343584 337068 343636 337074
rect 343584 337010 343636 337016
rect 343676 337068 343728 337074
rect 343676 337010 343728 337016
rect 342756 336932 342808 336938
rect 342756 336874 342808 336880
rect 343308 336932 343360 336938
rect 343308 336874 343360 336880
rect 342768 334694 342796 336874
rect 342756 334688 342808 334694
rect 342756 334630 342808 334636
rect 343398 320240 343454 320249
rect 343398 320175 343454 320184
rect 343412 319977 343440 320175
rect 343398 319968 343454 319977
rect 343398 319903 343454 319912
rect 342756 265668 342808 265674
rect 342756 265610 342808 265616
rect 342768 5114 342796 265610
rect 343398 7440 343454 7449
rect 343398 7375 343400 7384
rect 343452 7375 343454 7384
rect 343400 7346 343452 7352
rect 343596 5302 343624 337010
rect 343688 322250 343716 337010
rect 343676 322244 343728 322250
rect 343676 322186 343728 322192
rect 343780 304298 343808 337146
rect 343768 304292 343820 304298
rect 343768 304234 343820 304240
rect 343872 265674 343900 337742
rect 343860 265668 343912 265674
rect 343860 265610 343912 265616
rect 343584 5296 343636 5302
rect 343584 5238 343636 5244
rect 343964 5166 343992 340054
rect 344056 337074 344084 340068
rect 344332 337142 344360 340068
rect 344608 337210 344636 340068
rect 344806 340054 345004 340082
rect 345082 340054 345280 340082
rect 344976 337770 345004 340054
rect 344976 337742 345188 337770
rect 344596 337204 344648 337210
rect 344596 337146 344648 337152
rect 344320 337136 344372 337142
rect 344320 337078 344372 337084
rect 345056 337136 345108 337142
rect 345056 337078 345108 337084
rect 344044 337068 344096 337074
rect 344044 337010 344096 337016
rect 345068 324970 345096 337078
rect 345056 324964 345108 324970
rect 345056 324906 345108 324912
rect 345160 309806 345188 337742
rect 345148 309800 345200 309806
rect 345148 309742 345200 309748
rect 345252 262886 345280 340054
rect 345240 262880 345292 262886
rect 345240 262822 345292 262828
rect 345344 5273 345372 340068
rect 345424 337204 345476 337210
rect 345424 337146 345476 337152
rect 345436 5302 345464 337146
rect 345528 337074 345556 340068
rect 345516 337068 345568 337074
rect 345516 337010 345568 337016
rect 345804 337006 345832 340068
rect 346080 337142 346108 340068
rect 346264 337210 346292 340068
rect 346448 340054 346554 340082
rect 346724 340054 346830 340082
rect 346252 337204 346304 337210
rect 346252 337146 346304 337152
rect 346068 337136 346120 337142
rect 346068 337078 346120 337084
rect 345792 337000 345844 337006
rect 345792 336942 345844 336948
rect 346344 337000 346396 337006
rect 346344 336942 346396 336948
rect 346356 319462 346384 336942
rect 346344 319456 346396 319462
rect 346344 319398 346396 319404
rect 346448 301510 346476 340054
rect 346528 337204 346580 337210
rect 346528 337146 346580 337152
rect 346436 301504 346488 301510
rect 346436 301446 346488 301452
rect 346540 11218 346568 337146
rect 346620 337068 346672 337074
rect 346620 337010 346672 337016
rect 346528 11212 346580 11218
rect 346528 11154 346580 11160
rect 346632 9382 346660 337010
rect 346620 9376 346672 9382
rect 346620 9318 346672 9324
rect 345424 5296 345476 5302
rect 345330 5264 345386 5273
rect 345424 5238 345476 5244
rect 345330 5199 345386 5208
rect 345976 5228 346028 5234
rect 345976 5170 346028 5176
rect 343952 5160 344004 5166
rect 342768 5086 343624 5114
rect 343952 5102 344004 5108
rect 342662 4448 342718 4457
rect 342662 4383 342718 4392
rect 343596 480 343624 5086
rect 345332 5092 345384 5098
rect 345332 5034 345384 5040
rect 344780 4616 344832 4622
rect 345344 4593 345372 5034
rect 344780 4558 344832 4564
rect 345330 4584 345386 4593
rect 344792 480 344820 4558
rect 345330 4519 345386 4528
rect 345988 480 346016 5170
rect 346724 4690 346752 340054
rect 347000 337142 347028 340068
rect 346804 337136 346856 337142
rect 346804 337078 346856 337084
rect 346988 337136 347040 337142
rect 346988 337078 347040 337084
rect 346816 5166 346844 337078
rect 347276 337074 347304 340068
rect 347552 337210 347580 340068
rect 347540 337204 347592 337210
rect 347540 337146 347592 337152
rect 347264 337068 347316 337074
rect 347264 337010 347316 337016
rect 347736 337006 347764 340068
rect 347920 340054 348026 340082
rect 347816 337068 347868 337074
rect 347816 337010 347868 337016
rect 347724 337000 347776 337006
rect 347724 336942 347776 336948
rect 347828 300150 347856 337010
rect 347816 300144 347868 300150
rect 347816 300086 347868 300092
rect 347920 286346 347948 340054
rect 348288 337210 348316 340068
rect 348184 337204 348236 337210
rect 348184 337146 348236 337152
rect 348276 337204 348328 337210
rect 348276 337146 348328 337152
rect 348000 337136 348052 337142
rect 348000 337078 348052 337084
rect 347908 286340 347960 286346
rect 347908 286282 347960 286288
rect 346896 21412 346948 21418
rect 346896 21354 346948 21360
rect 346908 19310 346936 21354
rect 346896 19304 346948 19310
rect 346896 19246 346948 19252
rect 347080 19304 347132 19310
rect 347080 19246 347132 19252
rect 347092 9761 347120 19246
rect 347908 16584 347960 16590
rect 347908 16526 347960 16532
rect 346894 9752 346950 9761
rect 346894 9687 346950 9696
rect 347078 9752 347134 9761
rect 347078 9687 347134 9696
rect 346804 5160 346856 5166
rect 346804 5102 346856 5108
rect 346712 4684 346764 4690
rect 346712 4626 346764 4632
rect 346250 3360 346306 3369
rect 346250 3295 346306 3304
rect 346264 2961 346292 3295
rect 346342 3224 346398 3233
rect 346342 3159 346398 3168
rect 346250 2952 346306 2961
rect 346250 2887 346306 2896
rect 346356 2650 346384 3159
rect 346908 2802 346936 9687
rect 346986 7440 347042 7449
rect 346986 7375 346988 7384
rect 347040 7375 347042 7384
rect 346988 7346 347040 7352
rect 346986 6488 347042 6497
rect 346986 6423 347042 6432
rect 347000 6322 347028 6423
rect 346988 6316 347040 6322
rect 346988 6258 347040 6264
rect 347920 4758 347948 16526
rect 348012 9489 348040 337078
rect 348092 337000 348144 337006
rect 348092 336942 348144 336948
rect 348104 11286 348132 336942
rect 348196 16590 348224 337146
rect 348472 337074 348500 340068
rect 348748 337142 348776 340068
rect 348840 340054 349038 340082
rect 349222 340054 349420 340082
rect 348736 337136 348788 337142
rect 348736 337078 348788 337084
rect 348460 337068 348512 337074
rect 348460 337010 348512 337016
rect 348840 333266 348868 340054
rect 349196 337204 349248 337210
rect 349196 337146 349248 337152
rect 349288 337204 349340 337210
rect 349288 337146 349340 337152
rect 348828 333260 348880 333266
rect 348828 333202 348880 333208
rect 348184 16584 348236 16590
rect 348184 16526 348236 16532
rect 348092 11280 348144 11286
rect 348092 11222 348144 11228
rect 347998 9480 348054 9489
rect 347998 9415 348054 9424
rect 348366 4856 348422 4865
rect 348366 4791 348422 4800
rect 347908 4752 347960 4758
rect 347908 4694 347960 4700
rect 346908 2774 347120 2802
rect 347092 2666 347120 2774
rect 346344 2644 346396 2650
rect 347092 2638 347212 2666
rect 346344 2586 346396 2592
rect 347184 480 347212 2638
rect 348380 480 348408 4791
rect 349208 4729 349236 337146
rect 349300 283626 349328 337146
rect 349288 283620 349340 283626
rect 349288 283562 349340 283568
rect 349392 9450 349420 340054
rect 349484 337210 349512 340068
rect 349472 337204 349524 337210
rect 349472 337146 349524 337152
rect 349472 337068 349524 337074
rect 349472 337010 349524 337016
rect 349380 9444 349432 9450
rect 349380 9386 349432 9392
rect 349484 9382 349512 337010
rect 349760 337006 349788 340068
rect 349944 337210 349972 340068
rect 349932 337204 349984 337210
rect 349932 337146 349984 337152
rect 349748 337000 349800 337006
rect 349748 336942 349800 336948
rect 349656 253224 349708 253230
rect 349656 253166 349708 253172
rect 349288 9376 349340 9382
rect 349288 9318 349340 9324
rect 349472 9376 349524 9382
rect 349472 9318 349524 9324
rect 349300 9217 349328 9318
rect 349286 9208 349342 9217
rect 349286 9143 349342 9152
rect 349562 6352 349618 6361
rect 349562 6287 349618 6296
rect 349194 4720 349250 4729
rect 349194 4655 349250 4664
rect 349576 480 349604 6287
rect 349668 2446 349696 253166
rect 350036 26246 350064 459598
rect 350234 340054 350892 340082
rect 350760 337000 350812 337006
rect 350760 336942 350812 336948
rect 350772 312594 350800 336942
rect 350760 312588 350812 312594
rect 350760 312530 350812 312536
rect 350864 253230 350892 340054
rect 350944 337204 350996 337210
rect 350944 337146 350996 337152
rect 350852 253224 350904 253230
rect 350852 253166 350904 253172
rect 350024 26240 350076 26246
rect 350024 26182 350076 26188
rect 350850 9480 350906 9489
rect 350850 9415 350852 9424
rect 350904 9415 350906 9424
rect 350852 9386 350904 9392
rect 350956 8945 350984 337146
rect 351036 336320 351088 336326
rect 351036 336262 351088 336268
rect 351048 19310 351076 336262
rect 351692 148986 351720 461382
rect 353060 460148 353112 460154
rect 353060 460090 353112 460096
rect 351772 337136 351824 337142
rect 351772 337078 351824 337084
rect 351784 261526 351812 337078
rect 351772 261520 351824 261526
rect 351772 261462 351824 261468
rect 353072 195974 353100 460090
rect 354440 458924 354492 458930
rect 354440 458866 354492 458872
rect 353796 333396 353848 333402
rect 353796 333338 353848 333344
rect 353060 195968 353112 195974
rect 353060 195910 353112 195916
rect 351680 148980 351732 148986
rect 351680 148922 351732 148928
rect 351036 19304 351088 19310
rect 351036 19246 351088 19252
rect 351312 19304 351364 19310
rect 351312 19246 351364 19252
rect 351324 9761 351352 19246
rect 351310 9752 351366 9761
rect 351310 9687 351366 9696
rect 351586 9752 351642 9761
rect 351586 9687 351642 9696
rect 351128 9444 351180 9450
rect 351128 9386 351180 9392
rect 351140 9217 351168 9386
rect 351126 9208 351182 9217
rect 351126 9143 351182 9152
rect 351218 9072 351274 9081
rect 351218 9007 351220 9016
rect 351272 9007 351274 9016
rect 351220 8978 351272 8984
rect 351036 8968 351088 8974
rect 350942 8936 350998 8945
rect 351088 8916 351168 8922
rect 351036 8910 351168 8916
rect 351048 8894 351168 8910
rect 350942 8871 350998 8880
rect 351034 8392 351090 8401
rect 351140 8362 351168 8894
rect 351034 8327 351036 8336
rect 351088 8327 351090 8336
rect 351128 8356 351180 8362
rect 351036 8298 351088 8304
rect 351128 8298 351180 8304
rect 350852 8016 350904 8022
rect 350852 7958 350904 7964
rect 350668 7948 350720 7954
rect 350668 7890 350720 7896
rect 350680 7721 350708 7890
rect 350864 7857 350892 7958
rect 350850 7848 350906 7857
rect 350850 7783 350906 7792
rect 350666 7712 350722 7721
rect 350666 7647 350722 7656
rect 350942 5264 350998 5273
rect 350942 5199 350998 5208
rect 350956 5166 350984 5199
rect 350852 5160 350904 5166
rect 350850 5128 350852 5137
rect 350944 5160 350996 5166
rect 350904 5128 350906 5137
rect 350944 5102 350996 5108
rect 350850 5063 350906 5072
rect 350666 4992 350722 5001
rect 350666 4927 350722 4936
rect 350574 4856 350630 4865
rect 350574 4791 350630 4800
rect 350588 4758 350616 4791
rect 350576 4752 350628 4758
rect 350576 4694 350628 4700
rect 350680 4690 350708 4927
rect 351600 4842 351628 9687
rect 353060 8356 353112 8362
rect 353060 8298 353112 8304
rect 351600 4814 351904 4842
rect 350944 4752 350996 4758
rect 350944 4694 350996 4700
rect 350668 4684 350720 4690
rect 350668 4626 350720 4632
rect 350852 4684 350904 4690
rect 350852 4626 350904 4632
rect 350864 4457 350892 4626
rect 350956 4593 350984 4694
rect 350942 4584 350998 4593
rect 350942 4519 350998 4528
rect 350850 4448 350906 4457
rect 350850 4383 350906 4392
rect 351128 3528 351180 3534
rect 351128 3470 351180 3476
rect 351140 3233 351168 3470
rect 351126 3224 351182 3233
rect 351126 3159 351182 3168
rect 349656 2440 349708 2446
rect 349656 2382 349708 2388
rect 350760 2440 350812 2446
rect 350760 2382 350812 2388
rect 350772 480 350800 2382
rect 351876 480 351904 4814
rect 353072 480 353100 8298
rect 353808 1154 353836 333338
rect 354452 289814 354480 458866
rect 354544 368490 354572 463286
rect 355820 459944 355872 459950
rect 355820 459886 355872 459892
rect 354532 368484 354584 368490
rect 354532 368426 354584 368432
rect 355832 336666 355860 459886
rect 355924 415410 355952 463558
rect 358672 463412 358724 463418
rect 358672 463354 358724 463360
rect 357200 462868 357252 462874
rect 357200 462810 357252 462816
rect 355912 415404 355964 415410
rect 355912 415346 355964 415352
rect 357212 353258 357240 462810
rect 358580 459876 358632 459882
rect 358580 459818 358632 459824
rect 357200 353252 357252 353258
rect 357200 353194 357252 353200
rect 356556 338088 356608 338094
rect 356556 338030 356608 338036
rect 355820 336660 355872 336666
rect 355820 336602 355872 336608
rect 355176 330676 355228 330682
rect 355176 330618 355228 330624
rect 354440 289808 354492 289814
rect 354440 289750 354492 289756
rect 355188 2802 355216 330618
rect 356188 8424 356240 8430
rect 356188 8366 356240 8372
rect 356200 7721 356228 8366
rect 356186 7712 356242 7721
rect 356186 7647 356242 7656
rect 356462 7440 356518 7449
rect 356462 7375 356464 7384
rect 356516 7375 356518 7384
rect 356464 7346 356516 7352
rect 356462 6488 356518 6497
rect 356462 6423 356518 6432
rect 356476 6322 356504 6423
rect 356464 6316 356516 6322
rect 356464 6258 356516 6264
rect 355818 4856 355874 4865
rect 355818 4791 355874 4800
rect 355832 4593 355860 4791
rect 355818 4584 355874 4593
rect 355818 4519 355874 4528
rect 355268 2984 355320 2990
rect 355266 2952 355268 2961
rect 355320 2952 355322 2961
rect 355266 2887 355322 2896
rect 355188 2774 355308 2802
rect 355280 2666 355308 2774
rect 355280 2638 355492 2666
rect 353796 1148 353848 1154
rect 353796 1090 353848 1096
rect 354256 1148 354308 1154
rect 354256 1090 354308 1096
rect 354268 480 354296 1090
rect 355464 480 355492 2638
rect 356568 1426 356596 338030
rect 357936 336116 357988 336122
rect 357936 336058 357988 336064
rect 357948 309126 357976 336058
rect 357936 309120 357988 309126
rect 357936 309062 357988 309068
rect 357936 299532 357988 299538
rect 357936 299474 357988 299480
rect 357948 289746 357976 299474
rect 357936 289740 357988 289746
rect 357936 289682 357988 289688
rect 357936 280356 357988 280362
rect 357936 280298 357988 280304
rect 357948 270502 357976 280298
rect 358592 274650 358620 459818
rect 358684 400178 358712 463354
rect 359972 447098 360000 463626
rect 378832 463282 378860 470614
rect 378820 463276 378872 463282
rect 378820 463218 378872 463224
rect 508552 463146 508580 470614
rect 508540 463140 508592 463146
rect 508540 463082 508592 463088
rect 580666 461408 580722 461417
rect 580666 461343 580722 461352
rect 361340 461236 361392 461242
rect 361340 461178 361392 461184
rect 359960 447092 360012 447098
rect 359960 447034 360012 447040
rect 358672 400172 358724 400178
rect 358672 400114 358724 400120
rect 360602 320648 360658 320657
rect 360658 320606 360736 320634
rect 360602 320583 360658 320592
rect 360708 320385 360736 320606
rect 360694 320376 360750 320385
rect 360694 320311 360750 320320
rect 360696 314016 360748 314022
rect 360696 313958 360748 313964
rect 358580 274644 358632 274650
rect 358580 274586 358632 274592
rect 357936 270496 357988 270502
rect 357936 270438 357988 270444
rect 357936 260908 357988 260914
rect 357936 260850 357988 260856
rect 357948 251190 357976 260850
rect 357936 251184 357988 251190
rect 357936 251126 357988 251132
rect 357936 241664 357988 241670
rect 357936 241606 357988 241612
rect 357948 231849 357976 241606
rect 357934 231840 357990 231849
rect 357934 231775 357990 231784
rect 358118 231840 358174 231849
rect 358118 231775 358174 231784
rect 358132 222222 358160 231775
rect 360604 226568 360656 226574
rect 360602 226536 360604 226545
rect 360656 226536 360658 226545
rect 360602 226471 360658 226480
rect 357936 222216 357988 222222
rect 357936 222158 357988 222164
rect 358120 222216 358172 222222
rect 358120 222158 358172 222164
rect 357948 212498 357976 222158
rect 357936 212492 357988 212498
rect 357936 212434 357988 212440
rect 357936 203040 357988 203046
rect 357936 202982 357988 202988
rect 357948 193225 357976 202982
rect 357934 193216 357990 193225
rect 357934 193151 357990 193160
rect 358118 193216 358174 193225
rect 358118 193151 358174 193160
rect 358132 183598 358160 193151
rect 357936 183592 357988 183598
rect 357936 183534 357988 183540
rect 358120 183592 358172 183598
rect 358120 183534 358172 183540
rect 357948 173913 357976 183534
rect 357934 173904 357990 173913
rect 357934 173839 357990 173848
rect 357934 164384 357990 164393
rect 357934 164319 357990 164328
rect 357948 154465 357976 164319
rect 357934 154456 357990 154465
rect 357934 154391 357990 154400
rect 358210 154456 358266 154465
rect 358210 154391 358266 154400
rect 358224 144945 358252 154391
rect 357934 144936 357990 144945
rect 357934 144871 357990 144880
rect 358210 144936 358266 144945
rect 358210 144871 358266 144880
rect 357948 115802 357976 144871
rect 357936 115796 357988 115802
rect 357936 115738 357988 115744
rect 357936 106344 357988 106350
rect 357936 106286 357988 106292
rect 357948 96626 357976 106286
rect 360418 101008 360474 101017
rect 360418 100943 360420 100952
rect 360472 100943 360474 100952
rect 360420 100914 360472 100920
rect 357936 96620 357988 96626
rect 357936 96562 357988 96568
rect 358212 96620 358264 96626
rect 358212 96562 358264 96568
rect 358224 87145 358252 96562
rect 358210 87136 358266 87145
rect 358210 87071 358266 87080
rect 357934 87000 357990 87009
rect 357934 86935 357990 86944
rect 357948 77178 357976 86935
rect 357936 77172 357988 77178
rect 357936 77114 357988 77120
rect 357936 67652 357988 67658
rect 357936 67594 357988 67600
rect 357948 57934 357976 67594
rect 357936 57928 357988 57934
rect 357936 57870 357988 57876
rect 357936 48340 357988 48346
rect 357936 48282 357988 48288
rect 357948 38554 357976 48282
rect 357936 38548 357988 38554
rect 357936 38490 357988 38496
rect 357936 29028 357988 29034
rect 357936 28970 357988 28976
rect 356646 9072 356702 9081
rect 356646 9007 356702 9016
rect 356556 1420 356608 1426
rect 356556 1362 356608 1368
rect 356660 480 356688 9007
rect 357948 7562 357976 28970
rect 360234 8392 360290 8401
rect 360234 8327 360290 8336
rect 357948 7534 358068 7562
rect 358040 2650 358068 7534
rect 358028 2644 358080 2650
rect 358028 2586 358080 2592
rect 359040 2644 359092 2650
rect 359040 2586 359092 2592
rect 357844 1420 357896 1426
rect 357844 1362 357896 1368
rect 357856 480 357884 1362
rect 359052 480 359080 2586
rect 360248 480 360276 8327
rect 360512 3528 360564 3534
rect 360512 3470 360564 3476
rect 360604 3528 360656 3534
rect 360604 3470 360656 3476
rect 360524 3233 360552 3470
rect 360510 3224 360566 3233
rect 360510 3159 360566 3168
rect 360616 2961 360644 3470
rect 360602 2952 360658 2961
rect 360602 2887 360658 2896
rect 360708 2650 360736 313958
rect 361352 86970 361380 461178
rect 411020 461168 411072 461174
rect 411020 461110 411072 461116
rect 406880 458448 406932 458454
rect 406880 458390 406932 458396
rect 406892 383654 406920 458390
rect 411032 430574 411060 461110
rect 580680 460970 580708 461343
rect 580668 460964 580720 460970
rect 580668 460906 580720 460912
rect 580760 458244 580812 458250
rect 580760 458186 580812 458192
rect 580668 447092 580720 447098
rect 580668 447034 580720 447040
rect 580680 445777 580708 447034
rect 580666 445768 580722 445777
rect 580666 445703 580722 445712
rect 411020 430568 411072 430574
rect 411020 430510 411072 430516
rect 580668 430568 580720 430574
rect 580668 430510 580720 430516
rect 580680 430137 580708 430510
rect 580666 430128 580722 430137
rect 580666 430063 580722 430072
rect 580668 415404 580720 415410
rect 580668 415346 580720 415352
rect 580680 414497 580708 415346
rect 580666 414488 580722 414497
rect 580666 414423 580722 414432
rect 580668 400172 580720 400178
rect 580668 400114 580720 400120
rect 580680 398857 580708 400114
rect 580666 398848 580722 398857
rect 580666 398783 580722 398792
rect 406880 383648 406932 383654
rect 406880 383590 406932 383596
rect 580668 383648 580720 383654
rect 580668 383590 580720 383596
rect 580680 383217 580708 383590
rect 580666 383208 580722 383217
rect 580666 383143 580722 383152
rect 580668 368484 580720 368490
rect 580668 368426 580720 368432
rect 580680 367577 580708 368426
rect 580666 367568 580722 367577
rect 580666 367503 580722 367512
rect 580668 353252 580720 353258
rect 580668 353194 580720 353200
rect 580680 351937 580708 353194
rect 580666 351928 580722 351937
rect 580666 351863 580722 351872
rect 364836 338020 364888 338026
rect 364836 337962 364888 337968
rect 362076 327888 362128 327894
rect 362076 327830 362128 327836
rect 361340 86964 361392 86970
rect 361340 86906 361392 86912
rect 361154 8392 361210 8401
rect 361154 8327 361156 8336
rect 361208 8327 361210 8336
rect 361248 8356 361300 8362
rect 361156 8298 361208 8304
rect 361248 8298 361300 8304
rect 361260 7857 361288 8298
rect 361246 7848 361302 7857
rect 361246 7783 361302 7792
rect 360788 3528 360840 3534
rect 360788 3470 360840 3476
rect 360800 3233 360828 3470
rect 360786 3224 360842 3233
rect 360786 3159 360842 3168
rect 362088 2650 362116 327830
rect 362260 226568 362312 226574
rect 362258 226536 362260 226545
rect 362312 226536 362314 226545
rect 362258 226471 362314 226480
rect 363824 8492 363876 8498
rect 363824 8434 363876 8440
rect 363916 8492 363968 8498
rect 363916 8434 363968 8440
rect 360696 2644 360748 2650
rect 360696 2586 360748 2592
rect 361432 2644 361484 2650
rect 361432 2586 361484 2592
rect 362076 2644 362128 2650
rect 362076 2586 362128 2592
rect 362628 2644 362680 2650
rect 362628 2586 362680 2592
rect 361444 480 361472 2586
rect 362640 480 362668 2586
rect 363836 480 363864 8434
rect 363928 8401 363956 8434
rect 363914 8392 363970 8401
rect 363914 8327 363970 8336
rect 364848 7562 364876 337962
rect 378636 337748 378688 337754
rect 378636 337690 378688 337696
rect 366216 334756 366268 334762
rect 366216 334698 366268 334704
rect 366122 179616 366178 179625
rect 366122 179551 366178 179560
rect 366136 179353 366164 179551
rect 366122 179344 366178 179353
rect 366122 179279 366178 179288
rect 366124 100972 366176 100978
rect 366124 100914 366176 100920
rect 366136 100881 366164 100914
rect 366122 100872 366178 100881
rect 366122 100807 366178 100816
rect 366122 38856 366178 38865
rect 366122 38791 366178 38800
rect 366136 38593 366164 38791
rect 366122 38584 366178 38593
rect 366122 38519 366178 38528
rect 364848 7534 365060 7562
rect 364926 3496 364982 3505
rect 364926 3431 364982 3440
rect 364742 2952 364798 2961
rect 364742 2887 364798 2896
rect 364756 2854 364784 2887
rect 364940 2854 364968 3431
rect 364652 2848 364704 2854
rect 364650 2816 364652 2825
rect 364744 2848 364796 2854
rect 364704 2816 364706 2825
rect 364744 2790 364796 2796
rect 364928 2848 364980 2854
rect 364928 2790 364980 2796
rect 364650 2751 364706 2760
rect 365032 480 365060 7534
rect 366122 7032 366178 7041
rect 366122 6967 366178 6976
rect 366136 6633 366164 6967
rect 366122 6624 366178 6633
rect 366122 6559 366178 6568
rect 365294 3360 365350 3369
rect 365294 3295 365350 3304
rect 365308 2938 365336 3295
rect 365754 2952 365810 2961
rect 365308 2910 365754 2938
rect 365754 2887 365810 2896
rect 365112 2848 365164 2854
rect 365110 2816 365112 2825
rect 365164 2816 365166 2825
rect 365110 2751 365166 2760
rect 366228 480 366256 334698
rect 373024 332036 373076 332042
rect 373024 331978 373076 331984
rect 371920 331152 371972 331158
rect 371920 331094 371972 331100
rect 371932 328438 371960 331094
rect 371920 328432 371972 328438
rect 371920 328374 371972 328380
rect 373036 327078 373064 331978
rect 373024 327072 373076 327078
rect 373024 327014 373076 327020
rect 368976 325100 369028 325106
rect 368976 325042 369028 325048
rect 367596 311296 367648 311302
rect 367596 311238 367648 311244
rect 367608 22098 367636 311238
rect 368988 22098 369016 325042
rect 371920 321428 371972 321434
rect 371920 321370 371972 321376
rect 371932 318866 371960 321370
rect 371932 318838 372052 318866
rect 372024 311982 372052 318838
rect 373116 318708 373168 318714
rect 373116 318650 373168 318656
rect 372012 311976 372064 311982
rect 372012 311918 372064 311924
rect 371920 311840 371972 311846
rect 371920 311782 371972 311788
rect 371932 309126 371960 311782
rect 373128 309126 373156 318650
rect 371920 309120 371972 309126
rect 371920 309062 371972 309068
rect 373116 309120 373168 309126
rect 373116 309062 373168 309068
rect 373208 309120 373260 309126
rect 373208 309062 373260 309068
rect 373220 307766 373248 309062
rect 372932 307760 372984 307766
rect 372932 307702 372984 307708
rect 373208 307760 373260 307766
rect 373208 307702 373260 307708
rect 371828 302184 371880 302190
rect 371828 302126 371880 302132
rect 371840 292618 371868 302126
rect 372944 298217 372972 307702
rect 372930 298208 372986 298217
rect 372930 298143 372986 298152
rect 373114 298208 373170 298217
rect 373114 298143 373170 298152
rect 373128 298058 373156 298143
rect 373036 298030 373156 298058
rect 373036 296721 373064 298030
rect 374496 297492 374548 297498
rect 374496 297434 374548 297440
rect 372838 296712 372894 296721
rect 372838 296647 372894 296656
rect 373022 296712 373078 296721
rect 373022 296647 373078 296656
rect 371840 292590 371960 292618
rect 371932 289746 371960 292590
rect 371920 289740 371972 289746
rect 371920 289682 371972 289688
rect 372852 288250 372880 296647
rect 372840 288244 372892 288250
rect 372840 288186 372892 288192
rect 373116 288244 373168 288250
rect 373116 288186 373168 288192
rect 371920 282804 371972 282810
rect 371920 282746 371972 282752
rect 371932 280242 371960 282746
rect 373128 280294 373156 288186
rect 373116 280288 373168 280294
rect 371932 280214 372052 280242
rect 373116 280230 373168 280236
rect 372024 273358 372052 280214
rect 372932 278792 372984 278798
rect 372932 278734 372984 278740
rect 372012 273352 372064 273358
rect 372012 273294 372064 273300
rect 371920 273216 371972 273222
rect 371920 273158 371972 273164
rect 371932 264330 371960 273158
rect 372944 269142 372972 278734
rect 372932 269136 372984 269142
rect 372932 269078 372984 269084
rect 373116 269136 373168 269142
rect 373116 269078 373168 269084
rect 371932 264302 372144 264330
rect 372116 253978 372144 264302
rect 373128 264194 373156 269078
rect 372944 264166 373156 264194
rect 371920 253972 371972 253978
rect 371920 253914 371972 253920
rect 372104 253972 372156 253978
rect 372104 253914 372156 253920
rect 371932 244202 371960 253914
rect 372944 249830 372972 264166
rect 372932 249824 372984 249830
rect 372932 249766 372984 249772
rect 373116 249824 373168 249830
rect 373116 249766 373168 249772
rect 371840 244174 371960 244202
rect 371840 234734 371868 244174
rect 371828 234728 371880 234734
rect 371828 234670 371880 234676
rect 371736 234592 371788 234598
rect 371736 234534 371788 234540
rect 371748 231849 371776 234534
rect 373128 231849 373156 249766
rect 371550 231840 371606 231849
rect 371550 231775 371606 231784
rect 371734 231840 371790 231849
rect 371734 231775 371790 231784
rect 373114 231840 373170 231849
rect 373114 231775 373170 231784
rect 373298 231840 373354 231849
rect 373298 231775 373354 231784
rect 371564 222222 371592 231775
rect 371552 222216 371604 222222
rect 371552 222158 371604 222164
rect 371828 222216 371880 222222
rect 373312 222170 373340 231775
rect 371828 222158 371880 222164
rect 371840 217274 371868 222158
rect 373220 222142 373340 222170
rect 373220 220794 373248 222142
rect 373208 220788 373260 220794
rect 373208 220730 373260 220736
rect 371840 217246 371960 217274
rect 371932 206258 371960 217246
rect 373208 212492 373260 212498
rect 373208 212434 373260 212440
rect 371840 206230 371960 206258
rect 371840 201498 371868 206230
rect 373220 203538 373248 212434
rect 373128 203510 373248 203538
rect 371840 201470 372052 201498
rect 372024 200122 372052 201470
rect 373128 200122 373156 203510
rect 372012 200116 372064 200122
rect 372012 200058 372064 200064
rect 373116 200116 373168 200122
rect 373116 200058 373168 200064
rect 372012 191276 372064 191282
rect 372012 191218 372064 191224
rect 372024 180810 372052 191218
rect 373024 190596 373076 190602
rect 373024 190538 373076 190544
rect 373036 185586 373064 190538
rect 373036 185558 373248 185586
rect 373220 180826 373248 185558
rect 371920 180804 371972 180810
rect 371920 180746 371972 180752
rect 372012 180804 372064 180810
rect 373220 180798 373340 180826
rect 372012 180746 372064 180752
rect 370262 179616 370318 179625
rect 370318 179574 370488 179602
rect 370262 179551 370318 179560
rect 370460 179489 370488 179574
rect 370446 179480 370502 179489
rect 370446 179415 370502 179424
rect 371932 179382 371960 180746
rect 371920 179376 371972 179382
rect 371920 179318 371972 179324
rect 373312 172553 373340 180798
rect 373114 172544 373170 172553
rect 373114 172479 373170 172488
rect 373298 172544 373354 172553
rect 373298 172479 373354 172488
rect 372012 161492 372064 161498
rect 372012 161434 372064 161440
rect 372024 153270 372052 161434
rect 372012 153264 372064 153270
rect 372012 153206 372064 153212
rect 373128 153202 373156 172479
rect 371920 153196 371972 153202
rect 371920 153138 371972 153144
rect 373116 153196 373168 153202
rect 373116 153138 373168 153144
rect 371932 148322 371960 153138
rect 371840 148294 371960 148322
rect 371840 138038 371868 148294
rect 373116 145172 373168 145178
rect 373116 145114 373168 145120
rect 373128 143546 373156 145114
rect 373024 143540 373076 143546
rect 373024 143482 373076 143488
rect 373116 143540 373168 143546
rect 373116 143482 373168 143488
rect 371828 138032 371880 138038
rect 371828 137974 371880 137980
rect 371920 137964 371972 137970
rect 371920 137906 371972 137912
rect 371932 135250 371960 137906
rect 371920 135244 371972 135250
rect 371920 135186 371972 135192
rect 373036 133929 373064 143482
rect 373022 133920 373078 133929
rect 373022 133855 373078 133864
rect 373298 133920 373354 133929
rect 373298 133855 373354 133864
rect 371920 128308 371972 128314
rect 371920 128250 371972 128256
rect 371932 125610 371960 128250
rect 373312 125769 373340 133855
rect 373298 125760 373354 125769
rect 373298 125695 373354 125704
rect 373114 125624 373170 125633
rect 371932 125582 372052 125610
rect 372024 120578 372052 125582
rect 373114 125559 373170 125568
rect 373128 124166 373156 125559
rect 373116 124160 373168 124166
rect 373116 124102 373168 124108
rect 371932 120550 372052 120578
rect 371932 104922 371960 120550
rect 373116 114572 373168 114578
rect 373116 114514 373168 114520
rect 371828 104916 371880 104922
rect 371828 104858 371880 104864
rect 371920 104916 371972 104922
rect 371920 104858 371972 104864
rect 371840 104802 371868 104858
rect 373128 104854 373156 114514
rect 373116 104848 373168 104854
rect 371840 104774 372052 104802
rect 373116 104790 373168 104796
rect 372024 95334 372052 104774
rect 371920 95328 371972 95334
rect 371920 95270 371972 95276
rect 372012 95328 372064 95334
rect 372012 95270 372064 95276
rect 373116 95328 373168 95334
rect 373116 95270 373168 95276
rect 371932 95130 371960 95270
rect 371920 95124 371972 95130
rect 371920 95066 371972 95072
rect 372012 85604 372064 85610
rect 372012 85546 372064 85552
rect 372024 85513 372052 85546
rect 373128 85542 373156 95270
rect 373116 85536 373168 85542
rect 371826 85504 371882 85513
rect 371826 85439 371882 85448
rect 372010 85504 372066 85513
rect 373116 85478 373168 85484
rect 372010 85439 372066 85448
rect 371840 80050 371868 85439
rect 371840 80022 371960 80050
rect 371932 72214 371960 80022
rect 373116 75948 373168 75954
rect 373116 75890 373168 75896
rect 371920 72208 371972 72214
rect 371920 72150 371972 72156
rect 372104 72208 372156 72214
rect 372104 72150 372156 72156
rect 372116 66314 372144 72150
rect 373128 71482 373156 75890
rect 373128 71454 373248 71482
rect 372024 66286 372144 66314
rect 373220 66298 373248 71454
rect 373208 66292 373260 66298
rect 372024 64870 372052 66286
rect 373208 66234 373260 66240
rect 373300 66292 373352 66298
rect 373300 66234 373352 66240
rect 372012 64864 372064 64870
rect 372012 64806 372064 64812
rect 373312 56710 373340 66234
rect 373116 56704 373168 56710
rect 373116 56646 373168 56652
rect 373300 56704 373352 56710
rect 373300 56646 373352 56652
rect 371920 55276 371972 55282
rect 371920 55218 371972 55224
rect 371932 51762 371960 55218
rect 373128 51762 373156 56646
rect 371932 51734 372052 51762
rect 370262 38856 370318 38865
rect 370318 38814 370488 38842
rect 370262 38791 370318 38800
rect 370460 38729 370488 38814
rect 370446 38720 370502 38729
rect 370446 38655 370502 38664
rect 372024 37330 372052 51734
rect 373036 51734 373156 51762
rect 373036 37330 373064 51734
rect 371920 37324 371972 37330
rect 371920 37266 371972 37272
rect 372012 37324 372064 37330
rect 372012 37266 372064 37272
rect 373024 37324 373076 37330
rect 373024 37266 373076 37272
rect 373116 37324 373168 37330
rect 373116 37266 373168 37272
rect 371932 37210 371960 37266
rect 371932 37182 372052 37210
rect 372024 22114 372052 37182
rect 367596 22092 367648 22098
rect 367596 22034 367648 22040
rect 368332 22092 368384 22098
rect 368332 22034 368384 22040
rect 368976 22092 369028 22098
rect 368976 22034 369028 22040
rect 369528 22092 369580 22098
rect 369528 22034 369580 22040
rect 371840 22086 372052 22114
rect 368344 21978 368372 22034
rect 369540 21978 369568 22034
rect 371840 21978 371868 22086
rect 368344 21950 368464 21978
rect 369540 21950 369660 21978
rect 371840 21950 372052 21978
rect 367412 8492 367464 8498
rect 367412 8434 367464 8440
rect 367424 480 367452 8434
rect 368436 4162 368464 21950
rect 368436 4134 368556 4162
rect 368528 480 368556 4134
rect 369632 2530 369660 21950
rect 370816 8560 370868 8566
rect 370816 8502 370868 8508
rect 370356 8424 370408 8430
rect 370356 8366 370408 8372
rect 370368 7721 370396 8366
rect 370354 7712 370410 7721
rect 370354 7647 370410 7656
rect 370356 6180 370408 6186
rect 370356 6122 370408 6128
rect 370448 6180 370500 6186
rect 370448 6122 370500 6128
rect 370368 5953 370396 6122
rect 370460 6089 370488 6122
rect 370446 6080 370502 6089
rect 370446 6015 370502 6024
rect 370354 5944 370410 5953
rect 370354 5879 370410 5888
rect 370828 4978 370856 8502
rect 371000 5636 371052 5642
rect 371000 5578 371052 5584
rect 370908 5568 370960 5574
rect 370908 5510 370960 5516
rect 370920 5137 370948 5510
rect 370906 5128 370962 5137
rect 370906 5063 370962 5072
rect 371012 5001 371040 5578
rect 370998 4992 371054 5001
rect 370828 4950 370948 4978
rect 370632 3596 370684 3602
rect 370632 3538 370684 3544
rect 370172 3528 370224 3534
rect 370264 3528 370316 3534
rect 370172 3470 370224 3476
rect 370262 3496 370264 3505
rect 370540 3528 370592 3534
rect 370316 3496 370318 3505
rect 370184 3233 370212 3470
rect 370540 3470 370592 3476
rect 370262 3431 370318 3440
rect 370170 3224 370226 3233
rect 370170 3159 370226 3168
rect 370552 3097 370580 3470
rect 370644 3233 370672 3538
rect 370630 3224 370686 3233
rect 370630 3159 370686 3168
rect 370538 3088 370594 3097
rect 370538 3023 370594 3032
rect 369632 2502 369752 2530
rect 369724 480 369752 2502
rect 370920 480 370948 4950
rect 370998 4927 371054 4936
rect 372024 2530 372052 21950
rect 373128 17882 373156 37266
rect 373116 17876 373168 17882
rect 373116 17818 373168 17824
rect 374508 8430 374536 297434
rect 375876 132592 375928 132598
rect 375874 132560 375876 132569
rect 375928 132560 375930 132569
rect 375874 132495 375930 132504
rect 377348 38752 377400 38758
rect 377346 38720 377348 38729
rect 377400 38720 377402 38729
rect 377346 38655 377402 38664
rect 378084 8832 378136 8838
rect 378084 8774 378136 8780
rect 374588 8628 374640 8634
rect 374588 8570 374640 8576
rect 373116 8424 373168 8430
rect 373116 8366 373168 8372
rect 374496 8424 374548 8430
rect 374496 8366 374548 8372
rect 373128 2802 373156 8366
rect 374600 8242 374628 8570
rect 375692 8424 375744 8430
rect 375692 8366 375744 8372
rect 373036 2774 373156 2802
rect 374508 8214 374628 8242
rect 373036 2530 373064 2774
rect 372024 2502 372144 2530
rect 373036 2502 373340 2530
rect 372116 480 372144 2502
rect 373312 480 373340 2502
rect 374508 480 374536 8214
rect 375138 3496 375194 3505
rect 375138 3431 375194 3440
rect 375152 2961 375180 3431
rect 375138 2952 375194 2961
rect 375138 2887 375194 2896
rect 375704 480 375732 8366
rect 376886 5944 376942 5953
rect 376886 5879 376942 5888
rect 375782 3360 375838 3369
rect 375966 3360 376022 3369
rect 375838 3318 375966 3346
rect 375782 3295 375838 3304
rect 375966 3295 376022 3304
rect 376900 480 376928 5879
rect 378096 480 378124 8774
rect 378648 610 378676 337690
rect 385536 337680 385588 337686
rect 385536 337622 385588 337628
rect 385548 319161 385576 337622
rect 392436 337612 392488 337618
rect 392436 337554 392488 337560
rect 392448 336705 392476 337554
rect 400716 337544 400768 337550
rect 400716 337486 400768 337492
rect 392250 336696 392306 336705
rect 392250 336631 392306 336640
rect 392434 336696 392490 336705
rect 392434 336631 392490 336640
rect 392264 327146 392292 336631
rect 392252 327140 392304 327146
rect 392252 327082 392304 327088
rect 392436 327140 392488 327146
rect 392436 327082 392488 327088
rect 385534 319152 385590 319161
rect 385534 319087 385590 319096
rect 385534 318880 385590 318889
rect 385534 318815 385590 318824
rect 385548 317422 385576 318815
rect 392448 317422 392476 327082
rect 399336 323604 399388 323610
rect 399336 323546 399388 323552
rect 395196 319592 395248 319598
rect 395196 319534 395248 319540
rect 385536 317416 385588 317422
rect 385536 317358 385588 317364
rect 392436 317416 392488 317422
rect 392436 317358 392488 317364
rect 385536 307828 385588 307834
rect 385536 307770 385588 307776
rect 392436 307828 392488 307834
rect 392436 307770 392488 307776
rect 385548 298081 385576 307770
rect 392448 298081 392476 307770
rect 385534 298072 385590 298081
rect 385534 298007 385590 298016
rect 385718 298072 385774 298081
rect 385718 298007 385774 298016
rect 392434 298072 392490 298081
rect 392434 298007 392490 298016
rect 392618 298072 392674 298081
rect 392618 298007 392674 298016
rect 385732 288454 385760 298007
rect 392632 288454 392660 298007
rect 385536 288448 385588 288454
rect 385536 288390 385588 288396
rect 385720 288448 385772 288454
rect 385720 288390 385772 288396
rect 392436 288448 392488 288454
rect 392436 288390 392488 288396
rect 392620 288448 392672 288454
rect 392620 288390 392672 288396
rect 385548 278769 385576 288390
rect 392448 278769 392476 288390
rect 385534 278760 385590 278769
rect 385534 278695 385590 278704
rect 385718 278760 385774 278769
rect 385718 278695 385774 278704
rect 392434 278760 392490 278769
rect 392434 278695 392490 278704
rect 392618 278760 392674 278769
rect 392618 278695 392674 278704
rect 385732 269142 385760 278695
rect 392632 269142 392660 278695
rect 385536 269136 385588 269142
rect 385536 269078 385588 269084
rect 385720 269136 385772 269142
rect 385720 269078 385772 269084
rect 392436 269136 392488 269142
rect 392436 269078 392488 269084
rect 392620 269136 392672 269142
rect 392620 269078 392672 269084
rect 385548 259457 385576 269078
rect 392448 259457 392476 269078
rect 385534 259448 385590 259457
rect 385534 259383 385590 259392
rect 385718 259448 385774 259457
rect 385718 259383 385774 259392
rect 392434 259448 392490 259457
rect 392434 259383 392490 259392
rect 392618 259448 392674 259457
rect 392618 259383 392674 259392
rect 385732 249830 385760 259383
rect 392632 249830 392660 259383
rect 385536 249824 385588 249830
rect 385536 249766 385588 249772
rect 385720 249824 385772 249830
rect 385720 249766 385772 249772
rect 392436 249824 392488 249830
rect 392436 249766 392488 249772
rect 392620 249824 392672 249830
rect 392620 249766 392672 249772
rect 384062 242176 384118 242185
rect 384062 242111 384118 242120
rect 384076 241913 384104 242111
rect 384062 241904 384118 241913
rect 384062 241839 384118 241848
rect 385548 240145 385576 249766
rect 392448 240145 392476 249766
rect 385534 240136 385590 240145
rect 385534 240071 385590 240080
rect 385718 240136 385774 240145
rect 385718 240071 385774 240080
rect 392434 240136 392490 240145
rect 392434 240071 392490 240080
rect 392618 240136 392674 240145
rect 392618 240071 392674 240080
rect 385732 230518 385760 240071
rect 392632 230518 392660 240071
rect 385536 230512 385588 230518
rect 385536 230454 385588 230460
rect 385720 230512 385772 230518
rect 385720 230454 385772 230460
rect 392436 230512 392488 230518
rect 392436 230454 392488 230460
rect 392620 230512 392672 230518
rect 392620 230454 392672 230460
rect 385548 220833 385576 230454
rect 392448 220833 392476 230454
rect 385534 220824 385590 220833
rect 385534 220759 385590 220768
rect 385718 220824 385774 220833
rect 385718 220759 385774 220768
rect 392434 220824 392490 220833
rect 392434 220759 392490 220768
rect 392618 220824 392674 220833
rect 392618 220759 392674 220768
rect 385732 211206 385760 220759
rect 392632 211206 392660 220759
rect 385536 211200 385588 211206
rect 385536 211142 385588 211148
rect 385720 211200 385772 211206
rect 385720 211142 385772 211148
rect 392436 211200 392488 211206
rect 392436 211142 392488 211148
rect 392620 211200 392672 211206
rect 392620 211142 392672 211148
rect 385548 201482 385576 211142
rect 392448 201482 392476 211142
rect 385536 201476 385588 201482
rect 385536 201418 385588 201424
rect 385720 201476 385772 201482
rect 385720 201418 385772 201424
rect 392436 201476 392488 201482
rect 392436 201418 392488 201424
rect 392620 201476 392672 201482
rect 392620 201418 392672 201424
rect 385732 191865 385760 201418
rect 392632 191865 392660 201418
rect 385534 191856 385590 191865
rect 385534 191791 385590 191800
rect 385718 191856 385774 191865
rect 385718 191791 385774 191800
rect 392434 191856 392490 191865
rect 392434 191791 392490 191800
rect 392618 191856 392674 191865
rect 392618 191791 392674 191800
rect 385548 182170 385576 191791
rect 392448 182170 392476 191791
rect 385536 182164 385588 182170
rect 385536 182106 385588 182112
rect 385720 182164 385772 182170
rect 385720 182106 385772 182112
rect 392436 182164 392488 182170
rect 392436 182106 392488 182112
rect 392620 182164 392672 182170
rect 392620 182106 392672 182112
rect 380106 179616 380162 179625
rect 379936 179574 380106 179602
rect 379936 179489 379964 179574
rect 380106 179551 380162 179560
rect 379922 179480 379978 179489
rect 379922 179415 379978 179424
rect 385732 172553 385760 182106
rect 391698 179888 391754 179897
rect 391698 179823 391754 179832
rect 391712 179489 391740 179823
rect 391698 179480 391754 179489
rect 391698 179415 391754 179424
rect 392632 172553 392660 182106
rect 385534 172544 385590 172553
rect 385534 172479 385590 172488
rect 385718 172544 385774 172553
rect 385718 172479 385774 172488
rect 392434 172544 392490 172553
rect 392434 172479 392490 172488
rect 392618 172544 392674 172553
rect 392618 172479 392674 172488
rect 385548 164529 385576 172479
rect 392448 164529 392476 172479
rect 385534 164520 385590 164529
rect 385534 164455 385590 164464
rect 392434 164520 392490 164529
rect 392434 164455 392490 164464
rect 382040 164416 382092 164422
rect 382040 164358 382092 164364
rect 385812 164416 385864 164422
rect 385812 164358 385864 164364
rect 391700 164416 391752 164422
rect 391700 164358 391752 164364
rect 392712 164416 392764 164422
rect 392712 164358 392764 164364
rect 382052 164257 382080 164358
rect 385824 164257 385852 164358
rect 391712 164257 391740 164358
rect 392724 164257 392752 164358
rect 382038 164248 382094 164257
rect 382038 164183 382094 164192
rect 385534 164248 385590 164257
rect 385534 164183 385590 164192
rect 385810 164248 385866 164257
rect 385810 164183 385866 164192
rect 391698 164248 391754 164257
rect 391698 164183 391754 164192
rect 392434 164248 392490 164257
rect 392434 164183 392490 164192
rect 392710 164248 392766 164257
rect 392710 164183 392766 164192
rect 385548 162858 385576 164183
rect 392448 162858 392476 164183
rect 385536 162852 385588 162858
rect 385536 162794 385588 162800
rect 392436 162852 392488 162858
rect 392436 162794 392488 162800
rect 385536 153264 385588 153270
rect 385536 153206 385588 153212
rect 392436 153264 392488 153270
rect 392436 153206 392488 153212
rect 385548 143546 385576 153206
rect 392448 143546 392476 153206
rect 385536 143540 385588 143546
rect 385536 143482 385588 143488
rect 392436 143540 392488 143546
rect 392436 143482 392488 143488
rect 385536 133952 385588 133958
rect 385536 133894 385588 133900
rect 392436 133952 392488 133958
rect 392436 133894 392488 133900
rect 385442 132696 385498 132705
rect 385442 132631 385498 132640
rect 385456 132598 385484 132631
rect 385444 132592 385496 132598
rect 385444 132534 385496 132540
rect 385548 124166 385576 133894
rect 390318 132968 390374 132977
rect 390318 132903 390374 132912
rect 390332 132569 390360 132903
rect 390318 132560 390374 132569
rect 390318 132495 390374 132504
rect 392448 124166 392476 133894
rect 385536 124160 385588 124166
rect 385536 124102 385588 124108
rect 392436 124160 392488 124166
rect 392436 124102 392488 124108
rect 385536 114572 385588 114578
rect 385536 114514 385588 114520
rect 392436 114572 392488 114578
rect 392436 114514 392488 114520
rect 385548 104854 385576 114514
rect 392448 104854 392476 114514
rect 385536 104848 385588 104854
rect 385536 104790 385588 104796
rect 392436 104848 392488 104854
rect 392436 104790 392488 104796
rect 386822 101416 386878 101425
rect 386822 101351 386878 101360
rect 386836 101017 386864 101351
rect 391698 101280 391754 101289
rect 391698 101215 391754 101224
rect 386822 101008 386878 101017
rect 386822 100943 386878 100952
rect 391712 100881 391740 101215
rect 391698 100872 391754 100881
rect 391698 100807 391754 100816
rect 385536 95328 385588 95334
rect 385536 95270 385588 95276
rect 392436 95328 392488 95334
rect 392436 95270 392488 95276
rect 385548 85542 385576 95270
rect 392448 85542 392476 95270
rect 385536 85536 385588 85542
rect 385536 85478 385588 85484
rect 392436 85536 392488 85542
rect 392436 85478 392488 85484
rect 385536 75948 385588 75954
rect 385536 75890 385588 75896
rect 392436 75948 392488 75954
rect 392436 75890 392488 75896
rect 385548 66230 385576 75890
rect 392448 66230 392476 75890
rect 385536 66224 385588 66230
rect 385536 66166 385588 66172
rect 392436 66224 392488 66230
rect 392436 66166 392488 66172
rect 385536 56704 385588 56710
rect 385536 56646 385588 56652
rect 392436 56704 392488 56710
rect 392436 56646 392488 56652
rect 385548 46918 385576 56646
rect 392448 46918 392476 56646
rect 385536 46912 385588 46918
rect 385536 46854 385588 46860
rect 392436 46912 392488 46918
rect 392436 46854 392488 46860
rect 392528 46708 392580 46714
rect 392528 46650 392580 46656
rect 382038 38856 382094 38865
rect 382038 38791 382094 38800
rect 389582 38856 389638 38865
rect 389638 38814 389808 38842
rect 389582 38791 389638 38800
rect 382052 38758 382080 38791
rect 382040 38752 382092 38758
rect 389780 38729 389808 38814
rect 382040 38694 382092 38700
rect 389766 38720 389822 38729
rect 389766 38655 389822 38664
rect 385536 37324 385588 37330
rect 385536 37266 385588 37272
rect 385548 27606 385576 37266
rect 392540 29209 392568 46650
rect 392526 29200 392582 29209
rect 392526 29135 392582 29144
rect 392434 29064 392490 29073
rect 392434 28999 392490 29008
rect 392448 27606 392476 28999
rect 385536 27600 385588 27606
rect 385536 27542 385588 27548
rect 385996 27600 386048 27606
rect 385996 27542 386048 27548
rect 392436 27600 392488 27606
rect 392436 27542 392488 27548
rect 392620 27600 392672 27606
rect 392620 27542 392672 27548
rect 386008 9761 386036 27542
rect 392632 18057 392660 27542
rect 392342 18048 392398 18057
rect 392342 17983 392398 17992
rect 392618 18048 392674 18057
rect 392618 17983 392674 17992
rect 392356 15502 392384 17983
rect 392344 15496 392396 15502
rect 392344 15438 392396 15444
rect 393540 15496 393592 15502
rect 393540 15438 393592 15444
rect 385994 9752 386050 9761
rect 385994 9687 386050 9696
rect 386362 9752 386418 9761
rect 386362 9687 386418 9696
rect 385168 9648 385220 9654
rect 385168 9590 385220 9596
rect 381672 8900 381724 8906
rect 381672 8842 381724 8848
rect 380476 2508 380528 2514
rect 380476 2450 380528 2456
rect 378636 604 378688 610
rect 378636 546 378688 552
rect 379280 604 379332 610
rect 379280 546 379332 552
rect 379292 480 379320 546
rect 380488 480 380516 2450
rect 381684 480 381712 8842
rect 382868 2644 382920 2650
rect 382868 2586 382920 2592
rect 382880 480 382908 2586
rect 384064 2440 384116 2446
rect 384064 2382 384116 2388
rect 384076 480 384104 2382
rect 385180 480 385208 9590
rect 386376 480 386404 9687
rect 388756 9580 388808 9586
rect 388756 9522 388808 9528
rect 387560 5704 387612 5710
rect 387560 5646 387612 5652
rect 387572 480 387600 5646
rect 388768 480 388796 9522
rect 392344 9512 392396 9518
rect 392344 9454 392396 9460
rect 389858 7032 389914 7041
rect 389858 6967 389914 6976
rect 389872 6633 389900 6967
rect 389858 6624 389914 6633
rect 389858 6559 389914 6568
rect 391148 5772 391200 5778
rect 391148 5714 391200 5720
rect 389952 3460 390004 3466
rect 389952 3402 390004 3408
rect 389964 480 389992 3402
rect 391160 480 391188 5714
rect 392356 480 392384 9454
rect 392434 3360 392490 3369
rect 392434 3295 392490 3304
rect 392448 2961 392476 3295
rect 392434 2952 392490 2961
rect 392434 2887 392490 2896
rect 393552 480 393580 15438
rect 394736 5840 394788 5846
rect 394736 5782 394788 5788
rect 394748 480 394776 5782
rect 395208 610 395236 319534
rect 399244 132864 399296 132870
rect 399244 132806 399296 132812
rect 399256 132705 399284 132806
rect 399242 132696 399298 132705
rect 399242 132631 399298 132640
rect 399244 38888 399296 38894
rect 399242 38856 399244 38865
rect 399296 38856 399298 38865
rect 399242 38791 399298 38800
rect 398324 5908 398376 5914
rect 398324 5850 398376 5856
rect 397128 2848 397180 2854
rect 397128 2790 397180 2796
rect 395196 604 395248 610
rect 395196 546 395248 552
rect 395932 604 395984 610
rect 395932 546 395984 552
rect 395944 480 395972 546
rect 397140 480 397168 2790
rect 398336 480 398364 5850
rect 399348 626 399376 323546
rect 399428 8424 399480 8430
rect 399428 8366 399480 8372
rect 399440 7721 399468 8366
rect 399426 7712 399482 7721
rect 399426 7647 399482 7656
rect 399348 598 399560 626
rect 399532 480 399560 598
rect 400728 480 400756 337486
rect 407616 337476 407668 337482
rect 407616 337418 407668 337424
rect 406236 318164 406288 318170
rect 406236 318106 406288 318112
rect 402096 312656 402148 312662
rect 402096 312598 402148 312604
rect 401820 6112 401872 6118
rect 401820 6054 401872 6060
rect 401832 480 401860 6054
rect 402002 3224 402058 3233
rect 402002 3159 402058 3168
rect 402016 2961 402044 3159
rect 402002 2952 402058 2961
rect 402002 2887 402058 2896
rect 402108 610 402136 312598
rect 406144 132864 406196 132870
rect 406142 132832 406144 132841
rect 406196 132832 406198 132841
rect 406142 132767 406198 132776
rect 406142 38992 406198 39001
rect 406142 38927 406198 38936
rect 406156 38894 406184 38927
rect 406144 38888 406196 38894
rect 406144 38830 406196 38836
rect 405408 6860 405460 6866
rect 405408 6802 405460 6808
rect 404212 2848 404264 2854
rect 404212 2790 404264 2796
rect 402096 604 402148 610
rect 402096 546 402148 552
rect 403016 604 403068 610
rect 403016 546 403068 552
rect 403028 480 403056 546
rect 404224 480 404252 2790
rect 405420 480 405448 6802
rect 406248 610 406276 318106
rect 406878 3224 406934 3233
rect 406878 3159 406934 3168
rect 406892 2990 406920 3159
rect 406880 2984 406932 2990
rect 406880 2926 406932 2932
rect 407628 626 407656 337418
rect 414516 337408 414568 337414
rect 414516 337350 414568 337356
rect 413136 315376 413188 315382
rect 413136 315318 413188 315324
rect 408996 286408 409048 286414
rect 408996 286350 409048 286356
rect 409008 11218 409036 286350
rect 413148 14498 413176 315318
rect 414528 19310 414556 337350
rect 580392 336660 580444 336666
rect 580392 336602 580444 336608
rect 580404 336297 580432 336602
rect 580390 336288 580446 336297
rect 580390 336223 580446 336232
rect 454536 336048 454588 336054
rect 454536 335990 454588 335996
rect 447636 329248 447688 329254
rect 447636 329190 447688 329196
rect 425462 320512 425518 320521
rect 425462 320447 425518 320456
rect 444782 320512 444838 320521
rect 444782 320447 444838 320456
rect 418562 320376 418618 320385
rect 425476 320346 425504 320447
rect 437882 320376 437938 320385
rect 418562 320311 418564 320320
rect 418616 320311 418618 320320
rect 425464 320340 425516 320346
rect 418564 320282 418616 320288
rect 444796 320346 444824 320447
rect 437882 320311 437884 320320
rect 425464 320282 425516 320288
rect 437936 320311 437938 320320
rect 444784 320340 444836 320346
rect 437884 320282 437936 320288
rect 444784 320282 444836 320288
rect 420036 316736 420088 316742
rect 420036 316678 420088 316684
rect 417368 283688 417420 283694
rect 417368 283630 417420 283636
rect 414516 19304 414568 19310
rect 414516 19246 414568 19252
rect 414884 19304 414936 19310
rect 414884 19246 414936 19252
rect 413148 14470 413268 14498
rect 408996 11212 409048 11218
rect 408996 11154 409048 11160
rect 410192 11212 410244 11218
rect 410192 11154 410244 11160
rect 408994 10568 409050 10577
rect 408994 10503 408996 10512
rect 409048 10503 409050 10512
rect 408996 10474 409048 10480
rect 409180 8424 409232 8430
rect 409180 8366 409232 8372
rect 409192 7721 409220 8366
rect 409178 7712 409234 7721
rect 409178 7647 409234 7656
rect 408996 6792 409048 6798
rect 408996 6734 409048 6740
rect 406236 604 406288 610
rect 406236 546 406288 552
rect 406604 604 406656 610
rect 407628 598 407840 626
rect 406604 546 406656 552
rect 406616 480 406644 546
rect 407812 480 407840 598
rect 409008 480 409036 6734
rect 410204 480 410232 11154
rect 413240 9761 413268 14470
rect 414896 12322 414924 19246
rect 414896 12294 415016 12322
rect 413226 9752 413282 9761
rect 413226 9687 413282 9696
rect 413778 9752 413834 9761
rect 413778 9687 413834 9696
rect 411662 7440 411718 7449
rect 411662 7375 411718 7384
rect 413042 7440 413098 7449
rect 413042 7375 413098 7384
rect 411676 7177 411704 7375
rect 411662 7168 411718 7177
rect 411662 7103 411718 7112
rect 413056 7041 413084 7375
rect 413042 7032 413098 7041
rect 413042 6967 413098 6976
rect 412584 6724 412636 6730
rect 412584 6666 412636 6672
rect 411662 3360 411718 3369
rect 411662 3295 411718 3304
rect 411676 2990 411704 3295
rect 411664 2984 411716 2990
rect 411664 2926 411716 2932
rect 411388 2916 411440 2922
rect 411388 2858 411440 2864
rect 411400 480 411428 2858
rect 412596 480 412624 6666
rect 413792 480 413820 9687
rect 414528 3454 414648 3482
rect 414528 3369 414556 3454
rect 414514 3360 414570 3369
rect 414514 3295 414570 3304
rect 414620 2990 414648 3454
rect 414608 2984 414660 2990
rect 414608 2926 414660 2932
rect 414988 480 415016 12294
rect 416172 6656 416224 6662
rect 416172 6598 416224 6604
rect 416184 480 416212 6598
rect 417380 480 417408 283630
rect 418748 10464 418800 10470
rect 418746 10432 418748 10441
rect 418800 10432 418802 10441
rect 418746 10367 418802 10376
rect 419668 6452 419720 6458
rect 419668 6394 419720 6400
rect 418838 4720 418894 4729
rect 418838 4655 418894 4664
rect 418852 4146 418880 4655
rect 418840 4140 418892 4146
rect 418840 4082 418892 4088
rect 418472 3052 418524 3058
rect 418472 2994 418524 3000
rect 418484 480 418512 2994
rect 419680 480 419708 6394
rect 420048 2854 420076 316678
rect 440736 309868 440788 309874
rect 440736 309810 440788 309816
rect 424174 10568 424230 10577
rect 424174 10503 424230 10512
rect 424082 7032 424138 7041
rect 424082 6967 424138 6976
rect 424096 6798 424124 6967
rect 424084 6792 424136 6798
rect 424084 6734 424136 6740
rect 423256 6384 423308 6390
rect 423256 6326 423308 6332
rect 422060 3120 422112 3126
rect 422060 3062 422112 3068
rect 420036 2848 420088 2854
rect 420036 2790 420088 2796
rect 420864 604 420916 610
rect 420864 546 420916 552
rect 420876 480 420904 546
rect 422072 480 422100 3062
rect 423268 480 423296 6326
rect 424082 3224 424138 3233
rect 424082 3159 424138 3168
rect 424096 2990 424124 3159
rect 424084 2984 424136 2990
rect 424084 2926 424136 2932
rect 424188 610 424216 10503
rect 437976 9920 438028 9926
rect 437976 9862 438028 9868
rect 435124 9716 435176 9722
rect 435124 9658 435176 9664
rect 431076 9648 431128 9654
rect 431076 9590 431128 9596
rect 426936 9580 426988 9586
rect 426936 9522 426988 9528
rect 426844 6112 426896 6118
rect 426844 6054 426896 6060
rect 425648 3188 425700 3194
rect 425648 3130 425700 3136
rect 424176 604 424228 610
rect 424176 546 424228 552
rect 424452 604 424504 610
rect 424452 546 424504 552
rect 424464 480 424492 546
rect 425660 480 425688 3130
rect 426856 480 426884 6054
rect 426948 610 426976 9522
rect 428958 7168 429014 7177
rect 428958 7103 429014 7112
rect 428972 6798 429000 7103
rect 428960 6792 429012 6798
rect 428960 6734 429012 6740
rect 430432 6248 430484 6254
rect 430432 6190 430484 6196
rect 429236 3392 429288 3398
rect 429236 3334 429288 3340
rect 426936 604 426988 610
rect 426936 546 426988 552
rect 428040 604 428092 610
rect 428040 546 428092 552
rect 428052 480 428080 546
rect 429248 480 429276 3334
rect 430444 480 430472 6190
rect 431088 610 431116 9590
rect 434020 6180 434072 6186
rect 434020 6122 434072 6128
rect 433558 3496 433614 3505
rect 433558 3431 433614 3440
rect 433742 3496 433798 3505
rect 433742 3431 433798 3440
rect 433572 3380 433600 3431
rect 433756 3380 433784 3431
rect 433572 3352 433784 3380
rect 433836 3392 433888 3398
rect 433834 3360 433836 3369
rect 433888 3360 433890 3369
rect 433834 3295 433890 3304
rect 432824 3120 432876 3126
rect 432824 3062 432876 3068
rect 431076 604 431128 610
rect 431076 546 431128 552
rect 431628 604 431680 610
rect 431628 546 431680 552
rect 431640 480 431668 546
rect 432836 480 432864 3062
rect 434032 480 434060 6122
rect 435136 480 435164 9658
rect 437514 6216 437570 6225
rect 437514 6151 437570 6160
rect 436320 4072 436372 4078
rect 436320 4014 436372 4020
rect 436332 480 436360 4014
rect 437528 480 437556 6151
rect 437988 626 438016 9862
rect 438252 8424 438304 8430
rect 438252 8366 438304 8372
rect 438264 7721 438292 8366
rect 438250 7712 438306 7721
rect 438250 7647 438306 7656
rect 439908 4004 439960 4010
rect 439908 3946 439960 3952
rect 437988 598 438660 626
rect 438632 592 438660 598
rect 438632 564 438752 592
rect 438724 480 438752 564
rect 439920 480 439948 3946
rect 440748 626 440776 309810
rect 443588 307148 443640 307154
rect 443588 307090 443640 307096
rect 442116 9988 442168 9994
rect 442116 9930 442168 9936
rect 440748 598 441052 626
rect 442128 610 442156 9930
rect 443496 3936 443548 3942
rect 443496 3878 443548 3884
rect 441024 592 441052 598
rect 442116 604 442168 610
rect 441024 564 441144 592
rect 441116 480 441144 564
rect 442116 546 442168 552
rect 442300 604 442352 610
rect 442300 546 442352 552
rect 442312 480 442340 546
rect 443508 480 443536 3878
rect 443600 610 443628 307090
rect 444876 10056 444928 10062
rect 444876 9998 444928 10004
rect 444888 610 444916 9998
rect 447084 3732 447136 3738
rect 447084 3674 447136 3680
rect 443588 604 443640 610
rect 443588 546 443640 552
rect 444692 604 444744 610
rect 444692 546 444744 552
rect 444876 604 444928 610
rect 444876 546 444928 552
rect 445888 604 445940 610
rect 445888 546 445940 552
rect 444704 480 444732 546
rect 445900 480 445928 546
rect 447096 480 447124 3674
rect 447648 610 447676 329190
rect 451776 304360 451828 304366
rect 451776 304302 451828 304308
rect 449016 10124 449068 10130
rect 449016 10066 449068 10072
rect 449028 610 449056 10066
rect 450672 3664 450724 3670
rect 450672 3606 450724 3612
rect 447636 604 447688 610
rect 447636 546 447688 552
rect 448280 604 448332 610
rect 448280 546 448332 552
rect 449016 604 449068 610
rect 449016 546 449068 552
rect 449476 604 449528 610
rect 449476 546 449528 552
rect 448292 480 448320 546
rect 449488 480 449516 546
rect 450684 480 450712 3606
rect 451684 3392 451736 3398
rect 451684 3334 451736 3340
rect 451696 3233 451724 3334
rect 451682 3224 451738 3233
rect 451682 3159 451738 3168
rect 451788 480 451816 304302
rect 451868 10192 451920 10198
rect 451868 10134 451920 10140
rect 451880 610 451908 10134
rect 453246 7032 453302 7041
rect 453246 6967 453302 6976
rect 453260 6730 453288 6967
rect 453248 6724 453300 6730
rect 453248 6666 453300 6672
rect 454168 3596 454220 3602
rect 454168 3538 454220 3544
rect 451868 604 451920 610
rect 451868 546 451920 552
rect 452972 604 453024 610
rect 452972 546 453024 552
rect 452984 480 453012 546
rect 454180 480 454208 3538
rect 454548 610 454576 335990
rect 548376 334688 548428 334694
rect 548376 334630 548428 334636
rect 483516 333328 483568 333334
rect 483516 333270 483568 333276
rect 465576 326528 465628 326534
rect 465576 326470 465628 326476
rect 464102 320512 464158 320521
rect 464102 320447 464158 320456
rect 457202 320376 457258 320385
rect 464116 320346 464144 320447
rect 457202 320311 457204 320320
rect 457256 320311 457258 320320
rect 464104 320340 464156 320346
rect 457204 320282 457256 320288
rect 464104 320282 464156 320288
rect 458676 301572 458728 301578
rect 458676 301514 458728 301520
rect 455916 10260 455968 10266
rect 455916 10202 455968 10208
rect 455928 626 455956 10202
rect 457756 3528 457808 3534
rect 457756 3470 457808 3476
rect 454536 604 454588 610
rect 454536 546 454588 552
rect 455364 604 455416 610
rect 455928 598 456508 626
rect 456480 592 456508 598
rect 456480 564 456600 592
rect 455364 546 455416 552
rect 455376 480 455404 546
rect 456572 480 456600 564
rect 457768 480 457796 3470
rect 458688 626 458716 301514
rect 461436 300212 461488 300218
rect 461436 300154 461488 300160
rect 460148 11008 460200 11014
rect 460148 10950 460200 10956
rect 458688 598 458900 626
rect 458872 592 458900 598
rect 458872 564 458992 592
rect 458964 480 458992 564
rect 460160 480 460188 10950
rect 461344 3460 461396 3466
rect 461344 3402 461396 3408
rect 461356 480 461384 3402
rect 461448 610 461476 300154
rect 462816 10804 462868 10810
rect 462816 10746 462868 10752
rect 462722 7032 462778 7041
rect 462722 6967 462778 6976
rect 462736 6730 462764 6967
rect 462724 6724 462776 6730
rect 462724 6666 462776 6672
rect 462722 3224 462778 3233
rect 462722 3159 462778 3168
rect 462736 3097 462764 3159
rect 462722 3088 462778 3097
rect 462722 3023 462778 3032
rect 462828 610 462856 10746
rect 464930 4040 464986 4049
rect 464930 3975 464986 3984
rect 461436 604 461488 610
rect 461436 546 461488 552
rect 462540 604 462592 610
rect 462540 546 462592 552
rect 462816 604 462868 610
rect 462816 546 462868 552
rect 463736 604 463788 610
rect 463736 546 463788 552
rect 462552 480 462580 546
rect 463748 480 463776 546
rect 464944 480 464972 3975
rect 465588 610 465616 326470
rect 483422 320512 483478 320521
rect 483422 320447 483478 320456
rect 476522 320376 476578 320385
rect 483436 320346 483464 320447
rect 476522 320311 476524 320320
rect 476576 320311 476578 320320
rect 483424 320340 483476 320346
rect 476524 320282 476576 320288
rect 483424 320282 483476 320288
rect 483528 14618 483556 333270
rect 520776 331968 520828 331974
rect 520776 331910 520828 331916
rect 486276 330608 486328 330614
rect 486276 330550 486328 330556
rect 483516 14612 483568 14618
rect 483516 14554 483568 14560
rect 483976 14612 484028 14618
rect 483976 14554 484028 14560
rect 466956 10736 467008 10742
rect 466956 10678 467008 10684
rect 466588 3392 466640 3398
rect 466588 3334 466640 3340
rect 466600 3233 466628 3334
rect 466586 3224 466642 3233
rect 466586 3159 466642 3168
rect 466968 610 466996 10678
rect 469716 10668 469768 10674
rect 469716 10610 469768 10616
rect 469624 6860 469676 6866
rect 469624 6802 469676 6808
rect 468426 3904 468482 3913
rect 468426 3839 468482 3848
rect 465576 604 465628 610
rect 465576 546 465628 552
rect 466128 604 466180 610
rect 466128 546 466180 552
rect 466956 604 467008 610
rect 466956 546 467008 552
rect 467324 604 467376 610
rect 467324 546 467376 552
rect 466140 480 466168 546
rect 467336 480 467364 546
rect 468440 480 468468 3839
rect 469636 480 469664 6802
rect 469728 610 469756 10610
rect 474408 10600 474460 10606
rect 474408 10542 474460 10548
rect 473856 7200 473908 7206
rect 473854 7168 473856 7177
rect 474224 7200 474276 7206
rect 473908 7168 473910 7177
rect 473854 7103 473910 7112
rect 474222 7168 474224 7177
rect 474276 7168 474278 7177
rect 474222 7103 474278 7112
rect 473212 6792 473264 6798
rect 473212 6734 473264 6740
rect 472014 3768 472070 3777
rect 472014 3703 472070 3712
rect 469716 604 469768 610
rect 469716 546 469768 552
rect 470820 604 470872 610
rect 470820 546 470872 552
rect 470832 480 470860 546
rect 472028 480 472056 3703
rect 473224 480 473252 6734
rect 474420 480 474448 10542
rect 477996 10532 478048 10538
rect 477996 10474 478048 10480
rect 476800 6928 476852 6934
rect 476800 6870 476852 6876
rect 475602 3632 475658 3641
rect 475602 3567 475658 3576
rect 475616 480 475644 3567
rect 476812 480 476840 6870
rect 478008 480 478036 10474
rect 481584 10464 481636 10470
rect 481584 10406 481636 10412
rect 480768 7126 480888 7154
rect 480768 7041 480796 7126
rect 480754 7032 480810 7041
rect 480388 6996 480440 7002
rect 480860 7002 480888 7126
rect 480754 6967 480810 6976
rect 480848 6996 480900 7002
rect 480388 6938 480440 6944
rect 480848 6938 480900 6944
rect 479190 3496 479246 3505
rect 479190 3431 479246 3440
rect 479204 480 479232 3431
rect 480400 480 480428 6938
rect 480664 3392 480716 3398
rect 480664 3334 480716 3340
rect 480676 3233 480704 3334
rect 480662 3224 480718 3233
rect 480662 3159 480718 3168
rect 481596 480 481624 10406
rect 483514 7032 483570 7041
rect 483514 6967 483516 6976
rect 483568 6967 483570 6976
rect 483516 6938 483568 6944
rect 482778 3224 482834 3233
rect 482778 3159 482834 3168
rect 482792 480 482820 3159
rect 483988 480 484016 14554
rect 486288 7206 486316 330550
rect 490416 327820 490468 327826
rect 490416 327762 490468 327768
rect 488300 320544 488352 320550
rect 488298 320512 488300 320521
rect 488352 320512 488354 320521
rect 488298 320447 488354 320456
rect 489864 11688 489916 11694
rect 489864 11630 489916 11636
rect 486458 10296 486514 10305
rect 486458 10231 486514 10240
rect 485080 7200 485132 7206
rect 485080 7142 485132 7148
rect 486276 7200 486328 7206
rect 486276 7142 486328 7148
rect 485092 480 485120 7142
rect 486472 7018 486500 10231
rect 488668 7268 488720 7274
rect 488668 7210 488720 7216
rect 487472 7200 487524 7206
rect 487472 7142 487524 7148
rect 486288 6990 486500 7018
rect 486288 480 486316 6990
rect 487484 480 487512 7142
rect 488680 480 488708 7210
rect 489876 480 489904 11630
rect 490428 610 490456 327762
rect 494556 325032 494608 325038
rect 494556 324974 494608 324980
rect 493084 320544 493136 320550
rect 493082 320512 493084 320521
rect 493136 320512 493138 320521
rect 493082 320447 493138 320456
rect 493176 12436 493228 12442
rect 493176 12378 493228 12384
rect 492256 7336 492308 7342
rect 492256 7278 492308 7284
rect 490416 604 490468 610
rect 490416 546 490468 552
rect 491060 604 491112 610
rect 491060 546 491112 552
rect 491072 480 491100 546
rect 492268 480 492296 7278
rect 493188 626 493216 12378
rect 493188 598 493400 626
rect 493372 592 493400 598
rect 494568 592 494596 324974
rect 497316 322312 497368 322318
rect 497316 322254 497368 322260
rect 495936 12368 495988 12374
rect 495936 12310 495988 12316
rect 495844 7404 495896 7410
rect 495844 7346 495896 7352
rect 493372 564 493492 592
rect 494568 564 494688 592
rect 493464 480 493492 564
rect 494660 480 494688 564
rect 495856 480 495884 7346
rect 495948 610 495976 12310
rect 497328 610 497356 322254
rect 505594 320512 505650 320521
rect 505650 320470 505728 320498
rect 505594 320447 505650 320456
rect 505700 320249 505728 320470
rect 505686 320240 505742 320249
rect 505686 320175 505742 320184
rect 501456 319524 501508 319530
rect 501456 319466 501508 319472
rect 500076 12300 500128 12306
rect 500076 12242 500128 12248
rect 499432 7472 499484 7478
rect 499432 7414 499484 7420
rect 495936 604 495988 610
rect 495936 546 495988 552
rect 497040 604 497092 610
rect 497040 546 497092 552
rect 497316 604 497368 610
rect 497316 546 497368 552
rect 498236 604 498288 610
rect 498236 546 498288 552
rect 497052 480 497080 546
rect 498248 480 498276 546
rect 499444 480 499472 7414
rect 500088 610 500116 12242
rect 501468 610 501496 319466
rect 504216 318096 504268 318102
rect 504216 318038 504268 318044
rect 504124 12232 504176 12238
rect 504124 12174 504176 12180
rect 502928 7540 502980 7546
rect 502928 7482 502980 7488
rect 500076 604 500128 610
rect 500076 546 500128 552
rect 500628 604 500680 610
rect 500628 546 500680 552
rect 501456 604 501508 610
rect 501456 546 501508 552
rect 501732 604 501784 610
rect 501732 546 501784 552
rect 500640 480 500668 546
rect 501744 480 501772 546
rect 502940 480 502968 7482
rect 504136 480 504164 12174
rect 504228 610 504256 318038
rect 508356 315308 508408 315314
rect 508356 315250 508408 315256
rect 506976 279472 507028 279478
rect 506976 279414 507028 279420
rect 506516 8288 506568 8294
rect 506516 8230 506568 8236
rect 504216 604 504268 610
rect 504216 546 504268 552
rect 505320 604 505372 610
rect 505320 546 505372 552
rect 505332 480 505360 546
rect 506528 480 506556 8230
rect 506988 610 507016 279414
rect 508368 610 508396 315250
rect 513876 276684 513928 276690
rect 513876 276626 513928 276632
rect 513888 12442 513916 276626
rect 513876 12436 513928 12442
rect 513876 12378 513928 12384
rect 514888 12436 514940 12442
rect 514888 12378 514940 12384
rect 511300 12164 511352 12170
rect 511300 12106 511352 12112
rect 510104 8084 510156 8090
rect 510104 8026 510156 8032
rect 506976 604 507028 610
rect 506976 546 507028 552
rect 507712 604 507764 610
rect 507712 546 507764 552
rect 508356 604 508408 610
rect 508356 546 508408 552
rect 508908 604 508960 610
rect 508908 546 508960 552
rect 507724 480 507752 546
rect 508920 480 508948 546
rect 510116 480 510144 8026
rect 511022 7576 511078 7585
rect 511022 7511 511078 7520
rect 511036 7177 511064 7511
rect 511022 7168 511078 7177
rect 511022 7103 511078 7112
rect 511312 480 511340 12106
rect 513692 8016 513744 8022
rect 513692 7958 513744 7964
rect 512496 4072 512548 4078
rect 512496 4014 512548 4020
rect 512508 480 512536 4014
rect 513704 480 513732 7958
rect 514900 480 514928 12378
rect 518384 12096 518436 12102
rect 518384 12038 518436 12044
rect 517280 7948 517332 7954
rect 517280 7890 517332 7896
rect 515256 4820 515308 4826
rect 515256 4762 515308 4768
rect 515348 4820 515400 4826
rect 515348 4762 515400 4768
rect 515268 4729 515296 4762
rect 515254 4720 515310 4729
rect 515254 4655 515310 4664
rect 515360 4282 515388 4762
rect 515348 4276 515400 4282
rect 515348 4218 515400 4224
rect 516084 4004 516136 4010
rect 516084 3946 516136 3952
rect 516096 480 516124 3946
rect 517292 480 517320 7890
rect 518396 480 518424 12038
rect 520788 7546 520816 331910
rect 530436 330540 530488 330546
rect 530436 330482 530488 330488
rect 529056 307080 529108 307086
rect 529056 307022 529108 307028
rect 529068 298081 529096 307022
rect 528870 298072 528926 298081
rect 528870 298007 528926 298016
rect 529054 298072 529110 298081
rect 529054 298007 529110 298016
rect 528884 288454 528912 298007
rect 528872 288448 528924 288454
rect 528872 288390 528924 288396
rect 529056 288448 529108 288454
rect 529056 288390 529108 288396
rect 529068 278769 529096 288390
rect 528870 278760 528926 278769
rect 528870 278695 528926 278704
rect 529054 278760 529110 278769
rect 529054 278695 529110 278704
rect 528884 269142 528912 278695
rect 528872 269136 528924 269142
rect 528872 269078 528924 269084
rect 529056 269136 529108 269142
rect 529056 269078 529108 269084
rect 529068 259457 529096 269078
rect 528870 259448 528926 259457
rect 528870 259383 528926 259392
rect 529054 259448 529110 259457
rect 529054 259383 529110 259392
rect 528884 249830 528912 259383
rect 528872 249824 528924 249830
rect 528872 249766 528924 249772
rect 529056 249824 529108 249830
rect 529056 249766 529108 249772
rect 529068 240145 529096 249766
rect 528870 240136 528926 240145
rect 528870 240071 528926 240080
rect 529054 240136 529110 240145
rect 529054 240071 529110 240080
rect 528884 230518 528912 240071
rect 528872 230512 528924 230518
rect 528872 230454 528924 230460
rect 529056 230512 529108 230518
rect 529056 230454 529108 230460
rect 529068 220833 529096 230454
rect 528870 220824 528926 220833
rect 528870 220759 528926 220768
rect 529054 220824 529110 220833
rect 529054 220759 529110 220768
rect 528884 211206 528912 220759
rect 528872 211200 528924 211206
rect 528872 211142 528924 211148
rect 529056 211200 529108 211206
rect 529056 211142 529108 211148
rect 529068 201482 529096 211142
rect 528872 201476 528924 201482
rect 528872 201418 528924 201424
rect 529056 201476 529108 201482
rect 529056 201418 529108 201424
rect 528884 191865 528912 201418
rect 528870 191856 528926 191865
rect 528870 191791 528926 191800
rect 529054 191856 529110 191865
rect 529054 191791 529110 191800
rect 529068 182170 529096 191791
rect 528872 182164 528924 182170
rect 528872 182106 528924 182112
rect 529056 182164 529108 182170
rect 529056 182106 529108 182112
rect 528884 172553 528912 182106
rect 528870 172544 528926 172553
rect 528870 172479 528926 172488
rect 529054 172544 529110 172553
rect 529054 172479 529110 172488
rect 529068 164529 529096 172479
rect 529054 164520 529110 164529
rect 529054 164455 529110 164464
rect 526940 164416 526992 164422
rect 526940 164358 526992 164364
rect 529332 164416 529384 164422
rect 529332 164358 529384 164364
rect 526952 164257 526980 164358
rect 529344 164257 529372 164358
rect 526938 164248 526994 164257
rect 526938 164183 526994 164192
rect 529054 164248 529110 164257
rect 529054 164183 529110 164192
rect 529330 164248 529386 164257
rect 529330 164183 529386 164192
rect 529068 162858 529096 164183
rect 529056 162852 529108 162858
rect 529056 162794 529108 162800
rect 529056 153264 529108 153270
rect 529056 153206 529108 153212
rect 529068 143546 529096 153206
rect 529056 143540 529108 143546
rect 529056 143482 529108 143488
rect 529056 133952 529108 133958
rect 529056 133894 529108 133900
rect 529068 124166 529096 133894
rect 529056 124160 529108 124166
rect 529056 124102 529108 124108
rect 529056 114572 529108 114578
rect 529056 114514 529108 114520
rect 529068 104854 529096 114514
rect 529056 104848 529108 104854
rect 529056 104790 529108 104796
rect 529056 95328 529108 95334
rect 529056 95270 529108 95276
rect 529068 85542 529096 95270
rect 529056 85536 529108 85542
rect 529056 85478 529108 85484
rect 529056 75948 529108 75954
rect 529056 75890 529108 75896
rect 529068 66230 529096 75890
rect 529056 66224 529108 66230
rect 529056 66166 529108 66172
rect 529056 56704 529108 56710
rect 529056 56646 529108 56652
rect 529068 46918 529096 56646
rect 529056 46912 529108 46918
rect 529056 46854 529108 46860
rect 529056 37324 529108 37330
rect 529056 37266 529108 37272
rect 529068 27606 529096 37266
rect 529056 27600 529108 27606
rect 529056 27542 529108 27548
rect 530448 12442 530476 330482
rect 541476 327752 541528 327758
rect 541476 327694 541528 327700
rect 534576 297424 534628 297430
rect 534576 297366 534628 297372
rect 534588 12442 534616 297366
rect 537336 294636 537388 294642
rect 537336 294578 537388 294584
rect 535956 269136 536008 269142
rect 535956 269078 536008 269084
rect 535968 259457 535996 269078
rect 535954 259448 536010 259457
rect 535954 259383 536010 259392
rect 536138 259448 536194 259457
rect 536138 259383 536194 259392
rect 536152 249830 536180 259383
rect 535956 249824 536008 249830
rect 535956 249766 536008 249772
rect 536140 249824 536192 249830
rect 536140 249766 536192 249772
rect 535968 240145 535996 249766
rect 535954 240136 536010 240145
rect 535954 240071 536010 240080
rect 536138 240136 536194 240145
rect 536138 240071 536194 240080
rect 536152 230518 536180 240071
rect 535956 230512 536008 230518
rect 535956 230454 536008 230460
rect 536140 230512 536192 230518
rect 536140 230454 536192 230460
rect 535968 220833 535996 230454
rect 535954 220824 536010 220833
rect 535954 220759 536010 220768
rect 536138 220824 536194 220833
rect 536138 220759 536194 220768
rect 536152 211206 536180 220759
rect 535956 211200 536008 211206
rect 535956 211142 536008 211148
rect 536140 211200 536192 211206
rect 536140 211142 536192 211148
rect 535968 201482 535996 211142
rect 535956 201476 536008 201482
rect 535956 201418 536008 201424
rect 536140 201476 536192 201482
rect 536140 201418 536192 201424
rect 536152 191865 536180 201418
rect 535954 191856 536010 191865
rect 535954 191791 536010 191800
rect 536138 191856 536194 191865
rect 536138 191791 536194 191800
rect 535968 182170 535996 191791
rect 535956 182164 536008 182170
rect 535956 182106 536008 182112
rect 536140 182164 536192 182170
rect 536140 182106 536192 182112
rect 536152 172553 536180 182106
rect 535954 172544 536010 172553
rect 535954 172479 536010 172488
rect 536138 172544 536194 172553
rect 536138 172479 536194 172488
rect 535968 164529 535996 172479
rect 535954 164520 536010 164529
rect 535954 164455 536010 164464
rect 535680 164416 535732 164422
rect 535680 164358 535732 164364
rect 536600 164416 536652 164422
rect 536600 164358 536652 164364
rect 535692 164257 535720 164358
rect 536612 164257 536640 164358
rect 535678 164248 535734 164257
rect 535678 164183 535734 164192
rect 535954 164248 536010 164257
rect 535954 164183 536010 164192
rect 536598 164248 536654 164257
rect 536598 164183 536654 164192
rect 535968 162858 535996 164183
rect 535956 162852 536008 162858
rect 535956 162794 536008 162800
rect 535956 153264 536008 153270
rect 535956 153206 536008 153212
rect 535968 143546 535996 153206
rect 535956 143540 536008 143546
rect 535956 143482 536008 143488
rect 535956 133952 536008 133958
rect 535956 133894 536008 133900
rect 535968 124166 535996 133894
rect 535956 124160 536008 124166
rect 535956 124102 536008 124108
rect 535956 114572 536008 114578
rect 535956 114514 536008 114520
rect 535968 104854 535996 114514
rect 535956 104848 536008 104854
rect 535956 104790 536008 104796
rect 535956 95328 536008 95334
rect 535956 95270 536008 95276
rect 535968 85542 535996 95270
rect 535956 85536 536008 85542
rect 535956 85478 536008 85484
rect 535956 75948 536008 75954
rect 535956 75890 536008 75896
rect 535968 66230 535996 75890
rect 535956 66224 536008 66230
rect 535956 66166 536008 66172
rect 535956 56704 536008 56710
rect 535956 56646 536008 56652
rect 535968 46918 535996 56646
rect 535956 46912 536008 46918
rect 535956 46854 536008 46860
rect 535956 37324 536008 37330
rect 535956 37266 536008 37272
rect 535968 27606 535996 37266
rect 535956 27600 536008 27606
rect 535956 27542 536008 27548
rect 530436 12436 530488 12442
rect 530436 12378 530488 12384
rect 531540 12436 531592 12442
rect 531540 12378 531592 12384
rect 534576 12436 534628 12442
rect 534576 12378 534628 12384
rect 535036 12436 535088 12442
rect 535036 12378 535088 12384
rect 525560 11892 525612 11898
rect 525560 11834 525612 11840
rect 520868 7880 520920 7886
rect 520868 7822 520920 7828
rect 520776 7540 520828 7546
rect 520776 7482 520828 7488
rect 520682 7032 520738 7041
rect 520682 6967 520738 6976
rect 520696 6905 520724 6967
rect 520682 6896 520738 6905
rect 520682 6831 520738 6840
rect 519578 4720 519634 4729
rect 519578 4655 519634 4664
rect 519592 480 519620 4655
rect 520880 1442 520908 7822
rect 524364 7812 524416 7818
rect 524364 7754 524416 7760
rect 521972 7540 522024 7546
rect 521972 7482 522024 7488
rect 520788 1414 520908 1442
rect 520788 480 520816 1414
rect 521984 480 522012 7482
rect 523168 4208 523220 4214
rect 523168 4150 523220 4156
rect 523180 480 523208 4150
rect 524376 480 524404 7754
rect 525572 480 525600 11834
rect 529148 9716 529200 9722
rect 529148 9658 529200 9664
rect 529160 9602 529188 9658
rect 529160 9574 529280 9602
rect 527952 7744 528004 7750
rect 527952 7686 528004 7692
rect 526756 4820 526808 4826
rect 526756 4762 526808 4768
rect 526768 480 526796 4762
rect 527964 480 527992 7686
rect 529252 610 529280 9574
rect 530344 4480 530396 4486
rect 530344 4422 530396 4428
rect 529148 604 529200 610
rect 529148 546 529200 552
rect 529240 604 529292 610
rect 529240 546 529292 552
rect 529160 480 529188 546
rect 530356 480 530384 4422
rect 531552 480 531580 12378
rect 532736 11824 532788 11830
rect 532736 11766 532788 11772
rect 532748 480 532776 11766
rect 534666 7168 534722 7177
rect 534496 7126 534666 7154
rect 534496 7041 534524 7126
rect 534666 7103 534722 7112
rect 534482 7032 534538 7041
rect 534482 6967 534538 6976
rect 533932 4548 533984 4554
rect 533932 4490 533984 4496
rect 533944 480 533972 4490
rect 535048 480 535076 12378
rect 536232 9716 536284 9722
rect 536232 9658 536284 9664
rect 536244 480 536272 9658
rect 537348 7546 537376 294578
rect 541488 19310 541516 327694
rect 541566 320512 541622 320521
rect 541566 320447 541622 320456
rect 541580 320346 541608 320447
rect 541568 320340 541620 320346
rect 541568 320282 541620 320288
rect 544328 320340 544380 320346
rect 544328 320282 544380 320288
rect 544340 320249 544368 320282
rect 544326 320240 544382 320249
rect 544326 320175 544382 320184
rect 546996 304292 547048 304298
rect 546996 304234 547048 304240
rect 545616 291848 545668 291854
rect 545616 291790 545668 291796
rect 542856 268388 542908 268394
rect 542856 268330 542908 268336
rect 541476 19304 541528 19310
rect 541476 19246 541528 19252
rect 542868 12442 542896 268330
rect 545628 14498 545656 291790
rect 545536 14470 545656 14498
rect 542856 12436 542908 12442
rect 542856 12378 542908 12384
rect 543408 12436 543460 12442
rect 543408 12378 543460 12384
rect 539820 11756 539872 11762
rect 539820 11698 539872 11704
rect 537336 7540 537388 7546
rect 537336 7482 537388 7488
rect 538624 7540 538676 7546
rect 538624 7482 538676 7488
rect 537428 4276 537480 4282
rect 537428 4218 537480 4224
rect 537440 480 537468 4218
rect 538636 480 538664 7482
rect 539832 480 539860 11698
rect 542212 9716 542264 9722
rect 542212 9658 542264 9664
rect 541016 4616 541068 4622
rect 541016 4558 541068 4564
rect 541028 480 541056 4558
rect 542224 480 542252 9658
rect 543420 480 543448 12378
rect 545536 9722 545564 14470
rect 545524 9716 545576 9722
rect 545524 9658 545576 9664
rect 545800 9716 545852 9722
rect 545800 9658 545852 9664
rect 544604 4752 544656 4758
rect 544604 4694 544656 4700
rect 544616 480 544644 4694
rect 545812 480 545840 9658
rect 546902 7440 546958 7449
rect 546902 7375 546958 7384
rect 546916 7041 546944 7375
rect 546902 7032 546958 7041
rect 546902 6967 546958 6976
rect 547008 480 547036 304234
rect 548388 12442 548416 334630
rect 575976 333260 576028 333266
rect 575976 333202 576028 333208
rect 553896 324964 553948 324970
rect 553896 324906 553948 324912
rect 552516 322244 552568 322250
rect 552516 322186 552568 322192
rect 552528 309126 552556 322186
rect 553908 309346 553936 324906
rect 560796 319456 560848 319462
rect 560796 319398 560848 319404
rect 555276 309800 555328 309806
rect 555276 309742 555328 309748
rect 553816 309318 553936 309346
rect 553816 309210 553844 309318
rect 553816 309182 553936 309210
rect 552516 309120 552568 309126
rect 552516 309062 552568 309068
rect 552608 309120 552660 309126
rect 552608 309062 552660 309068
rect 552620 299554 552648 309062
rect 552528 299526 552648 299554
rect 552528 293298 552556 299526
rect 553908 299470 553936 309182
rect 553804 299464 553856 299470
rect 553804 299406 553856 299412
rect 553896 299464 553948 299470
rect 553896 299406 553948 299412
rect 552436 293270 552556 293298
rect 552436 288425 552464 293270
rect 553816 289898 553844 299406
rect 553816 289870 553936 289898
rect 553908 289746 553936 289870
rect 553896 289740 553948 289746
rect 553896 289682 553948 289688
rect 552422 288416 552478 288425
rect 552422 288351 552478 288360
rect 552606 288416 552662 288425
rect 552606 288351 552662 288360
rect 552528 278798 552556 278829
rect 552620 278798 552648 288351
rect 553896 280288 553948 280294
rect 553896 280230 553948 280236
rect 552516 278792 552568 278798
rect 552608 278792 552660 278798
rect 552606 278760 552608 278769
rect 552660 278760 552662 278769
rect 552568 278740 552606 278746
rect 552516 278734 552606 278740
rect 552528 278718 552606 278734
rect 552606 278695 552662 278704
rect 552790 278760 552846 278769
rect 552790 278695 552846 278704
rect 552804 269142 552832 278695
rect 553908 270722 553936 280230
rect 553816 270694 553936 270722
rect 553816 270586 553844 270694
rect 553816 270558 553936 270586
rect 553908 270502 553936 270558
rect 553896 270496 553948 270502
rect 553896 270438 553948 270444
rect 552608 269136 552660 269142
rect 552608 269078 552660 269084
rect 552792 269136 552844 269142
rect 552792 269078 552844 269084
rect 549756 265668 549808 265674
rect 549756 265610 549808 265616
rect 549768 12442 549796 265610
rect 552620 260930 552648 269078
rect 552528 260902 552648 260930
rect 553896 260976 553948 260982
rect 553896 260918 553948 260924
rect 552528 259457 552556 260902
rect 553908 260846 553936 260918
rect 553896 260840 553948 260846
rect 553896 260782 553948 260788
rect 553804 260772 553856 260778
rect 553804 260714 553856 260720
rect 552514 259448 552570 259457
rect 552514 259383 552570 259392
rect 552698 259448 552754 259457
rect 552698 259383 552754 259392
rect 552712 241641 552740 259383
rect 553816 251274 553844 260714
rect 553816 251246 553936 251274
rect 553908 251190 553936 251246
rect 553896 251184 553948 251190
rect 553896 251126 553948 251132
rect 553896 241664 553948 241670
rect 552514 241632 552570 241641
rect 552514 241567 552570 241576
rect 552698 241632 552754 241641
rect 553896 241606 553948 241612
rect 552698 241567 552754 241576
rect 552528 240122 552556 241567
rect 552436 240094 552556 240122
rect 552436 230518 552464 240094
rect 553908 231849 553936 241606
rect 553710 231840 553766 231849
rect 553710 231775 553766 231784
rect 553894 231840 553950 231849
rect 553894 231775 553950 231784
rect 552332 230512 552384 230518
rect 552332 230454 552384 230460
rect 552424 230512 552476 230518
rect 552424 230454 552476 230460
rect 552344 211206 552372 230454
rect 553724 222222 553752 231775
rect 553712 222216 553764 222222
rect 553710 222184 553712 222193
rect 553896 222216 553948 222222
rect 553764 222184 553766 222193
rect 553710 222119 553766 222128
rect 553894 222184 553896 222193
rect 553948 222184 553950 222193
rect 553894 222119 553950 222128
rect 553724 212566 553752 222119
rect 553712 212560 553764 212566
rect 553712 212502 553764 212508
rect 553896 212560 553948 212566
rect 553896 212502 553948 212508
rect 552332 211200 552384 211206
rect 552332 211142 552384 211148
rect 552516 211200 552568 211206
rect 552516 211142 552568 211148
rect 552528 201657 552556 211142
rect 553908 202881 553936 212502
rect 553710 202872 553766 202881
rect 553710 202807 553766 202816
rect 553894 202872 553950 202881
rect 553894 202807 553950 202816
rect 552514 201648 552570 201657
rect 552514 201583 552570 201592
rect 552422 201512 552478 201521
rect 552422 201447 552424 201456
rect 552476 201447 552478 201456
rect 552424 201418 552476 201424
rect 552424 196308 552476 196314
rect 552424 196250 552476 196256
rect 552436 191826 552464 196250
rect 553724 193254 553752 202807
rect 553712 193248 553764 193254
rect 553710 193216 553712 193225
rect 553896 193248 553948 193254
rect 553764 193216 553766 193225
rect 553710 193151 553766 193160
rect 553894 193216 553896 193225
rect 553948 193216 553950 193225
rect 553894 193151 553950 193160
rect 552424 191820 552476 191826
rect 552424 191762 552476 191768
rect 553724 183598 553752 193151
rect 553712 183592 553764 183598
rect 553896 183592 553948 183598
rect 553712 183534 553764 183540
rect 553894 183560 553896 183569
rect 553948 183560 553950 183569
rect 552424 183524 552476 183530
rect 553894 183495 553950 183504
rect 552424 183466 552476 183472
rect 552436 182186 552464 183466
rect 552344 182158 552464 182186
rect 552344 172553 552372 182158
rect 553894 174040 553950 174049
rect 553894 173975 553950 173984
rect 553908 173913 553936 173975
rect 553710 173904 553766 173913
rect 553710 173839 553766 173848
rect 553894 173904 553950 173913
rect 553894 173839 553950 173848
rect 552330 172544 552386 172553
rect 552330 172479 552386 172488
rect 552698 172544 552754 172553
rect 552698 172479 552754 172488
rect 552712 164422 552740 172479
rect 552516 164416 552568 164422
rect 552516 164358 552568 164364
rect 552700 164416 552752 164422
rect 552700 164358 552752 164364
rect 552528 162858 552556 164358
rect 553724 164234 553752 173839
rect 553724 164218 553936 164234
rect 553724 164212 553948 164218
rect 553724 164206 553896 164212
rect 553896 164154 553948 164160
rect 552516 162852 552568 162858
rect 552516 162794 552568 162800
rect 553896 154692 553948 154698
rect 553896 154634 553948 154640
rect 552516 153264 552568 153270
rect 552516 153206 552568 153212
rect 552528 143546 552556 153206
rect 553908 144906 553936 154634
rect 553896 144900 553948 144906
rect 553896 144842 553948 144848
rect 552516 143540 552568 143546
rect 552516 143482 552568 143488
rect 553896 135380 553948 135386
rect 553896 135322 553948 135328
rect 553908 135250 553936 135322
rect 553712 135244 553764 135250
rect 553712 135186 553764 135192
rect 553896 135244 553948 135250
rect 553896 135186 553948 135192
rect 552240 133952 552292 133958
rect 552240 133894 552292 133900
rect 552252 133754 552280 133894
rect 552240 133748 552292 133754
rect 552240 133690 552292 133696
rect 553724 125633 553752 135186
rect 553710 125624 553766 125633
rect 553710 125559 553766 125568
rect 553894 125624 553950 125633
rect 553894 125559 553950 125568
rect 552516 125452 552568 125458
rect 552516 125394 552568 125400
rect 552528 114510 552556 125394
rect 553908 122806 553936 125559
rect 553436 122800 553488 122806
rect 553436 122742 553488 122748
rect 553896 122800 553948 122806
rect 553896 122742 553948 122748
rect 552516 114504 552568 114510
rect 552516 114446 552568 114452
rect 552608 114504 552660 114510
rect 552608 114446 552660 114452
rect 552620 104961 552648 114446
rect 553448 113257 553476 122742
rect 553434 113248 553490 113257
rect 553434 113183 553490 113192
rect 553618 113248 553674 113257
rect 553618 113183 553674 113192
rect 553632 109750 553660 113183
rect 553620 109744 553672 109750
rect 553620 109686 553672 109692
rect 552422 104952 552478 104961
rect 552422 104887 552478 104896
rect 552606 104952 552662 104961
rect 552606 104887 552662 104896
rect 552436 103494 552464 104887
rect 552424 103488 552476 103494
rect 552424 103430 552476 103436
rect 553896 96756 553948 96762
rect 553896 96698 553948 96704
rect 553908 96626 553936 96698
rect 553712 96620 553764 96626
rect 553712 96562 553764 96568
rect 553896 96620 553948 96626
rect 553896 96562 553948 96568
rect 552424 93900 552476 93906
rect 552424 93842 552476 93848
rect 552436 87174 552464 93842
rect 552424 87168 552476 87174
rect 553724 87145 553752 96562
rect 552424 87110 552476 87116
rect 553710 87136 553766 87145
rect 553710 87071 553766 87080
rect 553894 87000 553950 87009
rect 553894 86935 553950 86944
rect 552424 86896 552476 86902
rect 552424 86838 552476 86844
rect 552436 85542 552464 86838
rect 552424 85536 552476 85542
rect 552424 85478 552476 85484
rect 553908 77194 553936 86935
rect 552332 77172 552384 77178
rect 553908 77166 554028 77194
rect 552332 77114 552384 77120
rect 552344 67697 552372 77114
rect 552330 67688 552386 67697
rect 552330 67623 552386 67632
rect 552514 67688 552570 67697
rect 554000 67658 554028 77166
rect 552514 67623 552570 67632
rect 553896 67652 553948 67658
rect 552528 66230 552556 67623
rect 553896 67594 553948 67600
rect 553988 67652 554040 67658
rect 553988 67594 554040 67600
rect 552516 66224 552568 66230
rect 552516 66166 552568 66172
rect 553908 58070 553936 67594
rect 553896 58064 553948 58070
rect 553896 58006 553948 58012
rect 553988 57928 554040 57934
rect 553988 57870 554040 57876
rect 552516 56704 552568 56710
rect 552516 56646 552568 56652
rect 554000 56658 554028 57870
rect 552528 46918 552556 56646
rect 554000 56630 554120 56658
rect 554092 48385 554120 56630
rect 553894 48376 553950 48385
rect 553894 48311 553950 48320
rect 554078 48376 554134 48385
rect 554078 48311 554134 48320
rect 553908 48278 553936 48311
rect 553804 48272 553856 48278
rect 553804 48214 553856 48220
rect 553896 48272 553948 48278
rect 553896 48214 553948 48220
rect 553816 46918 553844 48214
rect 552516 46912 552568 46918
rect 552516 46854 552568 46860
rect 553804 46912 553856 46918
rect 553804 46854 553856 46860
rect 553804 38412 553856 38418
rect 553804 38354 553856 38360
rect 552608 37324 552660 37330
rect 552608 37266 552660 37272
rect 552620 29050 552648 37266
rect 552528 29022 552648 29050
rect 553816 29034 553844 38354
rect 553804 29028 553856 29034
rect 552528 27606 552556 29022
rect 553804 28970 553856 28976
rect 553896 29028 553948 29034
rect 553896 28970 553948 28976
rect 552516 27600 552568 27606
rect 552516 27542 552568 27548
rect 553908 22930 553936 28970
rect 553908 22902 554120 22930
rect 548376 12436 548428 12442
rect 548376 12378 548428 12384
rect 549388 12436 549440 12442
rect 549388 12378 549440 12384
rect 549756 12436 549808 12442
rect 549756 12378 549808 12384
rect 550584 12436 550636 12442
rect 550584 12378 550636 12384
rect 548192 5364 548244 5370
rect 548192 5306 548244 5312
rect 548204 480 548232 5306
rect 549400 480 549428 12378
rect 550596 480 550624 12378
rect 552884 9716 552936 9722
rect 552884 9658 552936 9664
rect 551688 5296 551740 5302
rect 551688 5238 551740 5244
rect 551700 480 551728 5238
rect 552896 480 552924 9658
rect 554092 480 554120 22902
rect 555288 7546 555316 309742
rect 556656 262880 556708 262886
rect 556656 262822 556708 262828
rect 556668 12442 556696 262822
rect 560808 164506 560836 319398
rect 563556 301504 563608 301510
rect 563556 301446 563608 301452
rect 560808 164478 560928 164506
rect 560900 164234 560928 164478
rect 560808 164206 560928 164234
rect 560808 87281 560836 164206
rect 560794 87272 560850 87281
rect 560794 87207 560850 87216
rect 560794 87136 560850 87145
rect 560794 87071 560850 87080
rect 560808 48657 560836 87071
rect 560794 48648 560850 48657
rect 560794 48583 560850 48592
rect 560794 48512 560850 48521
rect 560794 48447 560850 48456
rect 560808 19310 560836 48447
rect 560796 19304 560848 19310
rect 560796 19246 560848 19252
rect 556656 12436 556708 12442
rect 556656 12378 556708 12384
rect 557668 12436 557720 12442
rect 557668 12378 557720 12384
rect 555276 7540 555328 7546
rect 555276 7482 555328 7488
rect 556472 7540 556524 7546
rect 556472 7482 556524 7488
rect 555276 5228 555328 5234
rect 555276 5170 555328 5176
rect 555288 480 555316 5170
rect 556484 480 556512 7482
rect 557680 480 557708 12378
rect 561256 9716 561308 9722
rect 561256 9658 561308 9664
rect 560060 9444 560112 9450
rect 560060 9386 560112 9392
rect 558034 7168 558090 7177
rect 558034 7103 558090 7112
rect 558048 7002 558076 7103
rect 558036 6996 558088 7002
rect 558036 6938 558088 6944
rect 558864 5160 558916 5166
rect 558864 5102 558916 5108
rect 558876 480 558904 5102
rect 560072 480 560100 9386
rect 561268 480 561296 9658
rect 563568 7546 563596 301446
rect 567696 300144 567748 300150
rect 567696 300086 567748 300092
rect 567708 12442 567736 300086
rect 571836 286340 571888 286346
rect 571836 286282 571888 286288
rect 571848 278769 571876 286282
rect 571834 278760 571890 278769
rect 571834 278695 571890 278704
rect 572018 278760 572074 278769
rect 572018 278695 572074 278704
rect 572032 269142 572060 278695
rect 571836 269136 571888 269142
rect 571836 269078 571888 269084
rect 572020 269136 572072 269142
rect 572020 269078 572072 269084
rect 571848 259457 571876 269078
rect 574596 261520 574648 261526
rect 574596 261462 574648 261468
rect 571834 259448 571890 259457
rect 571834 259383 571890 259392
rect 572018 259448 572074 259457
rect 572018 259383 572074 259392
rect 572032 249830 572060 259383
rect 571836 249824 571888 249830
rect 571836 249766 571888 249772
rect 572020 249824 572072 249830
rect 572020 249766 572072 249772
rect 571848 240145 571876 249766
rect 571834 240136 571890 240145
rect 571834 240071 571890 240080
rect 572018 240136 572074 240145
rect 572018 240071 572074 240080
rect 572032 230518 572060 240071
rect 571836 230512 571888 230518
rect 571836 230454 571888 230460
rect 572020 230512 572072 230518
rect 572020 230454 572072 230460
rect 571848 220833 571876 230454
rect 571834 220824 571890 220833
rect 571834 220759 571890 220768
rect 572018 220824 572074 220833
rect 572018 220759 572074 220768
rect 572032 211206 572060 220759
rect 571836 211200 571888 211206
rect 571836 211142 571888 211148
rect 572020 211200 572072 211206
rect 572020 211142 572072 211148
rect 571848 201482 571876 211142
rect 571836 201476 571888 201482
rect 571836 201418 571888 201424
rect 572020 201476 572072 201482
rect 572020 201418 572072 201424
rect 572032 191865 572060 201418
rect 571834 191856 571890 191865
rect 571834 191791 571890 191800
rect 572018 191856 572074 191865
rect 572018 191791 572074 191800
rect 571848 182170 571876 191791
rect 571836 182164 571888 182170
rect 571836 182106 571888 182112
rect 572020 182164 572072 182170
rect 572020 182106 572072 182112
rect 572032 172553 572060 182106
rect 571834 172544 571890 172553
rect 571834 172479 571890 172488
rect 572018 172544 572074 172553
rect 572018 172479 572074 172488
rect 570362 164656 570418 164665
rect 570362 164591 570418 164600
rect 570376 164257 570404 164591
rect 571848 164529 571876 172479
rect 571834 164520 571890 164529
rect 571834 164455 571890 164464
rect 571560 164416 571612 164422
rect 571560 164358 571612 164364
rect 572112 164416 572164 164422
rect 572112 164358 572164 164364
rect 571572 164257 571600 164358
rect 572124 164257 572152 164358
rect 570362 164248 570418 164257
rect 570362 164183 570418 164192
rect 571558 164248 571614 164257
rect 571558 164183 571614 164192
rect 571834 164248 571890 164257
rect 571834 164183 571890 164192
rect 572110 164248 572166 164257
rect 572110 164183 572166 164192
rect 571848 162858 571876 164183
rect 571836 162852 571888 162858
rect 571836 162794 571888 162800
rect 571836 153264 571888 153270
rect 571836 153206 571888 153212
rect 571848 143546 571876 153206
rect 571836 143540 571888 143546
rect 571836 143482 571888 143488
rect 571836 133952 571888 133958
rect 571836 133894 571888 133900
rect 571848 124166 571876 133894
rect 571836 124160 571888 124166
rect 571836 124102 571888 124108
rect 571836 114572 571888 114578
rect 571836 114514 571888 114520
rect 571848 104854 571876 114514
rect 571836 104848 571888 104854
rect 571836 104790 571888 104796
rect 571836 95328 571888 95334
rect 571836 95270 571888 95276
rect 571848 85542 571876 95270
rect 571836 85536 571888 85542
rect 571836 85478 571888 85484
rect 571836 75948 571888 75954
rect 571836 75890 571888 75896
rect 571848 66230 571876 75890
rect 571836 66224 571888 66230
rect 571836 66166 571888 66172
rect 571836 56704 571888 56710
rect 571836 56646 571888 56652
rect 571848 46918 571876 56646
rect 571836 46912 571888 46918
rect 571836 46854 571888 46860
rect 571836 37324 571888 37330
rect 571836 37266 571888 37272
rect 571848 27606 571876 37266
rect 571836 27600 571888 27606
rect 571836 27542 571888 27548
rect 574608 12442 574636 261462
rect 575988 12442 576016 333202
rect 579380 312588 579432 312594
rect 579380 312530 579432 312536
rect 578000 283620 578052 283626
rect 578000 283562 578052 283568
rect 567696 12436 567748 12442
rect 567696 12378 567748 12384
rect 568340 12436 568392 12442
rect 568340 12378 568392 12384
rect 574596 12436 574648 12442
rect 574596 12378 574648 12384
rect 575516 12436 575568 12442
rect 575516 12378 575568 12384
rect 575976 12436 576028 12442
rect 575976 12378 576028 12384
rect 576712 12436 576764 12442
rect 576712 12378 576764 12384
rect 563648 9376 563700 9382
rect 563648 9318 563700 9324
rect 563556 7540 563608 7546
rect 563556 7482 563608 7488
rect 562452 5092 562504 5098
rect 562452 5034 562504 5040
rect 562464 480 562492 5034
rect 563660 480 563688 9318
rect 567236 9172 567288 9178
rect 567236 9114 567288 9120
rect 564844 7540 564896 7546
rect 564844 7482 564896 7488
rect 564856 480 564884 7482
rect 566040 5024 566092 5030
rect 566040 4966 566092 4972
rect 566052 480 566080 4966
rect 567248 480 567276 9114
rect 567602 7032 567658 7041
rect 567602 6967 567604 6976
rect 567656 6967 567658 6976
rect 567604 6938 567656 6944
rect 568352 480 568380 12378
rect 571928 9716 571980 9722
rect 571928 9658 571980 9664
rect 570732 9104 570784 9110
rect 570732 9046 570784 9052
rect 569076 7200 569128 7206
rect 569076 7142 569128 7148
rect 569088 7041 569116 7142
rect 569074 7032 569130 7041
rect 569074 6967 569130 6976
rect 569536 4752 569588 4758
rect 569536 4694 569588 4700
rect 569548 480 569576 4694
rect 570744 480 570772 9046
rect 571940 480 571968 9658
rect 574320 9036 574372 9042
rect 574320 8978 574372 8984
rect 573122 4856 573178 4865
rect 573122 4791 573178 4800
rect 573136 480 573164 4791
rect 574332 480 574360 8978
rect 575528 480 575556 12378
rect 576724 480 576752 12378
rect 577908 8968 577960 8974
rect 577908 8910 577960 8916
rect 577920 480 577948 8910
rect 578012 4146 578040 283562
rect 578644 7200 578696 7206
rect 578642 7168 578644 7177
rect 578696 7168 578698 7177
rect 578642 7103 578698 7112
rect 579392 4146 579420 312530
rect 580668 289808 580720 289814
rect 580668 289750 580720 289756
rect 580680 289377 580708 289750
rect 580666 289368 580722 289377
rect 580666 289303 580722 289312
rect 580668 274644 580720 274650
rect 580668 274586 580720 274592
rect 580680 273737 580708 274586
rect 580666 273728 580722 273737
rect 580666 273663 580722 273672
rect 580668 195968 580720 195974
rect 580668 195910 580720 195916
rect 580680 195537 580708 195910
rect 580666 195528 580722 195537
rect 580666 195463 580722 195472
rect 580392 148980 580444 148986
rect 580392 148922 580444 148928
rect 580404 148617 580432 148922
rect 580390 148608 580446 148617
rect 580390 148543 580446 148552
rect 580668 86964 580720 86970
rect 580668 86906 580720 86912
rect 580680 86057 580708 86906
rect 580666 86048 580722 86057
rect 580666 85983 580722 85992
rect 580772 54777 580800 458186
rect 581496 253224 581548 253230
rect 581496 253166 581548 253172
rect 580758 54768 580814 54777
rect 580758 54703 580814 54712
rect 581508 7546 581536 253166
rect 581586 8936 581642 8945
rect 581586 8871 581642 8880
rect 581496 7540 581548 7546
rect 581496 7482 581548 7488
rect 578000 4140 578052 4146
rect 578000 4082 578052 4088
rect 579104 4140 579156 4146
rect 579104 4082 579156 4088
rect 579380 4140 579432 4146
rect 579380 4082 579432 4088
rect 580300 4140 580352 4146
rect 580300 4082 580352 4088
rect 579116 480 579144 4082
rect 580312 480 580340 4082
rect 581600 1442 581628 8871
rect 583886 7848 583942 7857
rect 583886 7783 583942 7792
rect 582692 7540 582744 7546
rect 582692 7482 582744 7488
rect 581508 1414 581628 1442
rect 581508 480 581536 1414
rect 582704 480 582732 7482
rect 583900 7177 583928 7783
rect 583886 7168 583942 7177
rect 583886 7103 583942 7112
rect 1066 0 1122 480
rect 2170 0 2226 480
rect 3366 0 3422 480
rect 4562 0 4618 480
rect 5758 0 5814 480
rect 6954 0 7010 480
rect 8150 0 8206 480
rect 9346 0 9402 480
rect 10542 0 10598 480
rect 11738 0 11794 480
rect 12934 0 12990 480
rect 14130 0 14186 480
rect 15326 0 15382 480
rect 16522 0 16578 480
rect 17718 0 17774 480
rect 18822 0 18878 480
rect 20018 0 20074 480
rect 21214 0 21270 480
rect 22410 0 22466 480
rect 23606 0 23662 480
rect 24802 0 24858 480
rect 25998 0 26054 480
rect 27194 0 27250 480
rect 28390 0 28446 480
rect 29586 0 29642 480
rect 30782 0 30838 480
rect 31978 0 32034 480
rect 33174 0 33230 480
rect 34370 0 34426 480
rect 35474 0 35530 480
rect 36670 0 36726 480
rect 37866 0 37922 480
rect 39062 0 39118 480
rect 40258 0 40314 480
rect 41454 0 41510 480
rect 42650 0 42706 480
rect 43846 0 43902 480
rect 45042 0 45098 480
rect 46238 0 46294 480
rect 47434 0 47490 480
rect 48630 0 48686 480
rect 49826 0 49882 480
rect 51022 0 51078 480
rect 52126 0 52182 480
rect 53322 0 53378 480
rect 54518 0 54574 480
rect 55714 0 55770 480
rect 56910 0 56966 480
rect 58106 0 58162 480
rect 59302 0 59358 480
rect 60498 0 60554 480
rect 61694 0 61750 480
rect 62890 0 62946 480
rect 64086 0 64142 480
rect 65282 0 65338 480
rect 66478 0 66534 480
rect 67674 0 67730 480
rect 68778 0 68834 480
rect 69974 0 70030 480
rect 71170 0 71226 480
rect 72366 0 72422 480
rect 73562 0 73618 480
rect 74758 0 74814 480
rect 75954 0 76010 480
rect 77150 0 77206 480
rect 78346 0 78402 480
rect 79542 0 79598 480
rect 80738 0 80794 480
rect 81934 0 81990 480
rect 83130 0 83186 480
rect 84326 0 84382 480
rect 85430 0 85486 480
rect 86626 0 86682 480
rect 87822 0 87878 480
rect 89018 0 89074 480
rect 90214 0 90270 480
rect 91410 0 91466 480
rect 92606 0 92662 480
rect 93802 0 93858 480
rect 94998 0 95054 480
rect 96194 0 96250 480
rect 97390 0 97446 480
rect 98586 0 98642 480
rect 99782 0 99838 480
rect 100978 0 101034 480
rect 102082 0 102138 480
rect 103278 0 103334 480
rect 104474 0 104530 480
rect 105670 0 105726 480
rect 106866 0 106922 480
rect 108062 0 108118 480
rect 109258 0 109314 480
rect 110454 0 110510 480
rect 111650 0 111706 480
rect 112846 0 112902 480
rect 114042 0 114098 480
rect 115238 0 115294 480
rect 116434 0 116490 480
rect 117630 0 117686 480
rect 118734 0 118790 480
rect 119930 0 119986 480
rect 121126 0 121182 480
rect 122322 0 122378 480
rect 123518 0 123574 480
rect 124714 0 124770 480
rect 125910 0 125966 480
rect 127106 0 127162 480
rect 128302 0 128358 480
rect 129498 0 129554 480
rect 130694 0 130750 480
rect 131890 0 131946 480
rect 133086 0 133142 480
rect 134282 0 134338 480
rect 135386 0 135442 480
rect 136582 0 136638 480
rect 137778 0 137834 480
rect 138974 0 139030 480
rect 140170 0 140226 480
rect 141366 0 141422 480
rect 142562 0 142618 480
rect 143758 0 143814 480
rect 144954 0 145010 480
rect 146150 0 146206 480
rect 147346 0 147402 480
rect 148542 0 148598 480
rect 149738 0 149794 480
rect 150934 0 150990 480
rect 152038 0 152094 480
rect 153234 0 153290 480
rect 154430 0 154486 480
rect 155626 0 155682 480
rect 156822 0 156878 480
rect 158018 0 158074 480
rect 159214 0 159270 480
rect 160410 0 160466 480
rect 161606 0 161662 480
rect 162802 0 162858 480
rect 163998 0 164054 480
rect 165194 0 165250 480
rect 166390 0 166446 480
rect 167586 0 167642 480
rect 168690 0 168746 480
rect 169886 0 169942 480
rect 171082 0 171138 480
rect 172278 0 172334 480
rect 173474 0 173530 480
rect 174670 0 174726 480
rect 175866 0 175922 480
rect 177062 0 177118 480
rect 178258 0 178314 480
rect 179454 0 179510 480
rect 180650 0 180706 480
rect 181846 0 181902 480
rect 183042 0 183098 480
rect 184238 0 184294 480
rect 185342 0 185398 480
rect 186538 0 186594 480
rect 187734 0 187790 480
rect 188930 0 188986 480
rect 190126 0 190182 480
rect 191322 0 191378 480
rect 192518 0 192574 480
rect 193714 0 193770 480
rect 194910 0 194966 480
rect 196106 0 196162 480
rect 197302 0 197358 480
rect 198498 0 198554 480
rect 199694 0 199750 480
rect 200890 0 200946 480
rect 201994 0 202050 480
rect 203190 0 203246 480
rect 204386 0 204442 480
rect 205582 0 205638 480
rect 206778 0 206834 480
rect 207974 0 208030 480
rect 209170 0 209226 480
rect 210366 0 210422 480
rect 211562 0 211618 480
rect 212758 0 212814 480
rect 213954 0 214010 480
rect 215150 0 215206 480
rect 216346 0 216402 480
rect 217542 0 217598 480
rect 218646 0 218702 480
rect 219842 0 219898 480
rect 221038 0 221094 480
rect 222234 0 222290 480
rect 223430 0 223486 480
rect 224626 0 224682 480
rect 225822 0 225878 480
rect 227018 0 227074 480
rect 228214 0 228270 480
rect 229410 0 229466 480
rect 230606 0 230662 480
rect 231802 0 231858 480
rect 232998 0 233054 480
rect 234194 0 234250 480
rect 235298 0 235354 480
rect 236494 0 236550 480
rect 237690 0 237746 480
rect 238886 0 238942 480
rect 240082 0 240138 480
rect 241278 0 241334 480
rect 242474 0 242530 480
rect 243670 0 243726 480
rect 244866 0 244922 480
rect 246062 0 246118 480
rect 247258 0 247314 480
rect 248454 0 248510 480
rect 249650 0 249706 480
rect 250846 0 250902 480
rect 251950 0 252006 480
rect 253146 0 253202 480
rect 254342 0 254398 480
rect 255538 0 255594 480
rect 256734 0 256790 480
rect 257930 0 257986 480
rect 259126 0 259182 480
rect 260322 0 260378 480
rect 261518 0 261574 480
rect 262714 0 262770 480
rect 263910 0 263966 480
rect 265106 0 265162 480
rect 266302 0 266358 480
rect 267498 0 267554 480
rect 268602 0 268658 480
rect 269798 0 269854 480
rect 270994 0 271050 480
rect 272190 0 272246 480
rect 273386 0 273442 480
rect 274582 0 274638 480
rect 275778 0 275834 480
rect 276974 0 277030 480
rect 278170 0 278226 480
rect 279366 0 279422 480
rect 280562 0 280618 480
rect 281758 0 281814 480
rect 282954 0 283010 480
rect 284150 0 284206 480
rect 285254 0 285310 480
rect 286450 0 286506 480
rect 287646 0 287702 480
rect 288842 0 288898 480
rect 290038 0 290094 480
rect 291234 0 291290 480
rect 292430 0 292486 480
rect 293626 0 293682 480
rect 294822 0 294878 480
rect 296018 0 296074 480
rect 297214 0 297270 480
rect 298410 0 298466 480
rect 299606 0 299662 480
rect 300802 0 300858 480
rect 301906 0 301962 480
rect 303102 0 303158 480
rect 304298 0 304354 480
rect 305494 0 305550 480
rect 306690 0 306746 480
rect 307886 0 307942 480
rect 309082 0 309138 480
rect 310278 0 310334 480
rect 311474 0 311530 480
rect 312670 0 312726 480
rect 313866 0 313922 480
rect 315062 0 315118 480
rect 316258 0 316314 480
rect 317454 0 317510 480
rect 318558 0 318614 480
rect 319754 0 319810 480
rect 320950 0 321006 480
rect 322146 0 322202 480
rect 323342 0 323398 480
rect 324538 0 324594 480
rect 325734 0 325790 480
rect 326930 0 326986 480
rect 328126 0 328182 480
rect 329322 0 329378 480
rect 330518 0 330574 480
rect 331714 0 331770 480
rect 332910 0 332966 480
rect 334106 0 334162 480
rect 335210 0 335266 480
rect 336406 0 336462 480
rect 337602 0 337658 480
rect 338798 0 338854 480
rect 339994 0 340050 480
rect 341190 0 341246 480
rect 342386 0 342442 480
rect 343582 0 343638 480
rect 344778 0 344834 480
rect 345974 0 346030 480
rect 347170 0 347226 480
rect 348366 0 348422 480
rect 349562 0 349618 480
rect 350758 0 350814 480
rect 351862 0 351918 480
rect 353058 0 353114 480
rect 354254 0 354310 480
rect 355450 0 355506 480
rect 356646 0 356702 480
rect 357842 0 357898 480
rect 359038 0 359094 480
rect 360234 0 360290 480
rect 361430 0 361486 480
rect 362626 0 362682 480
rect 363822 0 363878 480
rect 365018 0 365074 480
rect 366214 0 366270 480
rect 367410 0 367466 480
rect 368514 0 368570 480
rect 369710 0 369766 480
rect 370906 0 370962 480
rect 372102 0 372158 480
rect 373298 0 373354 480
rect 374494 0 374550 480
rect 375690 0 375746 480
rect 376886 0 376942 480
rect 378082 0 378138 480
rect 379278 0 379334 480
rect 380474 0 380530 480
rect 381670 0 381726 480
rect 382866 0 382922 480
rect 384062 0 384118 480
rect 385166 0 385222 480
rect 386362 0 386418 480
rect 387558 0 387614 480
rect 388754 0 388810 480
rect 389950 0 390006 480
rect 391146 0 391202 480
rect 392342 0 392398 480
rect 393538 0 393594 480
rect 394734 0 394790 480
rect 395930 0 395986 480
rect 397126 0 397182 480
rect 398322 0 398378 480
rect 399518 0 399574 480
rect 400714 0 400770 480
rect 401818 0 401874 480
rect 403014 0 403070 480
rect 404210 0 404266 480
rect 405406 0 405462 480
rect 406602 0 406658 480
rect 407798 0 407854 480
rect 408994 0 409050 480
rect 410190 0 410246 480
rect 411386 0 411442 480
rect 412582 0 412638 480
rect 413778 0 413834 480
rect 414974 0 415030 480
rect 416170 0 416226 480
rect 417366 0 417422 480
rect 418470 0 418526 480
rect 419666 0 419722 480
rect 420862 0 420918 480
rect 422058 0 422114 480
rect 423254 0 423310 480
rect 424450 0 424506 480
rect 425646 0 425702 480
rect 426842 0 426898 480
rect 428038 0 428094 480
rect 429234 0 429290 480
rect 430430 0 430486 480
rect 431626 0 431682 480
rect 432822 0 432878 480
rect 434018 0 434074 480
rect 435122 0 435178 480
rect 436318 0 436374 480
rect 437514 0 437570 480
rect 438710 0 438766 480
rect 439906 0 439962 480
rect 441102 0 441158 480
rect 442298 0 442354 480
rect 443494 0 443550 480
rect 444690 0 444746 480
rect 445886 0 445942 480
rect 447082 0 447138 480
rect 448278 0 448334 480
rect 449474 0 449530 480
rect 450670 0 450726 480
rect 451774 0 451830 480
rect 452970 0 453026 480
rect 454166 0 454222 480
rect 455362 0 455418 480
rect 456558 0 456614 480
rect 457754 0 457810 480
rect 458950 0 459006 480
rect 460146 0 460202 480
rect 461342 0 461398 480
rect 462538 0 462594 480
rect 463734 0 463790 480
rect 464930 0 464986 480
rect 466126 0 466182 480
rect 467322 0 467378 480
rect 468426 0 468482 480
rect 469622 0 469678 480
rect 470818 0 470874 480
rect 472014 0 472070 480
rect 473210 0 473266 480
rect 474406 0 474462 480
rect 475602 0 475658 480
rect 476798 0 476854 480
rect 477994 0 478050 480
rect 479190 0 479246 480
rect 480386 0 480442 480
rect 481582 0 481638 480
rect 482778 0 482834 480
rect 483974 0 484030 480
rect 485078 0 485134 480
rect 486274 0 486330 480
rect 487470 0 487526 480
rect 488666 0 488722 480
rect 489862 0 489918 480
rect 491058 0 491114 480
rect 492254 0 492310 480
rect 493450 0 493506 480
rect 494646 0 494702 480
rect 495842 0 495898 480
rect 497038 0 497094 480
rect 498234 0 498290 480
rect 499430 0 499486 480
rect 500626 0 500682 480
rect 501730 0 501786 480
rect 502926 0 502982 480
rect 504122 0 504178 480
rect 505318 0 505374 480
rect 506514 0 506570 480
rect 507710 0 507766 480
rect 508906 0 508962 480
rect 510102 0 510158 480
rect 511298 0 511354 480
rect 512494 0 512550 480
rect 513690 0 513746 480
rect 514886 0 514942 480
rect 516082 0 516138 480
rect 517278 0 517334 480
rect 518382 0 518438 480
rect 519578 0 519634 480
rect 520774 0 520830 480
rect 521970 0 522026 480
rect 523166 0 523222 480
rect 524362 0 524418 480
rect 525558 0 525614 480
rect 526754 0 526810 480
rect 527950 0 528006 480
rect 529146 0 529202 480
rect 530342 0 530398 480
rect 531538 0 531594 480
rect 532734 0 532790 480
rect 533930 0 533986 480
rect 535034 0 535090 480
rect 536230 0 536286 480
rect 537426 0 537482 480
rect 538622 0 538678 480
rect 539818 0 539874 480
rect 541014 0 541070 480
rect 542210 0 542266 480
rect 543406 0 543462 480
rect 544602 0 544658 480
rect 545798 0 545854 480
rect 546994 0 547050 480
rect 548190 0 548246 480
rect 549386 0 549442 480
rect 550582 0 550638 480
rect 551686 0 551742 480
rect 552882 0 552938 480
rect 554078 0 554134 480
rect 555274 0 555330 480
rect 556470 0 556526 480
rect 557666 0 557722 480
rect 558862 0 558918 480
rect 560058 0 560114 480
rect 561254 0 561310 480
rect 562450 0 562506 480
rect 563646 0 563702 480
rect 564842 0 564898 480
rect 566038 0 566094 480
rect 567234 0 567290 480
rect 568338 0 568394 480
rect 569534 0 569590 480
rect 570730 0 570786 480
rect 571926 0 571982 480
rect 573122 0 573178 480
rect 574318 0 574374 480
rect 575514 0 575570 480
rect 576710 0 576766 480
rect 577906 0 577962 480
rect 579102 0 579158 480
rect 580298 0 580354 480
rect 581494 0 581550 480
rect 582690 0 582746 480
rect 583886 0 583942 480
<< via2 >>
rect 11278 700304 11334 700360
rect 3734 695408 3790 695464
rect 3918 678680 3974 678736
rect 3918 661952 3974 662008
rect 3550 645224 3606 645280
rect 3918 628360 3974 628416
rect 3826 611632 3882 611688
rect 3918 594904 3974 594960
rect 3734 578176 3790 578232
rect 3918 561312 3974 561368
rect 3642 544584 3698 544640
rect 3642 527856 3698 527912
rect 4010 511128 4066 511184
rect 3734 494264 3790 494320
rect 3918 477556 3974 477592
rect 3918 477536 3920 477556
rect 3920 477536 3972 477556
rect 3972 477536 3974 477556
rect 3918 462440 3974 462496
rect 3642 460808 3698 460864
rect 3642 444116 3644 444136
rect 3644 444116 3696 444136
rect 3696 444116 3698 444136
rect 3642 444080 3698 444116
rect 3642 427216 3698 427272
rect 3826 410488 3882 410544
rect 3826 393760 3882 393816
rect 3550 377032 3606 377088
rect 3826 360304 3882 360360
rect 3826 343440 3882 343496
rect 3642 309984 3698 310040
rect 3550 293256 3606 293312
rect 3826 259664 3882 259720
rect 3826 242936 3882 242992
rect 3734 209344 3790 209400
rect 3826 192652 3828 192672
rect 3828 192652 3880 192672
rect 3880 192652 3882 192672
rect 3826 192616 3882 192652
rect 5942 337320 5998 337376
rect 4378 326712 4434 326768
rect 4286 276392 4342 276448
rect 4194 226208 4250 226264
rect 4102 175888 4158 175944
rect 4010 159160 4066 159216
rect 4010 142296 4066 142352
rect 4010 126928 4066 126984
rect 4010 125568 4066 125624
rect 3918 108840 3974 108896
rect 3642 58520 3698 58576
rect 3918 42744 3974 42800
rect 3918 41792 3974 41848
rect 3918 25064 3974 25120
rect 3918 9560 3974 9616
rect 3918 8336 3974 8392
rect 6954 3304 7010 3360
rect 16522 3576 16578 3632
rect 15326 3440 15382 3496
rect 25998 3848 26054 3904
rect 24802 3712 24858 3768
rect 30690 10240 30746 10296
rect 31978 3984 32034 4040
rect 48630 6160 48686 6216
rect 58198 3440 58254 3496
rect 58382 3440 58438 3496
rect 58198 3304 58254 3360
rect 58382 3304 58438 3360
rect 128854 337864 128910 337920
rect 119286 337728 119342 337784
rect 94354 337456 94410 337512
rect 103922 337456 103978 337512
rect 91318 231784 91374 231840
rect 91502 231784 91558 231840
rect 91318 212472 91374 212528
rect 91502 212472 91558 212528
rect 91318 193160 91374 193216
rect 91502 193160 91558 193216
rect 91502 173848 91558 173904
rect 91502 164192 91558 164248
rect 91502 154400 91558 154456
rect 91778 154400 91834 154456
rect 91502 144880 91558 144936
rect 91778 144880 91834 144936
rect 91318 125704 91374 125760
rect 91502 125568 91558 125624
rect 91318 87080 91374 87136
rect 91502 86944 91558 87000
rect 99690 3168 99746 3224
rect 103830 3168 103886 3224
rect 128578 337592 128634 337648
rect 123886 337456 123942 337512
rect 120482 10512 120538 10568
rect 123518 10548 123520 10568
rect 123520 10548 123572 10568
rect 123572 10548 123574 10568
rect 123518 10512 123574 10548
rect 113858 3168 113914 3224
rect 129038 337728 129094 337784
rect 128946 337592 129002 337648
rect 138422 337864 138478 337920
rect 142654 337728 142710 337784
rect 152222 337728 152278 337784
rect 161974 337728 162030 337784
rect 171542 337728 171598 337784
rect 128762 337456 128818 337512
rect 129222 337592 129278 337648
rect 138330 337628 138332 337648
rect 138332 337628 138384 337648
rect 138384 337628 138386 337648
rect 138330 337592 138386 337628
rect 142286 337456 142342 337512
rect 142470 337456 142526 337512
rect 142746 337456 142802 337512
rect 152130 337456 152186 337512
rect 152406 337456 152462 337512
rect 152590 337456 152646 337512
rect 161606 337456 161662 337512
rect 161790 337456 161846 337512
rect 162066 337456 162122 337512
rect 171450 337456 171506 337512
rect 171726 337456 171782 337512
rect 171910 337456 171966 337512
rect 138330 337184 138386 337240
rect 142562 337184 142618 337240
rect 152314 337184 152370 337240
rect 161882 337184 161938 337240
rect 171634 337184 171690 337240
rect 126094 3168 126150 3224
rect 135478 298016 135534 298072
rect 135662 298016 135718 298072
rect 135478 278704 135534 278760
rect 135662 278704 135718 278760
rect 135478 259392 135534 259448
rect 135662 259392 135718 259448
rect 135478 240080 135534 240136
rect 135662 240080 135718 240136
rect 135478 220768 135534 220824
rect 135662 220768 135718 220824
rect 135478 211112 135534 211168
rect 135662 211112 135718 211168
rect 135478 191800 135534 191856
rect 135662 191800 135718 191856
rect 135478 172488 135534 172544
rect 135662 172488 135718 172544
rect 135662 164464 135718 164520
rect 135570 164328 135626 164384
rect 135662 48592 135718 48648
rect 135662 48456 135718 48512
rect 135294 9696 135350 9752
rect 135478 9696 135534 9752
rect 138238 10124 138294 10160
rect 138238 10104 138240 10124
rect 138240 10104 138292 10124
rect 138292 10104 138294 10124
rect 138606 10140 138608 10160
rect 138608 10140 138660 10160
rect 138660 10140 138662 10160
rect 138606 10104 138662 10140
rect 147806 10512 147862 10568
rect 148450 10512 148506 10568
rect 152038 298016 152094 298072
rect 152222 298016 152278 298072
rect 152038 278704 152094 278760
rect 152222 278704 152278 278760
rect 152038 259392 152094 259448
rect 152222 259392 152278 259448
rect 152038 240080 152094 240136
rect 152222 240080 152278 240136
rect 152038 220768 152094 220824
rect 152222 220768 152278 220824
rect 152038 211112 152094 211168
rect 152222 211112 152278 211168
rect 152038 191800 152094 191856
rect 152222 191800 152278 191856
rect 152038 172488 152094 172544
rect 152222 172488 152278 172544
rect 151854 9696 151910 9752
rect 152038 9696 152094 9752
rect 148174 3304 148230 3360
rect 148082 3032 148138 3088
rect 157834 10376 157890 10432
rect 157466 10140 157468 10160
rect 157468 10140 157520 10160
rect 157520 10140 157522 10160
rect 157466 10104 157522 10140
rect 157834 10104 157890 10160
rect 157558 9968 157614 10024
rect 157650 3168 157706 3224
rect 158110 3168 158166 3224
rect 170162 298016 170218 298072
rect 170346 298016 170402 298072
rect 170162 278704 170218 278760
rect 170346 278704 170402 278760
rect 170162 259392 170218 259448
rect 170346 259392 170402 259448
rect 170162 240080 170218 240136
rect 170346 240080 170402 240136
rect 170162 220768 170218 220824
rect 170346 220768 170402 220824
rect 170162 211112 170218 211168
rect 170346 211112 170402 211168
rect 170162 191800 170218 191856
rect 170346 191800 170402 191856
rect 170162 172488 170218 172544
rect 170346 172488 170402 172544
rect 167862 10376 167918 10432
rect 167770 10124 167826 10160
rect 167770 10104 167772 10124
rect 167772 10104 167824 10124
rect 167824 10104 167826 10124
rect 167494 9968 167550 10024
rect 169702 9696 169758 9752
rect 169886 9696 169942 9752
rect 169518 9424 169574 9480
rect 170162 9424 170218 9480
rect 181294 337728 181350 337784
rect 190862 337728 190918 337784
rect 200614 337728 200670 337784
rect 210182 337728 210238 337784
rect 180926 337456 180982 337512
rect 181110 337456 181166 337512
rect 181386 337456 181442 337512
rect 190770 337456 190826 337512
rect 191046 337456 191102 337512
rect 191230 337456 191286 337512
rect 200246 337456 200302 337512
rect 200430 337456 200486 337512
rect 200706 337456 200762 337512
rect 210090 337456 210146 337512
rect 210366 337456 210422 337512
rect 210550 337456 210606 337512
rect 181202 337184 181258 337240
rect 190954 337184 191010 337240
rect 200522 337184 200578 337240
rect 210274 337184 210330 337240
rect 177246 10512 177302 10568
rect 186538 3168 186594 3224
rect 190678 298016 190734 298072
rect 190862 298016 190918 298072
rect 190678 278704 190734 278760
rect 190862 278704 190918 278760
rect 190678 259392 190734 259448
rect 190862 259392 190918 259448
rect 190678 240080 190734 240136
rect 190862 240080 190918 240136
rect 190678 220768 190734 220824
rect 190862 220768 190918 220824
rect 190678 211112 190734 211168
rect 190862 211112 190918 211168
rect 190678 191800 190734 191856
rect 190862 191800 190918 191856
rect 190678 172488 190734 172544
rect 190862 172488 190918 172544
rect 190218 17992 190274 18048
rect 190402 17992 190458 18048
rect 186814 10684 186816 10704
rect 186816 10684 186868 10704
rect 186868 10684 186870 10704
rect 186814 10648 186870 10684
rect 187090 10512 187146 10568
rect 191782 10104 191838 10160
rect 190402 9696 190458 9752
rect 190586 9696 190642 9752
rect 187734 4800 187790 4856
rect 187182 3188 187238 3224
rect 187182 3168 187184 3188
rect 187184 3168 187236 3188
rect 187236 3168 187238 3188
rect 196382 10648 196438 10704
rect 196474 10376 196530 10432
rect 195922 10140 195924 10160
rect 195924 10140 195976 10160
rect 195976 10140 195978 10160
rect 195922 10104 195978 10140
rect 196474 10104 196530 10160
rect 196014 9968 196070 10024
rect 196290 7828 196292 7848
rect 196292 7828 196344 7848
rect 196344 7828 196346 7848
rect 196290 7792 196346 7828
rect 193622 7692 193624 7712
rect 193624 7692 193676 7712
rect 193676 7692 193678 7712
rect 193622 7656 193678 7692
rect 196198 3188 196254 3224
rect 196198 3168 196200 3188
rect 196200 3168 196252 3188
rect 196252 3168 196254 3188
rect 195922 2932 195924 2952
rect 195924 2932 195976 2952
rect 195976 2932 195978 2952
rect 195922 2896 195978 2932
rect 196750 3188 196806 3224
rect 196750 3168 196752 3188
rect 196752 3168 196804 3188
rect 196804 3168 196806 3188
rect 214322 298016 214378 298072
rect 214506 298016 214562 298072
rect 214322 278704 214378 278760
rect 214506 278704 214562 278760
rect 214322 259392 214378 259448
rect 214506 259392 214562 259448
rect 214322 240080 214378 240136
rect 214506 240080 214562 240136
rect 214322 220768 214378 220824
rect 214506 220768 214562 220824
rect 214322 211112 214378 211168
rect 214506 211112 214562 211168
rect 214322 191800 214378 191856
rect 214506 191800 214562 191856
rect 214322 172488 214378 172544
rect 214506 172488 214562 172544
rect 206318 10376 206374 10432
rect 206318 10104 206374 10160
rect 215794 9968 215850 10024
rect 216162 10376 216218 10432
rect 216162 10104 216218 10160
rect 215978 9832 216034 9888
rect 213954 9696 214010 9752
rect 214506 9696 214562 9752
rect 206778 5888 206834 5944
rect 205858 3188 205914 3224
rect 205858 3168 205860 3188
rect 205860 3168 205912 3188
rect 205912 3168 205914 3188
rect 206226 3168 206282 3224
rect 207698 2896 207754 2952
rect 210366 5752 210422 5808
rect 208158 3304 208214 3360
rect 208158 2488 208214 2544
rect 210274 3032 210330 3088
rect 215794 7928 215850 7984
rect 215886 7656 215942 7712
rect 215794 6024 215850 6080
rect 215886 5888 215942 5944
rect 216346 4256 216402 4312
rect 215794 4120 215850 4176
rect 219934 337728 219990 337784
rect 219566 337456 219622 337512
rect 219750 337456 219806 337512
rect 220026 337456 220082 337512
rect 219842 337184 219898 337240
rect 219658 4664 219714 4720
rect 218646 4276 218702 4312
rect 218646 4256 218648 4276
rect 218648 4256 218700 4276
rect 218700 4256 218702 4276
rect 219750 4120 219806 4176
rect 226926 337592 226982 337648
rect 225362 212472 225418 212528
rect 225546 212472 225602 212528
rect 225362 173848 225418 173904
rect 225362 164192 225418 164248
rect 283598 463120 283654 463176
rect 282310 462984 282366 463040
rect 283414 462984 283470 463040
rect 288198 463140 288254 463176
rect 288198 463120 288200 463140
rect 288200 463120 288252 463140
rect 288252 463120 288254 463140
rect 288382 463120 288438 463176
rect 293166 463120 293222 463176
rect 304114 700304 304170 700360
rect 580114 695952 580170 696008
rect 580114 680348 580116 680368
rect 580116 680348 580168 680368
rect 580168 680348 580170 680368
rect 580114 680312 580170 680348
rect 580114 664672 580170 664728
rect 313774 618160 313830 618216
rect 314050 618160 314106 618216
rect 580114 649032 580170 649088
rect 443770 618160 443826 618216
rect 580114 633428 580116 633448
rect 580116 633428 580168 633448
rect 580168 633428 580170 633448
rect 580114 633392 580170 633428
rect 443678 608640 443734 608696
rect 580114 617752 580170 617808
rect 573398 608640 573454 608696
rect 573766 608640 573822 608696
rect 580114 602112 580170 602168
rect 580114 586508 580116 586528
rect 580116 586508 580168 586528
rect 580168 586508 580170 586528
rect 580114 586472 580170 586508
rect 313774 557504 313830 557560
rect 313774 518880 313830 518936
rect 580114 570832 580170 570888
rect 378726 560224 378782 560280
rect 378910 560224 378966 560280
rect 314050 557504 314106 557560
rect 508446 560224 508502 560280
rect 508630 560224 508686 560280
rect 580114 555192 580170 555248
rect 314050 518880 314106 518936
rect 580114 539552 580170 539608
rect 379002 529760 379058 529816
rect 508722 529760 508778 529816
rect 379186 520240 379242 520296
rect 508906 520240 508962 520296
rect 580114 523912 580170 523968
rect 443494 511944 443550 512000
rect 443678 511944 443734 512000
rect 573214 511944 573270 512000
rect 573398 511944 573454 512000
rect 580114 508272 580170 508328
rect 378542 502288 378598 502344
rect 378818 502324 378820 502344
rect 378820 502324 378872 502344
rect 378872 502324 378874 502344
rect 378818 502288 378874 502324
rect 378542 492632 378598 492688
rect 378726 492632 378782 492688
rect 508262 502288 508318 502344
rect 508538 502324 508540 502344
rect 508540 502324 508592 502344
rect 508592 502324 508594 502344
rect 508538 502288 508594 502324
rect 508262 492632 508318 492688
rect 508446 492632 508502 492688
rect 580114 492668 580116 492688
rect 580116 492668 580168 492688
rect 580168 492668 580170 492688
rect 580114 492632 580170 492668
rect 580114 476992 580170 477048
rect 342386 462440 342442 462496
rect 225178 48320 225234 48376
rect 225362 48320 225418 48376
rect 225454 10648 225510 10704
rect 225638 10376 225694 10432
rect 225638 9968 225694 10024
rect 225086 9696 225142 9752
rect 225270 9696 225326 9752
rect 229410 8880 229466 8936
rect 225822 8744 225878 8800
rect 224626 7928 224682 7984
rect 225270 7928 225326 7984
rect 225454 7928 225510 7984
rect 224534 3168 224590 3224
rect 225270 7656 225326 7712
rect 225546 7656 225602 7712
rect 225362 7520 225418 7576
rect 225454 6432 225510 6488
rect 225178 6296 225234 6352
rect 225454 5888 225510 5944
rect 225270 5752 225326 5808
rect 225270 5208 225326 5264
rect 225270 4664 225326 4720
rect 225454 4256 225510 4312
rect 225638 3168 225694 3224
rect 225178 3032 225234 3088
rect 226926 5208 226982 5264
rect 228122 3576 228178 3632
rect 232170 459584 232226 459640
rect 233182 459584 233238 459640
rect 236218 459584 236274 459640
rect 237414 459584 237470 459640
rect 238518 459584 238574 459640
rect 239622 459584 239678 459640
rect 241646 459584 241702 459640
rect 242750 459584 242806 459640
rect 244590 459584 244646 459640
rect 245878 459584 245934 459640
rect 246982 459584 247038 459640
rect 248822 459584 248878 459640
rect 251214 459584 251270 459640
rect 252134 459584 252190 459640
rect 343122 459584 343178 459640
rect 344226 459584 344282 459640
rect 346250 459584 346306 459640
rect 347354 459584 347410 459640
rect 348458 459584 348514 459640
rect 229594 7112 229650 7168
rect 229778 135224 229834 135280
rect 229962 135224 230018 135280
rect 231434 337320 231490 337376
rect 231342 7828 231344 7848
rect 231344 7828 231396 7848
rect 231396 7828 231398 7848
rect 231342 7792 231398 7828
rect 231526 6024 231582 6080
rect 232814 337748 232870 337784
rect 232814 337728 232816 337748
rect 232816 337728 232868 337748
rect 232868 337728 232870 337748
rect 232446 9968 232502 10024
rect 231894 9696 231950 9752
rect 232170 9696 232226 9752
rect 231618 5344 231674 5400
rect 231066 5208 231122 5264
rect 232446 7384 232502 7440
rect 232354 7112 232410 7168
rect 230146 4120 230202 4176
rect 230422 3576 230478 3632
rect 232906 3440 232962 3496
rect 232722 3304 232778 3360
rect 235390 278704 235446 278760
rect 235574 278704 235630 278760
rect 235574 244296 235630 244352
rect 235482 241576 235538 241632
rect 235666 221040 235722 221096
rect 235574 220904 235630 220960
rect 235390 220768 235446 220824
rect 235574 220768 235630 220824
rect 235574 182144 235630 182200
rect 235758 182144 235814 182200
rect 235574 154400 235630 154456
rect 235850 154400 235906 154456
rect 235482 144880 235538 144936
rect 235850 144880 235906 144936
rect 235574 125568 235630 125624
rect 235758 125568 235814 125624
rect 235390 48184 235446 48240
rect 235666 48048 235722 48104
rect 235022 10648 235078 10704
rect 234654 10512 234710 10568
rect 235022 10124 235078 10160
rect 235022 10104 235024 10124
rect 235024 10104 235076 10124
rect 235076 10104 235078 10124
rect 234930 8880 234986 8936
rect 235022 8744 235078 8800
rect 234010 7928 234066 7984
rect 235114 6568 235170 6624
rect 235390 10512 235446 10568
rect 234930 4120 234986 4176
rect 235114 4140 235170 4176
rect 235114 4120 235116 4140
rect 235116 4120 235168 4140
rect 235168 4120 235170 4140
rect 235206 3848 235262 3904
rect 235206 3576 235262 3632
rect 235114 3440 235170 3496
rect 234838 3304 234894 3360
rect 234746 3168 234802 3224
rect 235206 3168 235262 3224
rect 235666 4256 235722 4312
rect 236586 10240 236642 10296
rect 235574 3712 235630 3768
rect 235390 3304 235446 3360
rect 236954 3984 237010 4040
rect 236770 3576 236826 3632
rect 237782 9152 237838 9208
rect 237690 5208 237746 5264
rect 237138 3440 237194 3496
rect 239254 96600 239310 96656
rect 239254 51060 239310 51096
rect 239254 51040 239256 51060
rect 239256 51040 239308 51060
rect 239308 51040 239310 51060
rect 238058 4140 238114 4176
rect 238058 4120 238060 4140
rect 238060 4120 238112 4140
rect 238112 4120 238114 4140
rect 238518 10104 238574 10160
rect 239438 96600 239494 96656
rect 239438 51060 239494 51096
rect 239438 51040 239440 51060
rect 239440 51040 239492 51060
rect 239492 51040 239494 51060
rect 239438 6160 239494 6216
rect 240082 9288 240138 9344
rect 241002 6568 241058 6624
rect 240818 6296 240874 6352
rect 242198 318960 242254 319016
rect 242198 318824 242254 318880
rect 242014 153176 242070 153232
rect 242198 153176 242254 153232
rect 241830 134000 241886 134056
rect 242014 133864 242070 133920
rect 242198 133864 242254 133920
rect 241830 132776 241886 132832
rect 242198 125704 242254 125760
rect 242106 125568 242162 125624
rect 242198 106392 242254 106448
rect 242106 106256 242162 106312
rect 241922 9968 241978 10024
rect 242658 276120 242714 276176
rect 242750 275984 242806 276040
rect 242474 218048 242530 218104
rect 242842 218184 242898 218240
rect 242474 182144 242530 182200
rect 242658 164212 242714 164248
rect 242658 164192 242660 164212
rect 242660 164192 242712 164212
rect 242712 164192 242714 164212
rect 242842 164192 242898 164248
rect 242566 162968 242622 163024
rect 242474 157800 242530 157856
rect 242474 144880 242530 144936
rect 242474 96600 242530 96656
rect 242658 96600 242714 96656
rect 242750 77288 242806 77344
rect 242934 77288 242990 77344
rect 242566 17992 242622 18048
rect 242750 17992 242806 18048
rect 242198 6432 242254 6488
rect 244866 9324 244868 9344
rect 244868 9324 244920 9344
rect 244920 9324 244922 9344
rect 244866 9288 244922 9324
rect 244866 9172 244922 9208
rect 244866 9152 244868 9172
rect 244868 9152 244920 9172
rect 244920 9152 244922 9172
rect 244774 5480 244830 5536
rect 244866 5344 244922 5400
rect 244958 5228 245014 5264
rect 244958 5208 244960 5228
rect 244960 5208 245012 5228
rect 245012 5208 245014 5228
rect 246522 285776 246578 285832
rect 246614 285640 246670 285696
rect 246338 198736 246394 198792
rect 246430 198464 246486 198520
rect 246890 96736 246946 96792
rect 246798 96600 246854 96656
rect 251674 241748 251676 241768
rect 251676 241748 251728 241768
rect 251728 241748 251730 241768
rect 251674 241712 251730 241748
rect 251674 179560 251730 179616
rect 251766 132912 251822 132968
rect 251766 132640 251822 132696
rect 251674 100852 251676 100872
rect 251676 100852 251728 100872
rect 251728 100852 251730 100872
rect 251674 100816 251730 100852
rect 254158 320492 254160 320512
rect 254160 320492 254212 320512
rect 254212 320492 254214 320512
rect 254158 320456 254214 320492
rect 254250 9172 254306 9208
rect 254250 9152 254252 9172
rect 254252 9152 254304 9172
rect 254304 9152 254306 9172
rect 254526 9172 254582 9208
rect 254526 9152 254528 9172
rect 254528 9152 254580 9172
rect 254580 9152 254582 9172
rect 254434 8880 254490 8936
rect 254894 8880 254950 8936
rect 255078 7520 255134 7576
rect 255078 7112 255134 7168
rect 259862 179288 259918 179344
rect 261242 320320 261298 320376
rect 261150 241984 261206 242040
rect 261150 179696 261206 179752
rect 261150 179288 261206 179344
rect 261150 101088 261206 101144
rect 261058 38700 261060 38720
rect 261060 38700 261112 38720
rect 261112 38700 261114 38720
rect 261058 38664 261114 38700
rect 259954 7112 260010 7168
rect 259954 6704 260010 6760
rect 257746 5480 257802 5536
rect 257286 5344 257342 5400
rect 268142 38700 268144 38720
rect 268144 38700 268196 38720
rect 268196 38700 268198 38720
rect 268142 38664 268198 38700
rect 268510 191800 268566 191856
rect 268694 191800 268750 191856
rect 268510 183504 268566 183560
rect 268694 183504 268750 183560
rect 269522 6976 269578 7032
rect 269522 6704 269578 6760
rect 268694 4800 268750 4856
rect 264370 4548 264426 4584
rect 270902 226616 270958 226672
rect 270902 226208 270958 226264
rect 264370 4528 264372 4548
rect 264372 4528 264424 4548
rect 264424 4528 264426 4548
rect 269798 4548 269854 4584
rect 269798 4528 269800 4548
rect 269800 4528 269852 4548
rect 269852 4528 269854 4548
rect 271362 108976 271418 109032
rect 271638 108976 271694 109032
rect 264186 4428 264188 4448
rect 264188 4428 264240 4448
rect 264240 4428 264242 4448
rect 264186 4392 264242 4428
rect 273294 336912 273350 336968
rect 273294 336776 273350 336832
rect 272926 333920 272982 333976
rect 273294 333920 273350 333976
rect 273018 295296 273074 295352
rect 273202 295296 273258 295352
rect 272926 274760 272982 274816
rect 272834 274644 272890 274680
rect 272834 274624 272836 274644
rect 272836 274624 272888 274644
rect 272888 274624 272890 274644
rect 272834 264968 272890 265024
rect 273018 264968 273074 265024
rect 272926 52400 272982 52456
rect 273294 52400 273350 52456
rect 273018 33224 273074 33280
rect 273202 33224 273258 33280
rect 272926 4392 272982 4448
rect 275502 324264 275558 324320
rect 275686 324300 275688 324320
rect 275688 324300 275740 324320
rect 275740 324300 275742 324320
rect 275686 324264 275742 324300
rect 275594 187856 275650 187912
rect 275686 187720 275742 187776
rect 275502 118632 275558 118688
rect 275686 118632 275742 118688
rect 276514 295296 276570 295352
rect 276698 295316 276754 295352
rect 276698 295296 276700 295316
rect 276700 295296 276752 295316
rect 276752 295296 276754 295316
rect 276974 295296 277030 295352
rect 276790 227840 276846 227896
rect 276790 227704 276846 227760
rect 276514 221448 276570 221504
rect 276514 208392 276570 208448
rect 276974 227704 277030 227760
rect 276698 164464 276754 164520
rect 276790 164328 276846 164384
rect 276698 133864 276754 133920
rect 276422 62056 276478 62112
rect 276606 62056 276662 62112
rect 276882 133864 276938 133920
rect 277250 295432 277306 295488
rect 277250 227704 277306 227760
rect 278446 277480 278502 277536
rect 278446 277344 278502 277400
rect 278446 16496 278502 16552
rect 278722 306312 278778 306368
rect 278906 306312 278962 306368
rect 278630 277480 278686 277536
rect 278630 277344 278686 277400
rect 278814 267688 278870 267744
rect 278998 267688 279054 267744
rect 278814 162968 278870 163024
rect 278722 162832 278778 162888
rect 278630 16496 278686 16552
rect 279458 249736 279514 249792
rect 279734 278704 279790 278760
rect 279826 249736 279882 249792
rect 279826 100680 279882 100736
rect 280010 278704 280066 278760
rect 280010 100716 280012 100736
rect 280012 100716 280064 100736
rect 280064 100716 280066 100736
rect 280010 100680 280066 100716
rect 279734 64912 279790 64968
rect 280010 64912 280066 64968
rect 284794 164192 284850 164248
rect 285254 177248 285310 177304
rect 285162 164464 285218 164520
rect 285162 164328 285218 164384
rect 285346 164056 285402 164112
rect 285622 164192 285678 164248
rect 285070 28872 285126 28928
rect 285254 28872 285310 28928
rect 285070 19216 285126 19272
rect 285346 19216 285402 19272
rect 290314 320220 290316 320240
rect 290316 320220 290368 320240
rect 290368 320220 290370 320240
rect 290314 320184 290370 320220
rect 289946 241712 290002 241768
rect 290038 241576 290094 241632
rect 290314 241612 290316 241632
rect 290316 241612 290368 241632
rect 290368 241612 290370 241632
rect 290314 241576 290370 241612
rect 290314 132812 290316 132832
rect 290316 132812 290368 132832
rect 290368 132812 290370 132832
rect 290314 132776 290370 132812
rect 290222 101088 290278 101144
rect 290406 101088 290462 101144
rect 293626 179968 293682 180024
rect 293626 179696 293682 179752
rect 293258 132640 293314 132696
rect 294638 320456 294694 320512
rect 294822 241848 294878 241904
rect 298594 38820 298650 38856
rect 298594 38800 298596 38820
rect 298596 38800 298648 38820
rect 298648 38800 298650 38820
rect 300434 226636 300490 226672
rect 300434 226616 300436 226636
rect 300436 226616 300488 226636
rect 300488 226616 300490 226636
rect 304942 230424 304998 230480
rect 305126 230424 305182 230480
rect 304850 173848 304906 173904
rect 305126 173848 305182 173904
rect 307886 86944 307942 87000
rect 308162 226480 308218 226536
rect 309174 151680 309230 151736
rect 309174 142160 309230 142216
rect 308162 86944 308218 87000
rect 308162 38664 308218 38720
rect 308898 86944 308954 87000
rect 309082 86944 309138 87000
rect 302550 4800 302606 4856
rect 302550 4548 302606 4584
rect 302550 4528 302552 4548
rect 302552 4528 302604 4548
rect 302604 4528 302606 4548
rect 302458 4392 302514 4448
rect 302826 4936 302882 4992
rect 303102 4548 303158 4584
rect 303102 4528 303104 4548
rect 303104 4528 303156 4548
rect 303156 4528 303158 4548
rect 303010 4428 303012 4448
rect 303012 4428 303064 4448
rect 303064 4428 303066 4448
rect 303010 4392 303066 4428
rect 309634 242392 309690 242448
rect 309634 241712 309690 241768
rect 309634 227160 309690 227216
rect 309634 226480 309690 226536
rect 312210 4936 312266 4992
rect 312578 5244 312580 5264
rect 312580 5244 312632 5264
rect 312632 5244 312634 5264
rect 312578 5208 312634 5244
rect 317454 5208 317510 5264
rect 318650 335688 318706 335744
rect 319110 335688 319166 335744
rect 319018 318688 319074 318744
rect 318926 318416 318982 318472
rect 318926 6432 318982 6488
rect 318834 6332 318836 6352
rect 318836 6332 318888 6352
rect 318888 6332 318890 6352
rect 318834 6296 318890 6332
rect 320122 282920 320178 282976
rect 320030 278840 320086 278896
rect 320030 251096 320086 251152
rect 320030 241576 320086 241632
rect 320030 216008 320086 216064
rect 320030 206216 320086 206272
rect 319754 172488 319810 172544
rect 319938 172488 319994 172544
rect 319846 153176 319902 153232
rect 320030 153176 320086 153232
rect 319846 56480 319902 56536
rect 320122 56480 320178 56536
rect 320398 6160 320454 6216
rect 321962 6296 322018 6352
rect 321962 4664 322018 4720
rect 322238 6296 322294 6352
rect 322146 4664 322202 4720
rect 326010 3984 326066 4040
rect 327390 3848 327446 3904
rect 328218 288496 328274 288552
rect 328402 288496 328458 288552
rect 328218 266328 328274 266384
rect 328402 266328 328458 266384
rect 328218 115912 328274 115968
rect 328402 115912 328458 115968
rect 328494 95104 328550 95160
rect 328494 94968 328550 95024
rect 328218 77288 328274 77344
rect 328402 77288 328458 77344
rect 328402 58112 328458 58168
rect 328402 57976 328458 58032
rect 328402 9968 328458 10024
rect 328678 6432 328734 6488
rect 327482 3712 327538 3768
rect 328770 3576 328826 3632
rect 328862 3440 328918 3496
rect 329874 10512 329930 10568
rect 331070 241440 331126 241496
rect 331254 241440 331310 241496
rect 331070 222128 331126 222184
rect 331254 222128 331310 222184
rect 331070 202816 331126 202872
rect 331254 202816 331310 202872
rect 331070 183504 331126 183560
rect 331254 183504 331310 183560
rect 331070 154536 331126 154592
rect 331254 154536 331310 154592
rect 331070 135224 331126 135280
rect 331254 135224 331310 135280
rect 331070 115912 331126 115968
rect 331254 115912 331310 115968
rect 330978 100816 331034 100872
rect 330978 100544 331034 100600
rect 331070 96600 331126 96656
rect 331254 96600 331310 96656
rect 331070 77288 331126 77344
rect 331254 77288 331310 77344
rect 331254 10240 331310 10296
rect 331622 10512 331678 10568
rect 331622 10004 331624 10024
rect 331624 10004 331676 10024
rect 331676 10004 331678 10024
rect 331622 9968 331678 10004
rect 333370 338000 333426 338056
rect 333554 338000 333610 338056
rect 333738 320592 333794 320648
rect 333738 320184 333794 320240
rect 331714 6024 331770 6080
rect 329782 2896 329838 2952
rect 337234 39208 337290 39264
rect 337234 38936 337290 38992
rect 337234 6432 337290 6488
rect 338154 7384 338210 7440
rect 336682 3440 336738 3496
rect 338798 6432 338854 6488
rect 338522 3304 338578 3360
rect 338338 3168 338394 3224
rect 341098 290128 341154 290184
rect 341098 289856 341154 289912
rect 340914 270816 340970 270872
rect 341190 270544 341246 270600
rect 341190 173984 341246 174040
rect 341190 173848 341246 173904
rect 341098 164328 341154 164384
rect 341190 125568 341246 125624
rect 341190 115776 341246 115832
rect 341190 106256 341246 106312
rect 341190 86944 341246 87000
rect 340914 48320 340970 48376
rect 341098 48320 341154 48376
rect 340730 9696 340786 9752
rect 340914 9696 340970 9752
rect 340822 8200 340878 8256
rect 340730 8064 340786 8120
rect 341466 173984 341522 174040
rect 341374 173848 341430 173904
rect 341374 164328 341430 164384
rect 341374 125568 341430 125624
rect 341466 115776 341522 115832
rect 341466 106256 341522 106312
rect 341374 86944 341430 87000
rect 341466 10376 341522 10432
rect 341282 8236 341284 8256
rect 341284 8236 341336 8256
rect 341336 8236 341338 8256
rect 341282 8200 341338 8236
rect 341374 8084 341430 8120
rect 341374 8064 341376 8084
rect 341376 8064 341428 8084
rect 341428 8064 341430 8084
rect 341466 3476 341468 3496
rect 341468 3476 341520 3496
rect 341520 3476 341522 3496
rect 341466 3440 341522 3476
rect 343398 320184 343454 320240
rect 343398 319912 343454 319968
rect 343398 7404 343454 7440
rect 343398 7384 343400 7404
rect 343400 7384 343452 7404
rect 343452 7384 343454 7404
rect 345330 5208 345386 5264
rect 342662 4392 342718 4448
rect 345330 4528 345386 4584
rect 346894 9696 346950 9752
rect 347078 9696 347134 9752
rect 346250 3304 346306 3360
rect 346342 3168 346398 3224
rect 346250 2896 346306 2952
rect 346986 7404 347042 7440
rect 346986 7384 346988 7404
rect 346988 7384 347040 7404
rect 347040 7384 347042 7404
rect 346986 6432 347042 6488
rect 347998 9424 348054 9480
rect 348366 4800 348422 4856
rect 349286 9152 349342 9208
rect 349562 6296 349618 6352
rect 349194 4664 349250 4720
rect 350850 9444 350906 9480
rect 350850 9424 350852 9444
rect 350852 9424 350904 9444
rect 350904 9424 350906 9444
rect 351310 9696 351366 9752
rect 351586 9696 351642 9752
rect 351126 9152 351182 9208
rect 351218 9036 351274 9072
rect 351218 9016 351220 9036
rect 351220 9016 351272 9036
rect 351272 9016 351274 9036
rect 350942 8880 350998 8936
rect 351034 8356 351090 8392
rect 351034 8336 351036 8356
rect 351036 8336 351088 8356
rect 351088 8336 351090 8356
rect 350850 7792 350906 7848
rect 350666 7656 350722 7712
rect 350942 5208 350998 5264
rect 350850 5108 350852 5128
rect 350852 5108 350904 5128
rect 350904 5108 350906 5128
rect 350850 5072 350906 5108
rect 350666 4936 350722 4992
rect 350574 4800 350630 4856
rect 350942 4528 350998 4584
rect 350850 4392 350906 4448
rect 351126 3168 351182 3224
rect 356186 7656 356242 7712
rect 356462 7404 356518 7440
rect 356462 7384 356464 7404
rect 356464 7384 356516 7404
rect 356516 7384 356518 7404
rect 356462 6432 356518 6488
rect 355818 4800 355874 4856
rect 355818 4528 355874 4584
rect 355266 2932 355268 2952
rect 355268 2932 355320 2952
rect 355320 2932 355322 2952
rect 355266 2896 355322 2932
rect 580666 461352 580722 461408
rect 360602 320592 360658 320648
rect 360694 320320 360750 320376
rect 357934 231784 357990 231840
rect 358118 231784 358174 231840
rect 360602 226516 360604 226536
rect 360604 226516 360656 226536
rect 360656 226516 360658 226536
rect 360602 226480 360658 226516
rect 357934 193160 357990 193216
rect 358118 193160 358174 193216
rect 357934 173848 357990 173904
rect 357934 164328 357990 164384
rect 357934 154400 357990 154456
rect 358210 154400 358266 154456
rect 357934 144880 357990 144936
rect 358210 144880 358266 144936
rect 360418 100972 360474 101008
rect 360418 100952 360420 100972
rect 360420 100952 360472 100972
rect 360472 100952 360474 100972
rect 358210 87080 358266 87136
rect 357934 86944 357990 87000
rect 356646 9016 356702 9072
rect 360234 8336 360290 8392
rect 360510 3168 360566 3224
rect 360602 2896 360658 2952
rect 580666 445712 580722 445768
rect 580666 430072 580722 430128
rect 580666 414432 580722 414488
rect 580666 398792 580722 398848
rect 580666 383152 580722 383208
rect 580666 367512 580722 367568
rect 580666 351872 580722 351928
rect 361154 8356 361210 8392
rect 361154 8336 361156 8356
rect 361156 8336 361208 8356
rect 361208 8336 361210 8356
rect 361246 7792 361302 7848
rect 360786 3168 360842 3224
rect 362258 226516 362260 226536
rect 362260 226516 362312 226536
rect 362312 226516 362314 226536
rect 362258 226480 362314 226516
rect 363914 8336 363970 8392
rect 366122 179560 366178 179616
rect 366122 179288 366178 179344
rect 366122 100816 366178 100872
rect 366122 38800 366178 38856
rect 366122 38528 366178 38584
rect 364926 3440 364982 3496
rect 364742 2896 364798 2952
rect 364650 2796 364652 2816
rect 364652 2796 364704 2816
rect 364704 2796 364706 2816
rect 364650 2760 364706 2796
rect 366122 6976 366178 7032
rect 366122 6568 366178 6624
rect 365294 3304 365350 3360
rect 365754 2896 365810 2952
rect 365110 2796 365112 2816
rect 365112 2796 365164 2816
rect 365164 2796 365166 2816
rect 365110 2760 365166 2796
rect 372930 298152 372986 298208
rect 373114 298152 373170 298208
rect 372838 296656 372894 296712
rect 373022 296656 373078 296712
rect 371550 231784 371606 231840
rect 371734 231784 371790 231840
rect 373114 231784 373170 231840
rect 373298 231784 373354 231840
rect 370262 179560 370318 179616
rect 370446 179424 370502 179480
rect 373114 172488 373170 172544
rect 373298 172488 373354 172544
rect 373022 133864 373078 133920
rect 373298 133864 373354 133920
rect 373298 125704 373354 125760
rect 373114 125568 373170 125624
rect 371826 85448 371882 85504
rect 372010 85448 372066 85504
rect 370262 38800 370318 38856
rect 370446 38664 370502 38720
rect 370354 7656 370410 7712
rect 370446 6024 370502 6080
rect 370354 5888 370410 5944
rect 370906 5072 370962 5128
rect 370262 3476 370264 3496
rect 370264 3476 370316 3496
rect 370316 3476 370318 3496
rect 370262 3440 370318 3476
rect 370170 3168 370226 3224
rect 370630 3168 370686 3224
rect 370538 3032 370594 3088
rect 370998 4936 371054 4992
rect 375874 132540 375876 132560
rect 375876 132540 375928 132560
rect 375928 132540 375930 132560
rect 375874 132504 375930 132540
rect 377346 38700 377348 38720
rect 377348 38700 377400 38720
rect 377400 38700 377402 38720
rect 377346 38664 377402 38700
rect 375138 3440 375194 3496
rect 375138 2896 375194 2952
rect 376886 5888 376942 5944
rect 375782 3304 375838 3360
rect 375966 3304 376022 3360
rect 392250 336640 392306 336696
rect 392434 336640 392490 336696
rect 385534 319096 385590 319152
rect 385534 318824 385590 318880
rect 385534 298016 385590 298072
rect 385718 298016 385774 298072
rect 392434 298016 392490 298072
rect 392618 298016 392674 298072
rect 385534 278704 385590 278760
rect 385718 278704 385774 278760
rect 392434 278704 392490 278760
rect 392618 278704 392674 278760
rect 385534 259392 385590 259448
rect 385718 259392 385774 259448
rect 392434 259392 392490 259448
rect 392618 259392 392674 259448
rect 384062 242120 384118 242176
rect 384062 241848 384118 241904
rect 385534 240080 385590 240136
rect 385718 240080 385774 240136
rect 392434 240080 392490 240136
rect 392618 240080 392674 240136
rect 385534 220768 385590 220824
rect 385718 220768 385774 220824
rect 392434 220768 392490 220824
rect 392618 220768 392674 220824
rect 385534 191800 385590 191856
rect 385718 191800 385774 191856
rect 392434 191800 392490 191856
rect 392618 191800 392674 191856
rect 380106 179560 380162 179616
rect 379922 179424 379978 179480
rect 391698 179832 391754 179888
rect 391698 179424 391754 179480
rect 385534 172488 385590 172544
rect 385718 172488 385774 172544
rect 392434 172488 392490 172544
rect 392618 172488 392674 172544
rect 385534 164464 385590 164520
rect 392434 164464 392490 164520
rect 382038 164192 382094 164248
rect 385534 164192 385590 164248
rect 385810 164192 385866 164248
rect 391698 164192 391754 164248
rect 392434 164192 392490 164248
rect 392710 164192 392766 164248
rect 385442 132640 385498 132696
rect 390318 132912 390374 132968
rect 390318 132504 390374 132560
rect 386822 101360 386878 101416
rect 391698 101224 391754 101280
rect 386822 100952 386878 101008
rect 391698 100816 391754 100872
rect 382038 38800 382094 38856
rect 389582 38800 389638 38856
rect 389766 38664 389822 38720
rect 392526 29144 392582 29200
rect 392434 29008 392490 29064
rect 392342 17992 392398 18048
rect 392618 17992 392674 18048
rect 385994 9696 386050 9752
rect 386362 9696 386418 9752
rect 389858 6976 389914 7032
rect 389858 6568 389914 6624
rect 392434 3304 392490 3360
rect 392434 2896 392490 2952
rect 399242 132640 399298 132696
rect 399242 38836 399244 38856
rect 399244 38836 399296 38856
rect 399296 38836 399298 38856
rect 399242 38800 399298 38836
rect 399426 7656 399482 7712
rect 402002 3168 402058 3224
rect 402002 2896 402058 2952
rect 406142 132812 406144 132832
rect 406144 132812 406196 132832
rect 406196 132812 406198 132832
rect 406142 132776 406198 132812
rect 406142 38936 406198 38992
rect 406878 3168 406934 3224
rect 580390 336232 580446 336288
rect 425462 320456 425518 320512
rect 444782 320456 444838 320512
rect 418562 320340 418618 320376
rect 418562 320320 418564 320340
rect 418564 320320 418616 320340
rect 418616 320320 418618 320340
rect 437882 320340 437938 320376
rect 437882 320320 437884 320340
rect 437884 320320 437936 320340
rect 437936 320320 437938 320340
rect 408994 10532 409050 10568
rect 408994 10512 408996 10532
rect 408996 10512 409048 10532
rect 409048 10512 409050 10532
rect 409178 7656 409234 7712
rect 413226 9696 413282 9752
rect 413778 9696 413834 9752
rect 411662 7384 411718 7440
rect 413042 7384 413098 7440
rect 411662 7112 411718 7168
rect 413042 6976 413098 7032
rect 411662 3304 411718 3360
rect 414514 3304 414570 3360
rect 418746 10412 418748 10432
rect 418748 10412 418800 10432
rect 418800 10412 418802 10432
rect 418746 10376 418802 10412
rect 418838 4664 418894 4720
rect 424174 10512 424230 10568
rect 424082 6976 424138 7032
rect 424082 3168 424138 3224
rect 428958 7112 429014 7168
rect 433558 3440 433614 3496
rect 433742 3440 433798 3496
rect 433834 3340 433836 3360
rect 433836 3340 433888 3360
rect 433888 3340 433890 3360
rect 433834 3304 433890 3340
rect 437514 6160 437570 6216
rect 438250 7656 438306 7712
rect 451682 3168 451738 3224
rect 453246 6976 453302 7032
rect 464102 320456 464158 320512
rect 457202 320340 457258 320376
rect 457202 320320 457204 320340
rect 457204 320320 457256 320340
rect 457256 320320 457258 320340
rect 462722 6976 462778 7032
rect 462722 3168 462778 3224
rect 462722 3032 462778 3088
rect 464930 3984 464986 4040
rect 483422 320456 483478 320512
rect 476522 320340 476578 320376
rect 476522 320320 476524 320340
rect 476524 320320 476576 320340
rect 476576 320320 476578 320340
rect 466586 3168 466642 3224
rect 468426 3848 468482 3904
rect 473854 7148 473856 7168
rect 473856 7148 473908 7168
rect 473908 7148 473910 7168
rect 473854 7112 473910 7148
rect 474222 7148 474224 7168
rect 474224 7148 474276 7168
rect 474276 7148 474278 7168
rect 474222 7112 474278 7148
rect 472014 3712 472070 3768
rect 475602 3576 475658 3632
rect 480754 6976 480810 7032
rect 479190 3440 479246 3496
rect 480662 3168 480718 3224
rect 483514 6996 483570 7032
rect 483514 6976 483516 6996
rect 483516 6976 483568 6996
rect 483568 6976 483570 6996
rect 482778 3168 482834 3224
rect 488298 320492 488300 320512
rect 488300 320492 488352 320512
rect 488352 320492 488354 320512
rect 488298 320456 488354 320492
rect 486458 10240 486514 10296
rect 493082 320492 493084 320512
rect 493084 320492 493136 320512
rect 493136 320492 493138 320512
rect 493082 320456 493138 320492
rect 505594 320456 505650 320512
rect 505686 320184 505742 320240
rect 511022 7520 511078 7576
rect 511022 7112 511078 7168
rect 515254 4664 515310 4720
rect 528870 298016 528926 298072
rect 529054 298016 529110 298072
rect 528870 278704 528926 278760
rect 529054 278704 529110 278760
rect 528870 259392 528926 259448
rect 529054 259392 529110 259448
rect 528870 240080 528926 240136
rect 529054 240080 529110 240136
rect 528870 220768 528926 220824
rect 529054 220768 529110 220824
rect 528870 191800 528926 191856
rect 529054 191800 529110 191856
rect 528870 172488 528926 172544
rect 529054 172488 529110 172544
rect 529054 164464 529110 164520
rect 526938 164192 526994 164248
rect 529054 164192 529110 164248
rect 529330 164192 529386 164248
rect 535954 259392 536010 259448
rect 536138 259392 536194 259448
rect 535954 240080 536010 240136
rect 536138 240080 536194 240136
rect 535954 220768 536010 220824
rect 536138 220768 536194 220824
rect 535954 191800 536010 191856
rect 536138 191800 536194 191856
rect 535954 172488 536010 172544
rect 536138 172488 536194 172544
rect 535954 164464 536010 164520
rect 535678 164192 535734 164248
rect 535954 164192 536010 164248
rect 536598 164192 536654 164248
rect 520682 6976 520738 7032
rect 520682 6840 520738 6896
rect 519578 4664 519634 4720
rect 534666 7112 534722 7168
rect 534482 6976 534538 7032
rect 541566 320456 541622 320512
rect 544326 320184 544382 320240
rect 546902 7384 546958 7440
rect 546902 6976 546958 7032
rect 552422 288360 552478 288416
rect 552606 288360 552662 288416
rect 552606 278740 552608 278760
rect 552608 278740 552660 278760
rect 552660 278740 552662 278760
rect 552606 278704 552662 278740
rect 552790 278704 552846 278760
rect 552514 259392 552570 259448
rect 552698 259392 552754 259448
rect 552514 241576 552570 241632
rect 552698 241576 552754 241632
rect 553710 231784 553766 231840
rect 553894 231784 553950 231840
rect 553710 222164 553712 222184
rect 553712 222164 553764 222184
rect 553764 222164 553766 222184
rect 553710 222128 553766 222164
rect 553894 222164 553896 222184
rect 553896 222164 553948 222184
rect 553948 222164 553950 222184
rect 553894 222128 553950 222164
rect 553710 202816 553766 202872
rect 553894 202816 553950 202872
rect 552514 201592 552570 201648
rect 552422 201476 552478 201512
rect 552422 201456 552424 201476
rect 552424 201456 552476 201476
rect 552476 201456 552478 201476
rect 553710 193196 553712 193216
rect 553712 193196 553764 193216
rect 553764 193196 553766 193216
rect 553710 193160 553766 193196
rect 553894 193196 553896 193216
rect 553896 193196 553948 193216
rect 553948 193196 553950 193216
rect 553894 193160 553950 193196
rect 553894 183540 553896 183560
rect 553896 183540 553948 183560
rect 553948 183540 553950 183560
rect 553894 183504 553950 183540
rect 553894 173984 553950 174040
rect 553710 173848 553766 173904
rect 553894 173848 553950 173904
rect 552330 172488 552386 172544
rect 552698 172488 552754 172544
rect 553710 125568 553766 125624
rect 553894 125568 553950 125624
rect 553434 113192 553490 113248
rect 553618 113192 553674 113248
rect 552422 104896 552478 104952
rect 552606 104896 552662 104952
rect 553710 87080 553766 87136
rect 553894 86944 553950 87000
rect 552330 67632 552386 67688
rect 552514 67632 552570 67688
rect 553894 48320 553950 48376
rect 554078 48320 554134 48376
rect 560794 87216 560850 87272
rect 560794 87080 560850 87136
rect 560794 48592 560850 48648
rect 560794 48456 560850 48512
rect 558034 7112 558090 7168
rect 571834 278704 571890 278760
rect 572018 278704 572074 278760
rect 571834 259392 571890 259448
rect 572018 259392 572074 259448
rect 571834 240080 571890 240136
rect 572018 240080 572074 240136
rect 571834 220768 571890 220824
rect 572018 220768 572074 220824
rect 571834 191800 571890 191856
rect 572018 191800 572074 191856
rect 571834 172488 571890 172544
rect 572018 172488 572074 172544
rect 570362 164600 570418 164656
rect 571834 164464 571890 164520
rect 570362 164192 570418 164248
rect 571558 164192 571614 164248
rect 571834 164192 571890 164248
rect 572110 164192 572166 164248
rect 567602 6996 567658 7032
rect 567602 6976 567604 6996
rect 567604 6976 567656 6996
rect 567656 6976 567658 6996
rect 569074 6976 569130 7032
rect 573122 4800 573178 4856
rect 578642 7148 578644 7168
rect 578644 7148 578696 7168
rect 578696 7148 578698 7168
rect 578642 7112 578698 7148
rect 580666 289312 580722 289368
rect 580666 273672 580722 273728
rect 580666 195472 580722 195528
rect 580390 148552 580446 148608
rect 580666 85992 580722 86048
rect 580758 54712 580814 54768
rect 581586 8880 581642 8936
rect 583886 7792 583942 7848
rect 583886 7112 583942 7168
<< metal3 >>
rect 11273 700362 11339 700365
rect 304109 700362 304175 700365
rect 11273 700360 304175 700362
rect 11273 700304 11278 700360
rect 11334 700304 304114 700360
rect 304170 700304 304175 700360
rect 11273 700302 304175 700304
rect 11273 700299 11339 700302
rect 304109 700299 304175 700302
rect 580109 696010 580175 696013
rect 584016 696010 584496 696040
rect 580109 696008 584496 696010
rect 580109 695952 580114 696008
rect 580170 695952 584496 696008
rect 580109 695950 584496 695952
rect 580109 695947 580175 695950
rect 584016 695920 584496 695950
rect 496 695466 976 695496
rect 3729 695466 3795 695469
rect 496 695464 3795 695466
rect 496 695408 3734 695464
rect 3790 695408 3795 695464
rect 496 695406 3795 695408
rect 496 695376 976 695406
rect 3729 695403 3795 695406
rect 580109 680370 580175 680373
rect 584016 680370 584496 680400
rect 580109 680368 584496 680370
rect 580109 680312 580114 680368
rect 580170 680312 584496 680368
rect 580109 680310 584496 680312
rect 580109 680307 580175 680310
rect 584016 680280 584496 680310
rect 496 678738 976 678768
rect 3913 678738 3979 678741
rect 496 678736 3979 678738
rect 496 678680 3918 678736
rect 3974 678680 3979 678736
rect 496 678678 3979 678680
rect 496 678648 976 678678
rect 3913 678675 3979 678678
rect 580109 664730 580175 664733
rect 584016 664730 584496 664760
rect 580109 664728 584496 664730
rect 580109 664672 580114 664728
rect 580170 664672 584496 664728
rect 580109 664670 584496 664672
rect 580109 664667 580175 664670
rect 584016 664640 584496 664670
rect 496 662010 976 662040
rect 3913 662010 3979 662013
rect 496 662008 3979 662010
rect 496 661952 3918 662008
rect 3974 661952 3979 662008
rect 496 661950 3979 661952
rect 496 661920 976 661950
rect 3913 661947 3979 661950
rect 580109 649090 580175 649093
rect 584016 649090 584496 649120
rect 580109 649088 584496 649090
rect 580109 649032 580114 649088
rect 580170 649032 584496 649088
rect 580109 649030 584496 649032
rect 580109 649027 580175 649030
rect 584016 649000 584496 649030
rect 496 645282 976 645312
rect 3545 645282 3611 645285
rect 496 645280 3611 645282
rect 496 645224 3550 645280
rect 3606 645224 3611 645280
rect 496 645222 3611 645224
rect 496 645192 976 645222
rect 3545 645219 3611 645222
rect 580109 633450 580175 633453
rect 584016 633450 584496 633480
rect 580109 633448 584496 633450
rect 580109 633392 580114 633448
rect 580170 633392 584496 633448
rect 580109 633390 584496 633392
rect 580109 633387 580175 633390
rect 584016 633360 584496 633390
rect 496 628418 976 628448
rect 3913 628418 3979 628421
rect 496 628416 3979 628418
rect 496 628360 3918 628416
rect 3974 628360 3979 628416
rect 496 628358 3979 628360
rect 496 628328 976 628358
rect 3913 628355 3979 628358
rect 313769 618218 313835 618221
rect 314045 618218 314111 618221
rect 313769 618216 314111 618218
rect 313769 618160 313774 618216
rect 313830 618160 314050 618216
rect 314106 618160 314111 618216
rect 313769 618158 314111 618160
rect 313769 618155 313835 618158
rect 314045 618155 314111 618158
rect 443622 618156 443628 618220
rect 443692 618218 443698 618220
rect 443765 618218 443831 618221
rect 443692 618216 443831 618218
rect 443692 618160 443770 618216
rect 443826 618160 443831 618216
rect 443692 618158 443831 618160
rect 443692 618156 443698 618158
rect 443765 618155 443831 618158
rect 580109 617810 580175 617813
rect 584016 617810 584496 617840
rect 580109 617808 584496 617810
rect 580109 617752 580114 617808
rect 580170 617752 584496 617808
rect 580109 617750 584496 617752
rect 580109 617747 580175 617750
rect 584016 617720 584496 617750
rect 496 611690 976 611720
rect 3821 611690 3887 611693
rect 496 611688 3887 611690
rect 496 611632 3826 611688
rect 3882 611632 3887 611688
rect 496 611630 3887 611632
rect 496 611600 976 611630
rect 3821 611627 3887 611630
rect 443673 608700 443739 608701
rect 443622 608636 443628 608700
rect 443692 608698 443739 608700
rect 573393 608698 573459 608701
rect 573761 608698 573827 608701
rect 443692 608696 443784 608698
rect 443734 608640 443784 608696
rect 443692 608638 443784 608640
rect 573393 608696 573827 608698
rect 573393 608640 573398 608696
rect 573454 608640 573766 608696
rect 573822 608640 573827 608696
rect 573393 608638 573827 608640
rect 443692 608636 443739 608638
rect 443673 608635 443739 608636
rect 573393 608635 573459 608638
rect 573761 608635 573827 608638
rect 580109 602170 580175 602173
rect 584016 602170 584496 602200
rect 580109 602168 584496 602170
rect 580109 602112 580114 602168
rect 580170 602112 584496 602168
rect 580109 602110 584496 602112
rect 580109 602107 580175 602110
rect 584016 602080 584496 602110
rect 496 594962 976 594992
rect 3913 594962 3979 594965
rect 496 594960 3979 594962
rect 496 594904 3918 594960
rect 3974 594904 3979 594960
rect 496 594902 3979 594904
rect 496 594872 976 594902
rect 3913 594899 3979 594902
rect 580109 586530 580175 586533
rect 584016 586530 584496 586560
rect 580109 586528 584496 586530
rect 580109 586472 580114 586528
rect 580170 586472 584496 586528
rect 580109 586470 584496 586472
rect 580109 586467 580175 586470
rect 584016 586440 584496 586470
rect 496 578234 976 578264
rect 3729 578234 3795 578237
rect 496 578232 3795 578234
rect 496 578176 3734 578232
rect 3790 578176 3795 578232
rect 496 578174 3795 578176
rect 496 578144 976 578174
rect 3729 578171 3795 578174
rect 580109 570890 580175 570893
rect 584016 570890 584496 570920
rect 580109 570888 584496 570890
rect 580109 570832 580114 570888
rect 580170 570832 584496 570888
rect 580109 570830 584496 570832
rect 580109 570827 580175 570830
rect 584016 570800 584496 570830
rect 496 561370 976 561400
rect 3913 561370 3979 561373
rect 496 561368 3979 561370
rect 496 561312 3918 561368
rect 3974 561312 3979 561368
rect 496 561310 3979 561312
rect 496 561280 976 561310
rect 3913 561307 3979 561310
rect 378721 560282 378787 560285
rect 378905 560282 378971 560285
rect 378721 560280 378971 560282
rect 378721 560224 378726 560280
rect 378782 560224 378910 560280
rect 378966 560224 378971 560280
rect 378721 560222 378971 560224
rect 378721 560219 378787 560222
rect 378905 560219 378971 560222
rect 508441 560282 508507 560285
rect 508625 560282 508691 560285
rect 508441 560280 508691 560282
rect 508441 560224 508446 560280
rect 508502 560224 508630 560280
rect 508686 560224 508691 560280
rect 508441 560222 508691 560224
rect 508441 560219 508507 560222
rect 508625 560219 508691 560222
rect 313769 557562 313835 557565
rect 314045 557562 314111 557565
rect 313769 557560 314111 557562
rect 313769 557504 313774 557560
rect 313830 557504 314050 557560
rect 314106 557504 314111 557560
rect 313769 557502 314111 557504
rect 313769 557499 313835 557502
rect 314045 557499 314111 557502
rect 580109 555250 580175 555253
rect 584016 555250 584496 555280
rect 580109 555248 584496 555250
rect 580109 555192 580114 555248
rect 580170 555192 584496 555248
rect 580109 555190 584496 555192
rect 580109 555187 580175 555190
rect 584016 555160 584496 555190
rect 496 544642 976 544672
rect 3637 544642 3703 544645
rect 496 544640 3703 544642
rect 496 544584 3642 544640
rect 3698 544584 3703 544640
rect 496 544582 3703 544584
rect 496 544552 976 544582
rect 3637 544579 3703 544582
rect 580109 539610 580175 539613
rect 584016 539610 584496 539640
rect 580109 539608 584496 539610
rect 580109 539552 580114 539608
rect 580170 539552 584496 539608
rect 580109 539550 584496 539552
rect 580109 539547 580175 539550
rect 584016 539520 584496 539550
rect 378997 529820 379063 529821
rect 508717 529820 508783 529821
rect 378997 529818 379044 529820
rect 378952 529816 379044 529818
rect 378952 529760 379002 529816
rect 378952 529758 379044 529760
rect 378997 529756 379044 529758
rect 379108 529756 379114 529820
rect 508717 529818 508764 529820
rect 508672 529816 508764 529818
rect 508672 529760 508722 529816
rect 508672 529758 508764 529760
rect 508717 529756 508764 529758
rect 508828 529756 508834 529820
rect 378997 529755 379063 529756
rect 508717 529755 508783 529756
rect 496 527914 976 527944
rect 3637 527914 3703 527917
rect 496 527912 3703 527914
rect 496 527856 3642 527912
rect 3698 527856 3703 527912
rect 496 527854 3703 527856
rect 496 527824 976 527854
rect 3637 527851 3703 527854
rect 580109 523970 580175 523973
rect 584016 523970 584496 524000
rect 580109 523968 584496 523970
rect 580109 523912 580114 523968
rect 580170 523912 584496 523968
rect 580109 523910 584496 523912
rect 580109 523907 580175 523910
rect 584016 523880 584496 523910
rect 379038 520236 379044 520300
rect 379108 520298 379114 520300
rect 379181 520298 379247 520301
rect 379108 520296 379247 520298
rect 379108 520240 379186 520296
rect 379242 520240 379247 520296
rect 379108 520238 379247 520240
rect 379108 520236 379114 520238
rect 379181 520235 379247 520238
rect 508758 520236 508764 520300
rect 508828 520298 508834 520300
rect 508901 520298 508967 520301
rect 508828 520296 508967 520298
rect 508828 520240 508906 520296
rect 508962 520240 508967 520296
rect 508828 520238 508967 520240
rect 508828 520236 508834 520238
rect 508901 520235 508967 520238
rect 313769 518938 313835 518941
rect 314045 518938 314111 518941
rect 313769 518936 314111 518938
rect 313769 518880 313774 518936
rect 313830 518880 314050 518936
rect 314106 518880 314111 518936
rect 313769 518878 314111 518880
rect 313769 518875 313835 518878
rect 314045 518875 314111 518878
rect 443489 512002 443555 512005
rect 443673 512002 443739 512005
rect 443489 512000 443739 512002
rect 443489 511944 443494 512000
rect 443550 511944 443678 512000
rect 443734 511944 443739 512000
rect 443489 511942 443739 511944
rect 443489 511939 443555 511942
rect 443673 511939 443739 511942
rect 573209 512002 573275 512005
rect 573393 512002 573459 512005
rect 573209 512000 573459 512002
rect 573209 511944 573214 512000
rect 573270 511944 573398 512000
rect 573454 511944 573459 512000
rect 573209 511942 573459 511944
rect 573209 511939 573275 511942
rect 573393 511939 573459 511942
rect 496 511186 976 511216
rect 4005 511186 4071 511189
rect 496 511184 4071 511186
rect 496 511128 4010 511184
rect 4066 511128 4071 511184
rect 496 511126 4071 511128
rect 496 511096 976 511126
rect 4005 511123 4071 511126
rect 580109 508330 580175 508333
rect 584016 508330 584496 508360
rect 580109 508328 584496 508330
rect 580109 508272 580114 508328
rect 580170 508272 584496 508328
rect 580109 508270 584496 508272
rect 580109 508267 580175 508270
rect 584016 508240 584496 508270
rect 378537 502346 378603 502349
rect 378813 502346 378879 502349
rect 378537 502344 378879 502346
rect 378537 502288 378542 502344
rect 378598 502288 378818 502344
rect 378874 502288 378879 502344
rect 378537 502286 378879 502288
rect 378537 502283 378603 502286
rect 378813 502283 378879 502286
rect 508257 502346 508323 502349
rect 508533 502346 508599 502349
rect 508257 502344 508599 502346
rect 508257 502288 508262 502344
rect 508318 502288 508538 502344
rect 508594 502288 508599 502344
rect 508257 502286 508599 502288
rect 508257 502283 508323 502286
rect 508533 502283 508599 502286
rect 496 494322 976 494352
rect 3729 494322 3795 494325
rect 496 494320 3795 494322
rect 496 494264 3734 494320
rect 3790 494264 3795 494320
rect 496 494262 3795 494264
rect 496 494232 976 494262
rect 3729 494259 3795 494262
rect 378537 492690 378603 492693
rect 378721 492690 378787 492693
rect 378537 492688 378787 492690
rect 378537 492632 378542 492688
rect 378598 492632 378726 492688
rect 378782 492632 378787 492688
rect 378537 492630 378787 492632
rect 378537 492627 378603 492630
rect 378721 492627 378787 492630
rect 508257 492690 508323 492693
rect 508441 492690 508507 492693
rect 508257 492688 508507 492690
rect 508257 492632 508262 492688
rect 508318 492632 508446 492688
rect 508502 492632 508507 492688
rect 508257 492630 508507 492632
rect 508257 492627 508323 492630
rect 508441 492627 508507 492630
rect 580109 492690 580175 492693
rect 584016 492690 584496 492720
rect 580109 492688 584496 492690
rect 580109 492632 580114 492688
rect 580170 492632 584496 492688
rect 580109 492630 584496 492632
rect 580109 492627 580175 492630
rect 584016 492600 584496 492630
rect 496 477594 976 477624
rect 3913 477594 3979 477597
rect 496 477592 3979 477594
rect 496 477536 3918 477592
rect 3974 477536 3979 477592
rect 496 477534 3979 477536
rect 496 477504 976 477534
rect 3913 477531 3979 477534
rect 580109 477050 580175 477053
rect 584016 477050 584496 477080
rect 580109 477048 584496 477050
rect 580109 476992 580114 477048
rect 580170 476992 584496 477048
rect 580109 476990 584496 476992
rect 580109 476987 580175 476990
rect 584016 476960 584496 476990
rect 283593 463178 283659 463181
rect 288193 463178 288259 463181
rect 283593 463176 288259 463178
rect 283593 463120 283598 463176
rect 283654 463120 288198 463176
rect 288254 463120 288259 463176
rect 283593 463118 288259 463120
rect 283593 463115 283659 463118
rect 288193 463115 288259 463118
rect 288377 463178 288443 463181
rect 293161 463178 293227 463181
rect 288377 463176 293227 463178
rect 288377 463120 288382 463176
rect 288438 463120 293166 463176
rect 293222 463120 293227 463176
rect 288377 463118 293227 463120
rect 288377 463115 288443 463118
rect 293161 463115 293227 463118
rect 282305 463042 282371 463045
rect 283409 463042 283475 463045
rect 282305 463040 283475 463042
rect 282305 462984 282310 463040
rect 282366 462984 283414 463040
rect 283470 462984 283475 463040
rect 282305 462982 283475 462984
rect 282305 462979 282371 462982
rect 283409 462979 283475 462982
rect 3913 462498 3979 462501
rect 342381 462498 342447 462501
rect 3913 462496 342447 462498
rect 3913 462440 3918 462496
rect 3974 462440 342386 462496
rect 342442 462440 342447 462496
rect 3913 462438 342447 462440
rect 3913 462435 3979 462438
rect 342381 462435 342447 462438
rect 580661 461410 580727 461413
rect 584016 461410 584496 461440
rect 580661 461408 584496 461410
rect 580661 461352 580666 461408
rect 580722 461352 584496 461408
rect 580661 461350 584496 461352
rect 580661 461347 580727 461350
rect 584016 461320 584496 461350
rect 496 460866 976 460896
rect 3637 460866 3703 460869
rect 496 460864 3703 460866
rect 496 460808 3642 460864
rect 3698 460808 3703 460864
rect 496 460806 3703 460808
rect 496 460776 976 460806
rect 3637 460803 3703 460806
rect 232165 459644 232231 459645
rect 232165 459640 232212 459644
rect 232276 459642 232282 459644
rect 233177 459642 233243 459645
rect 236213 459644 236279 459645
rect 233494 459642 233500 459644
rect 232165 459584 232170 459640
rect 232165 459580 232212 459584
rect 232276 459582 232322 459642
rect 233177 459640 233500 459642
rect 233177 459584 233182 459640
rect 233238 459584 233500 459640
rect 233177 459582 233500 459584
rect 232276 459580 232282 459582
rect 232165 459579 232231 459580
rect 233177 459579 233243 459582
rect 233494 459580 233500 459582
rect 233564 459580 233570 459644
rect 236213 459640 236260 459644
rect 236324 459642 236330 459644
rect 237409 459642 237475 459645
rect 237726 459642 237732 459644
rect 236213 459584 236218 459640
rect 236213 459580 236260 459584
rect 236324 459582 236370 459642
rect 237409 459640 237732 459642
rect 237409 459584 237414 459640
rect 237470 459584 237732 459640
rect 237409 459582 237732 459584
rect 236324 459580 236330 459582
rect 236213 459579 236279 459580
rect 237409 459579 237475 459582
rect 237726 459580 237732 459582
rect 237796 459580 237802 459644
rect 238513 459642 238579 459645
rect 239014 459642 239020 459644
rect 238513 459640 239020 459642
rect 238513 459584 238518 459640
rect 238574 459584 239020 459640
rect 238513 459582 239020 459584
rect 238513 459579 238579 459582
rect 239014 459580 239020 459582
rect 239084 459580 239090 459644
rect 239617 459642 239683 459645
rect 240486 459642 240492 459644
rect 239617 459640 240492 459642
rect 239617 459584 239622 459640
rect 239678 459584 240492 459640
rect 239617 459582 240492 459584
rect 239617 459579 239683 459582
rect 240486 459580 240492 459582
rect 240556 459580 240562 459644
rect 241641 459642 241707 459645
rect 241774 459642 241780 459644
rect 241641 459640 241780 459642
rect 241641 459584 241646 459640
rect 241702 459584 241780 459640
rect 241641 459582 241780 459584
rect 241641 459579 241707 459582
rect 241774 459580 241780 459582
rect 241844 459580 241850 459644
rect 242745 459642 242811 459645
rect 244585 459644 244651 459645
rect 243246 459642 243252 459644
rect 242745 459640 243252 459642
rect 242745 459584 242750 459640
rect 242806 459584 243252 459640
rect 242745 459582 243252 459584
rect 242745 459579 242811 459582
rect 243246 459580 243252 459582
rect 243316 459580 243322 459644
rect 244534 459642 244540 459644
rect 244494 459582 244540 459642
rect 244604 459640 244651 459644
rect 244646 459584 244651 459640
rect 244534 459580 244540 459582
rect 244604 459580 244651 459584
rect 244585 459579 244651 459580
rect 245873 459642 245939 459645
rect 246006 459642 246012 459644
rect 245873 459640 246012 459642
rect 245873 459584 245878 459640
rect 245934 459584 246012 459640
rect 245873 459582 246012 459584
rect 245873 459579 245939 459582
rect 246006 459580 246012 459582
rect 246076 459580 246082 459644
rect 246977 459642 247043 459645
rect 248817 459644 248883 459645
rect 247294 459642 247300 459644
rect 246977 459640 247300 459642
rect 246977 459584 246982 459640
rect 247038 459584 247300 459640
rect 246977 459582 247300 459584
rect 246977 459579 247043 459582
rect 247294 459580 247300 459582
rect 247364 459580 247370 459644
rect 248766 459642 248772 459644
rect 248726 459582 248772 459642
rect 248836 459640 248883 459644
rect 248878 459584 248883 459640
rect 248766 459580 248772 459582
rect 248836 459580 248883 459584
rect 248817 459579 248883 459580
rect 251209 459642 251275 459645
rect 251526 459642 251532 459644
rect 251209 459640 251532 459642
rect 251209 459584 251214 459640
rect 251270 459584 251532 459640
rect 251209 459582 251532 459584
rect 251209 459579 251275 459582
rect 251526 459580 251532 459582
rect 251596 459580 251602 459644
rect 252129 459642 252195 459645
rect 252814 459642 252820 459644
rect 252129 459640 252820 459642
rect 252129 459584 252134 459640
rect 252190 459584 252820 459640
rect 252129 459582 252820 459584
rect 252129 459579 252195 459582
rect 252814 459580 252820 459582
rect 252884 459580 252890 459644
rect 342790 459580 342796 459644
rect 342860 459642 342866 459644
rect 343117 459642 343183 459645
rect 342860 459640 343183 459642
rect 342860 459584 343122 459640
rect 343178 459584 343183 459640
rect 342860 459582 343183 459584
rect 342860 459580 342866 459582
rect 343117 459579 343183 459582
rect 344078 459580 344084 459644
rect 344148 459642 344154 459644
rect 344221 459642 344287 459645
rect 344148 459640 344287 459642
rect 344148 459584 344226 459640
rect 344282 459584 344287 459640
rect 344148 459582 344287 459584
rect 344148 459580 344154 459582
rect 344221 459579 344287 459582
rect 345550 459580 345556 459644
rect 345620 459642 345626 459644
rect 346245 459642 346311 459645
rect 345620 459640 346311 459642
rect 345620 459584 346250 459640
rect 346306 459584 346311 459640
rect 345620 459582 346311 459584
rect 345620 459580 345626 459582
rect 346245 459579 346311 459582
rect 346838 459580 346844 459644
rect 346908 459642 346914 459644
rect 347349 459642 347415 459645
rect 346908 459640 347415 459642
rect 346908 459584 347354 459640
rect 347410 459584 347415 459640
rect 346908 459582 347415 459584
rect 346908 459580 346914 459582
rect 347349 459579 347415 459582
rect 348310 459580 348316 459644
rect 348380 459642 348386 459644
rect 348453 459642 348519 459645
rect 348380 459640 348519 459642
rect 348380 459584 348458 459640
rect 348514 459584 348519 459640
rect 348380 459582 348519 459584
rect 348380 459580 348386 459582
rect 348453 459579 348519 459582
rect 580661 445770 580727 445773
rect 584016 445770 584496 445800
rect 580661 445768 584496 445770
rect 580661 445712 580666 445768
rect 580722 445712 584496 445768
rect 580661 445710 584496 445712
rect 580661 445707 580727 445710
rect 584016 445680 584496 445710
rect 496 444138 976 444168
rect 3637 444138 3703 444141
rect 496 444136 3703 444138
rect 496 444080 3642 444136
rect 3698 444080 3703 444136
rect 496 444078 3703 444080
rect 496 444048 976 444078
rect 3637 444075 3703 444078
rect 580661 430130 580727 430133
rect 584016 430130 584496 430160
rect 580661 430128 584496 430130
rect 580661 430072 580666 430128
rect 580722 430072 584496 430128
rect 580661 430070 584496 430072
rect 580661 430067 580727 430070
rect 584016 430040 584496 430070
rect 496 427274 976 427304
rect 3637 427274 3703 427277
rect 496 427272 3703 427274
rect 496 427216 3642 427272
rect 3698 427216 3703 427272
rect 496 427214 3703 427216
rect 496 427184 976 427214
rect 3637 427211 3703 427214
rect 580661 414490 580727 414493
rect 584016 414490 584496 414520
rect 580661 414488 584496 414490
rect 580661 414432 580666 414488
rect 580722 414432 584496 414488
rect 580661 414430 584496 414432
rect 580661 414427 580727 414430
rect 584016 414400 584496 414430
rect 496 410546 976 410576
rect 3821 410546 3887 410549
rect 496 410544 3887 410546
rect 496 410488 3826 410544
rect 3882 410488 3887 410544
rect 496 410486 3887 410488
rect 496 410456 976 410486
rect 3821 410483 3887 410486
rect 580661 398850 580727 398853
rect 584016 398850 584496 398880
rect 580661 398848 584496 398850
rect 580661 398792 580666 398848
rect 580722 398792 584496 398848
rect 580661 398790 584496 398792
rect 580661 398787 580727 398790
rect 584016 398760 584496 398790
rect 496 393818 976 393848
rect 3821 393818 3887 393821
rect 496 393816 3887 393818
rect 496 393760 3826 393816
rect 3882 393760 3887 393816
rect 496 393758 3887 393760
rect 496 393728 976 393758
rect 3821 393755 3887 393758
rect 580661 383210 580727 383213
rect 584016 383210 584496 383240
rect 580661 383208 584496 383210
rect 580661 383152 580666 383208
rect 580722 383152 584496 383208
rect 580661 383150 584496 383152
rect 580661 383147 580727 383150
rect 584016 383120 584496 383150
rect 496 377090 976 377120
rect 3545 377090 3611 377093
rect 496 377088 3611 377090
rect 496 377032 3550 377088
rect 3606 377032 3611 377088
rect 496 377030 3611 377032
rect 496 377000 976 377030
rect 3545 377027 3611 377030
rect 580661 367570 580727 367573
rect 584016 367570 584496 367600
rect 580661 367568 584496 367570
rect 580661 367512 580666 367568
rect 580722 367512 584496 367568
rect 580661 367510 584496 367512
rect 580661 367507 580727 367510
rect 584016 367480 584496 367510
rect 496 360362 976 360392
rect 3821 360362 3887 360365
rect 496 360360 3887 360362
rect 496 360304 3826 360360
rect 3882 360304 3887 360360
rect 496 360302 3887 360304
rect 496 360272 976 360302
rect 3821 360299 3887 360302
rect 580661 351930 580727 351933
rect 584016 351930 584496 351960
rect 580661 351928 584496 351930
rect 580661 351872 580666 351928
rect 580722 351872 584496 351928
rect 580661 351870 584496 351872
rect 580661 351867 580727 351870
rect 584016 351840 584496 351870
rect 496 343498 976 343528
rect 3821 343498 3887 343501
rect 496 343496 3887 343498
rect 496 343440 3826 343496
rect 3882 343440 3887 343496
rect 496 343438 3887 343440
rect 496 343408 976 343438
rect 3821 343435 3887 343438
rect 333365 338058 333431 338061
rect 333549 338058 333615 338061
rect 333365 338056 333615 338058
rect 333365 338000 333370 338056
rect 333426 338000 333554 338056
rect 333610 338000 333615 338056
rect 333365 337998 333615 338000
rect 333365 337995 333431 337998
rect 333549 337995 333615 337998
rect 128849 337922 128915 337925
rect 138417 337922 138483 337925
rect 128849 337920 138483 337922
rect 128849 337864 128854 337920
rect 128910 337864 138422 337920
rect 138478 337864 138483 337920
rect 128849 337862 138483 337864
rect 128849 337859 128915 337862
rect 138417 337859 138483 337862
rect 119281 337786 119347 337789
rect 129033 337786 129099 337789
rect 119281 337784 129099 337786
rect 119281 337728 119286 337784
rect 119342 337728 129038 337784
rect 129094 337728 129099 337784
rect 119281 337726 129099 337728
rect 119281 337723 119347 337726
rect 129033 337723 129099 337726
rect 142649 337786 142715 337789
rect 152217 337786 152283 337789
rect 142649 337784 152283 337786
rect 142649 337728 142654 337784
rect 142710 337728 152222 337784
rect 152278 337728 152283 337784
rect 142649 337726 152283 337728
rect 142649 337723 142715 337726
rect 152217 337723 152283 337726
rect 161969 337786 162035 337789
rect 171537 337786 171603 337789
rect 161969 337784 171603 337786
rect 161969 337728 161974 337784
rect 162030 337728 171542 337784
rect 171598 337728 171603 337784
rect 161969 337726 171603 337728
rect 161969 337723 162035 337726
rect 171537 337723 171603 337726
rect 181289 337786 181355 337789
rect 190857 337786 190923 337789
rect 181289 337784 190923 337786
rect 181289 337728 181294 337784
rect 181350 337728 190862 337784
rect 190918 337728 190923 337784
rect 181289 337726 190923 337728
rect 181289 337723 181355 337726
rect 190857 337723 190923 337726
rect 200609 337786 200675 337789
rect 210177 337786 210243 337789
rect 200609 337784 210243 337786
rect 200609 337728 200614 337784
rect 200670 337728 210182 337784
rect 210238 337728 210243 337784
rect 200609 337726 210243 337728
rect 200609 337723 200675 337726
rect 210177 337723 210243 337726
rect 219929 337786 219995 337789
rect 232809 337786 232875 337789
rect 219929 337784 232875 337786
rect 219929 337728 219934 337784
rect 219990 337728 232814 337784
rect 232870 337728 232875 337784
rect 219929 337726 232875 337728
rect 219929 337723 219995 337726
rect 232809 337723 232875 337726
rect 128573 337650 128639 337653
rect 128941 337650 129007 337653
rect 128573 337648 129007 337650
rect 128573 337592 128578 337648
rect 128634 337592 128946 337648
rect 129002 337592 129007 337648
rect 128573 337590 129007 337592
rect 128573 337587 128639 337590
rect 128941 337587 129007 337590
rect 129217 337650 129283 337653
rect 138325 337650 138391 337653
rect 226921 337650 226987 337653
rect 129217 337648 131074 337650
rect 129217 337592 129222 337648
rect 129278 337592 131074 337648
rect 129217 337590 131074 337592
rect 129217 337587 129283 337590
rect 94349 337514 94415 337517
rect 103917 337514 103983 337517
rect 94349 337512 103983 337514
rect 94349 337456 94354 337512
rect 94410 337456 103922 337512
rect 103978 337456 103983 337512
rect 94349 337454 103983 337456
rect 94349 337451 94415 337454
rect 103917 337451 103983 337454
rect 123881 337514 123947 337517
rect 128757 337514 128823 337517
rect 123881 337512 128823 337514
rect 123881 337456 123886 337512
rect 123942 337456 128762 337512
rect 128818 337456 128823 337512
rect 123881 337454 128823 337456
rect 131014 337514 131074 337590
rect 138325 337648 226987 337650
rect 138325 337592 138330 337648
rect 138386 337592 226926 337648
rect 226982 337592 226987 337648
rect 138325 337590 226987 337592
rect 138325 337587 138391 337590
rect 226921 337587 226987 337590
rect 142281 337514 142347 337517
rect 131014 337512 142347 337514
rect 131014 337456 142286 337512
rect 142342 337456 142347 337512
rect 131014 337454 142347 337456
rect 123881 337451 123947 337454
rect 128757 337451 128823 337454
rect 142281 337451 142347 337454
rect 142465 337514 142531 337517
rect 142741 337514 142807 337517
rect 142465 337512 142807 337514
rect 142465 337456 142470 337512
rect 142526 337456 142746 337512
rect 142802 337456 142807 337512
rect 142465 337454 142807 337456
rect 142465 337451 142531 337454
rect 142741 337451 142807 337454
rect 152125 337514 152191 337517
rect 152401 337514 152467 337517
rect 152125 337512 152467 337514
rect 152125 337456 152130 337512
rect 152186 337456 152406 337512
rect 152462 337456 152467 337512
rect 152125 337454 152467 337456
rect 152125 337451 152191 337454
rect 152401 337451 152467 337454
rect 152585 337514 152651 337517
rect 161601 337514 161667 337517
rect 152585 337512 161667 337514
rect 152585 337456 152590 337512
rect 152646 337456 161606 337512
rect 161662 337456 161667 337512
rect 152585 337454 161667 337456
rect 152585 337451 152651 337454
rect 161601 337451 161667 337454
rect 161785 337514 161851 337517
rect 162061 337514 162127 337517
rect 161785 337512 162127 337514
rect 161785 337456 161790 337512
rect 161846 337456 162066 337512
rect 162122 337456 162127 337512
rect 161785 337454 162127 337456
rect 161785 337451 161851 337454
rect 162061 337451 162127 337454
rect 171445 337514 171511 337517
rect 171721 337514 171787 337517
rect 171445 337512 171787 337514
rect 171445 337456 171450 337512
rect 171506 337456 171726 337512
rect 171782 337456 171787 337512
rect 171445 337454 171787 337456
rect 171445 337451 171511 337454
rect 171721 337451 171787 337454
rect 171905 337514 171971 337517
rect 180921 337514 180987 337517
rect 171905 337512 180987 337514
rect 171905 337456 171910 337512
rect 171966 337456 180926 337512
rect 180982 337456 180987 337512
rect 171905 337454 180987 337456
rect 171905 337451 171971 337454
rect 180921 337451 180987 337454
rect 181105 337514 181171 337517
rect 181381 337514 181447 337517
rect 181105 337512 181447 337514
rect 181105 337456 181110 337512
rect 181166 337456 181386 337512
rect 181442 337456 181447 337512
rect 181105 337454 181447 337456
rect 181105 337451 181171 337454
rect 181381 337451 181447 337454
rect 190765 337514 190831 337517
rect 191041 337514 191107 337517
rect 190765 337512 191107 337514
rect 190765 337456 190770 337512
rect 190826 337456 191046 337512
rect 191102 337456 191107 337512
rect 190765 337454 191107 337456
rect 190765 337451 190831 337454
rect 191041 337451 191107 337454
rect 191225 337514 191291 337517
rect 200241 337514 200307 337517
rect 191225 337512 200307 337514
rect 191225 337456 191230 337512
rect 191286 337456 200246 337512
rect 200302 337456 200307 337512
rect 191225 337454 200307 337456
rect 191225 337451 191291 337454
rect 200241 337451 200307 337454
rect 200425 337514 200491 337517
rect 200701 337514 200767 337517
rect 200425 337512 200767 337514
rect 200425 337456 200430 337512
rect 200486 337456 200706 337512
rect 200762 337456 200767 337512
rect 200425 337454 200767 337456
rect 200425 337451 200491 337454
rect 200701 337451 200767 337454
rect 210085 337514 210151 337517
rect 210361 337514 210427 337517
rect 210085 337512 210427 337514
rect 210085 337456 210090 337512
rect 210146 337456 210366 337512
rect 210422 337456 210427 337512
rect 210085 337454 210427 337456
rect 210085 337451 210151 337454
rect 210361 337451 210427 337454
rect 210545 337514 210611 337517
rect 219561 337514 219627 337517
rect 210545 337512 219627 337514
rect 210545 337456 210550 337512
rect 210606 337456 219566 337512
rect 219622 337456 219627 337512
rect 210545 337454 219627 337456
rect 210545 337451 210611 337454
rect 219561 337451 219627 337454
rect 219745 337514 219811 337517
rect 220021 337514 220087 337517
rect 219745 337512 220087 337514
rect 219745 337456 219750 337512
rect 219806 337456 220026 337512
rect 220082 337456 220087 337512
rect 219745 337454 220087 337456
rect 219745 337451 219811 337454
rect 220021 337451 220087 337454
rect 5937 337378 6003 337381
rect 231429 337378 231495 337381
rect 5937 337376 231495 337378
rect 5937 337320 5942 337376
rect 5998 337320 231434 337376
rect 231490 337320 231495 337376
rect 5937 337318 231495 337320
rect 5937 337315 6003 337318
rect 231429 337315 231495 337318
rect 138325 337242 138391 337245
rect 142557 337242 142623 337245
rect 138325 337240 142623 337242
rect 138325 337184 138330 337240
rect 138386 337184 142562 337240
rect 142618 337184 142623 337240
rect 138325 337182 142623 337184
rect 138325 337179 138391 337182
rect 142557 337179 142623 337182
rect 152309 337242 152375 337245
rect 161877 337242 161943 337245
rect 152309 337240 161943 337242
rect 152309 337184 152314 337240
rect 152370 337184 161882 337240
rect 161938 337184 161943 337240
rect 152309 337182 161943 337184
rect 152309 337179 152375 337182
rect 161877 337179 161943 337182
rect 171629 337242 171695 337245
rect 181197 337242 181263 337245
rect 171629 337240 181263 337242
rect 171629 337184 171634 337240
rect 171690 337184 181202 337240
rect 181258 337184 181263 337240
rect 171629 337182 181263 337184
rect 171629 337179 171695 337182
rect 181197 337179 181263 337182
rect 190949 337242 191015 337245
rect 200517 337242 200583 337245
rect 190949 337240 200583 337242
rect 190949 337184 190954 337240
rect 191010 337184 200522 337240
rect 200578 337184 200583 337240
rect 190949 337182 200583 337184
rect 190949 337179 191015 337182
rect 200517 337179 200583 337182
rect 210269 337242 210335 337245
rect 219837 337242 219903 337245
rect 210269 337240 219903 337242
rect 210269 337184 210274 337240
rect 210330 337184 219842 337240
rect 219898 337184 219903 337240
rect 210269 337182 219903 337184
rect 210269 337179 210335 337182
rect 219837 337179 219903 337182
rect 273289 336970 273355 336973
rect 273289 336968 273490 336970
rect 273289 336912 273294 336968
rect 273350 336912 273490 336968
rect 273289 336910 273490 336912
rect 273289 336907 273355 336910
rect 273289 336834 273355 336837
rect 273430 336834 273490 336910
rect 273289 336832 273490 336834
rect 273289 336776 273294 336832
rect 273350 336776 273490 336832
rect 273289 336774 273490 336776
rect 273289 336771 273355 336774
rect 392245 336698 392311 336701
rect 392429 336698 392495 336701
rect 392245 336696 392495 336698
rect 392245 336640 392250 336696
rect 392306 336640 392434 336696
rect 392490 336640 392495 336696
rect 392245 336638 392495 336640
rect 392245 336635 392311 336638
rect 392429 336635 392495 336638
rect 580385 336290 580451 336293
rect 584016 336290 584496 336320
rect 580385 336288 584496 336290
rect 580385 336232 580390 336288
rect 580446 336232 584496 336288
rect 580385 336230 584496 336232
rect 580385 336227 580451 336230
rect 584016 336200 584496 336230
rect 318645 335746 318711 335749
rect 319105 335746 319171 335749
rect 318645 335744 319171 335746
rect 318645 335688 318650 335744
rect 318706 335688 319110 335744
rect 319166 335688 319171 335744
rect 318645 335686 319171 335688
rect 318645 335683 318711 335686
rect 319105 335683 319171 335686
rect 272921 333978 272987 333981
rect 273289 333978 273355 333981
rect 272921 333976 273355 333978
rect 272921 333920 272926 333976
rect 272982 333920 273294 333976
rect 273350 333920 273355 333976
rect 272921 333918 273355 333920
rect 272921 333915 272987 333918
rect 273289 333915 273355 333918
rect 496 326770 976 326800
rect 4373 326770 4439 326773
rect 496 326768 4439 326770
rect 496 326712 4378 326768
rect 4434 326712 4439 326768
rect 496 326710 4439 326712
rect 496 326680 976 326710
rect 4373 326707 4439 326710
rect 275497 324322 275563 324325
rect 275681 324322 275747 324325
rect 275497 324320 275747 324322
rect 275497 324264 275502 324320
rect 275558 324264 275686 324320
rect 275742 324264 275747 324320
rect 275497 324262 275747 324264
rect 275497 324259 275563 324262
rect 275681 324259 275747 324262
rect 280598 320588 280604 320652
rect 280668 320588 280674 320652
rect 333733 320650 333799 320653
rect 360597 320650 360663 320653
rect 584016 320650 584496 320680
rect 328998 320648 333799 320650
rect 328998 320592 333738 320648
rect 333794 320592 333799 320648
rect 328998 320590 333799 320592
rect 251526 320452 251532 320516
rect 251596 320514 251602 320516
rect 254153 320514 254219 320517
rect 280606 320514 280666 320588
rect 251596 320512 254219 320514
rect 251596 320456 254158 320512
rect 254214 320456 254219 320512
rect 251596 320454 254219 320456
rect 251596 320452 251602 320454
rect 254153 320451 254219 320454
rect 274350 320454 280666 320514
rect 294633 320514 294699 320517
rect 299918 320514 299924 320516
rect 294633 320512 299924 320514
rect 294633 320456 294638 320512
rect 294694 320456 299924 320512
rect 294633 320454 299924 320456
rect 261237 320378 261303 320381
rect 274350 320378 274410 320454
rect 294633 320451 294699 320454
rect 299918 320452 299924 320454
rect 299988 320452 299994 320516
rect 312254 320454 319122 320514
rect 261237 320376 274410 320378
rect 261237 320320 261242 320376
rect 261298 320320 274410 320376
rect 261237 320318 274410 320320
rect 261237 320315 261303 320318
rect 309486 320316 309492 320380
rect 309556 320378 309562 320380
rect 312254 320378 312314 320454
rect 309556 320318 312314 320378
rect 309556 320316 309562 320318
rect 280782 320180 280788 320244
rect 280852 320242 280858 320244
rect 290309 320242 290375 320245
rect 280852 320240 290375 320242
rect 280852 320184 290314 320240
rect 290370 320184 290375 320240
rect 280852 320182 290375 320184
rect 319062 320242 319122 320454
rect 328998 320378 329058 320590
rect 333733 320587 333799 320590
rect 351078 320648 360663 320650
rect 351078 320592 360602 320648
rect 360658 320592 360663 320648
rect 351078 320590 360663 320592
rect 351078 320378 351138 320590
rect 360597 320587 360663 320590
rect 583838 320590 584496 320650
rect 425457 320514 425523 320517
rect 444777 320514 444843 320517
rect 464097 320514 464163 320517
rect 483417 320514 483483 320517
rect 488293 320514 488359 320517
rect 399286 320454 409098 320514
rect 324030 320318 329058 320378
rect 348134 320318 351138 320378
rect 360689 320378 360755 320381
rect 360689 320376 370274 320378
rect 360689 320320 360694 320376
rect 360750 320320 370274 320376
rect 360689 320318 370274 320320
rect 324030 320242 324090 320318
rect 319062 320182 324090 320242
rect 333733 320242 333799 320245
rect 338558 320242 338564 320244
rect 333733 320240 338564 320242
rect 333733 320184 333738 320240
rect 333794 320184 338564 320240
rect 333733 320182 338564 320184
rect 280852 320180 280858 320182
rect 290309 320179 290375 320182
rect 333733 320179 333799 320182
rect 338558 320180 338564 320182
rect 338628 320180 338634 320244
rect 343393 320242 343459 320245
rect 348134 320242 348194 320318
rect 360689 320315 360755 320318
rect 343393 320240 348194 320242
rect 343393 320184 343398 320240
rect 343454 320184 348194 320240
rect 343393 320182 348194 320184
rect 370214 320242 370274 320318
rect 370398 320318 379842 320378
rect 370398 320242 370458 320318
rect 370214 320182 370458 320242
rect 379782 320242 379842 320318
rect 399286 320242 399346 320454
rect 409038 320378 409098 320454
rect 425457 320512 428418 320514
rect 425457 320456 425462 320512
rect 425518 320456 428418 320512
rect 425457 320454 428418 320456
rect 425457 320451 425523 320454
rect 418557 320378 418623 320381
rect 409038 320376 418623 320378
rect 409038 320320 418562 320376
rect 418618 320320 418623 320376
rect 409038 320318 418623 320320
rect 428358 320378 428418 320454
rect 444777 320512 447738 320514
rect 444777 320456 444782 320512
rect 444838 320456 447738 320512
rect 444777 320454 447738 320456
rect 444777 320451 444843 320454
rect 437877 320378 437943 320381
rect 428358 320376 437943 320378
rect 428358 320320 437882 320376
rect 437938 320320 437943 320376
rect 428358 320318 437943 320320
rect 447678 320378 447738 320454
rect 464097 320512 467058 320514
rect 464097 320456 464102 320512
rect 464158 320456 467058 320512
rect 464097 320454 467058 320456
rect 464097 320451 464163 320454
rect 457197 320378 457263 320381
rect 447678 320376 457263 320378
rect 447678 320320 457202 320376
rect 457258 320320 457263 320376
rect 447678 320318 457263 320320
rect 466998 320378 467058 320454
rect 483417 320512 488359 320514
rect 483417 320456 483422 320512
rect 483478 320456 488298 320512
rect 488354 320456 488359 320512
rect 483417 320454 488359 320456
rect 483417 320451 483483 320454
rect 488293 320451 488359 320454
rect 493077 320514 493143 320517
rect 505589 320514 505655 320517
rect 493077 320512 505655 320514
rect 493077 320456 493082 320512
rect 493138 320456 505594 320512
rect 505650 320456 505655 320512
rect 493077 320454 505655 320456
rect 493077 320451 493143 320454
rect 505589 320451 505655 320454
rect 512438 320452 512444 320516
rect 512508 320514 512514 320516
rect 541561 320514 541627 320517
rect 512508 320454 529066 320514
rect 512508 320452 512514 320454
rect 476517 320378 476583 320381
rect 466998 320376 476583 320378
rect 466998 320320 476522 320376
rect 476578 320320 476583 320376
rect 466998 320318 476583 320320
rect 529006 320378 529066 320454
rect 538758 320512 541627 320514
rect 538758 320456 541566 320512
rect 541622 320456 541627 320512
rect 538758 320454 541627 320456
rect 529006 320318 538634 320378
rect 418557 320315 418623 320318
rect 437877 320315 437943 320318
rect 457197 320315 457263 320318
rect 476517 320315 476583 320318
rect 379782 320182 399346 320242
rect 505681 320242 505747 320245
rect 512438 320242 512444 320244
rect 505681 320240 512444 320242
rect 505681 320184 505686 320240
rect 505742 320184 512444 320240
rect 505681 320182 512444 320184
rect 343393 320179 343459 320182
rect 505681 320179 505747 320182
rect 512438 320180 512444 320182
rect 512508 320180 512514 320244
rect 538574 320242 538634 320318
rect 538758 320242 538818 320454
rect 541561 320451 541627 320454
rect 551078 320452 551084 320516
rect 551148 320514 551154 320516
rect 551148 320454 567706 320514
rect 551148 320452 551154 320454
rect 567646 320378 567706 320454
rect 583838 320378 583898 320590
rect 584016 320560 584496 320590
rect 567646 320318 577274 320378
rect 538574 320182 538818 320242
rect 544321 320242 544387 320245
rect 551078 320242 551084 320244
rect 544321 320240 551084 320242
rect 544321 320184 544326 320240
rect 544382 320184 551084 320240
rect 544321 320182 551084 320184
rect 544321 320179 544387 320182
rect 551078 320180 551084 320182
rect 551148 320180 551154 320244
rect 577214 320242 577274 320318
rect 577398 320318 583898 320378
rect 577398 320242 577458 320318
rect 577214 320182 577458 320242
rect 299918 320044 299924 320108
rect 299988 320106 299994 320108
rect 309486 320106 309492 320108
rect 299988 320046 309492 320106
rect 299988 320044 299994 320046
rect 309486 320044 309492 320046
rect 309556 320044 309562 320108
rect 338558 319908 338564 319972
rect 338628 319970 338634 319972
rect 343393 319970 343459 319973
rect 338628 319968 343459 319970
rect 338628 319912 343398 319968
rect 343454 319912 343459 319968
rect 338628 319910 343459 319912
rect 338628 319908 338634 319910
rect 343393 319907 343459 319910
rect 385529 319156 385595 319157
rect 385478 319154 385484 319156
rect 385438 319094 385484 319154
rect 385548 319152 385595 319156
rect 385590 319096 385595 319152
rect 385478 319092 385484 319094
rect 385548 319092 385595 319096
rect 385529 319091 385595 319092
rect 242193 319018 242259 319021
rect 242193 319016 242394 319018
rect 242193 318960 242198 319016
rect 242254 318960 242394 319016
rect 242193 318958 242394 318960
rect 242193 318955 242259 318958
rect 242193 318882 242259 318885
rect 242334 318882 242394 318958
rect 385529 318884 385595 318885
rect 242193 318880 242394 318882
rect 242193 318824 242198 318880
rect 242254 318824 242394 318880
rect 242193 318822 242394 318824
rect 242193 318819 242259 318822
rect 385478 318820 385484 318884
rect 385548 318882 385595 318884
rect 385548 318880 385640 318882
rect 385590 318824 385640 318880
rect 385548 318822 385640 318824
rect 385548 318820 385595 318822
rect 385529 318819 385595 318820
rect 319013 318746 319079 318749
rect 318694 318744 319079 318746
rect 318694 318688 319018 318744
rect 319074 318688 319079 318744
rect 318694 318686 319079 318688
rect 318694 318474 318754 318686
rect 319013 318683 319079 318686
rect 318921 318474 318987 318477
rect 318694 318472 318987 318474
rect 318694 318416 318926 318472
rect 318982 318416 318987 318472
rect 318694 318414 318987 318416
rect 318921 318411 318987 318414
rect 496 310042 976 310072
rect 3637 310042 3703 310045
rect 496 310040 3703 310042
rect 496 309984 3642 310040
rect 3698 309984 3703 310040
rect 496 309982 3703 309984
rect 496 309952 976 309982
rect 3637 309979 3703 309982
rect 278717 306370 278783 306373
rect 278901 306370 278967 306373
rect 278717 306368 278967 306370
rect 278717 306312 278722 306368
rect 278778 306312 278906 306368
rect 278962 306312 278967 306368
rect 278717 306310 278967 306312
rect 278717 306307 278783 306310
rect 278901 306307 278967 306310
rect 252814 304948 252820 305012
rect 252884 305010 252890 305012
rect 584016 305010 584496 305040
rect 252884 304950 584496 305010
rect 252884 304948 252890 304950
rect 584016 304920 584496 304950
rect 372925 298210 372991 298213
rect 373109 298210 373175 298213
rect 372925 298208 373175 298210
rect 372925 298152 372930 298208
rect 372986 298152 373114 298208
rect 373170 298152 373175 298208
rect 372925 298150 373175 298152
rect 372925 298147 372991 298150
rect 373109 298147 373175 298150
rect 135473 298074 135539 298077
rect 135657 298074 135723 298077
rect 135473 298072 135723 298074
rect 135473 298016 135478 298072
rect 135534 298016 135662 298072
rect 135718 298016 135723 298072
rect 135473 298014 135723 298016
rect 135473 298011 135539 298014
rect 135657 298011 135723 298014
rect 152033 298074 152099 298077
rect 152217 298074 152283 298077
rect 152033 298072 152283 298074
rect 152033 298016 152038 298072
rect 152094 298016 152222 298072
rect 152278 298016 152283 298072
rect 152033 298014 152283 298016
rect 152033 298011 152099 298014
rect 152217 298011 152283 298014
rect 170157 298074 170223 298077
rect 170341 298074 170407 298077
rect 170157 298072 170407 298074
rect 170157 298016 170162 298072
rect 170218 298016 170346 298072
rect 170402 298016 170407 298072
rect 170157 298014 170407 298016
rect 170157 298011 170223 298014
rect 170341 298011 170407 298014
rect 190673 298074 190739 298077
rect 190857 298074 190923 298077
rect 190673 298072 190923 298074
rect 190673 298016 190678 298072
rect 190734 298016 190862 298072
rect 190918 298016 190923 298072
rect 190673 298014 190923 298016
rect 190673 298011 190739 298014
rect 190857 298011 190923 298014
rect 214317 298074 214383 298077
rect 214501 298074 214567 298077
rect 214317 298072 214567 298074
rect 214317 298016 214322 298072
rect 214378 298016 214506 298072
rect 214562 298016 214567 298072
rect 214317 298014 214567 298016
rect 214317 298011 214383 298014
rect 214501 298011 214567 298014
rect 385529 298074 385595 298077
rect 385713 298074 385779 298077
rect 385529 298072 385779 298074
rect 385529 298016 385534 298072
rect 385590 298016 385718 298072
rect 385774 298016 385779 298072
rect 385529 298014 385779 298016
rect 385529 298011 385595 298014
rect 385713 298011 385779 298014
rect 392429 298074 392495 298077
rect 392613 298074 392679 298077
rect 392429 298072 392679 298074
rect 392429 298016 392434 298072
rect 392490 298016 392618 298072
rect 392674 298016 392679 298072
rect 392429 298014 392679 298016
rect 392429 298011 392495 298014
rect 392613 298011 392679 298014
rect 528865 298074 528931 298077
rect 529049 298074 529115 298077
rect 528865 298072 529115 298074
rect 528865 298016 528870 298072
rect 528926 298016 529054 298072
rect 529110 298016 529115 298072
rect 528865 298014 529115 298016
rect 528865 298011 528931 298014
rect 529049 298011 529115 298014
rect 372833 296714 372899 296717
rect 373017 296714 373083 296717
rect 372833 296712 373083 296714
rect 372833 296656 372838 296712
rect 372894 296656 373022 296712
rect 373078 296656 373083 296712
rect 372833 296654 373083 296656
rect 372833 296651 372899 296654
rect 373017 296651 373083 296654
rect 277245 295490 277311 295493
rect 276558 295488 277311 295490
rect 276558 295432 277250 295488
rect 277306 295432 277311 295488
rect 276558 295430 277311 295432
rect 276558 295357 276618 295430
rect 277245 295427 277311 295430
rect 273013 295354 273079 295357
rect 273197 295354 273263 295357
rect 273013 295352 273263 295354
rect 273013 295296 273018 295352
rect 273074 295296 273202 295352
rect 273258 295296 273263 295352
rect 273013 295294 273263 295296
rect 273013 295291 273079 295294
rect 273197 295291 273263 295294
rect 276509 295352 276618 295357
rect 276509 295296 276514 295352
rect 276570 295296 276618 295352
rect 276509 295294 276618 295296
rect 276693 295354 276759 295357
rect 276969 295354 277035 295357
rect 276693 295352 277035 295354
rect 276693 295296 276698 295352
rect 276754 295296 276974 295352
rect 277030 295296 277035 295352
rect 276693 295294 277035 295296
rect 276509 295291 276575 295294
rect 276693 295291 276759 295294
rect 276969 295291 277035 295294
rect 496 293314 976 293344
rect 3545 293314 3611 293317
rect 496 293312 3611 293314
rect 496 293256 3550 293312
rect 3606 293256 3611 293312
rect 496 293254 3611 293256
rect 496 293224 976 293254
rect 3545 293251 3611 293254
rect 341093 290188 341159 290189
rect 341093 290184 341140 290188
rect 341204 290186 341210 290188
rect 341093 290128 341098 290184
rect 341093 290124 341140 290128
rect 341204 290126 341250 290186
rect 341204 290124 341210 290126
rect 341093 290123 341159 290124
rect 341093 289916 341159 289917
rect 341093 289914 341140 289916
rect 341048 289912 341140 289914
rect 341048 289856 341098 289912
rect 341048 289854 341140 289856
rect 341093 289852 341140 289854
rect 341204 289852 341210 289916
rect 341093 289851 341159 289852
rect 580661 289370 580727 289373
rect 584016 289370 584496 289400
rect 580661 289368 584496 289370
rect 580661 289312 580666 289368
rect 580722 289312 584496 289368
rect 580661 289310 584496 289312
rect 580661 289307 580727 289310
rect 584016 289280 584496 289310
rect 328213 288554 328279 288557
rect 328397 288554 328463 288557
rect 328213 288552 328463 288554
rect 328213 288496 328218 288552
rect 328274 288496 328402 288552
rect 328458 288496 328463 288552
rect 328213 288494 328463 288496
rect 328213 288491 328279 288494
rect 328397 288491 328463 288494
rect 552417 288418 552483 288421
rect 552601 288418 552667 288421
rect 552417 288416 552667 288418
rect 552417 288360 552422 288416
rect 552478 288360 552606 288416
rect 552662 288360 552667 288416
rect 552417 288358 552667 288360
rect 552417 288355 552483 288358
rect 552601 288355 552667 288358
rect 246517 285834 246583 285837
rect 246517 285832 246626 285834
rect 246517 285776 246522 285832
rect 246578 285776 246626 285832
rect 246517 285771 246626 285776
rect 246566 285701 246626 285771
rect 246566 285696 246675 285701
rect 246566 285640 246614 285696
rect 246670 285640 246675 285696
rect 246566 285638 246675 285640
rect 246609 285635 246675 285638
rect 319974 282916 319980 282980
rect 320044 282978 320050 282980
rect 320117 282978 320183 282981
rect 320044 282976 320183 282978
rect 320044 282920 320122 282976
rect 320178 282920 320183 282976
rect 320044 282918 320183 282920
rect 320044 282916 320050 282918
rect 320117 282915 320183 282918
rect 320025 278900 320091 278901
rect 319974 278836 319980 278900
rect 320044 278898 320091 278900
rect 320044 278896 320136 278898
rect 320086 278840 320136 278896
rect 320044 278838 320136 278840
rect 320044 278836 320091 278838
rect 320025 278835 320091 278836
rect 135473 278762 135539 278765
rect 135657 278762 135723 278765
rect 135473 278760 135723 278762
rect 135473 278704 135478 278760
rect 135534 278704 135662 278760
rect 135718 278704 135723 278760
rect 135473 278702 135723 278704
rect 135473 278699 135539 278702
rect 135657 278699 135723 278702
rect 152033 278762 152099 278765
rect 152217 278762 152283 278765
rect 152033 278760 152283 278762
rect 152033 278704 152038 278760
rect 152094 278704 152222 278760
rect 152278 278704 152283 278760
rect 152033 278702 152283 278704
rect 152033 278699 152099 278702
rect 152217 278699 152283 278702
rect 170157 278762 170223 278765
rect 170341 278762 170407 278765
rect 170157 278760 170407 278762
rect 170157 278704 170162 278760
rect 170218 278704 170346 278760
rect 170402 278704 170407 278760
rect 170157 278702 170407 278704
rect 170157 278699 170223 278702
rect 170341 278699 170407 278702
rect 190673 278762 190739 278765
rect 190857 278762 190923 278765
rect 190673 278760 190923 278762
rect 190673 278704 190678 278760
rect 190734 278704 190862 278760
rect 190918 278704 190923 278760
rect 190673 278702 190923 278704
rect 190673 278699 190739 278702
rect 190857 278699 190923 278702
rect 214317 278762 214383 278765
rect 214501 278762 214567 278765
rect 214317 278760 214567 278762
rect 214317 278704 214322 278760
rect 214378 278704 214506 278760
rect 214562 278704 214567 278760
rect 214317 278702 214567 278704
rect 214317 278699 214383 278702
rect 214501 278699 214567 278702
rect 235385 278762 235451 278765
rect 235569 278762 235635 278765
rect 235385 278760 235635 278762
rect 235385 278704 235390 278760
rect 235446 278704 235574 278760
rect 235630 278704 235635 278760
rect 235385 278702 235635 278704
rect 235385 278699 235451 278702
rect 235569 278699 235635 278702
rect 279729 278762 279795 278765
rect 280005 278762 280071 278765
rect 279729 278760 280071 278762
rect 279729 278704 279734 278760
rect 279790 278704 280010 278760
rect 280066 278704 280071 278760
rect 279729 278702 280071 278704
rect 279729 278699 279795 278702
rect 280005 278699 280071 278702
rect 385529 278762 385595 278765
rect 385713 278762 385779 278765
rect 385529 278760 385779 278762
rect 385529 278704 385534 278760
rect 385590 278704 385718 278760
rect 385774 278704 385779 278760
rect 385529 278702 385779 278704
rect 385529 278699 385595 278702
rect 385713 278699 385779 278702
rect 392429 278762 392495 278765
rect 392613 278762 392679 278765
rect 392429 278760 392679 278762
rect 392429 278704 392434 278760
rect 392490 278704 392618 278760
rect 392674 278704 392679 278760
rect 392429 278702 392679 278704
rect 392429 278699 392495 278702
rect 392613 278699 392679 278702
rect 528865 278762 528931 278765
rect 529049 278762 529115 278765
rect 528865 278760 529115 278762
rect 528865 278704 528870 278760
rect 528926 278704 529054 278760
rect 529110 278704 529115 278760
rect 528865 278702 529115 278704
rect 528865 278699 528931 278702
rect 529049 278699 529115 278702
rect 552601 278762 552667 278765
rect 552785 278762 552851 278765
rect 552601 278760 552851 278762
rect 552601 278704 552606 278760
rect 552662 278704 552790 278760
rect 552846 278704 552851 278760
rect 552601 278702 552851 278704
rect 552601 278699 552667 278702
rect 552785 278699 552851 278702
rect 571829 278762 571895 278765
rect 572013 278762 572079 278765
rect 571829 278760 572079 278762
rect 571829 278704 571834 278760
rect 571890 278704 572018 278760
rect 572074 278704 572079 278760
rect 571829 278702 572079 278704
rect 571829 278699 571895 278702
rect 572013 278699 572079 278702
rect 278441 277538 278507 277541
rect 278625 277538 278691 277541
rect 278441 277536 278691 277538
rect 278441 277480 278446 277536
rect 278502 277480 278630 277536
rect 278686 277480 278691 277536
rect 278441 277478 278691 277480
rect 278441 277475 278507 277478
rect 278625 277475 278691 277478
rect 278441 277402 278507 277405
rect 278625 277402 278691 277405
rect 278441 277400 278691 277402
rect 278441 277344 278446 277400
rect 278502 277344 278630 277400
rect 278686 277344 278691 277400
rect 278441 277342 278691 277344
rect 278441 277339 278507 277342
rect 278625 277339 278691 277342
rect 496 276450 976 276480
rect 4281 276450 4347 276453
rect 496 276448 4347 276450
rect 496 276392 4286 276448
rect 4342 276392 4347 276448
rect 496 276390 4347 276392
rect 496 276360 976 276390
rect 4281 276387 4347 276390
rect 242653 276178 242719 276181
rect 242653 276176 242762 276178
rect 242653 276120 242658 276176
rect 242714 276120 242762 276176
rect 242653 276115 242762 276120
rect 242702 276045 242762 276115
rect 242702 276040 242811 276045
rect 242702 275984 242750 276040
rect 242806 275984 242811 276040
rect 242702 275982 242811 275984
rect 242745 275979 242811 275982
rect 272921 274818 272987 274821
rect 272878 274816 272987 274818
rect 272878 274760 272926 274816
rect 272982 274760 272987 274816
rect 272878 274755 272987 274760
rect 272878 274685 272938 274755
rect 272829 274680 272938 274685
rect 272829 274624 272834 274680
rect 272890 274624 272938 274680
rect 272829 274622 272938 274624
rect 272829 274619 272895 274622
rect 580661 273730 580727 273733
rect 584016 273730 584496 273760
rect 580661 273728 584496 273730
rect 580661 273672 580666 273728
rect 580722 273672 584496 273728
rect 580661 273670 584496 273672
rect 580661 273667 580727 273670
rect 584016 273640 584496 273670
rect 340909 270874 340975 270877
rect 340909 270872 341386 270874
rect 340909 270816 340914 270872
rect 340970 270816 341386 270872
rect 340909 270814 341386 270816
rect 340909 270811 340975 270814
rect 341185 270602 341251 270605
rect 341326 270602 341386 270814
rect 341185 270600 341386 270602
rect 341185 270544 341190 270600
rect 341246 270544 341386 270600
rect 341185 270542 341386 270544
rect 341185 270539 341251 270542
rect 278809 267746 278875 267749
rect 278993 267746 279059 267749
rect 278809 267744 279059 267746
rect 278809 267688 278814 267744
rect 278870 267688 278998 267744
rect 279054 267688 279059 267744
rect 278809 267686 279059 267688
rect 278809 267683 278875 267686
rect 278993 267683 279059 267686
rect 328213 266386 328279 266389
rect 328397 266386 328463 266389
rect 328213 266384 328463 266386
rect 328213 266328 328218 266384
rect 328274 266328 328402 266384
rect 328458 266328 328463 266384
rect 328213 266326 328463 266328
rect 328213 266323 328279 266326
rect 328397 266323 328463 266326
rect 272829 265026 272895 265029
rect 273013 265026 273079 265029
rect 272829 265024 273079 265026
rect 272829 264968 272834 265024
rect 272890 264968 273018 265024
rect 273074 264968 273079 265024
rect 272829 264966 273079 264968
rect 272829 264963 272895 264966
rect 273013 264963 273079 264966
rect 496 259722 976 259752
rect 3821 259722 3887 259725
rect 496 259720 3887 259722
rect 496 259664 3826 259720
rect 3882 259664 3887 259720
rect 496 259662 3887 259664
rect 496 259632 976 259662
rect 3821 259659 3887 259662
rect 135473 259450 135539 259453
rect 135657 259450 135723 259453
rect 135473 259448 135723 259450
rect 135473 259392 135478 259448
rect 135534 259392 135662 259448
rect 135718 259392 135723 259448
rect 135473 259390 135723 259392
rect 135473 259387 135539 259390
rect 135657 259387 135723 259390
rect 152033 259450 152099 259453
rect 152217 259450 152283 259453
rect 152033 259448 152283 259450
rect 152033 259392 152038 259448
rect 152094 259392 152222 259448
rect 152278 259392 152283 259448
rect 152033 259390 152283 259392
rect 152033 259387 152099 259390
rect 152217 259387 152283 259390
rect 170157 259450 170223 259453
rect 170341 259450 170407 259453
rect 170157 259448 170407 259450
rect 170157 259392 170162 259448
rect 170218 259392 170346 259448
rect 170402 259392 170407 259448
rect 170157 259390 170407 259392
rect 170157 259387 170223 259390
rect 170341 259387 170407 259390
rect 190673 259450 190739 259453
rect 190857 259450 190923 259453
rect 190673 259448 190923 259450
rect 190673 259392 190678 259448
rect 190734 259392 190862 259448
rect 190918 259392 190923 259448
rect 190673 259390 190923 259392
rect 190673 259387 190739 259390
rect 190857 259387 190923 259390
rect 214317 259450 214383 259453
rect 214501 259450 214567 259453
rect 214317 259448 214567 259450
rect 214317 259392 214322 259448
rect 214378 259392 214506 259448
rect 214562 259392 214567 259448
rect 214317 259390 214567 259392
rect 214317 259387 214383 259390
rect 214501 259387 214567 259390
rect 385529 259450 385595 259453
rect 385713 259450 385779 259453
rect 385529 259448 385779 259450
rect 385529 259392 385534 259448
rect 385590 259392 385718 259448
rect 385774 259392 385779 259448
rect 385529 259390 385779 259392
rect 385529 259387 385595 259390
rect 385713 259387 385779 259390
rect 392429 259450 392495 259453
rect 392613 259450 392679 259453
rect 392429 259448 392679 259450
rect 392429 259392 392434 259448
rect 392490 259392 392618 259448
rect 392674 259392 392679 259448
rect 392429 259390 392679 259392
rect 392429 259387 392495 259390
rect 392613 259387 392679 259390
rect 528865 259450 528931 259453
rect 529049 259450 529115 259453
rect 528865 259448 529115 259450
rect 528865 259392 528870 259448
rect 528926 259392 529054 259448
rect 529110 259392 529115 259448
rect 528865 259390 529115 259392
rect 528865 259387 528931 259390
rect 529049 259387 529115 259390
rect 535949 259450 536015 259453
rect 536133 259450 536199 259453
rect 535949 259448 536199 259450
rect 535949 259392 535954 259448
rect 536010 259392 536138 259448
rect 536194 259392 536199 259448
rect 535949 259390 536199 259392
rect 535949 259387 536015 259390
rect 536133 259387 536199 259390
rect 552509 259450 552575 259453
rect 552693 259450 552759 259453
rect 552509 259448 552759 259450
rect 552509 259392 552514 259448
rect 552570 259392 552698 259448
rect 552754 259392 552759 259448
rect 552509 259390 552759 259392
rect 552509 259387 552575 259390
rect 552693 259387 552759 259390
rect 571829 259450 571895 259453
rect 572013 259450 572079 259453
rect 571829 259448 572079 259450
rect 571829 259392 571834 259448
rect 571890 259392 572018 259448
rect 572074 259392 572079 259448
rect 571829 259390 572079 259392
rect 571829 259387 571895 259390
rect 572013 259387 572079 259390
rect 248766 258028 248772 258092
rect 248836 258090 248842 258092
rect 584016 258090 584496 258120
rect 248836 258030 584496 258090
rect 248836 258028 248842 258030
rect 584016 258000 584496 258030
rect 320025 251156 320091 251157
rect 319974 251154 319980 251156
rect 319934 251094 319980 251154
rect 320044 251152 320091 251156
rect 320086 251096 320091 251152
rect 319974 251092 319980 251094
rect 320044 251092 320091 251096
rect 320025 251091 320091 251092
rect 279453 249794 279519 249797
rect 279821 249794 279887 249797
rect 279453 249792 279887 249794
rect 279453 249736 279458 249792
rect 279514 249736 279826 249792
rect 279882 249736 279887 249792
rect 279453 249734 279887 249736
rect 279453 249731 279519 249734
rect 279821 249731 279887 249734
rect 235569 244356 235635 244357
rect 235518 244354 235524 244356
rect 235478 244294 235524 244354
rect 235588 244352 235635 244356
rect 235630 244296 235635 244352
rect 235518 244292 235524 244294
rect 235588 244292 235635 244296
rect 235569 244291 235635 244292
rect 496 242994 976 243024
rect 3821 242994 3887 242997
rect 496 242992 3887 242994
rect 496 242936 3826 242992
rect 3882 242936 3887 242992
rect 496 242934 3887 242936
rect 496 242904 976 242934
rect 3821 242931 3887 242934
rect 309629 242450 309695 242453
rect 319054 242450 319060 242452
rect 309629 242448 319060 242450
rect 309629 242392 309634 242448
rect 309690 242392 319060 242448
rect 309629 242390 319060 242392
rect 309629 242387 309695 242390
rect 319054 242388 319060 242390
rect 319124 242388 319130 242452
rect 584016 242450 584496 242480
rect 583838 242390 584496 242450
rect 377198 242116 377204 242180
rect 377268 242178 377274 242180
rect 384057 242178 384123 242181
rect 377268 242176 384123 242178
rect 377268 242120 384062 242176
rect 384118 242120 384123 242176
rect 377268 242118 384123 242120
rect 377268 242116 377274 242118
rect 384057 242115 384123 242118
rect 261145 242042 261211 242045
rect 261145 242040 264290 242042
rect 261145 241984 261150 242040
rect 261206 241984 264290 242040
rect 261145 241982 264290 241984
rect 261145 241979 261211 241982
rect 247294 241708 247300 241772
rect 247364 241770 247370 241772
rect 251669 241770 251735 241773
rect 247364 241768 251735 241770
rect 247364 241712 251674 241768
rect 251730 241712 251735 241768
rect 247364 241710 251735 241712
rect 264230 241770 264290 241982
rect 319054 241980 319060 242044
rect 319124 242042 319130 242044
rect 319124 241982 322250 242042
rect 319124 241980 319130 241982
rect 294817 241906 294883 241909
rect 299918 241906 299924 241908
rect 294817 241904 299924 241906
rect 294817 241848 294822 241904
rect 294878 241848 299924 241904
rect 294817 241846 299924 241848
rect 294817 241843 294883 241846
rect 299918 241844 299924 241846
rect 299988 241844 299994 241908
rect 289941 241770 290007 241773
rect 264230 241768 290007 241770
rect 264230 241712 289946 241768
rect 290002 241712 290007 241768
rect 264230 241710 290007 241712
rect 247364 241708 247370 241710
rect 251669 241707 251735 241710
rect 289941 241707 290007 241710
rect 300102 241708 300108 241772
rect 300172 241770 300178 241772
rect 309629 241770 309695 241773
rect 300172 241768 309695 241770
rect 300172 241712 309634 241768
rect 309690 241712 309695 241768
rect 300172 241710 309695 241712
rect 322190 241770 322250 241982
rect 384057 241906 384123 241909
rect 336542 241846 341386 241906
rect 336542 241770 336602 241846
rect 322190 241710 336602 241770
rect 300172 241708 300178 241710
rect 309629 241707 309695 241710
rect 235477 241636 235543 241637
rect 235477 241632 235524 241636
rect 235588 241634 235594 241636
rect 290033 241634 290099 241637
rect 290309 241634 290375 241637
rect 320025 241636 320091 241637
rect 235477 241576 235482 241632
rect 235477 241572 235524 241576
rect 235588 241574 235634 241634
rect 290033 241632 290375 241634
rect 290033 241576 290038 241632
rect 290094 241576 290314 241632
rect 290370 241576 290375 241632
rect 290033 241574 290375 241576
rect 235588 241572 235594 241574
rect 235477 241571 235543 241572
rect 290033 241571 290099 241574
rect 290309 241571 290375 241574
rect 319974 241572 319980 241636
rect 320044 241634 320091 241636
rect 341326 241634 341386 241846
rect 360462 241846 367514 241906
rect 360462 241770 360522 241846
rect 351078 241710 360522 241770
rect 367454 241770 367514 241846
rect 384057 241904 393826 241906
rect 384057 241848 384062 241904
rect 384118 241848 393826 241904
rect 384057 241846 393826 241848
rect 384057 241843 384123 241846
rect 377198 241770 377204 241772
rect 367454 241710 377204 241770
rect 351078 241634 351138 241710
rect 377198 241708 377204 241710
rect 377268 241708 377274 241772
rect 393766 241770 393826 241846
rect 403518 241846 413146 241906
rect 393766 241710 403394 241770
rect 320044 241632 320136 241634
rect 320086 241576 320136 241632
rect 320044 241574 320136 241576
rect 341326 241574 351138 241634
rect 403334 241634 403394 241710
rect 403518 241634 403578 241846
rect 413086 241770 413146 241846
rect 422838 241846 432466 241906
rect 413086 241710 422714 241770
rect 403334 241574 403578 241634
rect 422654 241634 422714 241710
rect 422838 241634 422898 241846
rect 432406 241770 432466 241846
rect 442158 241846 451786 241906
rect 432406 241710 442034 241770
rect 422654 241574 422898 241634
rect 441974 241634 442034 241710
rect 442158 241634 442218 241846
rect 451726 241770 451786 241846
rect 461478 241846 471106 241906
rect 451726 241710 461354 241770
rect 441974 241574 442218 241634
rect 461294 241634 461354 241710
rect 461478 241634 461538 241846
rect 471046 241770 471106 241846
rect 480798 241846 490426 241906
rect 471046 241710 480674 241770
rect 461294 241574 461538 241634
rect 480614 241634 480674 241710
rect 480798 241634 480858 241846
rect 490366 241770 490426 241846
rect 500118 241846 509746 241906
rect 490366 241710 499994 241770
rect 480614 241574 480858 241634
rect 499934 241634 499994 241710
rect 500118 241634 500178 241846
rect 509686 241770 509746 241846
rect 519438 241846 529066 241906
rect 509686 241710 519314 241770
rect 499934 241574 500178 241634
rect 519254 241634 519314 241710
rect 519438 241634 519498 241846
rect 529006 241770 529066 241846
rect 538758 241846 544338 241906
rect 529006 241710 538634 241770
rect 519254 241574 519498 241634
rect 538574 241634 538634 241710
rect 538758 241634 538818 241846
rect 538574 241574 538818 241634
rect 544278 241634 544338 241846
rect 551078 241844 551084 241908
rect 551148 241906 551154 241908
rect 551148 241846 567706 241906
rect 551148 241844 551154 241846
rect 567646 241770 567706 241846
rect 583838 241770 583898 242390
rect 584016 242360 584496 242390
rect 567646 241710 577274 241770
rect 551078 241634 551084 241636
rect 544278 241574 551084 241634
rect 320044 241572 320091 241574
rect 551078 241572 551084 241574
rect 551148 241572 551154 241636
rect 552509 241634 552575 241637
rect 552693 241634 552759 241637
rect 552509 241632 552759 241634
rect 552509 241576 552514 241632
rect 552570 241576 552698 241632
rect 552754 241576 552759 241632
rect 552509 241574 552759 241576
rect 577214 241634 577274 241710
rect 577398 241710 583898 241770
rect 577398 241634 577458 241710
rect 577214 241574 577458 241634
rect 320025 241571 320091 241572
rect 552509 241571 552575 241574
rect 552693 241571 552759 241574
rect 331065 241498 331131 241501
rect 331249 241498 331315 241501
rect 331065 241496 331315 241498
rect 331065 241440 331070 241496
rect 331126 241440 331254 241496
rect 331310 241440 331315 241496
rect 331065 241438 331315 241440
rect 331065 241435 331131 241438
rect 331249 241435 331315 241438
rect 135473 240138 135539 240141
rect 135657 240138 135723 240141
rect 135473 240136 135723 240138
rect 135473 240080 135478 240136
rect 135534 240080 135662 240136
rect 135718 240080 135723 240136
rect 135473 240078 135723 240080
rect 135473 240075 135539 240078
rect 135657 240075 135723 240078
rect 152033 240138 152099 240141
rect 152217 240138 152283 240141
rect 152033 240136 152283 240138
rect 152033 240080 152038 240136
rect 152094 240080 152222 240136
rect 152278 240080 152283 240136
rect 152033 240078 152283 240080
rect 152033 240075 152099 240078
rect 152217 240075 152283 240078
rect 170157 240138 170223 240141
rect 170341 240138 170407 240141
rect 170157 240136 170407 240138
rect 170157 240080 170162 240136
rect 170218 240080 170346 240136
rect 170402 240080 170407 240136
rect 170157 240078 170407 240080
rect 170157 240075 170223 240078
rect 170341 240075 170407 240078
rect 190673 240138 190739 240141
rect 190857 240138 190923 240141
rect 190673 240136 190923 240138
rect 190673 240080 190678 240136
rect 190734 240080 190862 240136
rect 190918 240080 190923 240136
rect 190673 240078 190923 240080
rect 190673 240075 190739 240078
rect 190857 240075 190923 240078
rect 214317 240138 214383 240141
rect 214501 240138 214567 240141
rect 214317 240136 214567 240138
rect 214317 240080 214322 240136
rect 214378 240080 214506 240136
rect 214562 240080 214567 240136
rect 214317 240078 214567 240080
rect 214317 240075 214383 240078
rect 214501 240075 214567 240078
rect 385529 240138 385595 240141
rect 385713 240138 385779 240141
rect 385529 240136 385779 240138
rect 385529 240080 385534 240136
rect 385590 240080 385718 240136
rect 385774 240080 385779 240136
rect 385529 240078 385779 240080
rect 385529 240075 385595 240078
rect 385713 240075 385779 240078
rect 392429 240138 392495 240141
rect 392613 240138 392679 240141
rect 392429 240136 392679 240138
rect 392429 240080 392434 240136
rect 392490 240080 392618 240136
rect 392674 240080 392679 240136
rect 392429 240078 392679 240080
rect 392429 240075 392495 240078
rect 392613 240075 392679 240078
rect 528865 240138 528931 240141
rect 529049 240138 529115 240141
rect 528865 240136 529115 240138
rect 528865 240080 528870 240136
rect 528926 240080 529054 240136
rect 529110 240080 529115 240136
rect 528865 240078 529115 240080
rect 528865 240075 528931 240078
rect 529049 240075 529115 240078
rect 535949 240138 536015 240141
rect 536133 240138 536199 240141
rect 535949 240136 536199 240138
rect 535949 240080 535954 240136
rect 536010 240080 536138 240136
rect 536194 240080 536199 240136
rect 535949 240078 536199 240080
rect 535949 240075 536015 240078
rect 536133 240075 536199 240078
rect 571829 240138 571895 240141
rect 572013 240138 572079 240141
rect 571829 240136 572079 240138
rect 571829 240080 571834 240136
rect 571890 240080 572018 240136
rect 572074 240080 572079 240136
rect 571829 240078 572079 240080
rect 571829 240075 571895 240078
rect 572013 240075 572079 240078
rect 91313 231842 91379 231845
rect 91497 231842 91563 231845
rect 91313 231840 91563 231842
rect 91313 231784 91318 231840
rect 91374 231784 91502 231840
rect 91558 231784 91563 231840
rect 91313 231782 91563 231784
rect 91313 231779 91379 231782
rect 91497 231779 91563 231782
rect 357929 231842 357995 231845
rect 358113 231842 358179 231845
rect 357929 231840 358179 231842
rect 357929 231784 357934 231840
rect 357990 231784 358118 231840
rect 358174 231784 358179 231840
rect 357929 231782 358179 231784
rect 357929 231779 357995 231782
rect 358113 231779 358179 231782
rect 371545 231842 371611 231845
rect 371729 231842 371795 231845
rect 371545 231840 371795 231842
rect 371545 231784 371550 231840
rect 371606 231784 371734 231840
rect 371790 231784 371795 231840
rect 371545 231782 371795 231784
rect 371545 231779 371611 231782
rect 371729 231779 371795 231782
rect 373109 231842 373175 231845
rect 373293 231842 373359 231845
rect 373109 231840 373359 231842
rect 373109 231784 373114 231840
rect 373170 231784 373298 231840
rect 373354 231784 373359 231840
rect 373109 231782 373359 231784
rect 373109 231779 373175 231782
rect 373293 231779 373359 231782
rect 553705 231842 553771 231845
rect 553889 231842 553955 231845
rect 553705 231840 553955 231842
rect 553705 231784 553710 231840
rect 553766 231784 553894 231840
rect 553950 231784 553955 231840
rect 553705 231782 553955 231784
rect 553705 231779 553771 231782
rect 553889 231779 553955 231782
rect 304937 230482 305003 230485
rect 305121 230482 305187 230485
rect 304937 230480 305187 230482
rect 304937 230424 304942 230480
rect 304998 230424 305126 230480
rect 305182 230424 305187 230480
rect 304937 230422 305187 230424
rect 304937 230419 305003 230422
rect 305121 230419 305187 230422
rect 276785 227898 276851 227901
rect 276742 227896 276851 227898
rect 276742 227840 276790 227896
rect 276846 227840 276851 227896
rect 276742 227835 276851 227840
rect 276742 227765 276802 227835
rect 276742 227760 276851 227765
rect 276742 227704 276790 227760
rect 276846 227704 276851 227760
rect 276742 227702 276851 227704
rect 276785 227699 276851 227702
rect 276969 227762 277035 227765
rect 277245 227762 277311 227765
rect 276969 227760 277311 227762
rect 276969 227704 276974 227760
rect 277030 227704 277250 227760
rect 277306 227704 277311 227760
rect 276969 227702 277311 227704
rect 276969 227699 277035 227702
rect 277245 227699 277311 227702
rect 309629 227218 309695 227221
rect 319054 227218 319060 227220
rect 309629 227216 319060 227218
rect 309629 227160 309634 227216
rect 309690 227160 319060 227216
rect 309629 227158 319060 227160
rect 309629 227155 309695 227158
rect 319054 227156 319060 227158
rect 319124 227156 319130 227220
rect 319054 226748 319060 226812
rect 319124 226810 319130 226812
rect 584016 226810 584496 226840
rect 319124 226750 322250 226810
rect 319124 226748 319130 226750
rect 244534 226612 244540 226676
rect 244604 226674 244610 226676
rect 270897 226674 270963 226677
rect 244604 226614 254538 226674
rect 244604 226612 244610 226614
rect 254478 226538 254538 226614
rect 270897 226672 283426 226674
rect 270897 226616 270902 226672
rect 270958 226616 283426 226672
rect 270897 226614 283426 226616
rect 270897 226611 270963 226614
rect 261278 226538 261284 226540
rect 254478 226478 261284 226538
rect 261278 226476 261284 226478
rect 261348 226476 261354 226540
rect 283366 226402 283426 226614
rect 288878 226612 288884 226676
rect 288948 226674 288954 226676
rect 300429 226674 300495 226677
rect 288948 226672 300495 226674
rect 288948 226616 300434 226672
rect 300490 226616 300495 226672
rect 288948 226614 300495 226616
rect 288948 226612 288954 226614
rect 300429 226611 300495 226614
rect 308157 226538 308223 226541
rect 309629 226538 309695 226541
rect 308157 226536 309695 226538
rect 308157 226480 308162 226536
rect 308218 226480 309634 226536
rect 309690 226480 309695 226536
rect 308157 226478 309695 226480
rect 322190 226538 322250 226750
rect 583838 226750 584496 226810
rect 336542 226614 341386 226674
rect 336542 226538 336602 226614
rect 322190 226478 336602 226538
rect 308157 226475 308223 226478
rect 309629 226475 309695 226478
rect 288878 226402 288884 226404
rect 283366 226342 288884 226402
rect 288878 226340 288884 226342
rect 288948 226340 288954 226404
rect 341326 226402 341386 226614
rect 374446 226614 384074 226674
rect 360597 226538 360663 226541
rect 351078 226536 360663 226538
rect 351078 226480 360602 226536
rect 360658 226480 360663 226536
rect 351078 226478 360663 226480
rect 351078 226402 351138 226478
rect 360597 226475 360663 226478
rect 362253 226538 362319 226541
rect 362253 226536 370274 226538
rect 362253 226480 362258 226536
rect 362314 226480 370274 226536
rect 362253 226478 370274 226480
rect 362253 226475 362319 226478
rect 341326 226342 351138 226402
rect 370214 226402 370274 226478
rect 374446 226402 374506 226614
rect 370214 226342 374506 226402
rect 384014 226402 384074 226614
rect 384198 226614 393826 226674
rect 384198 226402 384258 226614
rect 393766 226538 393826 226614
rect 403518 226614 413146 226674
rect 393766 226478 403394 226538
rect 384014 226342 384258 226402
rect 403334 226402 403394 226478
rect 403518 226402 403578 226614
rect 413086 226538 413146 226614
rect 422838 226614 432466 226674
rect 413086 226478 422714 226538
rect 403334 226342 403578 226402
rect 422654 226402 422714 226478
rect 422838 226402 422898 226614
rect 432406 226538 432466 226614
rect 442158 226614 451786 226674
rect 432406 226478 442034 226538
rect 422654 226342 422898 226402
rect 441974 226402 442034 226478
rect 442158 226402 442218 226614
rect 451726 226538 451786 226614
rect 461478 226614 471106 226674
rect 451726 226478 461354 226538
rect 441974 226342 442218 226402
rect 461294 226402 461354 226478
rect 461478 226402 461538 226614
rect 471046 226538 471106 226614
rect 480798 226614 490426 226674
rect 471046 226478 480674 226538
rect 461294 226342 461538 226402
rect 480614 226402 480674 226478
rect 480798 226402 480858 226614
rect 490366 226538 490426 226614
rect 500118 226614 509746 226674
rect 490366 226478 499994 226538
rect 480614 226342 480858 226402
rect 499934 226402 499994 226478
rect 500118 226402 500178 226614
rect 509686 226538 509746 226614
rect 519438 226614 529066 226674
rect 509686 226478 519314 226538
rect 499934 226342 500178 226402
rect 519254 226402 519314 226478
rect 519438 226402 519498 226614
rect 529006 226538 529066 226614
rect 538758 226614 544338 226674
rect 529006 226478 538634 226538
rect 519254 226342 519498 226402
rect 538574 226402 538634 226478
rect 538758 226402 538818 226614
rect 538574 226342 538818 226402
rect 544278 226402 544338 226614
rect 551078 226612 551084 226676
rect 551148 226674 551154 226676
rect 551148 226614 567706 226674
rect 551148 226612 551154 226614
rect 567646 226538 567706 226614
rect 583838 226538 583898 226750
rect 584016 226720 584496 226750
rect 567646 226478 577274 226538
rect 551078 226402 551084 226404
rect 544278 226342 551084 226402
rect 551078 226340 551084 226342
rect 551148 226340 551154 226404
rect 577214 226402 577274 226478
rect 577398 226478 583898 226538
rect 577398 226402 577458 226478
rect 577214 226342 577458 226402
rect 496 226266 976 226296
rect 4189 226266 4255 226269
rect 496 226264 4255 226266
rect 496 226208 4194 226264
rect 4250 226208 4255 226264
rect 496 226206 4255 226208
rect 496 226176 976 226206
rect 4189 226203 4255 226206
rect 261278 226204 261284 226268
rect 261348 226266 261354 226268
rect 270897 226266 270963 226269
rect 261348 226264 270963 226266
rect 261348 226208 270902 226264
rect 270958 226208 270963 226264
rect 261348 226206 270963 226208
rect 261348 226204 261354 226206
rect 270897 226203 270963 226206
rect 331065 222186 331131 222189
rect 331249 222186 331315 222189
rect 331065 222184 331315 222186
rect 331065 222128 331070 222184
rect 331126 222128 331254 222184
rect 331310 222128 331315 222184
rect 331065 222126 331315 222128
rect 331065 222123 331131 222126
rect 331249 222123 331315 222126
rect 553705 222186 553771 222189
rect 553889 222186 553955 222189
rect 553705 222184 553955 222186
rect 553705 222128 553710 222184
rect 553766 222128 553894 222184
rect 553950 222128 553955 222184
rect 553705 222126 553955 222128
rect 553705 222123 553771 222126
rect 553889 222123 553955 222126
rect 276509 221508 276575 221509
rect 276509 221506 276556 221508
rect 276464 221504 276556 221506
rect 276464 221448 276514 221504
rect 276464 221446 276556 221448
rect 276509 221444 276556 221446
rect 276620 221444 276626 221508
rect 276509 221443 276575 221444
rect 235661 221098 235727 221101
rect 235526 221096 235727 221098
rect 235526 221040 235666 221096
rect 235722 221040 235727 221096
rect 235526 221038 235727 221040
rect 235526 220965 235586 221038
rect 235661 221035 235727 221038
rect 235526 220960 235635 220965
rect 235526 220904 235574 220960
rect 235630 220904 235635 220960
rect 235526 220902 235635 220904
rect 235569 220899 235635 220902
rect 135473 220826 135539 220829
rect 135657 220826 135723 220829
rect 135473 220824 135723 220826
rect 135473 220768 135478 220824
rect 135534 220768 135662 220824
rect 135718 220768 135723 220824
rect 135473 220766 135723 220768
rect 135473 220763 135539 220766
rect 135657 220763 135723 220766
rect 152033 220826 152099 220829
rect 152217 220826 152283 220829
rect 152033 220824 152283 220826
rect 152033 220768 152038 220824
rect 152094 220768 152222 220824
rect 152278 220768 152283 220824
rect 152033 220766 152283 220768
rect 152033 220763 152099 220766
rect 152217 220763 152283 220766
rect 170157 220826 170223 220829
rect 170341 220826 170407 220829
rect 170157 220824 170407 220826
rect 170157 220768 170162 220824
rect 170218 220768 170346 220824
rect 170402 220768 170407 220824
rect 170157 220766 170407 220768
rect 170157 220763 170223 220766
rect 170341 220763 170407 220766
rect 190673 220826 190739 220829
rect 190857 220826 190923 220829
rect 190673 220824 190923 220826
rect 190673 220768 190678 220824
rect 190734 220768 190862 220824
rect 190918 220768 190923 220824
rect 190673 220766 190923 220768
rect 190673 220763 190739 220766
rect 190857 220763 190923 220766
rect 214317 220826 214383 220829
rect 214501 220826 214567 220829
rect 214317 220824 214567 220826
rect 214317 220768 214322 220824
rect 214378 220768 214506 220824
rect 214562 220768 214567 220824
rect 214317 220766 214567 220768
rect 214317 220763 214383 220766
rect 214501 220763 214567 220766
rect 235385 220826 235451 220829
rect 235569 220826 235635 220829
rect 235385 220824 235635 220826
rect 235385 220768 235390 220824
rect 235446 220768 235574 220824
rect 235630 220768 235635 220824
rect 235385 220766 235635 220768
rect 235385 220763 235451 220766
rect 235569 220763 235635 220766
rect 385529 220826 385595 220829
rect 385713 220826 385779 220829
rect 385529 220824 385779 220826
rect 385529 220768 385534 220824
rect 385590 220768 385718 220824
rect 385774 220768 385779 220824
rect 385529 220766 385779 220768
rect 385529 220763 385595 220766
rect 385713 220763 385779 220766
rect 392429 220826 392495 220829
rect 392613 220826 392679 220829
rect 392429 220824 392679 220826
rect 392429 220768 392434 220824
rect 392490 220768 392618 220824
rect 392674 220768 392679 220824
rect 392429 220766 392679 220768
rect 392429 220763 392495 220766
rect 392613 220763 392679 220766
rect 528865 220826 528931 220829
rect 529049 220826 529115 220829
rect 528865 220824 529115 220826
rect 528865 220768 528870 220824
rect 528926 220768 529054 220824
rect 529110 220768 529115 220824
rect 528865 220766 529115 220768
rect 528865 220763 528931 220766
rect 529049 220763 529115 220766
rect 535949 220826 536015 220829
rect 536133 220826 536199 220829
rect 535949 220824 536199 220826
rect 535949 220768 535954 220824
rect 536010 220768 536138 220824
rect 536194 220768 536199 220824
rect 535949 220766 536199 220768
rect 535949 220763 536015 220766
rect 536133 220763 536199 220766
rect 571829 220826 571895 220829
rect 572013 220826 572079 220829
rect 571829 220824 572079 220826
rect 571829 220768 571834 220824
rect 571890 220768 572018 220824
rect 572074 220768 572079 220824
rect 571829 220766 572079 220768
rect 571829 220763 571895 220766
rect 572013 220763 572079 220766
rect 242837 218242 242903 218245
rect 242334 218240 242903 218242
rect 242334 218184 242842 218240
rect 242898 218184 242903 218240
rect 242334 218182 242903 218184
rect 242334 218106 242394 218182
rect 242837 218179 242903 218182
rect 242469 218106 242535 218109
rect 242334 218104 242535 218106
rect 242334 218048 242474 218104
rect 242530 218048 242535 218104
rect 242334 218046 242535 218048
rect 242469 218043 242535 218046
rect 320025 216068 320091 216069
rect 319974 216066 319980 216068
rect 319934 216006 319980 216066
rect 320044 216064 320091 216068
rect 320086 216008 320091 216064
rect 319974 216004 319980 216006
rect 320044 216004 320091 216008
rect 320025 216003 320091 216004
rect 91313 212530 91379 212533
rect 91497 212530 91563 212533
rect 91313 212528 91563 212530
rect 91313 212472 91318 212528
rect 91374 212472 91502 212528
rect 91558 212472 91563 212528
rect 91313 212470 91563 212472
rect 91313 212467 91379 212470
rect 91497 212467 91563 212470
rect 225357 212530 225423 212533
rect 225541 212530 225607 212533
rect 225357 212528 225607 212530
rect 225357 212472 225362 212528
rect 225418 212472 225546 212528
rect 225602 212472 225607 212528
rect 225357 212470 225607 212472
rect 225357 212467 225423 212470
rect 225541 212467 225607 212470
rect 135473 211170 135539 211173
rect 135657 211170 135723 211173
rect 135473 211168 135723 211170
rect 135473 211112 135478 211168
rect 135534 211112 135662 211168
rect 135718 211112 135723 211168
rect 135473 211110 135723 211112
rect 135473 211107 135539 211110
rect 135657 211107 135723 211110
rect 152033 211170 152099 211173
rect 152217 211170 152283 211173
rect 152033 211168 152283 211170
rect 152033 211112 152038 211168
rect 152094 211112 152222 211168
rect 152278 211112 152283 211168
rect 152033 211110 152283 211112
rect 152033 211107 152099 211110
rect 152217 211107 152283 211110
rect 170157 211170 170223 211173
rect 170341 211170 170407 211173
rect 170157 211168 170407 211170
rect 170157 211112 170162 211168
rect 170218 211112 170346 211168
rect 170402 211112 170407 211168
rect 170157 211110 170407 211112
rect 170157 211107 170223 211110
rect 170341 211107 170407 211110
rect 190673 211170 190739 211173
rect 190857 211170 190923 211173
rect 190673 211168 190923 211170
rect 190673 211112 190678 211168
rect 190734 211112 190862 211168
rect 190918 211112 190923 211168
rect 190673 211110 190923 211112
rect 190673 211107 190739 211110
rect 190857 211107 190923 211110
rect 214317 211170 214383 211173
rect 214501 211170 214567 211173
rect 214317 211168 214567 211170
rect 214317 211112 214322 211168
rect 214378 211112 214506 211168
rect 214562 211112 214567 211168
rect 214317 211110 214567 211112
rect 214317 211107 214383 211110
rect 214501 211107 214567 211110
rect 246006 211108 246012 211172
rect 246076 211170 246082 211172
rect 584016 211170 584496 211200
rect 246076 211110 584496 211170
rect 246076 211108 246082 211110
rect 584016 211080 584496 211110
rect 496 209402 976 209432
rect 3729 209402 3795 209405
rect 496 209400 3795 209402
rect 496 209344 3734 209400
rect 3790 209344 3795 209400
rect 496 209342 3795 209344
rect 496 209312 976 209342
rect 3729 209339 3795 209342
rect 276509 208452 276575 208453
rect 276509 208448 276556 208452
rect 276620 208450 276626 208452
rect 276509 208392 276514 208448
rect 276509 208388 276556 208392
rect 276620 208390 276666 208450
rect 276620 208388 276626 208390
rect 276509 208387 276575 208388
rect 320025 206276 320091 206277
rect 319974 206274 319980 206276
rect 319934 206214 319980 206274
rect 320044 206272 320091 206276
rect 320086 206216 320091 206272
rect 319974 206212 319980 206214
rect 320044 206212 320091 206216
rect 320025 206211 320091 206212
rect 331065 202874 331131 202877
rect 331249 202874 331315 202877
rect 331065 202872 331315 202874
rect 331065 202816 331070 202872
rect 331126 202816 331254 202872
rect 331310 202816 331315 202872
rect 331065 202814 331315 202816
rect 331065 202811 331131 202814
rect 331249 202811 331315 202814
rect 553705 202874 553771 202877
rect 553889 202874 553955 202877
rect 553705 202872 553955 202874
rect 553705 202816 553710 202872
rect 553766 202816 553894 202872
rect 553950 202816 553955 202872
rect 553705 202814 553955 202816
rect 553705 202811 553771 202814
rect 553889 202811 553955 202814
rect 552509 201650 552575 201653
rect 552374 201648 552575 201650
rect 552374 201592 552514 201648
rect 552570 201592 552575 201648
rect 552374 201590 552575 201592
rect 552374 201517 552434 201590
rect 552509 201587 552575 201590
rect 552374 201512 552483 201517
rect 552374 201456 552422 201512
rect 552478 201456 552483 201512
rect 552374 201454 552483 201456
rect 552417 201451 552483 201454
rect 246333 198794 246399 198797
rect 246333 198792 246626 198794
rect 246333 198736 246338 198792
rect 246394 198736 246626 198792
rect 246333 198734 246626 198736
rect 246333 198731 246399 198734
rect 246425 198522 246491 198525
rect 246566 198522 246626 198734
rect 246425 198520 246626 198522
rect 246425 198464 246430 198520
rect 246486 198464 246626 198520
rect 246425 198462 246626 198464
rect 246425 198459 246491 198462
rect 580661 195530 580727 195533
rect 584016 195530 584496 195560
rect 580661 195528 584496 195530
rect 580661 195472 580666 195528
rect 580722 195472 584496 195528
rect 580661 195470 584496 195472
rect 580661 195467 580727 195470
rect 584016 195440 584496 195470
rect 91313 193218 91379 193221
rect 91497 193218 91563 193221
rect 91313 193216 91563 193218
rect 91313 193160 91318 193216
rect 91374 193160 91502 193216
rect 91558 193160 91563 193216
rect 91313 193158 91563 193160
rect 91313 193155 91379 193158
rect 91497 193155 91563 193158
rect 357929 193218 357995 193221
rect 358113 193218 358179 193221
rect 357929 193216 358179 193218
rect 357929 193160 357934 193216
rect 357990 193160 358118 193216
rect 358174 193160 358179 193216
rect 357929 193158 358179 193160
rect 357929 193155 357995 193158
rect 358113 193155 358179 193158
rect 553705 193218 553771 193221
rect 553889 193218 553955 193221
rect 553705 193216 553955 193218
rect 553705 193160 553710 193216
rect 553766 193160 553894 193216
rect 553950 193160 553955 193216
rect 553705 193158 553955 193160
rect 553705 193155 553771 193158
rect 553889 193155 553955 193158
rect 496 192674 976 192704
rect 3821 192674 3887 192677
rect 496 192672 3887 192674
rect 496 192616 3826 192672
rect 3882 192616 3887 192672
rect 496 192614 3887 192616
rect 496 192584 976 192614
rect 3821 192611 3887 192614
rect 135473 191858 135539 191861
rect 135657 191858 135723 191861
rect 135473 191856 135723 191858
rect 135473 191800 135478 191856
rect 135534 191800 135662 191856
rect 135718 191800 135723 191856
rect 135473 191798 135723 191800
rect 135473 191795 135539 191798
rect 135657 191795 135723 191798
rect 152033 191858 152099 191861
rect 152217 191858 152283 191861
rect 152033 191856 152283 191858
rect 152033 191800 152038 191856
rect 152094 191800 152222 191856
rect 152278 191800 152283 191856
rect 152033 191798 152283 191800
rect 152033 191795 152099 191798
rect 152217 191795 152283 191798
rect 170157 191858 170223 191861
rect 170341 191858 170407 191861
rect 170157 191856 170407 191858
rect 170157 191800 170162 191856
rect 170218 191800 170346 191856
rect 170402 191800 170407 191856
rect 170157 191798 170407 191800
rect 170157 191795 170223 191798
rect 170341 191795 170407 191798
rect 190673 191858 190739 191861
rect 190857 191858 190923 191861
rect 190673 191856 190923 191858
rect 190673 191800 190678 191856
rect 190734 191800 190862 191856
rect 190918 191800 190923 191856
rect 190673 191798 190923 191800
rect 190673 191795 190739 191798
rect 190857 191795 190923 191798
rect 214317 191858 214383 191861
rect 214501 191858 214567 191861
rect 214317 191856 214567 191858
rect 214317 191800 214322 191856
rect 214378 191800 214506 191856
rect 214562 191800 214567 191856
rect 214317 191798 214567 191800
rect 214317 191795 214383 191798
rect 214501 191795 214567 191798
rect 268505 191858 268571 191861
rect 268689 191858 268755 191861
rect 268505 191856 268755 191858
rect 268505 191800 268510 191856
rect 268566 191800 268694 191856
rect 268750 191800 268755 191856
rect 268505 191798 268755 191800
rect 268505 191795 268571 191798
rect 268689 191795 268755 191798
rect 385529 191858 385595 191861
rect 385713 191858 385779 191861
rect 385529 191856 385779 191858
rect 385529 191800 385534 191856
rect 385590 191800 385718 191856
rect 385774 191800 385779 191856
rect 385529 191798 385779 191800
rect 385529 191795 385595 191798
rect 385713 191795 385779 191798
rect 392429 191858 392495 191861
rect 392613 191858 392679 191861
rect 392429 191856 392679 191858
rect 392429 191800 392434 191856
rect 392490 191800 392618 191856
rect 392674 191800 392679 191856
rect 392429 191798 392679 191800
rect 392429 191795 392495 191798
rect 392613 191795 392679 191798
rect 528865 191858 528931 191861
rect 529049 191858 529115 191861
rect 528865 191856 529115 191858
rect 528865 191800 528870 191856
rect 528926 191800 529054 191856
rect 529110 191800 529115 191856
rect 528865 191798 529115 191800
rect 528865 191795 528931 191798
rect 529049 191795 529115 191798
rect 535949 191858 536015 191861
rect 536133 191858 536199 191861
rect 535949 191856 536199 191858
rect 535949 191800 535954 191856
rect 536010 191800 536138 191856
rect 536194 191800 536199 191856
rect 535949 191798 536199 191800
rect 535949 191795 536015 191798
rect 536133 191795 536199 191798
rect 571829 191858 571895 191861
rect 572013 191858 572079 191861
rect 571829 191856 572079 191858
rect 571829 191800 571834 191856
rect 571890 191800 572018 191856
rect 572074 191800 572079 191856
rect 571829 191798 572079 191800
rect 571829 191795 571895 191798
rect 572013 191795 572079 191798
rect 275589 187914 275655 187917
rect 275589 187912 275882 187914
rect 275589 187856 275594 187912
rect 275650 187856 275882 187912
rect 275589 187854 275882 187856
rect 275589 187851 275655 187854
rect 275681 187778 275747 187781
rect 275822 187778 275882 187854
rect 275681 187776 275882 187778
rect 275681 187720 275686 187776
rect 275742 187720 275882 187776
rect 275681 187718 275882 187720
rect 275681 187715 275747 187718
rect 268505 183562 268571 183565
rect 268689 183562 268755 183565
rect 268505 183560 268755 183562
rect 268505 183504 268510 183560
rect 268566 183504 268694 183560
rect 268750 183504 268755 183560
rect 268505 183502 268755 183504
rect 268505 183499 268571 183502
rect 268689 183499 268755 183502
rect 331065 183562 331131 183565
rect 331249 183562 331315 183565
rect 553889 183564 553955 183565
rect 553838 183562 553844 183564
rect 331065 183560 331315 183562
rect 331065 183504 331070 183560
rect 331126 183504 331254 183560
rect 331310 183504 331315 183560
rect 331065 183502 331315 183504
rect 553798 183502 553844 183562
rect 553908 183560 553955 183564
rect 553950 183504 553955 183560
rect 331065 183499 331131 183502
rect 331249 183499 331315 183502
rect 553838 183500 553844 183502
rect 553908 183500 553955 183504
rect 553889 183499 553955 183500
rect 235569 182202 235635 182205
rect 235753 182202 235819 182205
rect 235569 182200 235819 182202
rect 235569 182144 235574 182200
rect 235630 182144 235758 182200
rect 235814 182144 235819 182200
rect 235569 182142 235819 182144
rect 235569 182139 235635 182142
rect 235753 182139 235819 182142
rect 242469 182202 242535 182205
rect 242469 182200 242762 182202
rect 242469 182144 242474 182200
rect 242530 182144 242762 182200
rect 242469 182142 242762 182144
rect 242469 182139 242535 182142
rect 242510 182004 242516 182068
rect 242580 182066 242586 182068
rect 242702 182066 242762 182142
rect 242580 182006 242762 182066
rect 242580 182004 242586 182006
rect 288878 179964 288884 180028
rect 288948 180026 288954 180028
rect 293621 180026 293687 180029
rect 288948 180024 293687 180026
rect 288948 179968 293626 180024
rect 293682 179968 293687 180024
rect 288948 179966 293687 179968
rect 288948 179964 288954 179966
rect 293621 179963 293687 179966
rect 391693 179890 391759 179893
rect 584016 179890 584496 179920
rect 386958 179888 391759 179890
rect 386958 179832 391698 179888
rect 391754 179832 391759 179888
rect 386958 179830 391759 179832
rect 261145 179754 261211 179757
rect 261145 179752 264290 179754
rect 261145 179696 261150 179752
rect 261206 179696 264290 179752
rect 261145 179694 264290 179696
rect 261145 179691 261211 179694
rect 241774 179556 241780 179620
rect 241844 179618 241850 179620
rect 251669 179618 251735 179621
rect 241844 179616 251735 179618
rect 241844 179560 251674 179616
rect 251730 179560 251735 179616
rect 241844 179558 251735 179560
rect 241844 179556 241850 179558
rect 251669 179555 251735 179558
rect 264230 179482 264290 179694
rect 269558 179692 269564 179756
rect 269628 179754 269634 179756
rect 288878 179754 288884 179756
rect 269628 179694 288884 179754
rect 269628 179692 269634 179694
rect 288878 179692 288884 179694
rect 288948 179692 288954 179756
rect 293621 179754 293687 179757
rect 293621 179752 298514 179754
rect 293621 179696 293626 179752
rect 293682 179696 298514 179752
rect 293621 179694 298514 179696
rect 293621 179691 293687 179694
rect 298454 179618 298514 179694
rect 327518 179692 327524 179756
rect 327588 179754 327594 179756
rect 356590 179754 356596 179756
rect 327588 179694 341386 179754
rect 327588 179692 327594 179694
rect 299918 179618 299924 179620
rect 298454 179558 299924 179618
rect 299918 179556 299924 179558
rect 299988 179556 299994 179620
rect 269558 179482 269564 179484
rect 264230 179422 269564 179482
rect 269558 179420 269564 179422
rect 269628 179420 269634 179484
rect 308198 179420 308204 179484
rect 308268 179482 308274 179484
rect 327518 179482 327524 179484
rect 308268 179422 327524 179482
rect 308268 179420 308274 179422
rect 327518 179420 327524 179422
rect 327588 179420 327594 179484
rect 341326 179482 341386 179694
rect 351262 179694 356596 179754
rect 351262 179618 351322 179694
rect 356590 179692 356596 179694
rect 356660 179692 356666 179756
rect 346846 179558 351322 179618
rect 366117 179618 366183 179621
rect 370257 179618 370323 179621
rect 366117 179616 370323 179618
rect 366117 179560 366122 179616
rect 366178 179560 370262 179616
rect 370318 179560 370323 179616
rect 366117 179558 370323 179560
rect 346846 179482 346906 179558
rect 366117 179555 366183 179558
rect 370257 179555 370323 179558
rect 380101 179618 380167 179621
rect 386958 179618 387018 179830
rect 391693 179827 391759 179830
rect 583838 179830 584496 179890
rect 396518 179692 396524 179756
rect 396588 179754 396594 179756
rect 396588 179694 413146 179754
rect 396588 179692 396594 179694
rect 380101 179616 387018 179618
rect 380101 179560 380106 179616
rect 380162 179560 387018 179616
rect 380101 179558 387018 179560
rect 413086 179618 413146 179694
rect 422838 179694 432466 179754
rect 413086 179558 422714 179618
rect 380101 179555 380167 179558
rect 341326 179422 346906 179482
rect 370441 179482 370507 179485
rect 379917 179482 379983 179485
rect 370441 179480 379983 179482
rect 370441 179424 370446 179480
rect 370502 179424 379922 179480
rect 379978 179424 379983 179480
rect 370441 179422 379983 179424
rect 370441 179419 370507 179422
rect 379917 179419 379983 179422
rect 391693 179482 391759 179485
rect 396518 179482 396524 179484
rect 391693 179480 396524 179482
rect 391693 179424 391698 179480
rect 391754 179424 396524 179480
rect 391693 179422 396524 179424
rect 391693 179419 391759 179422
rect 396518 179420 396524 179422
rect 396588 179420 396594 179484
rect 422654 179482 422714 179558
rect 422838 179482 422898 179694
rect 432406 179618 432466 179694
rect 442158 179694 451786 179754
rect 432406 179558 442034 179618
rect 422654 179422 422898 179482
rect 441974 179482 442034 179558
rect 442158 179482 442218 179694
rect 451726 179618 451786 179694
rect 461478 179694 471106 179754
rect 451726 179558 461354 179618
rect 441974 179422 442218 179482
rect 461294 179482 461354 179558
rect 461478 179482 461538 179694
rect 471046 179618 471106 179694
rect 480798 179694 490426 179754
rect 471046 179558 480674 179618
rect 461294 179422 461538 179482
rect 480614 179482 480674 179558
rect 480798 179482 480858 179694
rect 490366 179618 490426 179694
rect 500118 179694 509746 179754
rect 490366 179558 499994 179618
rect 480614 179422 480858 179482
rect 499934 179482 499994 179558
rect 500118 179482 500178 179694
rect 509686 179618 509746 179694
rect 519438 179694 529066 179754
rect 509686 179558 519314 179618
rect 499934 179422 500178 179482
rect 519254 179482 519314 179558
rect 519438 179482 519498 179694
rect 529006 179618 529066 179694
rect 538758 179694 544338 179754
rect 529006 179558 538634 179618
rect 519254 179422 519498 179482
rect 538574 179482 538634 179558
rect 538758 179482 538818 179694
rect 538574 179422 538818 179482
rect 544278 179482 544338 179694
rect 551078 179692 551084 179756
rect 551148 179754 551154 179756
rect 551148 179694 567706 179754
rect 551148 179692 551154 179694
rect 567646 179618 567706 179694
rect 583838 179618 583898 179830
rect 584016 179800 584496 179830
rect 567646 179558 577274 179618
rect 551078 179482 551084 179484
rect 544278 179422 551084 179482
rect 551078 179420 551084 179422
rect 551148 179420 551154 179484
rect 577214 179482 577274 179558
rect 577398 179558 583898 179618
rect 577398 179482 577458 179558
rect 577214 179422 577458 179482
rect 259857 179346 259923 179349
rect 261145 179346 261211 179349
rect 259857 179344 261211 179346
rect 259857 179288 259862 179344
rect 259918 179288 261150 179344
rect 261206 179288 261211 179344
rect 259857 179286 261211 179288
rect 259857 179283 259923 179286
rect 261145 179283 261211 179286
rect 356590 179284 356596 179348
rect 356660 179346 356666 179348
rect 366117 179346 366183 179349
rect 356660 179344 366183 179346
rect 356660 179288 366122 179344
rect 366178 179288 366183 179344
rect 356660 179286 366183 179288
rect 356660 179284 356666 179286
rect 366117 179283 366183 179286
rect 299918 179148 299924 179212
rect 299988 179210 299994 179212
rect 308198 179210 308204 179212
rect 299988 179150 308204 179210
rect 299988 179148 299994 179150
rect 308198 179148 308204 179150
rect 308268 179148 308274 179212
rect 285249 177306 285315 177309
rect 285382 177306 285388 177308
rect 285249 177304 285388 177306
rect 285249 177248 285254 177304
rect 285310 177248 285388 177304
rect 285249 177246 285388 177248
rect 285249 177243 285315 177246
rect 285382 177244 285388 177246
rect 285452 177244 285458 177308
rect 496 175946 976 175976
rect 4097 175946 4163 175949
rect 496 175944 4163 175946
rect 496 175888 4102 175944
rect 4158 175888 4163 175944
rect 496 175886 4163 175888
rect 496 175856 976 175886
rect 4097 175883 4163 175886
rect 341185 174042 341251 174045
rect 341461 174042 341527 174045
rect 553889 174044 553955 174045
rect 341185 174040 341527 174042
rect 341185 173984 341190 174040
rect 341246 173984 341466 174040
rect 341522 173984 341527 174040
rect 341185 173982 341527 173984
rect 341185 173979 341251 173982
rect 341461 173979 341527 173982
rect 553838 173980 553844 174044
rect 553908 174042 553955 174044
rect 553908 174040 554000 174042
rect 553950 173984 554000 174040
rect 553908 173982 554000 173984
rect 553908 173980 553955 173982
rect 553889 173979 553955 173980
rect 91497 173908 91563 173909
rect 91446 173906 91452 173908
rect 91406 173846 91452 173906
rect 91516 173904 91563 173908
rect 91558 173848 91563 173904
rect 91446 173844 91452 173846
rect 91516 173844 91563 173848
rect 91497 173843 91563 173844
rect 225357 173908 225423 173909
rect 225357 173904 225404 173908
rect 225468 173906 225474 173908
rect 304845 173906 304911 173909
rect 305121 173906 305187 173909
rect 225357 173848 225362 173904
rect 225357 173844 225404 173848
rect 225468 173846 225514 173906
rect 304845 173904 305187 173906
rect 304845 173848 304850 173904
rect 304906 173848 305126 173904
rect 305182 173848 305187 173904
rect 304845 173846 305187 173848
rect 225468 173844 225474 173846
rect 225357 173843 225423 173844
rect 304845 173843 304911 173846
rect 305121 173843 305187 173846
rect 341185 173906 341251 173909
rect 341369 173906 341435 173909
rect 357929 173908 357995 173909
rect 341185 173904 341435 173906
rect 341185 173848 341190 173904
rect 341246 173848 341374 173904
rect 341430 173848 341435 173904
rect 341185 173846 341435 173848
rect 341185 173843 341251 173846
rect 341369 173843 341435 173846
rect 357878 173844 357884 173908
rect 357948 173906 357995 173908
rect 553705 173906 553771 173909
rect 553889 173906 553955 173909
rect 357948 173904 358040 173906
rect 357990 173848 358040 173904
rect 357948 173846 358040 173848
rect 553705 173904 553955 173906
rect 553705 173848 553710 173904
rect 553766 173848 553894 173904
rect 553950 173848 553955 173904
rect 553705 173846 553955 173848
rect 357948 173844 357995 173846
rect 357929 173843 357995 173844
rect 553705 173843 553771 173846
rect 553889 173843 553955 173846
rect 135473 172546 135539 172549
rect 135657 172546 135723 172549
rect 135473 172544 135723 172546
rect 135473 172488 135478 172544
rect 135534 172488 135662 172544
rect 135718 172488 135723 172544
rect 135473 172486 135723 172488
rect 135473 172483 135539 172486
rect 135657 172483 135723 172486
rect 152033 172546 152099 172549
rect 152217 172546 152283 172549
rect 152033 172544 152283 172546
rect 152033 172488 152038 172544
rect 152094 172488 152222 172544
rect 152278 172488 152283 172544
rect 152033 172486 152283 172488
rect 152033 172483 152099 172486
rect 152217 172483 152283 172486
rect 170157 172546 170223 172549
rect 170341 172546 170407 172549
rect 170157 172544 170407 172546
rect 170157 172488 170162 172544
rect 170218 172488 170346 172544
rect 170402 172488 170407 172544
rect 170157 172486 170407 172488
rect 170157 172483 170223 172486
rect 170341 172483 170407 172486
rect 190673 172546 190739 172549
rect 190857 172546 190923 172549
rect 190673 172544 190923 172546
rect 190673 172488 190678 172544
rect 190734 172488 190862 172544
rect 190918 172488 190923 172544
rect 190673 172486 190923 172488
rect 190673 172483 190739 172486
rect 190857 172483 190923 172486
rect 214317 172546 214383 172549
rect 214501 172546 214567 172549
rect 214317 172544 214567 172546
rect 214317 172488 214322 172544
rect 214378 172488 214506 172544
rect 214562 172488 214567 172544
rect 214317 172486 214567 172488
rect 214317 172483 214383 172486
rect 214501 172483 214567 172486
rect 319749 172546 319815 172549
rect 319933 172546 319999 172549
rect 319749 172544 319999 172546
rect 319749 172488 319754 172544
rect 319810 172488 319938 172544
rect 319994 172488 319999 172544
rect 319749 172486 319999 172488
rect 319749 172483 319815 172486
rect 319933 172483 319999 172486
rect 373109 172546 373175 172549
rect 373293 172546 373359 172549
rect 373109 172544 373359 172546
rect 373109 172488 373114 172544
rect 373170 172488 373298 172544
rect 373354 172488 373359 172544
rect 373109 172486 373359 172488
rect 373109 172483 373175 172486
rect 373293 172483 373359 172486
rect 385529 172546 385595 172549
rect 385713 172546 385779 172549
rect 385529 172544 385779 172546
rect 385529 172488 385534 172544
rect 385590 172488 385718 172544
rect 385774 172488 385779 172544
rect 385529 172486 385779 172488
rect 385529 172483 385595 172486
rect 385713 172483 385779 172486
rect 392429 172546 392495 172549
rect 392613 172546 392679 172549
rect 392429 172544 392679 172546
rect 392429 172488 392434 172544
rect 392490 172488 392618 172544
rect 392674 172488 392679 172544
rect 392429 172486 392679 172488
rect 392429 172483 392495 172486
rect 392613 172483 392679 172486
rect 528865 172546 528931 172549
rect 529049 172546 529115 172549
rect 528865 172544 529115 172546
rect 528865 172488 528870 172544
rect 528926 172488 529054 172544
rect 529110 172488 529115 172544
rect 528865 172486 529115 172488
rect 528865 172483 528931 172486
rect 529049 172483 529115 172486
rect 535949 172546 536015 172549
rect 536133 172546 536199 172549
rect 535949 172544 536199 172546
rect 535949 172488 535954 172544
rect 536010 172488 536138 172544
rect 536194 172488 536199 172544
rect 535949 172486 536199 172488
rect 535949 172483 536015 172486
rect 536133 172483 536199 172486
rect 552325 172546 552391 172549
rect 552693 172546 552759 172549
rect 552325 172544 552759 172546
rect 552325 172488 552330 172544
rect 552386 172488 552698 172544
rect 552754 172488 552759 172544
rect 552325 172486 552759 172488
rect 552325 172483 552391 172486
rect 552693 172483 552759 172486
rect 571829 172546 571895 172549
rect 572013 172546 572079 172549
rect 571829 172544 572079 172546
rect 571829 172488 571834 172544
rect 571890 172488 572018 172544
rect 572074 172488 572079 172544
rect 571829 172486 572079 172488
rect 571829 172483 571895 172486
rect 572013 172483 572079 172486
rect 560830 164596 560836 164660
rect 560900 164658 560906 164660
rect 570357 164658 570423 164661
rect 560900 164656 570423 164658
rect 560900 164600 570362 164656
rect 570418 164600 570423 164656
rect 560900 164598 570423 164600
rect 560900 164596 560906 164598
rect 570357 164595 570423 164598
rect 135657 164522 135723 164525
rect 135614 164520 135723 164522
rect 135614 164464 135662 164520
rect 135718 164464 135723 164520
rect 135614 164459 135723 164464
rect 276693 164522 276759 164525
rect 285157 164522 285223 164525
rect 385529 164522 385595 164525
rect 276693 164520 276802 164522
rect 276693 164464 276698 164520
rect 276754 164464 276802 164520
rect 276693 164459 276802 164464
rect 285157 164520 285266 164522
rect 285157 164464 285162 164520
rect 285218 164464 285266 164520
rect 285157 164459 285266 164464
rect 135614 164389 135674 164459
rect 135565 164384 135674 164389
rect 135565 164328 135570 164384
rect 135626 164328 135674 164384
rect 135565 164326 135674 164328
rect 276742 164389 276802 164459
rect 285206 164389 285266 164459
rect 385486 164520 385595 164522
rect 385486 164464 385534 164520
rect 385590 164464 385595 164520
rect 385486 164459 385595 164464
rect 392429 164522 392495 164525
rect 529049 164522 529115 164525
rect 392429 164520 392538 164522
rect 392429 164464 392434 164520
rect 392490 164464 392538 164520
rect 392429 164459 392538 164464
rect 276742 164384 276851 164389
rect 276742 164328 276790 164384
rect 276846 164328 276851 164384
rect 276742 164326 276851 164328
rect 135565 164323 135631 164326
rect 276785 164323 276851 164326
rect 285157 164384 285266 164389
rect 285157 164328 285162 164384
rect 285218 164328 285266 164384
rect 285157 164326 285266 164328
rect 341093 164386 341159 164389
rect 341369 164386 341435 164389
rect 357929 164388 357995 164389
rect 341093 164384 341435 164386
rect 341093 164328 341098 164384
rect 341154 164328 341374 164384
rect 341430 164328 341435 164384
rect 341093 164326 341435 164328
rect 285157 164323 285223 164326
rect 341093 164323 341159 164326
rect 341369 164323 341435 164326
rect 357878 164324 357884 164388
rect 357948 164386 357995 164388
rect 357948 164384 358040 164386
rect 357990 164328 358040 164384
rect 357948 164326 358040 164328
rect 357948 164324 357995 164326
rect 357929 164323 357995 164324
rect 385486 164253 385546 164459
rect 392478 164253 392538 164459
rect 529006 164520 529115 164522
rect 529006 164464 529054 164520
rect 529110 164464 529115 164520
rect 529006 164459 529115 164464
rect 535949 164522 536015 164525
rect 571829 164522 571895 164525
rect 535949 164520 536058 164522
rect 535949 164464 535954 164520
rect 536010 164464 536058 164520
rect 535949 164459 536058 164464
rect 571829 164520 571938 164522
rect 571829 164464 571834 164520
rect 571890 164464 571938 164520
rect 571829 164459 571938 164464
rect 529006 164253 529066 164459
rect 535998 164253 536058 164459
rect 571878 164253 571938 164459
rect 91497 164252 91563 164253
rect 91446 164188 91452 164252
rect 91516 164250 91563 164252
rect 225357 164252 225423 164253
rect 91516 164248 91608 164250
rect 91558 164192 91608 164248
rect 91516 164190 91608 164192
rect 225357 164248 225404 164252
rect 225468 164250 225474 164252
rect 242653 164250 242719 164253
rect 242837 164250 242903 164253
rect 225357 164192 225362 164248
rect 91516 164188 91563 164190
rect 91497 164187 91563 164188
rect 225357 164188 225404 164192
rect 225468 164190 225514 164250
rect 242653 164248 242903 164250
rect 242653 164192 242658 164248
rect 242714 164192 242842 164248
rect 242898 164192 242903 164248
rect 242653 164190 242903 164192
rect 225468 164188 225474 164190
rect 225357 164187 225423 164188
rect 242653 164187 242719 164190
rect 242837 164187 242903 164190
rect 243246 164188 243252 164252
rect 243316 164250 243322 164252
rect 284789 164250 284855 164253
rect 243316 164248 284855 164250
rect 243316 164192 284794 164248
rect 284850 164192 284855 164248
rect 243316 164190 284855 164192
rect 243316 164188 243322 164190
rect 284789 164187 284855 164190
rect 285617 164250 285683 164253
rect 382033 164250 382099 164253
rect 285617 164248 382099 164250
rect 285617 164192 285622 164248
rect 285678 164192 382038 164248
rect 382094 164192 382099 164248
rect 285617 164190 382099 164192
rect 385486 164248 385595 164253
rect 385486 164192 385534 164248
rect 385590 164192 385595 164248
rect 385486 164190 385595 164192
rect 285617 164187 285683 164190
rect 382033 164187 382099 164190
rect 385529 164187 385595 164190
rect 385805 164250 385871 164253
rect 391693 164250 391759 164253
rect 385805 164248 391759 164250
rect 385805 164192 385810 164248
rect 385866 164192 391698 164248
rect 391754 164192 391759 164248
rect 385805 164190 391759 164192
rect 385805 164187 385871 164190
rect 391693 164187 391759 164190
rect 392429 164248 392538 164253
rect 392429 164192 392434 164248
rect 392490 164192 392538 164248
rect 392429 164190 392538 164192
rect 392705 164250 392771 164253
rect 526933 164250 526999 164253
rect 392705 164248 526999 164250
rect 392705 164192 392710 164248
rect 392766 164192 526938 164248
rect 526994 164192 526999 164248
rect 392705 164190 526999 164192
rect 529006 164248 529115 164253
rect 529006 164192 529054 164248
rect 529110 164192 529115 164248
rect 529006 164190 529115 164192
rect 392429 164187 392495 164190
rect 392705 164187 392771 164190
rect 526933 164187 526999 164190
rect 529049 164187 529115 164190
rect 529325 164250 529391 164253
rect 535673 164250 535739 164253
rect 529325 164248 535739 164250
rect 529325 164192 529330 164248
rect 529386 164192 535678 164248
rect 535734 164192 535739 164248
rect 529325 164190 535739 164192
rect 529325 164187 529391 164190
rect 535673 164187 535739 164190
rect 535949 164248 536058 164253
rect 535949 164192 535954 164248
rect 536010 164192 536058 164248
rect 535949 164190 536058 164192
rect 536593 164250 536659 164253
rect 560830 164250 560836 164252
rect 536593 164248 560836 164250
rect 536593 164192 536598 164248
rect 536654 164192 560836 164248
rect 536593 164190 560836 164192
rect 535949 164187 536015 164190
rect 536593 164187 536659 164190
rect 560830 164188 560836 164190
rect 560900 164188 560906 164252
rect 570357 164250 570423 164253
rect 571553 164250 571619 164253
rect 570357 164248 571619 164250
rect 570357 164192 570362 164248
rect 570418 164192 571558 164248
rect 571614 164192 571619 164248
rect 570357 164190 571619 164192
rect 570357 164187 570423 164190
rect 571553 164187 571619 164190
rect 571829 164248 571938 164253
rect 571829 164192 571834 164248
rect 571890 164192 571938 164248
rect 571829 164190 571938 164192
rect 572105 164250 572171 164253
rect 584016 164250 584496 164280
rect 572105 164248 584496 164250
rect 572105 164192 572110 164248
rect 572166 164192 584496 164248
rect 572105 164190 584496 164192
rect 571829 164187 571895 164190
rect 572105 164187 572171 164190
rect 584016 164160 584496 164190
rect 285341 164116 285407 164117
rect 285341 164114 285388 164116
rect 285296 164112 285388 164114
rect 285296 164056 285346 164112
rect 285296 164054 285388 164056
rect 285341 164052 285388 164054
rect 285452 164052 285458 164116
rect 285341 164051 285407 164052
rect 242561 163028 242627 163029
rect 242510 162964 242516 163028
rect 242580 163026 242627 163028
rect 278809 163026 278875 163029
rect 242580 163024 242672 163026
rect 242622 162968 242672 163024
rect 242580 162966 242672 162968
rect 278766 163024 278875 163026
rect 278766 162968 278814 163024
rect 278870 162968 278875 163024
rect 242580 162964 242627 162966
rect 242561 162963 242627 162964
rect 278766 162963 278875 162968
rect 278766 162893 278826 162963
rect 278717 162888 278826 162893
rect 278717 162832 278722 162888
rect 278778 162832 278826 162888
rect 278717 162830 278826 162832
rect 278717 162827 278783 162830
rect 496 159218 976 159248
rect 4005 159218 4071 159221
rect 496 159216 4071 159218
rect 496 159160 4010 159216
rect 4066 159160 4071 159216
rect 496 159158 4071 159160
rect 496 159128 976 159158
rect 4005 159155 4071 159158
rect 242469 157860 242535 157861
rect 242469 157858 242516 157860
rect 242424 157856 242516 157858
rect 242424 157800 242474 157856
rect 242424 157798 242516 157800
rect 242469 157796 242516 157798
rect 242580 157796 242586 157860
rect 242469 157795 242535 157796
rect 331065 154594 331131 154597
rect 331249 154594 331315 154597
rect 331065 154592 331315 154594
rect 331065 154536 331070 154592
rect 331126 154536 331254 154592
rect 331310 154536 331315 154592
rect 331065 154534 331315 154536
rect 331065 154531 331131 154534
rect 331249 154531 331315 154534
rect 91497 154458 91563 154461
rect 91773 154458 91839 154461
rect 91497 154456 91839 154458
rect 91497 154400 91502 154456
rect 91558 154400 91778 154456
rect 91834 154400 91839 154456
rect 91497 154398 91839 154400
rect 91497 154395 91563 154398
rect 91773 154395 91839 154398
rect 235569 154458 235635 154461
rect 235845 154458 235911 154461
rect 235569 154456 235911 154458
rect 235569 154400 235574 154456
rect 235630 154400 235850 154456
rect 235906 154400 235911 154456
rect 235569 154398 235911 154400
rect 235569 154395 235635 154398
rect 235845 154395 235911 154398
rect 357929 154458 357995 154461
rect 358205 154458 358271 154461
rect 357929 154456 358271 154458
rect 357929 154400 357934 154456
rect 357990 154400 358210 154456
rect 358266 154400 358271 154456
rect 357929 154398 358271 154400
rect 357929 154395 357995 154398
rect 358205 154395 358271 154398
rect 242009 153234 242075 153237
rect 242193 153234 242259 153237
rect 242009 153232 242259 153234
rect 242009 153176 242014 153232
rect 242070 153176 242198 153232
rect 242254 153176 242259 153232
rect 242009 153174 242259 153176
rect 242009 153171 242075 153174
rect 242193 153171 242259 153174
rect 319841 153234 319907 153237
rect 320025 153234 320091 153237
rect 319841 153232 320091 153234
rect 319841 153176 319846 153232
rect 319902 153176 320030 153232
rect 320086 153176 320091 153232
rect 319841 153174 320091 153176
rect 319841 153171 319907 153174
rect 320025 153171 320091 153174
rect 309169 151738 309235 151741
rect 309302 151738 309308 151740
rect 309169 151736 309308 151738
rect 309169 151680 309174 151736
rect 309230 151680 309308 151736
rect 309169 151678 309308 151680
rect 309169 151675 309235 151678
rect 309302 151676 309308 151678
rect 309372 151676 309378 151740
rect 580385 148610 580451 148613
rect 584016 148610 584496 148640
rect 580385 148608 584496 148610
rect 580385 148552 580390 148608
rect 580446 148552 584496 148608
rect 580385 148550 584496 148552
rect 580385 148547 580451 148550
rect 584016 148520 584496 148550
rect 91497 144938 91563 144941
rect 91773 144938 91839 144941
rect 91497 144936 91839 144938
rect 91497 144880 91502 144936
rect 91558 144880 91778 144936
rect 91834 144880 91839 144936
rect 91497 144878 91839 144880
rect 91497 144875 91563 144878
rect 91773 144875 91839 144878
rect 235477 144938 235543 144941
rect 235845 144938 235911 144941
rect 242469 144940 242535 144941
rect 242469 144938 242516 144940
rect 235477 144936 235911 144938
rect 235477 144880 235482 144936
rect 235538 144880 235850 144936
rect 235906 144880 235911 144936
rect 235477 144878 235911 144880
rect 242424 144936 242516 144938
rect 242424 144880 242474 144936
rect 242424 144878 242516 144880
rect 235477 144875 235543 144878
rect 235845 144875 235911 144878
rect 242469 144876 242516 144878
rect 242580 144876 242586 144940
rect 357929 144938 357995 144941
rect 358205 144938 358271 144941
rect 357929 144936 358271 144938
rect 357929 144880 357934 144936
rect 357990 144880 358210 144936
rect 358266 144880 358271 144936
rect 357929 144878 358271 144880
rect 242469 144875 242535 144876
rect 357929 144875 357995 144878
rect 358205 144875 358271 144878
rect 496 142354 976 142384
rect 4005 142354 4071 142357
rect 496 142352 4071 142354
rect 496 142296 4010 142352
rect 4066 142296 4071 142352
rect 496 142294 4071 142296
rect 496 142264 976 142294
rect 4005 142291 4071 142294
rect 309169 142218 309235 142221
rect 309302 142218 309308 142220
rect 309169 142216 309308 142218
rect 309169 142160 309174 142216
rect 309230 142160 309308 142216
rect 309169 142158 309308 142160
rect 309169 142155 309235 142158
rect 309302 142156 309308 142158
rect 309372 142156 309378 142220
rect 229773 135282 229839 135285
rect 229957 135282 230023 135285
rect 229773 135280 230023 135282
rect 229773 135224 229778 135280
rect 229834 135224 229962 135280
rect 230018 135224 230023 135280
rect 229773 135222 230023 135224
rect 229773 135219 229839 135222
rect 229957 135219 230023 135222
rect 331065 135282 331131 135285
rect 331249 135282 331315 135285
rect 331065 135280 331315 135282
rect 331065 135224 331070 135280
rect 331126 135224 331254 135280
rect 331310 135224 331315 135280
rect 331065 135222 331315 135224
rect 331065 135219 331131 135222
rect 331249 135219 331315 135222
rect 239014 133996 239020 134060
rect 239084 134058 239090 134060
rect 241825 134058 241891 134061
rect 239084 134056 241891 134058
rect 239084 134000 241830 134056
rect 241886 134000 241891 134056
rect 239084 133998 241891 134000
rect 239084 133996 239090 133998
rect 241825 133995 241891 133998
rect 242009 133922 242075 133925
rect 242193 133922 242259 133925
rect 242009 133920 242259 133922
rect 242009 133864 242014 133920
rect 242070 133864 242198 133920
rect 242254 133864 242259 133920
rect 242009 133862 242259 133864
rect 242009 133859 242075 133862
rect 242193 133859 242259 133862
rect 276693 133922 276759 133925
rect 276877 133922 276943 133925
rect 276693 133920 276943 133922
rect 276693 133864 276698 133920
rect 276754 133864 276882 133920
rect 276938 133864 276943 133920
rect 276693 133862 276943 133864
rect 276693 133859 276759 133862
rect 276877 133859 276943 133862
rect 373017 133922 373083 133925
rect 373293 133922 373359 133925
rect 373017 133920 373359 133922
rect 373017 133864 373022 133920
rect 373078 133864 373298 133920
rect 373354 133864 373359 133920
rect 373017 133862 373359 133864
rect 373017 133859 373083 133862
rect 373293 133859 373359 133862
rect 357878 133044 357884 133108
rect 357948 133106 357954 133108
rect 366158 133106 366164 133108
rect 357948 133046 366164 133106
rect 357948 133044 357954 133046
rect 366158 133044 366164 133046
rect 366228 133044 366234 133108
rect 251761 132970 251827 132973
rect 390313 132970 390379 132973
rect 584016 132970 584496 133000
rect 251761 132968 275146 132970
rect 251761 132912 251766 132968
rect 251822 132912 275146 132968
rect 251761 132910 275146 132912
rect 251761 132907 251827 132910
rect 241825 132834 241891 132837
rect 275086 132834 275146 132910
rect 385486 132968 390379 132970
rect 385486 132912 390318 132968
rect 390374 132912 390379 132968
rect 385486 132910 390379 132912
rect 290309 132834 290375 132837
rect 241825 132832 246810 132834
rect 241825 132776 241830 132832
rect 241886 132776 246810 132832
rect 241825 132774 246810 132776
rect 275086 132832 290375 132834
rect 275086 132776 290314 132832
rect 290370 132776 290375 132832
rect 275086 132774 290375 132776
rect 241825 132771 241891 132774
rect 246750 132698 246810 132774
rect 290309 132771 290375 132774
rect 308198 132772 308204 132836
rect 308268 132834 308274 132836
rect 317766 132834 317772 132836
rect 308268 132774 317772 132834
rect 308268 132772 308274 132774
rect 317766 132772 317772 132774
rect 317836 132772 317842 132836
rect 327518 132772 327524 132836
rect 327588 132834 327594 132836
rect 357878 132834 357884 132836
rect 327588 132774 341386 132834
rect 327588 132772 327594 132774
rect 251761 132698 251827 132701
rect 246750 132696 251827 132698
rect 246750 132640 251766 132696
rect 251822 132640 251827 132696
rect 246750 132638 251827 132640
rect 251761 132635 251827 132638
rect 293253 132698 293319 132701
rect 293253 132696 302562 132698
rect 293253 132640 293258 132696
rect 293314 132640 302562 132696
rect 293253 132638 302562 132640
rect 293253 132635 293319 132638
rect 302502 132562 302562 132638
rect 308198 132562 308204 132564
rect 302502 132502 308204 132562
rect 308198 132500 308204 132502
rect 308268 132500 308274 132564
rect 317766 132500 317772 132564
rect 317836 132562 317842 132564
rect 327518 132562 327524 132564
rect 317836 132502 327524 132562
rect 317836 132500 317842 132502
rect 327518 132500 327524 132502
rect 327588 132500 327594 132564
rect 341326 132562 341386 132774
rect 351078 132774 357884 132834
rect 351078 132562 351138 132774
rect 357878 132772 357884 132774
rect 357948 132772 357954 132836
rect 385486 132701 385546 132910
rect 390313 132907 390379 132910
rect 583838 132910 584496 132970
rect 406137 132834 406203 132837
rect 406137 132832 413146 132834
rect 406137 132776 406142 132832
rect 406198 132776 413146 132832
rect 406137 132774 413146 132776
rect 406137 132771 406203 132774
rect 366158 132636 366164 132700
rect 366228 132698 366234 132700
rect 385437 132698 385546 132701
rect 399237 132698 399303 132701
rect 366228 132638 368250 132698
rect 385356 132696 385546 132698
rect 385356 132640 385442 132696
rect 385498 132640 385546 132696
rect 385356 132638 385546 132640
rect 396526 132696 399303 132698
rect 396526 132640 399242 132696
rect 399298 132640 399303 132696
rect 396526 132638 399303 132640
rect 413086 132698 413146 132774
rect 422838 132774 432466 132834
rect 413086 132638 422714 132698
rect 366228 132636 366234 132638
rect 341326 132502 351138 132562
rect 368190 132562 368250 132638
rect 385437 132635 385503 132638
rect 375869 132562 375935 132565
rect 368190 132560 375935 132562
rect 368190 132504 375874 132560
rect 375930 132504 375935 132560
rect 368190 132502 375935 132504
rect 375869 132499 375935 132502
rect 390313 132562 390379 132565
rect 396526 132562 396586 132638
rect 399237 132635 399303 132638
rect 390313 132560 396586 132562
rect 390313 132504 390318 132560
rect 390374 132504 396586 132560
rect 390313 132502 396586 132504
rect 422654 132562 422714 132638
rect 422838 132562 422898 132774
rect 432406 132698 432466 132774
rect 442158 132774 451786 132834
rect 432406 132638 442034 132698
rect 422654 132502 422898 132562
rect 441974 132562 442034 132638
rect 442158 132562 442218 132774
rect 451726 132698 451786 132774
rect 461478 132774 471106 132834
rect 451726 132638 461354 132698
rect 441974 132502 442218 132562
rect 461294 132562 461354 132638
rect 461478 132562 461538 132774
rect 471046 132698 471106 132774
rect 480798 132774 490426 132834
rect 471046 132638 480674 132698
rect 461294 132502 461538 132562
rect 480614 132562 480674 132638
rect 480798 132562 480858 132774
rect 490366 132698 490426 132774
rect 500118 132774 509746 132834
rect 490366 132638 499994 132698
rect 480614 132502 480858 132562
rect 499934 132562 499994 132638
rect 500118 132562 500178 132774
rect 509686 132698 509746 132774
rect 519438 132774 529066 132834
rect 509686 132638 519314 132698
rect 499934 132502 500178 132562
rect 519254 132562 519314 132638
rect 519438 132562 519498 132774
rect 529006 132698 529066 132774
rect 538758 132774 544338 132834
rect 529006 132638 538634 132698
rect 519254 132502 519498 132562
rect 538574 132562 538634 132638
rect 538758 132562 538818 132774
rect 538574 132502 538818 132562
rect 544278 132562 544338 132774
rect 551078 132772 551084 132836
rect 551148 132834 551154 132836
rect 551148 132774 567706 132834
rect 551148 132772 551154 132774
rect 567646 132698 567706 132774
rect 583838 132698 583898 132910
rect 584016 132880 584496 132910
rect 567646 132638 577274 132698
rect 551078 132562 551084 132564
rect 544278 132502 551084 132562
rect 390313 132499 390379 132502
rect 551078 132500 551084 132502
rect 551148 132500 551154 132564
rect 577214 132562 577274 132638
rect 577398 132638 583898 132698
rect 577398 132562 577458 132638
rect 577214 132502 577458 132562
rect 4005 126986 4071 126989
rect 342790 126986 342796 126988
rect 4005 126984 342796 126986
rect 4005 126928 4010 126984
rect 4066 126928 342796 126984
rect 4005 126926 342796 126928
rect 4005 126923 4071 126926
rect 342790 126924 342796 126926
rect 342860 126924 342866 126988
rect 91313 125762 91379 125765
rect 242193 125762 242259 125765
rect 373293 125762 373359 125765
rect 91313 125760 91514 125762
rect 91313 125704 91318 125760
rect 91374 125704 91514 125760
rect 91313 125702 91514 125704
rect 91313 125699 91379 125702
rect 496 125626 976 125656
rect 91454 125629 91514 125702
rect 242150 125760 242259 125762
rect 242150 125704 242198 125760
rect 242254 125704 242259 125760
rect 242150 125699 242259 125704
rect 372974 125760 373359 125762
rect 372974 125704 373298 125760
rect 373354 125704 373359 125760
rect 372974 125702 373359 125704
rect 242150 125629 242210 125699
rect 4005 125626 4071 125629
rect 496 125624 4071 125626
rect 496 125568 4010 125624
rect 4066 125568 4071 125624
rect 496 125566 4071 125568
rect 91454 125624 91563 125629
rect 91454 125568 91502 125624
rect 91558 125568 91563 125624
rect 91454 125566 91563 125568
rect 496 125536 976 125566
rect 4005 125563 4071 125566
rect 91497 125563 91563 125566
rect 235569 125626 235635 125629
rect 235753 125626 235819 125629
rect 235569 125624 235819 125626
rect 235569 125568 235574 125624
rect 235630 125568 235758 125624
rect 235814 125568 235819 125624
rect 235569 125566 235819 125568
rect 235569 125563 235635 125566
rect 235753 125563 235819 125566
rect 242101 125624 242210 125629
rect 242101 125568 242106 125624
rect 242162 125568 242210 125624
rect 242101 125566 242210 125568
rect 341185 125626 341251 125629
rect 341369 125626 341435 125629
rect 341185 125624 341435 125626
rect 341185 125568 341190 125624
rect 341246 125568 341374 125624
rect 341430 125568 341435 125624
rect 341185 125566 341435 125568
rect 372974 125626 373034 125702
rect 373293 125699 373359 125702
rect 373109 125626 373175 125629
rect 372974 125624 373175 125626
rect 372974 125568 373114 125624
rect 373170 125568 373175 125624
rect 372974 125566 373175 125568
rect 242101 125563 242167 125566
rect 341185 125563 341251 125566
rect 341369 125563 341435 125566
rect 373109 125563 373175 125566
rect 553705 125626 553771 125629
rect 553889 125626 553955 125629
rect 553705 125624 553955 125626
rect 553705 125568 553710 125624
rect 553766 125568 553894 125624
rect 553950 125568 553955 125624
rect 553705 125566 553955 125568
rect 553705 125563 553771 125566
rect 553889 125563 553955 125566
rect 275497 118690 275563 118693
rect 275681 118690 275747 118693
rect 275497 118688 275747 118690
rect 275497 118632 275502 118688
rect 275558 118632 275686 118688
rect 275742 118632 275747 118688
rect 275497 118630 275747 118632
rect 275497 118627 275563 118630
rect 275681 118627 275747 118630
rect 240486 117268 240492 117332
rect 240556 117330 240562 117332
rect 584016 117330 584496 117360
rect 240556 117270 584496 117330
rect 240556 117268 240562 117270
rect 584016 117240 584496 117270
rect 328213 115970 328279 115973
rect 328397 115970 328463 115973
rect 328213 115968 328463 115970
rect 328213 115912 328218 115968
rect 328274 115912 328402 115968
rect 328458 115912 328463 115968
rect 328213 115910 328463 115912
rect 328213 115907 328279 115910
rect 328397 115907 328463 115910
rect 331065 115970 331131 115973
rect 331249 115970 331315 115973
rect 331065 115968 331315 115970
rect 331065 115912 331070 115968
rect 331126 115912 331254 115968
rect 331310 115912 331315 115968
rect 331065 115910 331315 115912
rect 331065 115907 331131 115910
rect 331249 115907 331315 115910
rect 341185 115834 341251 115837
rect 341461 115834 341527 115837
rect 341185 115832 341527 115834
rect 341185 115776 341190 115832
rect 341246 115776 341466 115832
rect 341522 115776 341527 115832
rect 341185 115774 341527 115776
rect 341185 115771 341251 115774
rect 341461 115771 341527 115774
rect 553429 113250 553495 113253
rect 553613 113250 553679 113253
rect 553429 113248 553679 113250
rect 553429 113192 553434 113248
rect 553490 113192 553618 113248
rect 553674 113192 553679 113248
rect 553429 113190 553679 113192
rect 553429 113187 553495 113190
rect 553613 113187 553679 113190
rect 271357 109034 271423 109037
rect 271633 109034 271699 109037
rect 271357 109032 271699 109034
rect 271357 108976 271362 109032
rect 271418 108976 271638 109032
rect 271694 108976 271699 109032
rect 271357 108974 271699 108976
rect 271357 108971 271423 108974
rect 271633 108971 271699 108974
rect 496 108898 976 108928
rect 3913 108898 3979 108901
rect 496 108896 3979 108898
rect 496 108840 3918 108896
rect 3974 108840 3979 108896
rect 496 108838 3979 108840
rect 496 108808 976 108838
rect 3913 108835 3979 108838
rect 242193 106450 242259 106453
rect 242150 106448 242259 106450
rect 242150 106392 242198 106448
rect 242254 106392 242259 106448
rect 242150 106387 242259 106392
rect 242150 106317 242210 106387
rect 242101 106312 242210 106317
rect 242101 106256 242106 106312
rect 242162 106256 242210 106312
rect 242101 106254 242210 106256
rect 341185 106314 341251 106317
rect 341461 106314 341527 106317
rect 341185 106312 341527 106314
rect 341185 106256 341190 106312
rect 341246 106256 341466 106312
rect 341522 106256 341527 106312
rect 341185 106254 341527 106256
rect 242101 106251 242167 106254
rect 341185 106251 341251 106254
rect 341461 106251 341527 106254
rect 552417 104954 552483 104957
rect 552601 104954 552667 104957
rect 552417 104952 552667 104954
rect 552417 104896 552422 104952
rect 552478 104896 552606 104952
rect 552662 104896 552667 104952
rect 552417 104894 552667 104896
rect 552417 104891 552483 104894
rect 552601 104891 552667 104894
rect 584016 101690 584496 101720
rect 583838 101630 584496 101690
rect 377198 101356 377204 101420
rect 377268 101418 377274 101420
rect 386817 101418 386883 101421
rect 377268 101416 386883 101418
rect 377268 101360 386822 101416
rect 386878 101360 386883 101416
rect 377268 101358 386883 101360
rect 377268 101356 377274 101358
rect 386817 101355 386883 101358
rect 391693 101282 391759 101285
rect 386958 101280 391759 101282
rect 386958 101224 391698 101280
rect 391754 101224 391759 101280
rect 386958 101222 391759 101224
rect 237726 101084 237732 101148
rect 237796 101146 237802 101148
rect 261145 101146 261211 101149
rect 290217 101146 290283 101149
rect 237796 101086 244970 101146
rect 237796 101084 237802 101086
rect 244910 100874 244970 101086
rect 261145 101144 264290 101146
rect 261145 101088 261150 101144
rect 261206 101088 264290 101144
rect 261145 101086 264290 101088
rect 261145 101083 261211 101086
rect 251669 100874 251735 100877
rect 244910 100872 251735 100874
rect 244910 100816 251674 100872
rect 251730 100816 251735 100872
rect 244910 100814 251735 100816
rect 264230 100874 264290 101086
rect 275822 101144 290283 101146
rect 275822 101088 290222 101144
rect 290278 101088 290283 101144
rect 275822 101086 290283 101088
rect 275822 100874 275882 101086
rect 290217 101083 290283 101086
rect 290401 101146 290467 101149
rect 377198 101146 377204 101148
rect 290401 101144 293730 101146
rect 290401 101088 290406 101144
rect 290462 101088 293730 101144
rect 290401 101086 293730 101088
rect 290401 101083 290467 101086
rect 293670 101010 293730 101086
rect 335622 101086 341386 101146
rect 293670 100950 302562 101010
rect 264230 100814 275882 100874
rect 251669 100811 251735 100814
rect 279821 100738 279887 100741
rect 280005 100738 280071 100741
rect 279821 100736 280071 100738
rect 279821 100680 279826 100736
rect 279882 100680 280010 100736
rect 280066 100680 280071 100736
rect 279821 100678 280071 100680
rect 302502 100738 302562 100950
rect 316478 100874 316484 100876
rect 316302 100814 316484 100874
rect 302502 100678 308082 100738
rect 279821 100675 279887 100678
rect 280005 100675 280071 100678
rect 308022 100602 308082 100678
rect 316302 100602 316362 100814
rect 316478 100812 316484 100814
rect 316548 100812 316554 100876
rect 330973 100874 331039 100877
rect 335622 100874 335682 101086
rect 330973 100872 335682 100874
rect 330973 100816 330978 100872
rect 331034 100816 335682 100872
rect 330973 100814 335682 100816
rect 341326 100874 341386 101086
rect 370398 101086 377204 101146
rect 360413 101010 360479 101013
rect 351078 101008 360479 101010
rect 351078 100952 360418 101008
rect 360474 100952 360479 101008
rect 351078 100950 360479 100952
rect 351078 100874 351138 100950
rect 360413 100947 360479 100950
rect 341326 100814 351138 100874
rect 366117 100874 366183 100877
rect 370398 100874 370458 101086
rect 377198 101084 377204 101086
rect 377268 101084 377274 101148
rect 386817 101010 386883 101013
rect 386958 101010 387018 101222
rect 391693 101219 391759 101222
rect 396518 101084 396524 101148
rect 396588 101146 396594 101148
rect 396588 101086 413146 101146
rect 396588 101084 396594 101086
rect 386817 101008 387018 101010
rect 386817 100952 386822 101008
rect 386878 100952 387018 101008
rect 386817 100950 387018 100952
rect 413086 101010 413146 101086
rect 422838 101086 432466 101146
rect 413086 100950 422714 101010
rect 386817 100947 386883 100950
rect 366117 100872 370458 100874
rect 366117 100816 366122 100872
rect 366178 100816 370458 100872
rect 366117 100814 370458 100816
rect 391693 100874 391759 100877
rect 396518 100874 396524 100876
rect 391693 100872 396524 100874
rect 391693 100816 391698 100872
rect 391754 100816 396524 100872
rect 391693 100814 396524 100816
rect 330973 100811 331039 100814
rect 366117 100811 366183 100814
rect 391693 100811 391759 100814
rect 396518 100812 396524 100814
rect 396588 100812 396594 100876
rect 422654 100874 422714 100950
rect 422838 100874 422898 101086
rect 432406 101010 432466 101086
rect 442158 101086 451786 101146
rect 432406 100950 442034 101010
rect 422654 100814 422898 100874
rect 441974 100874 442034 100950
rect 442158 100874 442218 101086
rect 451726 101010 451786 101086
rect 461478 101086 471106 101146
rect 451726 100950 461354 101010
rect 441974 100814 442218 100874
rect 461294 100874 461354 100950
rect 461478 100874 461538 101086
rect 471046 101010 471106 101086
rect 480798 101086 490426 101146
rect 471046 100950 480674 101010
rect 461294 100814 461538 100874
rect 480614 100874 480674 100950
rect 480798 100874 480858 101086
rect 490366 101010 490426 101086
rect 500118 101086 509746 101146
rect 490366 100950 499994 101010
rect 480614 100814 480858 100874
rect 499934 100874 499994 100950
rect 500118 100874 500178 101086
rect 509686 101010 509746 101086
rect 519438 101086 529066 101146
rect 509686 100950 519314 101010
rect 499934 100814 500178 100874
rect 519254 100874 519314 100950
rect 519438 100874 519498 101086
rect 529006 101010 529066 101086
rect 538758 101086 544338 101146
rect 529006 100950 538634 101010
rect 519254 100814 519498 100874
rect 538574 100874 538634 100950
rect 538758 100874 538818 101086
rect 538574 100814 538818 100874
rect 544278 100874 544338 101086
rect 551078 101084 551084 101148
rect 551148 101146 551154 101148
rect 551148 101086 567706 101146
rect 551148 101084 551154 101086
rect 567646 101010 567706 101086
rect 583838 101010 583898 101630
rect 584016 101600 584496 101630
rect 567646 100950 577274 101010
rect 551078 100874 551084 100876
rect 544278 100814 551084 100874
rect 551078 100812 551084 100814
rect 551148 100812 551154 100876
rect 577214 100874 577274 100950
rect 577398 100950 583898 101010
rect 577398 100874 577458 100950
rect 577214 100814 577458 100874
rect 308022 100542 316362 100602
rect 316478 100540 316484 100604
rect 316548 100602 316554 100604
rect 330973 100602 331039 100605
rect 316548 100600 331039 100602
rect 316548 100544 330978 100600
rect 331034 100544 331039 100600
rect 316548 100542 331039 100544
rect 316548 100540 316554 100542
rect 330973 100539 331039 100542
rect 246885 96794 246951 96797
rect 246750 96792 246951 96794
rect 246750 96736 246890 96792
rect 246946 96736 246951 96792
rect 246750 96734 246951 96736
rect 246750 96661 246810 96734
rect 246885 96731 246951 96734
rect 239249 96658 239315 96661
rect 239433 96658 239499 96661
rect 239249 96656 239499 96658
rect 239249 96600 239254 96656
rect 239310 96600 239438 96656
rect 239494 96600 239499 96656
rect 239249 96598 239499 96600
rect 239249 96595 239315 96598
rect 239433 96595 239499 96598
rect 242469 96658 242535 96661
rect 242653 96658 242719 96661
rect 242469 96656 242719 96658
rect 242469 96600 242474 96656
rect 242530 96600 242658 96656
rect 242714 96600 242719 96656
rect 242469 96598 242719 96600
rect 246750 96656 246859 96661
rect 246750 96600 246798 96656
rect 246854 96600 246859 96656
rect 246750 96598 246859 96600
rect 242469 96595 242535 96598
rect 242653 96595 242719 96598
rect 246793 96595 246859 96598
rect 331065 96658 331131 96661
rect 331249 96658 331315 96661
rect 331065 96656 331315 96658
rect 331065 96600 331070 96656
rect 331126 96600 331254 96656
rect 331310 96600 331315 96656
rect 331065 96598 331315 96600
rect 331065 96595 331131 96598
rect 331249 96595 331315 96598
rect 328489 95162 328555 95165
rect 328446 95160 328555 95162
rect 328446 95104 328494 95160
rect 328550 95104 328555 95160
rect 328446 95099 328555 95104
rect 328446 95029 328506 95099
rect 328446 95024 328555 95029
rect 328446 94968 328494 95024
rect 328550 94968 328555 95024
rect 328446 94966 328555 94968
rect 328489 94963 328555 94966
rect 344078 92442 344084 92444
rect 1110 92382 344084 92442
rect 496 92170 976 92200
rect 1110 92170 1170 92382
rect 344078 92380 344084 92382
rect 344148 92380 344154 92444
rect 496 92110 1170 92170
rect 496 92080 976 92110
rect 560789 87274 560855 87277
rect 560789 87272 560898 87274
rect 560789 87216 560794 87272
rect 560850 87216 560898 87272
rect 560789 87211 560898 87216
rect 560838 87141 560898 87211
rect 91313 87138 91379 87141
rect 358205 87138 358271 87141
rect 91313 87136 91514 87138
rect 91313 87080 91318 87136
rect 91374 87080 91514 87136
rect 91313 87078 91514 87080
rect 91313 87075 91379 87078
rect 91454 87005 91514 87078
rect 357886 87136 358271 87138
rect 357886 87080 358210 87136
rect 358266 87080 358271 87136
rect 357886 87078 358271 87080
rect 357886 87005 357946 87078
rect 358205 87075 358271 87078
rect 553705 87138 553771 87141
rect 553705 87136 553906 87138
rect 553705 87080 553710 87136
rect 553766 87080 553906 87136
rect 553705 87078 553906 87080
rect 553705 87075 553771 87078
rect 553846 87005 553906 87078
rect 560789 87136 560898 87141
rect 560789 87080 560794 87136
rect 560850 87080 560898 87136
rect 560789 87078 560898 87080
rect 560789 87075 560855 87078
rect 91454 87000 91563 87005
rect 91454 86944 91502 87000
rect 91558 86944 91563 87000
rect 91454 86942 91563 86944
rect 91497 86939 91563 86942
rect 307881 87002 307947 87005
rect 308157 87002 308223 87005
rect 307881 87000 308223 87002
rect 307881 86944 307886 87000
rect 307942 86944 308162 87000
rect 308218 86944 308223 87000
rect 307881 86942 308223 86944
rect 307881 86939 307947 86942
rect 308157 86939 308223 86942
rect 308893 87002 308959 87005
rect 309077 87002 309143 87005
rect 308893 87000 309143 87002
rect 308893 86944 308898 87000
rect 308954 86944 309082 87000
rect 309138 86944 309143 87000
rect 308893 86942 309143 86944
rect 308893 86939 308959 86942
rect 309077 86939 309143 86942
rect 341185 87002 341251 87005
rect 341369 87002 341435 87005
rect 341185 87000 341435 87002
rect 341185 86944 341190 87000
rect 341246 86944 341374 87000
rect 341430 86944 341435 87000
rect 341185 86942 341435 86944
rect 357886 87000 357995 87005
rect 357886 86944 357934 87000
rect 357990 86944 357995 87000
rect 357886 86942 357995 86944
rect 553846 87000 553955 87005
rect 553846 86944 553894 87000
rect 553950 86944 553955 87000
rect 553846 86942 553955 86944
rect 341185 86939 341251 86942
rect 341369 86939 341435 86942
rect 357929 86939 357995 86942
rect 553889 86939 553955 86942
rect 580661 86050 580727 86053
rect 584016 86050 584496 86080
rect 580661 86048 584496 86050
rect 580661 85992 580666 86048
rect 580722 85992 584496 86048
rect 580661 85990 584496 85992
rect 580661 85987 580727 85990
rect 584016 85960 584496 85990
rect 371821 85506 371887 85509
rect 372005 85506 372071 85509
rect 371821 85504 372071 85506
rect 371821 85448 371826 85504
rect 371882 85448 372010 85504
rect 372066 85448 372071 85504
rect 371821 85446 372071 85448
rect 371821 85443 371887 85446
rect 372005 85443 372071 85446
rect 242745 77346 242811 77349
rect 242929 77346 242995 77349
rect 242745 77344 242995 77346
rect 242745 77288 242750 77344
rect 242806 77288 242934 77344
rect 242990 77288 242995 77344
rect 242745 77286 242995 77288
rect 242745 77283 242811 77286
rect 242929 77283 242995 77286
rect 328213 77346 328279 77349
rect 328397 77346 328463 77349
rect 328213 77344 328463 77346
rect 328213 77288 328218 77344
rect 328274 77288 328402 77344
rect 328458 77288 328463 77344
rect 328213 77286 328463 77288
rect 328213 77283 328279 77286
rect 328397 77283 328463 77286
rect 331065 77346 331131 77349
rect 331249 77346 331315 77349
rect 331065 77344 331315 77346
rect 331065 77288 331070 77344
rect 331126 77288 331254 77344
rect 331310 77288 331315 77344
rect 331065 77286 331315 77288
rect 331065 77283 331131 77286
rect 331249 77283 331315 77286
rect 345550 75850 345556 75852
rect 1110 75790 345556 75850
rect 496 75306 976 75336
rect 1110 75306 1170 75790
rect 345550 75788 345556 75790
rect 345620 75788 345626 75852
rect 496 75246 1170 75306
rect 496 75216 976 75246
rect 236254 70348 236260 70412
rect 236324 70410 236330 70412
rect 584016 70410 584496 70440
rect 236324 70350 584496 70410
rect 236324 70348 236330 70350
rect 584016 70320 584496 70350
rect 552325 67690 552391 67693
rect 552509 67690 552575 67693
rect 552325 67688 552575 67690
rect 552325 67632 552330 67688
rect 552386 67632 552514 67688
rect 552570 67632 552575 67688
rect 552325 67630 552575 67632
rect 552325 67627 552391 67630
rect 552509 67627 552575 67630
rect 279729 64970 279795 64973
rect 280005 64970 280071 64973
rect 279729 64968 280071 64970
rect 279729 64912 279734 64968
rect 279790 64912 280010 64968
rect 280066 64912 280071 64968
rect 279729 64910 280071 64912
rect 279729 64907 279795 64910
rect 280005 64907 280071 64910
rect 276417 62114 276483 62117
rect 276601 62114 276667 62117
rect 276417 62112 276667 62114
rect 276417 62056 276422 62112
rect 276478 62056 276606 62112
rect 276662 62056 276667 62112
rect 276417 62054 276667 62056
rect 276417 62051 276483 62054
rect 276601 62051 276667 62054
rect 496 58578 976 58608
rect 3637 58578 3703 58581
rect 496 58576 3703 58578
rect 496 58520 3642 58576
rect 3698 58520 3703 58576
rect 496 58518 3703 58520
rect 496 58488 976 58518
rect 3637 58515 3703 58518
rect 328397 58170 328463 58173
rect 328262 58168 328463 58170
rect 328262 58112 328402 58168
rect 328458 58112 328463 58168
rect 328262 58110 328463 58112
rect 328262 58034 328322 58110
rect 328397 58107 328463 58110
rect 328397 58034 328463 58037
rect 328262 58032 328463 58034
rect 328262 57976 328402 58032
rect 328458 57976 328463 58032
rect 328262 57974 328463 57976
rect 328397 57971 328463 57974
rect 319841 56538 319907 56541
rect 320117 56538 320183 56541
rect 319841 56536 320183 56538
rect 319841 56480 319846 56536
rect 319902 56480 320122 56536
rect 320178 56480 320183 56536
rect 319841 56478 320183 56480
rect 319841 56475 319907 56478
rect 320117 56475 320183 56478
rect 580753 54770 580819 54773
rect 584016 54770 584496 54800
rect 580753 54768 584496 54770
rect 580753 54712 580758 54768
rect 580814 54712 584496 54768
rect 580753 54710 584496 54712
rect 580753 54707 580819 54710
rect 584016 54680 584496 54710
rect 272921 52458 272987 52461
rect 273289 52458 273355 52461
rect 272921 52456 273355 52458
rect 272921 52400 272926 52456
rect 272982 52400 273294 52456
rect 273350 52400 273355 52456
rect 272921 52398 273355 52400
rect 272921 52395 272987 52398
rect 273289 52395 273355 52398
rect 239249 51098 239315 51101
rect 239433 51098 239499 51101
rect 239249 51096 239499 51098
rect 239249 51040 239254 51096
rect 239310 51040 239438 51096
rect 239494 51040 239499 51096
rect 239249 51038 239499 51040
rect 239249 51035 239315 51038
rect 239433 51035 239499 51038
rect 135657 48650 135723 48653
rect 135614 48648 135723 48650
rect 135614 48592 135662 48648
rect 135718 48592 135723 48648
rect 135614 48587 135723 48592
rect 560789 48650 560855 48653
rect 560789 48648 560898 48650
rect 560789 48592 560794 48648
rect 560850 48592 560898 48648
rect 560789 48587 560898 48592
rect 135614 48517 135674 48587
rect 560838 48517 560898 48587
rect 135614 48512 135723 48517
rect 135614 48456 135662 48512
rect 135718 48456 135723 48512
rect 135614 48454 135723 48456
rect 135657 48451 135723 48454
rect 560789 48512 560898 48517
rect 560789 48456 560794 48512
rect 560850 48456 560898 48512
rect 560789 48454 560898 48456
rect 560789 48451 560855 48454
rect 225173 48378 225239 48381
rect 225357 48378 225423 48381
rect 225173 48376 225423 48378
rect 225173 48320 225178 48376
rect 225234 48320 225362 48376
rect 225418 48320 225423 48376
rect 225173 48318 225423 48320
rect 225173 48315 225239 48318
rect 225357 48315 225423 48318
rect 340909 48378 340975 48381
rect 341093 48378 341159 48381
rect 340909 48376 341159 48378
rect 340909 48320 340914 48376
rect 340970 48320 341098 48376
rect 341154 48320 341159 48376
rect 340909 48318 341159 48320
rect 340909 48315 340975 48318
rect 341093 48315 341159 48318
rect 553889 48378 553955 48381
rect 554073 48378 554139 48381
rect 553889 48376 554139 48378
rect 553889 48320 553894 48376
rect 553950 48320 554078 48376
rect 554134 48320 554139 48376
rect 553889 48318 554139 48320
rect 553889 48315 553955 48318
rect 554073 48315 554139 48318
rect 235385 48242 235451 48245
rect 235342 48240 235451 48242
rect 235342 48184 235390 48240
rect 235446 48184 235451 48240
rect 235342 48179 235451 48184
rect 235342 48106 235402 48179
rect 235661 48106 235727 48109
rect 235342 48104 235727 48106
rect 235342 48048 235666 48104
rect 235722 48048 235727 48104
rect 235342 48046 235727 48048
rect 235661 48043 235727 48046
rect 3913 42802 3979 42805
rect 346838 42802 346844 42804
rect 3913 42800 346844 42802
rect 3913 42744 3918 42800
rect 3974 42744 346844 42800
rect 3913 42742 346844 42744
rect 3913 42739 3979 42742
rect 346838 42740 346844 42742
rect 346908 42740 346914 42804
rect 496 41850 976 41880
rect 3913 41850 3979 41853
rect 496 41848 3979 41850
rect 496 41792 3918 41848
rect 3974 41792 3979 41848
rect 496 41790 3979 41792
rect 496 41760 976 41790
rect 3913 41787 3979 41790
rect 337229 39266 337295 39269
rect 346654 39266 346660 39268
rect 327526 39206 337154 39266
rect 327526 39132 327586 39206
rect 327518 39068 327524 39132
rect 327588 39068 327594 39132
rect 232206 38932 232212 38996
rect 232276 38994 232282 38996
rect 317766 38994 317772 38996
rect 232276 38934 244970 38994
rect 232276 38932 232282 38934
rect 244910 38722 244970 38934
rect 284102 38934 288946 38994
rect 261053 38722 261119 38725
rect 244910 38720 261119 38722
rect 244910 38664 261058 38720
rect 261114 38664 261119 38720
rect 244910 38662 261119 38664
rect 261053 38659 261119 38662
rect 268137 38722 268203 38725
rect 284102 38722 284162 38934
rect 288886 38858 288946 38934
rect 308206 38934 317772 38994
rect 298589 38858 298655 38861
rect 288886 38856 298655 38858
rect 288886 38800 298594 38856
rect 298650 38800 298655 38856
rect 288886 38798 298655 38800
rect 298589 38795 298655 38798
rect 308206 38725 308266 38934
rect 317766 38932 317772 38934
rect 317836 38932 317842 38996
rect 337094 38994 337154 39206
rect 337229 39264 346660 39266
rect 337229 39208 337234 39264
rect 337290 39208 346660 39264
rect 337229 39206 346660 39208
rect 337229 39203 337295 39206
rect 346654 39204 346660 39206
rect 346724 39204 346730 39268
rect 584016 39130 584496 39160
rect 583838 39070 584496 39130
rect 337229 38994 337295 38997
rect 337094 38992 337295 38994
rect 337094 38936 337234 38992
rect 337290 38936 337295 38992
rect 337094 38934 337295 38936
rect 337229 38931 337295 38934
rect 346838 38932 346844 38996
rect 346908 38994 346914 38996
rect 356590 38994 356596 38996
rect 346908 38934 356596 38994
rect 346908 38932 346914 38934
rect 356590 38932 356596 38934
rect 356660 38932 356666 38996
rect 406137 38994 406203 38997
rect 406137 38992 413146 38994
rect 406137 38936 406142 38992
rect 406198 38936 413146 38992
rect 406137 38934 413146 38936
rect 406137 38931 406203 38934
rect 366117 38858 366183 38861
rect 370257 38858 370323 38861
rect 366117 38856 370323 38858
rect 366117 38800 366122 38856
rect 366178 38800 370262 38856
rect 370318 38800 370323 38856
rect 366117 38798 370323 38800
rect 366117 38795 366183 38798
rect 370257 38795 370323 38798
rect 382033 38858 382099 38861
rect 389577 38858 389643 38861
rect 399237 38858 399303 38861
rect 382033 38856 389643 38858
rect 382033 38800 382038 38856
rect 382094 38800 389582 38856
rect 389638 38800 389643 38856
rect 382033 38798 389643 38800
rect 382033 38795 382099 38798
rect 389577 38795 389643 38798
rect 396526 38856 399303 38858
rect 396526 38800 399242 38856
rect 399298 38800 399303 38856
rect 396526 38798 399303 38800
rect 413086 38858 413146 38934
rect 422838 38934 432466 38994
rect 413086 38798 422714 38858
rect 308157 38722 308266 38725
rect 268137 38720 284162 38722
rect 268137 38664 268142 38720
rect 268198 38664 284162 38720
rect 268137 38662 284162 38664
rect 308076 38720 308266 38722
rect 308076 38664 308162 38720
rect 308218 38664 308266 38720
rect 308076 38662 308266 38664
rect 268137 38659 268203 38662
rect 308157 38659 308223 38662
rect 317766 38660 317772 38724
rect 317836 38722 317842 38724
rect 327518 38722 327524 38724
rect 317836 38662 327524 38722
rect 317836 38660 317842 38662
rect 327518 38660 327524 38662
rect 327588 38660 327594 38724
rect 346654 38660 346660 38724
rect 346724 38722 346730 38724
rect 346838 38722 346844 38724
rect 346724 38662 346844 38722
rect 346724 38660 346730 38662
rect 346838 38660 346844 38662
rect 346908 38660 346914 38724
rect 370441 38722 370507 38725
rect 377341 38722 377407 38725
rect 370441 38720 377407 38722
rect 370441 38664 370446 38720
rect 370502 38664 377346 38720
rect 377402 38664 377407 38720
rect 370441 38662 377407 38664
rect 370441 38659 370507 38662
rect 377341 38659 377407 38662
rect 389761 38722 389827 38725
rect 396526 38722 396586 38798
rect 399237 38795 399303 38798
rect 389761 38720 396586 38722
rect 389761 38664 389766 38720
rect 389822 38664 396586 38720
rect 389761 38662 396586 38664
rect 422654 38722 422714 38798
rect 422838 38722 422898 38934
rect 432406 38858 432466 38934
rect 442158 38934 451786 38994
rect 432406 38798 442034 38858
rect 422654 38662 422898 38722
rect 441974 38722 442034 38798
rect 442158 38722 442218 38934
rect 451726 38858 451786 38934
rect 461478 38934 471106 38994
rect 451726 38798 461354 38858
rect 441974 38662 442218 38722
rect 461294 38722 461354 38798
rect 461478 38722 461538 38934
rect 471046 38858 471106 38934
rect 480798 38934 490426 38994
rect 471046 38798 480674 38858
rect 461294 38662 461538 38722
rect 480614 38722 480674 38798
rect 480798 38722 480858 38934
rect 490366 38858 490426 38934
rect 500118 38934 509746 38994
rect 490366 38798 499994 38858
rect 480614 38662 480858 38722
rect 499934 38722 499994 38798
rect 500118 38722 500178 38934
rect 509686 38858 509746 38934
rect 519438 38934 529066 38994
rect 509686 38798 519314 38858
rect 499934 38662 500178 38722
rect 519254 38722 519314 38798
rect 519438 38722 519498 38934
rect 529006 38858 529066 38934
rect 538758 38934 544338 38994
rect 529006 38798 538634 38858
rect 519254 38662 519498 38722
rect 538574 38722 538634 38798
rect 538758 38722 538818 38934
rect 538574 38662 538818 38722
rect 544278 38722 544338 38934
rect 551078 38932 551084 38996
rect 551148 38994 551154 38996
rect 551148 38934 567706 38994
rect 551148 38932 551154 38934
rect 567646 38858 567706 38934
rect 583838 38858 583898 39070
rect 584016 39040 584496 39070
rect 567646 38798 577274 38858
rect 551078 38722 551084 38724
rect 544278 38662 551084 38722
rect 389761 38659 389827 38662
rect 551078 38660 551084 38662
rect 551148 38660 551154 38724
rect 577214 38722 577274 38798
rect 577398 38798 583898 38858
rect 577398 38722 577458 38798
rect 577214 38662 577458 38722
rect 356590 38524 356596 38588
rect 356660 38586 356666 38588
rect 366117 38586 366183 38589
rect 356660 38584 366183 38586
rect 356660 38528 366122 38584
rect 366178 38528 366183 38584
rect 356660 38526 366183 38528
rect 356660 38524 356666 38526
rect 366117 38523 366183 38526
rect 273013 33282 273079 33285
rect 273197 33282 273263 33285
rect 273013 33280 273263 33282
rect 273013 33224 273018 33280
rect 273074 33224 273202 33280
rect 273258 33224 273263 33280
rect 273013 33222 273263 33224
rect 273013 33219 273079 33222
rect 273197 33219 273263 33222
rect 392521 29202 392587 29205
rect 392294 29200 392587 29202
rect 392294 29144 392526 29200
rect 392582 29144 392587 29200
rect 392294 29142 392587 29144
rect 392294 29066 392354 29142
rect 392521 29139 392587 29142
rect 392429 29066 392495 29069
rect 392294 29064 392495 29066
rect 392294 29008 392434 29064
rect 392490 29008 392495 29064
rect 392294 29006 392495 29008
rect 392429 29003 392495 29006
rect 285065 28930 285131 28933
rect 285249 28930 285315 28933
rect 285065 28928 285315 28930
rect 285065 28872 285070 28928
rect 285126 28872 285254 28928
rect 285310 28872 285315 28928
rect 285065 28870 285315 28872
rect 285065 28867 285131 28870
rect 285249 28867 285315 28870
rect 496 25122 976 25152
rect 3913 25122 3979 25125
rect 496 25120 3979 25122
rect 496 25064 3918 25120
rect 3974 25064 3979 25120
rect 496 25062 3979 25064
rect 496 25032 976 25062
rect 3913 25059 3979 25062
rect 233494 23428 233500 23492
rect 233564 23490 233570 23492
rect 584016 23490 584496 23520
rect 233564 23430 584496 23490
rect 233564 23428 233570 23430
rect 584016 23400 584496 23430
rect 285065 19274 285131 19277
rect 285341 19274 285407 19277
rect 285065 19272 285407 19274
rect 285065 19216 285070 19272
rect 285126 19216 285346 19272
rect 285402 19216 285407 19272
rect 285065 19214 285407 19216
rect 285065 19211 285131 19214
rect 285341 19211 285407 19214
rect 190213 18050 190279 18053
rect 190397 18050 190463 18053
rect 190213 18048 190463 18050
rect 190213 17992 190218 18048
rect 190274 17992 190402 18048
rect 190458 17992 190463 18048
rect 190213 17990 190463 17992
rect 190213 17987 190279 17990
rect 190397 17987 190463 17990
rect 242561 18050 242627 18053
rect 242745 18050 242811 18053
rect 242561 18048 242811 18050
rect 242561 17992 242566 18048
rect 242622 17992 242750 18048
rect 242806 17992 242811 18048
rect 242561 17990 242811 17992
rect 242561 17987 242627 17990
rect 242745 17987 242811 17990
rect 392337 18050 392403 18053
rect 392613 18050 392679 18053
rect 392337 18048 392679 18050
rect 392337 17992 392342 18048
rect 392398 17992 392618 18048
rect 392674 17992 392679 18048
rect 392337 17990 392679 17992
rect 392337 17987 392403 17990
rect 392613 17987 392679 17990
rect 278441 16554 278507 16557
rect 278625 16554 278691 16557
rect 278441 16552 278691 16554
rect 278441 16496 278446 16552
rect 278502 16496 278630 16552
rect 278686 16496 278691 16552
rect 278441 16494 278691 16496
rect 278441 16491 278507 16494
rect 278625 16491 278691 16494
rect 186809 10706 186875 10709
rect 196377 10706 196443 10709
rect 186809 10704 196443 10706
rect 186809 10648 186814 10704
rect 186870 10648 196382 10704
rect 196438 10648 196443 10704
rect 186809 10646 196443 10648
rect 186809 10643 186875 10646
rect 196377 10643 196443 10646
rect 225449 10706 225515 10709
rect 235017 10706 235083 10709
rect 225449 10704 235083 10706
rect 225449 10648 225454 10704
rect 225510 10648 235022 10704
rect 235078 10648 235083 10704
rect 225449 10646 235083 10648
rect 225449 10643 225515 10646
rect 235017 10643 235083 10646
rect 120477 10570 120543 10573
rect 123513 10570 123579 10573
rect 120477 10568 123579 10570
rect 120477 10512 120482 10568
rect 120538 10512 123518 10568
rect 123574 10512 123579 10568
rect 120477 10510 123579 10512
rect 120477 10507 120543 10510
rect 123513 10507 123579 10510
rect 147801 10570 147867 10573
rect 148445 10570 148511 10573
rect 147801 10568 148511 10570
rect 147801 10512 147806 10568
rect 147862 10512 148450 10568
rect 148506 10512 148511 10568
rect 147801 10510 148511 10512
rect 147801 10507 147867 10510
rect 148445 10507 148511 10510
rect 177241 10570 177307 10573
rect 187085 10570 187151 10573
rect 177241 10568 187151 10570
rect 177241 10512 177246 10568
rect 177302 10512 187090 10568
rect 187146 10512 187151 10568
rect 177241 10510 187151 10512
rect 177241 10507 177307 10510
rect 187085 10507 187151 10510
rect 234649 10570 234715 10573
rect 235385 10570 235451 10573
rect 234649 10568 235451 10570
rect 234649 10512 234654 10568
rect 234710 10512 235390 10568
rect 235446 10512 235451 10568
rect 234649 10510 235451 10512
rect 234649 10507 234715 10510
rect 235385 10507 235451 10510
rect 329869 10570 329935 10573
rect 331617 10570 331683 10573
rect 329869 10568 331683 10570
rect 329869 10512 329874 10568
rect 329930 10512 331622 10568
rect 331678 10512 331683 10568
rect 329869 10510 331683 10512
rect 329869 10507 329935 10510
rect 331617 10507 331683 10510
rect 408989 10570 409055 10573
rect 424169 10570 424235 10573
rect 408989 10568 424235 10570
rect 408989 10512 408994 10568
rect 409050 10512 424174 10568
rect 424230 10512 424235 10568
rect 408989 10510 424235 10512
rect 408989 10507 409055 10510
rect 424169 10507 424235 10510
rect 157829 10434 157895 10437
rect 167857 10434 167923 10437
rect 157829 10432 167923 10434
rect 157829 10376 157834 10432
rect 157890 10376 167862 10432
rect 167918 10376 167923 10432
rect 157829 10374 167923 10376
rect 157829 10371 157895 10374
rect 167857 10371 167923 10374
rect 196469 10434 196535 10437
rect 206313 10434 206379 10437
rect 196469 10432 206379 10434
rect 196469 10376 196474 10432
rect 196530 10376 206318 10432
rect 206374 10376 206379 10432
rect 196469 10374 206379 10376
rect 196469 10371 196535 10374
rect 206313 10371 206379 10374
rect 216157 10434 216223 10437
rect 225633 10434 225699 10437
rect 216157 10432 225699 10434
rect 216157 10376 216162 10432
rect 216218 10376 225638 10432
rect 225694 10376 225699 10432
rect 216157 10374 225699 10376
rect 216157 10371 216223 10374
rect 225633 10371 225699 10374
rect 341461 10434 341527 10437
rect 418741 10434 418807 10437
rect 341461 10432 418807 10434
rect 341461 10376 341466 10432
rect 341522 10376 418746 10432
rect 418802 10376 418807 10432
rect 341461 10374 418807 10376
rect 341461 10371 341527 10374
rect 418741 10371 418807 10374
rect 30685 10298 30751 10301
rect 236581 10298 236647 10301
rect 30685 10296 236647 10298
rect 30685 10240 30690 10296
rect 30746 10240 236586 10296
rect 236642 10240 236647 10296
rect 30685 10238 236647 10240
rect 30685 10235 30751 10238
rect 236581 10235 236647 10238
rect 331249 10298 331315 10301
rect 486453 10298 486519 10301
rect 331249 10296 486519 10298
rect 331249 10240 331254 10296
rect 331310 10240 486458 10296
rect 486514 10240 486519 10296
rect 331249 10238 486519 10240
rect 331249 10235 331315 10238
rect 486453 10235 486519 10238
rect 138233 10162 138299 10165
rect 138601 10162 138667 10165
rect 138233 10160 138667 10162
rect 138233 10104 138238 10160
rect 138294 10104 138606 10160
rect 138662 10104 138667 10160
rect 138233 10102 138667 10104
rect 138233 10099 138299 10102
rect 138601 10099 138667 10102
rect 157461 10162 157527 10165
rect 157829 10162 157895 10165
rect 167765 10162 167831 10165
rect 157461 10160 157895 10162
rect 157461 10104 157466 10160
rect 157522 10104 157834 10160
rect 157890 10104 157895 10160
rect 157461 10102 157895 10104
rect 157461 10099 157527 10102
rect 157829 10099 157895 10102
rect 158246 10160 167831 10162
rect 158246 10104 167770 10160
rect 167826 10104 167831 10160
rect 158246 10102 167831 10104
rect 157553 10026 157619 10029
rect 158246 10026 158306 10102
rect 167765 10099 167831 10102
rect 177190 10100 177196 10164
rect 177260 10162 177266 10164
rect 191777 10162 191843 10165
rect 177260 10160 191843 10162
rect 177260 10104 191782 10160
rect 191838 10104 191843 10160
rect 177260 10102 191843 10104
rect 177260 10100 177266 10102
rect 191777 10099 191843 10102
rect 195917 10162 195983 10165
rect 196469 10162 196535 10165
rect 206313 10162 206379 10165
rect 216157 10162 216223 10165
rect 195917 10160 196535 10162
rect 195917 10104 195922 10160
rect 195978 10104 196474 10160
rect 196530 10104 196535 10160
rect 195917 10102 196535 10104
rect 195917 10099 195983 10102
rect 196469 10099 196535 10102
rect 196702 10102 206146 10162
rect 157553 10024 158306 10026
rect 157553 9968 157558 10024
rect 157614 9968 158306 10024
rect 157553 9966 158306 9968
rect 167489 10026 167555 10029
rect 177006 10026 177012 10028
rect 167489 10024 177012 10026
rect 167489 9968 167494 10024
rect 167550 9968 177012 10024
rect 167489 9966 177012 9968
rect 157553 9963 157619 9966
rect 167489 9963 167555 9966
rect 177006 9964 177012 9966
rect 177076 9964 177082 10028
rect 196009 10026 196075 10029
rect 196702 10026 196762 10102
rect 196009 10024 196762 10026
rect 196009 9968 196014 10024
rect 196070 9968 196762 10024
rect 196009 9966 196762 9968
rect 196009 9963 196075 9966
rect 206086 9890 206146 10102
rect 206313 10160 216223 10162
rect 206313 10104 206318 10160
rect 206374 10104 216162 10160
rect 216218 10104 216223 10160
rect 206313 10102 216223 10104
rect 206313 10099 206379 10102
rect 216157 10099 216223 10102
rect 235017 10162 235083 10165
rect 238513 10162 238579 10165
rect 235017 10160 238579 10162
rect 235017 10104 235022 10160
rect 235078 10104 238518 10160
rect 238574 10104 238579 10160
rect 235017 10102 238579 10104
rect 235017 10099 235083 10102
rect 238513 10099 238579 10102
rect 215789 10026 215855 10029
rect 225633 10026 225699 10029
rect 215789 10024 225699 10026
rect 215789 9968 215794 10024
rect 215850 9968 225638 10024
rect 225694 9968 225699 10024
rect 215789 9966 225699 9968
rect 215789 9963 215855 9966
rect 225633 9963 225699 9966
rect 232441 10026 232507 10029
rect 241917 10026 241983 10029
rect 232441 10024 241983 10026
rect 232441 9968 232446 10024
rect 232502 9968 241922 10024
rect 241978 9968 241983 10024
rect 232441 9966 241983 9968
rect 232441 9963 232507 9966
rect 241917 9963 241983 9966
rect 328397 10026 328463 10029
rect 331617 10026 331683 10029
rect 328397 10024 331683 10026
rect 328397 9968 328402 10024
rect 328458 9968 331622 10024
rect 331678 9968 331683 10024
rect 328397 9966 331683 9968
rect 328397 9963 328463 9966
rect 331617 9963 331683 9966
rect 215973 9890 216039 9893
rect 206086 9888 216039 9890
rect 206086 9832 215978 9888
rect 216034 9832 216039 9888
rect 206086 9830 216039 9832
rect 215973 9827 216039 9830
rect 135289 9754 135355 9757
rect 135473 9754 135539 9757
rect 135289 9752 135539 9754
rect 135289 9696 135294 9752
rect 135350 9696 135478 9752
rect 135534 9696 135539 9752
rect 135289 9694 135539 9696
rect 135289 9691 135355 9694
rect 135473 9691 135539 9694
rect 151849 9754 151915 9757
rect 152033 9754 152099 9757
rect 151849 9752 152099 9754
rect 151849 9696 151854 9752
rect 151910 9696 152038 9752
rect 152094 9696 152099 9752
rect 151849 9694 152099 9696
rect 151849 9691 151915 9694
rect 152033 9691 152099 9694
rect 169697 9754 169763 9757
rect 169881 9754 169947 9757
rect 169697 9752 169947 9754
rect 169697 9696 169702 9752
rect 169758 9696 169886 9752
rect 169942 9696 169947 9752
rect 169697 9694 169947 9696
rect 169697 9691 169763 9694
rect 169881 9691 169947 9694
rect 190397 9754 190463 9757
rect 190581 9754 190647 9757
rect 190397 9752 190647 9754
rect 190397 9696 190402 9752
rect 190458 9696 190586 9752
rect 190642 9696 190647 9752
rect 190397 9694 190647 9696
rect 190397 9691 190463 9694
rect 190581 9691 190647 9694
rect 213949 9754 214015 9757
rect 214501 9754 214567 9757
rect 213949 9752 214567 9754
rect 213949 9696 213954 9752
rect 214010 9696 214506 9752
rect 214562 9696 214567 9752
rect 213949 9694 214567 9696
rect 213949 9691 214015 9694
rect 214501 9691 214567 9694
rect 225081 9754 225147 9757
rect 225265 9754 225331 9757
rect 225081 9752 225331 9754
rect 225081 9696 225086 9752
rect 225142 9696 225270 9752
rect 225326 9696 225331 9752
rect 225081 9694 225331 9696
rect 225081 9691 225147 9694
rect 225265 9691 225331 9694
rect 231889 9754 231955 9757
rect 232165 9754 232231 9757
rect 231889 9752 232231 9754
rect 231889 9696 231894 9752
rect 231950 9696 232170 9752
rect 232226 9696 232231 9752
rect 231889 9694 232231 9696
rect 231889 9691 231955 9694
rect 232165 9691 232231 9694
rect 340725 9754 340791 9757
rect 340909 9754 340975 9757
rect 340725 9752 340975 9754
rect 340725 9696 340730 9752
rect 340786 9696 340914 9752
rect 340970 9696 340975 9752
rect 340725 9694 340975 9696
rect 340725 9691 340791 9694
rect 340909 9691 340975 9694
rect 346889 9754 346955 9757
rect 347073 9754 347139 9757
rect 346889 9752 347139 9754
rect 346889 9696 346894 9752
rect 346950 9696 347078 9752
rect 347134 9696 347139 9752
rect 346889 9694 347139 9696
rect 346889 9691 346955 9694
rect 347073 9691 347139 9694
rect 351305 9754 351371 9757
rect 351581 9754 351647 9757
rect 351305 9752 351647 9754
rect 351305 9696 351310 9752
rect 351366 9696 351586 9752
rect 351642 9696 351647 9752
rect 351305 9694 351647 9696
rect 351305 9691 351371 9694
rect 351581 9691 351647 9694
rect 385989 9754 386055 9757
rect 386357 9754 386423 9757
rect 385989 9752 386423 9754
rect 385989 9696 385994 9752
rect 386050 9696 386362 9752
rect 386418 9696 386423 9752
rect 385989 9694 386423 9696
rect 385989 9691 386055 9694
rect 386357 9691 386423 9694
rect 413221 9754 413287 9757
rect 413773 9754 413839 9757
rect 413221 9752 413839 9754
rect 413221 9696 413226 9752
rect 413282 9696 413778 9752
rect 413834 9696 413839 9752
rect 413221 9694 413839 9696
rect 413221 9691 413287 9694
rect 413773 9691 413839 9694
rect 3913 9618 3979 9621
rect 348310 9618 348316 9620
rect 3913 9616 348316 9618
rect 3913 9560 3918 9616
rect 3974 9560 348316 9616
rect 3913 9558 348316 9560
rect 3913 9555 3979 9558
rect 348310 9556 348316 9558
rect 348380 9556 348386 9620
rect 169513 9482 169579 9485
rect 170157 9482 170223 9485
rect 169513 9480 170223 9482
rect 169513 9424 169518 9480
rect 169574 9424 170162 9480
rect 170218 9424 170223 9480
rect 169513 9422 170223 9424
rect 169513 9419 169579 9422
rect 170157 9419 170223 9422
rect 347993 9482 348059 9485
rect 350845 9482 350911 9485
rect 347993 9480 350911 9482
rect 347993 9424 347998 9480
rect 348054 9424 350850 9480
rect 350906 9424 350911 9480
rect 347993 9422 350911 9424
rect 347993 9419 348059 9422
rect 350845 9419 350911 9422
rect 240077 9346 240143 9349
rect 244861 9346 244927 9349
rect 240077 9344 244927 9346
rect 240077 9288 240082 9344
rect 240138 9288 244866 9344
rect 244922 9288 244927 9344
rect 240077 9286 244927 9288
rect 240077 9283 240143 9286
rect 244861 9283 244927 9286
rect 237777 9210 237843 9213
rect 244861 9210 244927 9213
rect 237777 9208 244927 9210
rect 237777 9152 237782 9208
rect 237838 9152 244866 9208
rect 244922 9152 244927 9208
rect 237777 9150 244927 9152
rect 237777 9147 237843 9150
rect 244861 9147 244927 9150
rect 254245 9210 254311 9213
rect 254521 9210 254587 9213
rect 254245 9208 254587 9210
rect 254245 9152 254250 9208
rect 254306 9152 254526 9208
rect 254582 9152 254587 9208
rect 254245 9150 254587 9152
rect 254245 9147 254311 9150
rect 254521 9147 254587 9150
rect 349281 9210 349347 9213
rect 351121 9210 351187 9213
rect 349281 9208 351187 9210
rect 349281 9152 349286 9208
rect 349342 9152 351126 9208
rect 351182 9152 351187 9208
rect 349281 9150 351187 9152
rect 349281 9147 349347 9150
rect 351121 9147 351187 9150
rect 351213 9074 351279 9077
rect 356641 9074 356707 9077
rect 351213 9072 356707 9074
rect 351213 9016 351218 9072
rect 351274 9016 356646 9072
rect 356702 9016 356707 9072
rect 351213 9014 356707 9016
rect 351213 9011 351279 9014
rect 356641 9011 356707 9014
rect 229405 8938 229471 8941
rect 234925 8938 234991 8941
rect 229405 8936 234991 8938
rect 229405 8880 229410 8936
rect 229466 8880 234930 8936
rect 234986 8880 234991 8936
rect 229405 8878 234991 8880
rect 229405 8875 229471 8878
rect 234925 8875 234991 8878
rect 254429 8938 254495 8941
rect 254889 8938 254955 8941
rect 254429 8936 254955 8938
rect 254429 8880 254434 8936
rect 254490 8880 254894 8936
rect 254950 8880 254955 8936
rect 254429 8878 254955 8880
rect 254429 8875 254495 8878
rect 254889 8875 254955 8878
rect 350937 8938 351003 8941
rect 581581 8938 581647 8941
rect 350937 8936 581647 8938
rect 350937 8880 350942 8936
rect 350998 8880 581586 8936
rect 581642 8880 581647 8936
rect 350937 8878 581647 8880
rect 350937 8875 351003 8878
rect 581581 8875 581647 8878
rect 225817 8802 225883 8805
rect 235017 8802 235083 8805
rect 225817 8800 235083 8802
rect 225817 8744 225822 8800
rect 225878 8744 235022 8800
rect 235078 8744 235083 8800
rect 225817 8742 235083 8744
rect 225817 8739 225883 8742
rect 235017 8739 235083 8742
rect 496 8394 976 8424
rect 3913 8394 3979 8397
rect 496 8392 3979 8394
rect 496 8336 3918 8392
rect 3974 8336 3979 8392
rect 496 8334 3979 8336
rect 496 8304 976 8334
rect 3913 8331 3979 8334
rect 351029 8394 351095 8397
rect 360229 8394 360295 8397
rect 351029 8392 360295 8394
rect 351029 8336 351034 8392
rect 351090 8336 360234 8392
rect 360290 8336 360295 8392
rect 351029 8334 360295 8336
rect 351029 8331 351095 8334
rect 360229 8331 360295 8334
rect 361149 8394 361215 8397
rect 363909 8394 363975 8397
rect 361149 8392 363975 8394
rect 361149 8336 361154 8392
rect 361210 8336 363914 8392
rect 363970 8336 363975 8392
rect 361149 8334 363975 8336
rect 361149 8331 361215 8334
rect 363909 8331 363975 8334
rect 340817 8258 340883 8261
rect 341277 8258 341343 8261
rect 340817 8256 341343 8258
rect 340817 8200 340822 8256
rect 340878 8200 341282 8256
rect 341338 8200 341343 8256
rect 340817 8198 341343 8200
rect 340817 8195 340883 8198
rect 341277 8195 341343 8198
rect 340725 8122 340791 8125
rect 341369 8122 341435 8125
rect 340725 8120 341435 8122
rect 340725 8064 340730 8120
rect 340786 8064 341374 8120
rect 341430 8064 341435 8120
rect 340725 8062 341435 8064
rect 340725 8059 340791 8062
rect 341369 8059 341435 8062
rect 215789 7986 215855 7989
rect 224621 7986 224687 7989
rect 225265 7986 225331 7989
rect 215789 7984 216450 7986
rect 215789 7928 215794 7984
rect 215850 7928 216450 7984
rect 215789 7926 216450 7928
rect 215789 7923 215855 7926
rect 196285 7850 196351 7853
rect 216390 7850 216450 7926
rect 224621 7984 225331 7986
rect 224621 7928 224626 7984
rect 224682 7928 225270 7984
rect 225326 7928 225331 7984
rect 224621 7926 225331 7928
rect 224621 7923 224687 7926
rect 225265 7923 225331 7926
rect 225449 7986 225515 7989
rect 234005 7986 234071 7989
rect 225449 7984 234071 7986
rect 225449 7928 225454 7984
rect 225510 7928 234010 7984
rect 234066 7928 234071 7984
rect 225449 7926 234071 7928
rect 225449 7923 225515 7926
rect 234005 7923 234071 7926
rect 231337 7850 231403 7853
rect 196285 7848 216082 7850
rect 196285 7792 196290 7848
rect 196346 7792 216082 7848
rect 196285 7790 216082 7792
rect 216390 7848 231403 7850
rect 216390 7792 231342 7848
rect 231398 7792 231403 7848
rect 216390 7790 231403 7792
rect 196285 7787 196351 7790
rect 193617 7714 193683 7717
rect 215881 7714 215947 7717
rect 193617 7712 215947 7714
rect 193617 7656 193622 7712
rect 193678 7656 215886 7712
rect 215942 7656 215947 7712
rect 193617 7654 215947 7656
rect 193617 7651 193683 7654
rect 215881 7651 215947 7654
rect 216022 7578 216082 7790
rect 231337 7787 231403 7790
rect 350845 7850 350911 7853
rect 361241 7850 361307 7853
rect 350845 7848 361307 7850
rect 350845 7792 350850 7848
rect 350906 7792 361246 7848
rect 361302 7792 361307 7848
rect 350845 7790 361307 7792
rect 350845 7787 350911 7790
rect 361241 7787 361307 7790
rect 583881 7850 583947 7853
rect 584016 7850 584496 7880
rect 583881 7848 584496 7850
rect 583881 7792 583886 7848
rect 583942 7792 584496 7848
rect 583881 7790 584496 7792
rect 583881 7787 583947 7790
rect 584016 7760 584496 7790
rect 225265 7714 225331 7717
rect 225541 7714 225607 7717
rect 225265 7712 225607 7714
rect 225265 7656 225270 7712
rect 225326 7656 225546 7712
rect 225602 7656 225607 7712
rect 225265 7654 225607 7656
rect 225265 7651 225331 7654
rect 225541 7651 225607 7654
rect 350661 7714 350727 7717
rect 356181 7714 356247 7717
rect 350661 7712 356247 7714
rect 350661 7656 350666 7712
rect 350722 7656 356186 7712
rect 356242 7656 356247 7712
rect 350661 7654 356247 7656
rect 350661 7651 350727 7654
rect 356181 7651 356247 7654
rect 370349 7714 370415 7717
rect 399421 7714 399487 7717
rect 370349 7712 399487 7714
rect 370349 7656 370354 7712
rect 370410 7656 399426 7712
rect 399482 7656 399487 7712
rect 370349 7654 399487 7656
rect 370349 7651 370415 7654
rect 399421 7651 399487 7654
rect 409173 7714 409239 7717
rect 438245 7714 438311 7717
rect 409173 7712 438311 7714
rect 409173 7656 409178 7712
rect 409234 7656 438250 7712
rect 438306 7656 438311 7712
rect 409173 7654 438311 7656
rect 409173 7651 409239 7654
rect 438245 7651 438311 7654
rect 225357 7578 225423 7581
rect 216022 7576 225423 7578
rect 216022 7520 225362 7576
rect 225418 7520 225423 7576
rect 216022 7518 225423 7520
rect 225357 7515 225423 7518
rect 250238 7516 250244 7580
rect 250308 7578 250314 7580
rect 255073 7578 255139 7581
rect 250308 7576 255139 7578
rect 250308 7520 255078 7576
rect 255134 7520 255139 7576
rect 250308 7518 255139 7520
rect 250308 7516 250314 7518
rect 255073 7515 255139 7518
rect 501398 7516 501404 7580
rect 501468 7578 501474 7580
rect 511017 7578 511083 7581
rect 501468 7576 511083 7578
rect 501468 7520 511022 7576
rect 511078 7520 511083 7576
rect 501468 7518 511083 7520
rect 501468 7516 501474 7518
rect 511017 7515 511083 7518
rect 232441 7442 232507 7445
rect 338149 7442 338215 7445
rect 343393 7442 343459 7445
rect 232441 7440 242026 7442
rect 232441 7384 232446 7440
rect 232502 7384 242026 7440
rect 232441 7382 242026 7384
rect 232441 7379 232507 7382
rect 241966 7306 242026 7382
rect 338149 7440 343459 7442
rect 338149 7384 338154 7440
rect 338210 7384 343398 7440
rect 343454 7384 343459 7440
rect 338149 7382 343459 7384
rect 338149 7379 338215 7382
rect 343393 7379 343459 7382
rect 346981 7442 347047 7445
rect 356457 7442 356523 7445
rect 346981 7440 356523 7442
rect 346981 7384 346986 7440
rect 347042 7384 356462 7440
rect 356518 7384 356523 7440
rect 346981 7382 356523 7384
rect 346981 7379 347047 7382
rect 356457 7379 356523 7382
rect 393758 7380 393764 7444
rect 393828 7442 393834 7444
rect 411657 7442 411723 7445
rect 413037 7442 413103 7445
rect 393828 7382 403210 7442
rect 393828 7380 393834 7382
rect 250238 7306 250244 7308
rect 241966 7246 250244 7306
rect 250238 7244 250244 7246
rect 250308 7244 250314 7308
rect 308198 7244 308204 7308
rect 308268 7306 308274 7308
rect 308268 7246 317834 7306
rect 308268 7244 308274 7246
rect 229589 7170 229655 7173
rect 232349 7170 232415 7173
rect 229589 7168 232415 7170
rect 229589 7112 229594 7168
rect 229650 7112 232354 7168
rect 232410 7112 232415 7168
rect 229589 7110 232415 7112
rect 229589 7107 229655 7110
rect 232349 7107 232415 7110
rect 255073 7170 255139 7173
rect 259949 7170 260015 7173
rect 292926 7170 292932 7172
rect 255073 7168 260015 7170
rect 255073 7112 255078 7168
rect 255134 7112 259954 7168
rect 260010 7112 260015 7168
rect 255073 7110 260015 7112
rect 255073 7107 255139 7110
rect 259949 7107 260015 7110
rect 288886 7110 292932 7170
rect 269517 7034 269583 7037
rect 288886 7034 288946 7110
rect 292926 7108 292932 7110
rect 292996 7108 293002 7172
rect 293110 7108 293116 7172
rect 293180 7170 293186 7172
rect 299918 7170 299924 7172
rect 293180 7110 299924 7170
rect 293180 7108 293186 7110
rect 299918 7108 299924 7110
rect 299988 7108 299994 7172
rect 269517 7032 288946 7034
rect 269517 6976 269522 7032
rect 269578 6976 288946 7032
rect 269517 6974 288946 6976
rect 317774 7034 317834 7246
rect 319246 7246 328920 7306
rect 319246 7034 319306 7246
rect 317774 6974 319306 7034
rect 328860 7034 328920 7246
rect 366166 7246 375794 7306
rect 366166 7037 366226 7246
rect 375734 7172 375794 7246
rect 375726 7108 375732 7172
rect 375796 7108 375802 7172
rect 403150 7170 403210 7382
rect 411657 7440 413103 7442
rect 411657 7384 411662 7440
rect 411718 7384 413042 7440
rect 413098 7384 413103 7440
rect 411657 7382 413103 7384
rect 411657 7379 411723 7382
rect 413037 7379 413103 7382
rect 537278 7380 537284 7444
rect 537348 7442 537354 7444
rect 546897 7442 546963 7445
rect 537348 7440 546963 7442
rect 537348 7384 546902 7440
rect 546958 7384 546963 7440
rect 537348 7382 546963 7384
rect 537348 7380 537354 7382
rect 546897 7379 546963 7382
rect 501398 7306 501404 7308
rect 495886 7246 501404 7306
rect 411657 7170 411723 7173
rect 403150 7168 411723 7170
rect 403150 7112 411662 7168
rect 411718 7112 411723 7168
rect 403150 7110 411723 7112
rect 411657 7107 411723 7110
rect 428953 7170 429019 7173
rect 443438 7170 443444 7172
rect 428953 7168 443444 7170
rect 428953 7112 428958 7168
rect 429014 7112 443444 7168
rect 428953 7110 443444 7112
rect 428953 7107 429019 7110
rect 443438 7108 443444 7110
rect 443508 7108 443514 7172
rect 473849 7170 473915 7173
rect 474217 7170 474283 7173
rect 473849 7168 474283 7170
rect 473849 7112 473854 7168
rect 473910 7112 474222 7168
rect 474278 7112 474283 7168
rect 473849 7110 474283 7112
rect 473849 7107 473915 7110
rect 474217 7107 474283 7110
rect 346654 7034 346660 7036
rect 328860 6974 346660 7034
rect 269517 6971 269583 6974
rect 346654 6972 346660 6974
rect 346724 6972 346730 7036
rect 346838 6972 346844 7036
rect 346908 7034 346914 7036
rect 366117 7034 366226 7037
rect 346908 6974 356474 7034
rect 366036 7032 366226 7034
rect 366036 6976 366122 7032
rect 366178 6976 366226 7032
rect 366036 6974 366226 6976
rect 389853 7034 389919 7037
rect 393758 7034 393764 7036
rect 389853 7032 393764 7034
rect 389853 6976 389858 7032
rect 389914 6976 393764 7032
rect 389853 6974 393764 6976
rect 346908 6972 346914 6974
rect 300102 6836 300108 6900
rect 300172 6898 300178 6900
rect 308198 6898 308204 6900
rect 300172 6838 308204 6898
rect 300172 6836 300178 6838
rect 308198 6836 308204 6838
rect 308268 6836 308274 6900
rect 356414 6898 356474 6974
rect 366117 6971 366183 6974
rect 389853 6971 389919 6974
rect 393758 6972 393764 6974
rect 393828 6972 393834 7036
rect 413037 7034 413103 7037
rect 424077 7034 424143 7037
rect 453241 7034 453307 7037
rect 413037 7032 424143 7034
rect 413037 6976 413042 7032
rect 413098 6976 424082 7032
rect 424138 6976 424143 7032
rect 413037 6974 424143 6976
rect 413037 6971 413103 6974
rect 424077 6971 424143 6974
rect 453014 7032 453307 7034
rect 453014 6976 453246 7032
rect 453302 6976 453307 7032
rect 453014 6974 453307 6976
rect 356414 6838 356658 6898
rect 259949 6762 260015 6765
rect 269517 6762 269583 6765
rect 259949 6760 269583 6762
rect 259949 6704 259954 6760
rect 260010 6704 269522 6760
rect 269578 6704 269583 6760
rect 259949 6702 269583 6704
rect 259949 6699 260015 6702
rect 269517 6699 269583 6702
rect 346654 6700 346660 6764
rect 346724 6762 346730 6764
rect 346838 6762 346844 6764
rect 346724 6702 346844 6762
rect 346724 6700 346730 6702
rect 346838 6700 346844 6702
rect 346908 6700 346914 6764
rect 235109 6626 235175 6629
rect 240997 6626 241063 6629
rect 235109 6624 241063 6626
rect 235109 6568 235114 6624
rect 235170 6568 241002 6624
rect 241058 6568 241063 6624
rect 235109 6566 241063 6568
rect 356598 6626 356658 6838
rect 375910 6836 375916 6900
rect 375980 6898 375986 6900
rect 382718 6898 382724 6900
rect 375980 6838 382724 6898
rect 375980 6836 375986 6838
rect 382718 6836 382724 6838
rect 382788 6836 382794 6900
rect 443438 6836 443444 6900
rect 443508 6898 443514 6900
rect 453014 6898 453074 6974
rect 453241 6971 453307 6974
rect 462717 7034 462783 7037
rect 480749 7034 480815 7037
rect 462717 7032 480815 7034
rect 462717 6976 462722 7032
rect 462778 6976 480754 7032
rect 480810 6976 480815 7032
rect 462717 6974 480815 6976
rect 462717 6971 462783 6974
rect 480749 6971 480815 6974
rect 483509 7034 483575 7037
rect 495886 7034 495946 7246
rect 501398 7244 501404 7246
rect 501468 7244 501474 7308
rect 511017 7170 511083 7173
rect 534661 7170 534727 7173
rect 537278 7170 537284 7172
rect 511017 7168 511218 7170
rect 511017 7112 511022 7168
rect 511078 7112 511218 7168
rect 511017 7110 511218 7112
rect 511017 7107 511083 7110
rect 483509 7032 495946 7034
rect 483509 6976 483514 7032
rect 483570 6976 495946 7032
rect 483509 6974 495946 6976
rect 483509 6971 483575 6974
rect 443508 6838 453074 6898
rect 511158 6898 511218 7110
rect 534661 7168 537284 7170
rect 534661 7112 534666 7168
rect 534722 7112 537284 7168
rect 534661 7110 537284 7112
rect 534661 7107 534727 7110
rect 537278 7108 537284 7110
rect 537348 7108 537354 7172
rect 558029 7170 558095 7173
rect 553662 7168 558095 7170
rect 553662 7112 558034 7168
rect 558090 7112 558095 7168
rect 553662 7110 558095 7112
rect 520677 7034 520743 7037
rect 534477 7034 534543 7037
rect 520677 7032 534543 7034
rect 520677 6976 520682 7032
rect 520738 6976 534482 7032
rect 534538 6976 534543 7032
rect 520677 6974 534543 6976
rect 520677 6971 520743 6974
rect 534477 6971 534543 6974
rect 546897 7034 546963 7037
rect 553662 7034 553722 7110
rect 558029 7107 558095 7110
rect 578637 7170 578703 7173
rect 583881 7170 583947 7173
rect 578637 7168 583947 7170
rect 578637 7112 578642 7168
rect 578698 7112 583886 7168
rect 583942 7112 583947 7168
rect 578637 7110 583947 7112
rect 578637 7107 578703 7110
rect 583881 7107 583947 7110
rect 546897 7032 553722 7034
rect 546897 6976 546902 7032
rect 546958 6976 553722 7032
rect 546897 6974 553722 6976
rect 567597 7034 567663 7037
rect 569069 7034 569135 7037
rect 567597 7032 569135 7034
rect 567597 6976 567602 7032
rect 567658 6976 569074 7032
rect 569130 6976 569135 7032
rect 567597 6974 569135 6976
rect 546897 6971 546963 6974
rect 567597 6971 567663 6974
rect 569069 6971 569135 6974
rect 520677 6898 520743 6901
rect 511158 6896 520743 6898
rect 511158 6840 520682 6896
rect 520738 6840 520743 6896
rect 511158 6838 520743 6840
rect 443508 6836 443514 6838
rect 520677 6835 520743 6838
rect 366117 6626 366183 6629
rect 356598 6624 366183 6626
rect 356598 6568 366122 6624
rect 366178 6568 366183 6624
rect 356598 6566 366183 6568
rect 235109 6563 235175 6566
rect 240997 6563 241063 6566
rect 366117 6563 366183 6566
rect 382718 6564 382724 6628
rect 382788 6626 382794 6628
rect 389853 6626 389919 6629
rect 382788 6624 389919 6626
rect 382788 6568 389858 6624
rect 389914 6568 389919 6624
rect 382788 6566 389919 6568
rect 382788 6564 382794 6566
rect 389853 6563 389919 6566
rect 225449 6490 225515 6493
rect 242193 6490 242259 6493
rect 225449 6488 242259 6490
rect 225449 6432 225454 6488
rect 225510 6432 242198 6488
rect 242254 6432 242259 6488
rect 225449 6430 242259 6432
rect 225449 6427 225515 6430
rect 242193 6427 242259 6430
rect 318921 6490 318987 6493
rect 328673 6490 328739 6493
rect 318921 6488 328739 6490
rect 318921 6432 318926 6488
rect 318982 6432 328678 6488
rect 328734 6432 328739 6488
rect 318921 6430 328739 6432
rect 318921 6427 318987 6430
rect 328673 6427 328739 6430
rect 337229 6490 337295 6493
rect 338793 6490 338859 6493
rect 337229 6488 338859 6490
rect 337229 6432 337234 6488
rect 337290 6432 338798 6488
rect 338854 6432 338859 6488
rect 337229 6430 338859 6432
rect 337229 6427 337295 6430
rect 338793 6427 338859 6430
rect 346981 6490 347047 6493
rect 356457 6490 356523 6493
rect 346981 6488 356523 6490
rect 346981 6432 346986 6488
rect 347042 6432 356462 6488
rect 356518 6432 356523 6488
rect 346981 6430 356523 6432
rect 346981 6427 347047 6430
rect 356457 6427 356523 6430
rect 225173 6354 225239 6357
rect 240813 6354 240879 6357
rect 225173 6352 240879 6354
rect 225173 6296 225178 6352
rect 225234 6296 240818 6352
rect 240874 6296 240879 6352
rect 225173 6294 240879 6296
rect 225173 6291 225239 6294
rect 240813 6291 240879 6294
rect 318829 6354 318895 6357
rect 321957 6354 322023 6357
rect 318829 6352 322023 6354
rect 318829 6296 318834 6352
rect 318890 6296 321962 6352
rect 322018 6296 322023 6352
rect 318829 6294 322023 6296
rect 318829 6291 318895 6294
rect 321957 6291 322023 6294
rect 322233 6354 322299 6357
rect 349557 6354 349623 6357
rect 322233 6352 349623 6354
rect 322233 6296 322238 6352
rect 322294 6296 349562 6352
rect 349618 6296 349623 6352
rect 322233 6294 349623 6296
rect 322233 6291 322299 6294
rect 349557 6291 349623 6294
rect 48625 6218 48691 6221
rect 239433 6218 239499 6221
rect 48625 6216 239499 6218
rect 48625 6160 48630 6216
rect 48686 6160 239438 6216
rect 239494 6160 239499 6216
rect 48625 6158 239499 6160
rect 48625 6155 48691 6158
rect 239433 6155 239499 6158
rect 320393 6218 320459 6221
rect 437509 6218 437575 6221
rect 320393 6216 437575 6218
rect 320393 6160 320398 6216
rect 320454 6160 437514 6216
rect 437570 6160 437575 6216
rect 320393 6158 437575 6160
rect 320393 6155 320459 6158
rect 437509 6155 437575 6158
rect 215789 6082 215855 6085
rect 215789 6080 217002 6082
rect 215789 6024 215794 6080
rect 215850 6024 217002 6080
rect 215789 6022 217002 6024
rect 215789 6019 215855 6022
rect 206773 5946 206839 5949
rect 215881 5946 215947 5949
rect 206773 5944 215947 5946
rect 206773 5888 206778 5944
rect 206834 5888 215886 5944
rect 215942 5888 215947 5944
rect 206773 5886 215947 5888
rect 216942 5946 217002 6022
rect 222638 6020 222644 6084
rect 222708 6082 222714 6084
rect 231521 6082 231587 6085
rect 222708 6080 231587 6082
rect 222708 6024 231526 6080
rect 231582 6024 231587 6080
rect 222708 6022 231587 6024
rect 222708 6020 222714 6022
rect 231521 6019 231587 6022
rect 331709 6082 331775 6085
rect 370441 6082 370507 6085
rect 331709 6080 370507 6082
rect 331709 6024 331714 6080
rect 331770 6024 370446 6080
rect 370502 6024 370507 6080
rect 331709 6022 370507 6024
rect 331709 6019 331775 6022
rect 370441 6019 370507 6022
rect 225449 5946 225515 5949
rect 216942 5944 225515 5946
rect 216942 5888 225454 5944
rect 225510 5888 225515 5944
rect 216942 5886 225515 5888
rect 206773 5883 206839 5886
rect 215881 5883 215947 5886
rect 225449 5883 225515 5886
rect 370349 5946 370415 5949
rect 376881 5946 376947 5949
rect 370349 5944 376947 5946
rect 370349 5888 370354 5944
rect 370410 5888 376886 5944
rect 376942 5888 376947 5944
rect 370349 5886 376947 5888
rect 370349 5883 370415 5886
rect 376881 5883 376947 5886
rect 210361 5810 210427 5813
rect 225265 5810 225331 5813
rect 210361 5808 225331 5810
rect 210361 5752 210366 5808
rect 210422 5752 225270 5808
rect 225326 5752 225331 5808
rect 210361 5750 225331 5752
rect 210361 5747 210427 5750
rect 225265 5747 225331 5750
rect 244769 5538 244835 5541
rect 257741 5538 257807 5541
rect 244769 5536 257807 5538
rect 244769 5480 244774 5536
rect 244830 5480 257746 5536
rect 257802 5480 257807 5536
rect 244769 5478 257807 5480
rect 244769 5475 244835 5478
rect 257741 5475 257807 5478
rect 231613 5402 231679 5405
rect 225590 5400 231679 5402
rect 225590 5344 231618 5400
rect 231674 5344 231679 5400
rect 225590 5342 231679 5344
rect 225265 5266 225331 5269
rect 225590 5266 225650 5342
rect 231613 5339 231679 5342
rect 244861 5402 244927 5405
rect 257281 5402 257347 5405
rect 244861 5400 257347 5402
rect 244861 5344 244866 5400
rect 244922 5344 257286 5400
rect 257342 5344 257347 5400
rect 244861 5342 257347 5344
rect 244861 5339 244927 5342
rect 257281 5339 257347 5342
rect 225265 5264 225650 5266
rect 225265 5208 225270 5264
rect 225326 5208 225650 5264
rect 225265 5206 225650 5208
rect 226921 5266 226987 5269
rect 231061 5266 231127 5269
rect 226921 5264 231127 5266
rect 226921 5208 226926 5264
rect 226982 5208 231066 5264
rect 231122 5208 231127 5264
rect 226921 5206 231127 5208
rect 225265 5203 225331 5206
rect 226921 5203 226987 5206
rect 231061 5203 231127 5206
rect 237685 5266 237751 5269
rect 244953 5266 245019 5269
rect 237685 5264 245019 5266
rect 237685 5208 237690 5264
rect 237746 5208 244958 5264
rect 245014 5208 245019 5264
rect 237685 5206 245019 5208
rect 237685 5203 237751 5206
rect 244953 5203 245019 5206
rect 312573 5266 312639 5269
rect 317449 5266 317515 5269
rect 312573 5264 317515 5266
rect 312573 5208 312578 5264
rect 312634 5208 317454 5264
rect 317510 5208 317515 5264
rect 312573 5206 317515 5208
rect 312573 5203 312639 5206
rect 317449 5203 317515 5206
rect 345325 5266 345391 5269
rect 350937 5266 351003 5269
rect 345325 5264 351003 5266
rect 345325 5208 345330 5264
rect 345386 5208 350942 5264
rect 350998 5208 351003 5264
rect 345325 5206 351003 5208
rect 345325 5203 345391 5206
rect 350937 5203 351003 5206
rect 350845 5130 350911 5133
rect 370901 5130 370967 5133
rect 350845 5128 370967 5130
rect 350845 5072 350850 5128
rect 350906 5072 370906 5128
rect 370962 5072 370967 5128
rect 350845 5070 370967 5072
rect 350845 5067 350911 5070
rect 370901 5067 370967 5070
rect 302821 4994 302887 4997
rect 312205 4994 312271 4997
rect 302821 4992 312271 4994
rect 302821 4936 302826 4992
rect 302882 4936 312210 4992
rect 312266 4936 312271 4992
rect 302821 4934 312271 4936
rect 302821 4931 302887 4934
rect 312205 4931 312271 4934
rect 350661 4994 350727 4997
rect 370993 4994 371059 4997
rect 350661 4992 371059 4994
rect 350661 4936 350666 4992
rect 350722 4936 370998 4992
rect 371054 4936 371059 4992
rect 350661 4934 371059 4936
rect 350661 4931 350727 4934
rect 370993 4931 371059 4934
rect 187729 4858 187795 4861
rect 268689 4858 268755 4861
rect 187729 4856 268755 4858
rect 187729 4800 187734 4856
rect 187790 4800 268694 4856
rect 268750 4800 268755 4856
rect 187729 4798 268755 4800
rect 187729 4795 187795 4798
rect 268689 4795 268755 4798
rect 302545 4858 302611 4861
rect 348361 4858 348427 4861
rect 302545 4856 348427 4858
rect 302545 4800 302550 4856
rect 302606 4800 348366 4856
rect 348422 4800 348427 4856
rect 302545 4798 348427 4800
rect 302545 4795 302611 4798
rect 348361 4795 348427 4798
rect 350569 4858 350635 4861
rect 355813 4858 355879 4861
rect 573117 4858 573183 4861
rect 350569 4856 351874 4858
rect 350569 4800 350574 4856
rect 350630 4800 351874 4856
rect 350569 4798 351874 4800
rect 350569 4795 350635 4798
rect 219653 4722 219719 4725
rect 225265 4722 225331 4725
rect 219653 4720 225331 4722
rect 219653 4664 219658 4720
rect 219714 4664 225270 4720
rect 225326 4664 225331 4720
rect 219653 4662 225331 4664
rect 219653 4659 219719 4662
rect 225265 4659 225331 4662
rect 321957 4722 322023 4725
rect 322141 4722 322207 4725
rect 321957 4720 322207 4722
rect 321957 4664 321962 4720
rect 322018 4664 322146 4720
rect 322202 4664 322207 4720
rect 321957 4662 322207 4664
rect 321957 4659 322023 4662
rect 322141 4659 322207 4662
rect 349189 4722 349255 4725
rect 351814 4722 351874 4798
rect 355813 4856 573183 4858
rect 355813 4800 355818 4856
rect 355874 4800 573122 4856
rect 573178 4800 573183 4856
rect 355813 4798 573183 4800
rect 355813 4795 355879 4798
rect 573117 4795 573183 4798
rect 418833 4722 418899 4725
rect 349189 4720 351690 4722
rect 349189 4664 349194 4720
rect 349250 4664 351690 4720
rect 349189 4662 351690 4664
rect 351814 4720 418899 4722
rect 351814 4664 418838 4720
rect 418894 4664 418899 4720
rect 351814 4662 418899 4664
rect 349189 4659 349255 4662
rect 264365 4586 264431 4589
rect 269793 4586 269859 4589
rect 264365 4584 269859 4586
rect 264365 4528 264370 4584
rect 264426 4528 269798 4584
rect 269854 4528 269859 4584
rect 264365 4526 269859 4528
rect 264365 4523 264431 4526
rect 269793 4523 269859 4526
rect 302545 4586 302611 4589
rect 303097 4586 303163 4589
rect 302545 4584 303163 4586
rect 302545 4528 302550 4584
rect 302606 4528 303102 4584
rect 303158 4528 303163 4584
rect 302545 4526 303163 4528
rect 302545 4523 302611 4526
rect 303097 4523 303163 4526
rect 345325 4586 345391 4589
rect 350937 4586 351003 4589
rect 345325 4584 351003 4586
rect 345325 4528 345330 4584
rect 345386 4528 350942 4584
rect 350998 4528 351003 4584
rect 345325 4526 351003 4528
rect 351630 4586 351690 4662
rect 418833 4659 418899 4662
rect 515249 4722 515315 4725
rect 519573 4722 519639 4725
rect 515249 4720 519639 4722
rect 515249 4664 515254 4720
rect 515310 4664 519578 4720
rect 519634 4664 519639 4720
rect 515249 4662 519639 4664
rect 515249 4659 515315 4662
rect 519573 4659 519639 4662
rect 355813 4586 355879 4589
rect 351630 4584 355879 4586
rect 351630 4528 355818 4584
rect 355874 4528 355879 4584
rect 351630 4526 355879 4528
rect 345325 4523 345391 4526
rect 350937 4523 351003 4526
rect 355813 4523 355879 4526
rect 264181 4450 264247 4453
rect 272921 4450 272987 4453
rect 264181 4448 272987 4450
rect 264181 4392 264186 4448
rect 264242 4392 272926 4448
rect 272982 4392 272987 4448
rect 264181 4390 272987 4392
rect 264181 4387 264247 4390
rect 272921 4387 272987 4390
rect 302453 4450 302519 4453
rect 303005 4450 303071 4453
rect 302453 4448 303071 4450
rect 302453 4392 302458 4448
rect 302514 4392 303010 4448
rect 303066 4392 303071 4448
rect 302453 4390 303071 4392
rect 302453 4387 302519 4390
rect 303005 4387 303071 4390
rect 342657 4450 342723 4453
rect 350845 4450 350911 4453
rect 342657 4448 350911 4450
rect 342657 4392 342662 4448
rect 342718 4392 350850 4448
rect 350906 4392 350911 4448
rect 342657 4390 350911 4392
rect 342657 4387 342723 4390
rect 350845 4387 350911 4390
rect 216341 4314 216407 4317
rect 218641 4314 218707 4317
rect 216341 4312 218707 4314
rect 216341 4256 216346 4312
rect 216402 4256 218646 4312
rect 218702 4256 218707 4312
rect 216341 4254 218707 4256
rect 216341 4251 216407 4254
rect 218641 4251 218707 4254
rect 225449 4314 225515 4317
rect 235661 4314 235727 4317
rect 225449 4312 235727 4314
rect 225449 4256 225454 4312
rect 225510 4256 235666 4312
rect 235722 4256 235727 4312
rect 225449 4254 235727 4256
rect 225449 4251 225515 4254
rect 235661 4251 235727 4254
rect 215789 4178 215855 4181
rect 219745 4178 219811 4181
rect 215789 4176 219811 4178
rect 215789 4120 215794 4176
rect 215850 4120 219750 4176
rect 219806 4120 219811 4176
rect 215789 4118 219811 4120
rect 215789 4115 215855 4118
rect 219745 4115 219811 4118
rect 230141 4178 230207 4181
rect 234925 4178 234991 4181
rect 230141 4176 234991 4178
rect 230141 4120 230146 4176
rect 230202 4120 234930 4176
rect 234986 4120 234991 4176
rect 230141 4118 234991 4120
rect 230141 4115 230207 4118
rect 234925 4115 234991 4118
rect 235109 4178 235175 4181
rect 238053 4178 238119 4181
rect 235109 4176 238119 4178
rect 235109 4120 235114 4176
rect 235170 4120 238058 4176
rect 238114 4120 238119 4176
rect 235109 4118 238119 4120
rect 235109 4115 235175 4118
rect 238053 4115 238119 4118
rect 31973 4042 32039 4045
rect 236949 4042 237015 4045
rect 31973 4040 237015 4042
rect 31973 3984 31978 4040
rect 32034 3984 236954 4040
rect 237010 3984 237015 4040
rect 31973 3982 237015 3984
rect 31973 3979 32039 3982
rect 236949 3979 237015 3982
rect 326005 4042 326071 4045
rect 464925 4042 464991 4045
rect 326005 4040 464991 4042
rect 326005 3984 326010 4040
rect 326066 3984 464930 4040
rect 464986 3984 464991 4040
rect 326005 3982 464991 3984
rect 326005 3979 326071 3982
rect 464925 3979 464991 3982
rect 25993 3906 26059 3909
rect 235201 3906 235267 3909
rect 25993 3904 235267 3906
rect 25993 3848 25998 3904
rect 26054 3848 235206 3904
rect 235262 3848 235267 3904
rect 25993 3846 235267 3848
rect 25993 3843 26059 3846
rect 235201 3843 235267 3846
rect 327385 3906 327451 3909
rect 468421 3906 468487 3909
rect 327385 3904 468487 3906
rect 327385 3848 327390 3904
rect 327446 3848 468426 3904
rect 468482 3848 468487 3904
rect 327385 3846 468487 3848
rect 327385 3843 327451 3846
rect 468421 3843 468487 3846
rect 24797 3770 24863 3773
rect 235569 3770 235635 3773
rect 24797 3768 235635 3770
rect 24797 3712 24802 3768
rect 24858 3712 235574 3768
rect 235630 3712 235635 3768
rect 24797 3710 235635 3712
rect 24797 3707 24863 3710
rect 235569 3707 235635 3710
rect 327477 3770 327543 3773
rect 472009 3770 472075 3773
rect 327477 3768 472075 3770
rect 327477 3712 327482 3768
rect 327538 3712 472014 3768
rect 472070 3712 472075 3768
rect 327477 3710 472075 3712
rect 327477 3707 327543 3710
rect 472009 3707 472075 3710
rect 16517 3634 16583 3637
rect 228117 3634 228183 3637
rect 230417 3634 230483 3637
rect 16517 3632 228042 3634
rect 16517 3576 16522 3632
rect 16578 3576 228042 3632
rect 16517 3574 228042 3576
rect 16517 3571 16583 3574
rect 15321 3498 15387 3501
rect 58193 3498 58259 3501
rect 15321 3496 58259 3498
rect 15321 3440 15326 3496
rect 15382 3440 58198 3496
rect 58254 3440 58259 3496
rect 15321 3438 58259 3440
rect 15321 3435 15387 3438
rect 58193 3435 58259 3438
rect 58377 3498 58443 3501
rect 227982 3498 228042 3574
rect 228117 3632 230483 3634
rect 228117 3576 228122 3632
rect 228178 3576 230422 3632
rect 230478 3576 230483 3632
rect 228117 3574 230483 3576
rect 228117 3571 228183 3574
rect 230417 3571 230483 3574
rect 235201 3634 235267 3637
rect 236765 3634 236831 3637
rect 235201 3632 236831 3634
rect 235201 3576 235206 3632
rect 235262 3576 236770 3632
rect 236826 3576 236831 3632
rect 235201 3574 236831 3576
rect 235201 3571 235267 3574
rect 236765 3571 236831 3574
rect 328765 3634 328831 3637
rect 347942 3634 347948 3636
rect 328765 3632 347948 3634
rect 328765 3576 328770 3632
rect 328826 3576 347948 3632
rect 328765 3574 347948 3576
rect 328765 3571 328831 3574
rect 347942 3572 347948 3574
rect 348012 3572 348018 3636
rect 348494 3572 348500 3636
rect 348564 3634 348570 3636
rect 475597 3634 475663 3637
rect 348564 3632 475663 3634
rect 348564 3576 475602 3632
rect 475658 3576 475663 3632
rect 348564 3574 475663 3576
rect 348564 3572 348570 3574
rect 475597 3571 475663 3574
rect 232901 3498 232967 3501
rect 58377 3496 227858 3498
rect 58377 3440 58382 3496
rect 58438 3440 227858 3496
rect 58377 3438 227858 3440
rect 227982 3496 232967 3498
rect 227982 3440 232906 3496
rect 232962 3440 232967 3496
rect 227982 3438 232967 3440
rect 58377 3435 58443 3438
rect 6949 3362 7015 3365
rect 58193 3362 58259 3365
rect 6949 3360 58259 3362
rect 6949 3304 6954 3360
rect 7010 3304 58198 3360
rect 58254 3304 58259 3360
rect 6949 3302 58259 3304
rect 6949 3299 7015 3302
rect 58193 3299 58259 3302
rect 58377 3362 58443 3365
rect 145358 3362 145364 3364
rect 58377 3360 145364 3362
rect 58377 3304 58382 3360
rect 58438 3304 145364 3360
rect 58377 3302 145364 3304
rect 58377 3299 58443 3302
rect 145358 3300 145364 3302
rect 145428 3300 145434 3364
rect 148169 3362 148235 3365
rect 208153 3362 208219 3365
rect 148169 3360 208219 3362
rect 148169 3304 148174 3360
rect 148230 3304 208158 3360
rect 208214 3304 208219 3360
rect 148169 3302 208219 3304
rect 227798 3362 227858 3438
rect 232901 3435 232967 3438
rect 235109 3498 235175 3501
rect 237133 3498 237199 3501
rect 235109 3496 237199 3498
rect 235109 3440 235114 3496
rect 235170 3440 237138 3496
rect 237194 3440 237199 3496
rect 235109 3438 237199 3440
rect 235109 3435 235175 3438
rect 237133 3435 237199 3438
rect 328857 3498 328923 3501
rect 336677 3498 336743 3501
rect 341461 3498 341527 3501
rect 348180 3498 348424 3532
rect 364921 3498 364987 3501
rect 370257 3498 370323 3501
rect 328857 3496 333658 3498
rect 328857 3440 328862 3496
rect 328918 3440 333658 3496
rect 328857 3438 333658 3440
rect 328857 3435 328923 3438
rect 232717 3362 232783 3365
rect 227798 3360 232783 3362
rect 227798 3304 232722 3360
rect 232778 3304 232783 3360
rect 227798 3302 232783 3304
rect 148169 3299 148235 3302
rect 208153 3299 208219 3302
rect 232717 3299 232783 3302
rect 234833 3362 234899 3365
rect 235385 3362 235451 3365
rect 234833 3360 235451 3362
rect 234833 3304 234838 3360
rect 234894 3304 235390 3360
rect 235446 3304 235451 3360
rect 234833 3302 235451 3304
rect 234833 3299 234899 3302
rect 235385 3299 235451 3302
rect 99685 3226 99751 3229
rect 103825 3226 103891 3229
rect 99685 3224 103891 3226
rect 99685 3168 99690 3224
rect 99746 3168 103830 3224
rect 103886 3168 103891 3224
rect 99685 3166 103891 3168
rect 99685 3163 99751 3166
rect 103825 3163 103891 3166
rect 113853 3226 113919 3229
rect 126089 3226 126155 3229
rect 113853 3224 126155 3226
rect 113853 3168 113858 3224
rect 113914 3168 126094 3224
rect 126150 3168 126155 3224
rect 113853 3166 126155 3168
rect 113853 3163 113919 3166
rect 126089 3163 126155 3166
rect 157645 3226 157711 3229
rect 158105 3226 158171 3229
rect 157645 3224 158171 3226
rect 157645 3168 157650 3224
rect 157706 3168 158110 3224
rect 158166 3168 158171 3224
rect 157645 3166 158171 3168
rect 157645 3163 157711 3166
rect 158105 3163 158171 3166
rect 186533 3226 186599 3229
rect 187177 3226 187243 3229
rect 186533 3224 187243 3226
rect 186533 3168 186538 3224
rect 186594 3168 187182 3224
rect 187238 3168 187243 3224
rect 186533 3166 187243 3168
rect 186533 3163 186599 3166
rect 187177 3163 187243 3166
rect 196193 3226 196259 3229
rect 196745 3226 196811 3229
rect 196193 3224 196811 3226
rect 196193 3168 196198 3224
rect 196254 3168 196750 3224
rect 196806 3168 196811 3224
rect 196193 3166 196811 3168
rect 196193 3163 196259 3166
rect 196745 3163 196811 3166
rect 205853 3226 205919 3229
rect 206221 3226 206287 3229
rect 205853 3224 206287 3226
rect 205853 3168 205858 3224
rect 205914 3168 206226 3224
rect 206282 3168 206287 3224
rect 205853 3166 206287 3168
rect 205853 3163 205919 3166
rect 206221 3163 206287 3166
rect 224529 3226 224595 3229
rect 225633 3226 225699 3229
rect 224529 3224 225699 3226
rect 224529 3168 224534 3224
rect 224590 3168 225638 3224
rect 225694 3168 225699 3224
rect 224529 3166 225699 3168
rect 224529 3163 224595 3166
rect 225633 3163 225699 3166
rect 234741 3226 234807 3229
rect 235201 3226 235267 3229
rect 234741 3224 235267 3226
rect 234741 3168 234746 3224
rect 234802 3168 235206 3224
rect 235262 3168 235267 3224
rect 234741 3166 235267 3168
rect 333598 3226 333658 3438
rect 336677 3496 341527 3498
rect 336677 3440 336682 3496
rect 336738 3440 341466 3496
rect 341522 3440 341527 3496
rect 336677 3438 341527 3440
rect 336677 3435 336743 3438
rect 341461 3435 341527 3438
rect 343350 3472 362730 3498
rect 343350 3438 348240 3472
rect 348364 3438 362730 3472
rect 338517 3362 338583 3365
rect 343350 3362 343410 3438
rect 338517 3360 343410 3362
rect 338517 3304 338522 3360
rect 338578 3304 343410 3360
rect 338517 3302 343410 3304
rect 346245 3362 346311 3365
rect 362670 3362 362730 3438
rect 364921 3496 370323 3498
rect 364921 3440 364926 3496
rect 364982 3440 370262 3496
rect 370318 3440 370323 3496
rect 364921 3438 370323 3440
rect 364921 3435 364987 3438
rect 370257 3435 370323 3438
rect 375133 3498 375199 3501
rect 433553 3498 433619 3501
rect 375133 3496 433619 3498
rect 375133 3440 375138 3496
rect 375194 3440 433558 3496
rect 433614 3440 433619 3496
rect 375133 3438 433619 3440
rect 375133 3435 375199 3438
rect 433553 3435 433619 3438
rect 433737 3498 433803 3501
rect 479185 3498 479251 3501
rect 433737 3496 479251 3498
rect 433737 3440 433742 3496
rect 433798 3440 479190 3496
rect 479246 3440 479251 3496
rect 433737 3438 479251 3440
rect 433737 3435 433803 3438
rect 479185 3435 479251 3438
rect 365289 3362 365355 3365
rect 375777 3362 375843 3365
rect 346245 3360 355922 3362
rect 346245 3304 346250 3360
rect 346306 3304 355922 3360
rect 346245 3302 355922 3304
rect 362670 3360 365355 3362
rect 362670 3304 365294 3360
rect 365350 3304 365355 3360
rect 362670 3302 365355 3304
rect 338517 3299 338583 3302
rect 346245 3299 346311 3302
rect 338333 3226 338399 3229
rect 333598 3224 338399 3226
rect 333598 3168 338338 3224
rect 338394 3168 338399 3224
rect 333598 3166 338399 3168
rect 234741 3163 234807 3166
rect 235201 3163 235267 3166
rect 338333 3163 338399 3166
rect 346337 3226 346403 3229
rect 351121 3226 351187 3229
rect 346337 3224 351187 3226
rect 346337 3168 346342 3224
rect 346398 3168 351126 3224
rect 351182 3168 351187 3224
rect 346337 3166 351187 3168
rect 346337 3163 346403 3166
rect 351121 3163 351187 3166
rect 145358 3028 145364 3092
rect 145428 3090 145434 3092
rect 148077 3090 148143 3093
rect 145428 3088 148143 3090
rect 145428 3032 148082 3088
rect 148138 3032 148143 3088
rect 145428 3030 148143 3032
rect 145428 3028 145434 3030
rect 148077 3027 148143 3030
rect 210269 3090 210335 3093
rect 225173 3090 225239 3093
rect 210269 3088 225239 3090
rect 210269 3032 210274 3088
rect 210330 3032 225178 3088
rect 225234 3032 225239 3088
rect 210269 3030 225239 3032
rect 355862 3090 355922 3302
rect 365289 3299 365355 3302
rect 365430 3360 375843 3362
rect 365430 3304 375782 3360
rect 375838 3304 375843 3360
rect 365430 3302 375843 3304
rect 360505 3226 360571 3229
rect 360781 3226 360847 3229
rect 360505 3224 360847 3226
rect 360505 3168 360510 3224
rect 360566 3168 360786 3224
rect 360842 3168 360847 3224
rect 360505 3166 360847 3168
rect 360505 3163 360571 3166
rect 360781 3163 360847 3166
rect 365430 3090 365490 3302
rect 375777 3299 375843 3302
rect 375961 3362 376027 3365
rect 392429 3362 392495 3365
rect 375961 3360 392495 3362
rect 375961 3304 375966 3360
rect 376022 3304 392434 3360
rect 392490 3304 392495 3360
rect 375961 3302 392495 3304
rect 375961 3299 376027 3302
rect 392429 3299 392495 3302
rect 411657 3362 411723 3365
rect 414509 3362 414575 3365
rect 433829 3362 433895 3365
rect 411657 3360 414575 3362
rect 411657 3304 411662 3360
rect 411718 3304 414514 3360
rect 414570 3304 414575 3360
rect 411657 3302 414575 3304
rect 411657 3299 411723 3302
rect 414509 3299 414575 3302
rect 433694 3360 433895 3362
rect 433694 3304 433834 3360
rect 433890 3304 433895 3360
rect 433694 3302 433895 3304
rect 370165 3226 370231 3229
rect 370625 3226 370691 3229
rect 370165 3224 370691 3226
rect 370165 3168 370170 3224
rect 370226 3168 370630 3224
rect 370686 3168 370691 3224
rect 370165 3166 370691 3168
rect 370165 3163 370231 3166
rect 370625 3163 370691 3166
rect 401997 3226 402063 3229
rect 406873 3226 406939 3229
rect 401997 3224 406939 3226
rect 401997 3168 402002 3224
rect 402058 3168 406878 3224
rect 406934 3168 406939 3224
rect 401997 3166 406939 3168
rect 401997 3163 402063 3166
rect 406873 3163 406939 3166
rect 424077 3226 424143 3229
rect 424077 3224 428050 3226
rect 424077 3168 424082 3224
rect 424138 3168 428050 3224
rect 424077 3166 428050 3168
rect 424077 3163 424143 3166
rect 370533 3090 370599 3093
rect 355862 3030 365490 3090
rect 365614 3088 370599 3090
rect 365614 3032 370538 3088
rect 370594 3032 370599 3088
rect 365614 3030 370599 3032
rect 427990 3090 428050 3166
rect 433694 3090 433754 3302
rect 433829 3299 433895 3302
rect 451677 3226 451743 3229
rect 462717 3226 462783 3229
rect 466581 3226 466647 3229
rect 451677 3224 453258 3226
rect 451677 3168 451682 3224
rect 451738 3168 453258 3224
rect 451677 3166 453258 3168
rect 451677 3163 451743 3166
rect 427990 3030 433754 3090
rect 453198 3090 453258 3166
rect 462717 3224 466647 3226
rect 462717 3168 462722 3224
rect 462778 3168 466586 3224
rect 466642 3168 466647 3224
rect 462717 3166 466647 3168
rect 462717 3163 462783 3166
rect 466581 3163 466647 3166
rect 480657 3226 480723 3229
rect 482773 3226 482839 3229
rect 480657 3224 482839 3226
rect 480657 3168 480662 3224
rect 480718 3168 482778 3224
rect 482834 3168 482839 3224
rect 480657 3166 482839 3168
rect 480657 3163 480723 3166
rect 482773 3163 482839 3166
rect 462717 3090 462783 3093
rect 453198 3088 462783 3090
rect 453198 3032 462722 3088
rect 462778 3032 462783 3088
rect 453198 3030 462783 3032
rect 210269 3027 210335 3030
rect 225173 3027 225239 3030
rect 195917 2954 195983 2957
rect 207693 2954 207759 2957
rect 195917 2952 207759 2954
rect 195917 2896 195922 2952
rect 195978 2896 207698 2952
rect 207754 2896 207759 2952
rect 195917 2894 207759 2896
rect 195917 2891 195983 2894
rect 207693 2891 207759 2894
rect 329777 2954 329843 2957
rect 346245 2954 346311 2957
rect 329777 2952 346311 2954
rect 329777 2896 329782 2952
rect 329838 2896 346250 2952
rect 346306 2896 346311 2952
rect 329777 2894 346311 2896
rect 329777 2891 329843 2894
rect 346245 2891 346311 2894
rect 355261 2954 355327 2957
rect 360597 2954 360663 2957
rect 355261 2952 360663 2954
rect 355261 2896 355266 2952
rect 355322 2896 360602 2952
rect 360658 2896 360663 2952
rect 355261 2894 360663 2896
rect 355261 2891 355327 2894
rect 360597 2891 360663 2894
rect 364737 2954 364803 2957
rect 365614 2954 365674 3030
rect 370533 3027 370599 3030
rect 462717 3027 462783 3030
rect 364737 2952 365674 2954
rect 364737 2896 364742 2952
rect 364798 2896 365674 2952
rect 364737 2894 365674 2896
rect 365749 2954 365815 2957
rect 375133 2954 375199 2957
rect 365749 2952 375199 2954
rect 365749 2896 365754 2952
rect 365810 2896 375138 2952
rect 375194 2896 375199 2952
rect 365749 2894 375199 2896
rect 364737 2891 364803 2894
rect 365749 2891 365815 2894
rect 375133 2891 375199 2894
rect 392429 2954 392495 2957
rect 401997 2954 402063 2957
rect 392429 2952 402063 2954
rect 392429 2896 392434 2952
rect 392490 2896 402002 2952
rect 402058 2896 402063 2952
rect 392429 2894 402063 2896
rect 392429 2891 392495 2894
rect 401997 2891 402063 2894
rect 222638 2818 222644 2820
rect 212894 2758 222644 2818
rect 208153 2546 208219 2549
rect 212894 2546 212954 2758
rect 222638 2756 222644 2758
rect 222708 2756 222714 2820
rect 364645 2818 364711 2821
rect 365105 2818 365171 2821
rect 364645 2816 365171 2818
rect 364645 2760 364650 2816
rect 364706 2760 365110 2816
rect 365166 2760 365171 2816
rect 364645 2758 365171 2760
rect 364645 2755 364711 2758
rect 365105 2755 365171 2758
rect 208153 2544 212954 2546
rect 208153 2488 208158 2544
rect 208214 2488 212954 2544
rect 208153 2486 212954 2488
rect 208153 2483 208219 2486
<< via3 >>
rect 443628 618156 443692 618220
rect 443628 608696 443692 608700
rect 443628 608640 443678 608696
rect 443678 608640 443692 608696
rect 443628 608636 443692 608640
rect 379044 529816 379108 529820
rect 379044 529760 379058 529816
rect 379058 529760 379108 529816
rect 379044 529756 379108 529760
rect 508764 529816 508828 529820
rect 508764 529760 508778 529816
rect 508778 529760 508828 529816
rect 508764 529756 508828 529760
rect 379044 520236 379108 520300
rect 508764 520236 508828 520300
rect 232212 459640 232276 459644
rect 232212 459584 232226 459640
rect 232226 459584 232276 459640
rect 232212 459580 232276 459584
rect 233500 459580 233564 459644
rect 236260 459640 236324 459644
rect 236260 459584 236274 459640
rect 236274 459584 236324 459640
rect 236260 459580 236324 459584
rect 237732 459580 237796 459644
rect 239020 459580 239084 459644
rect 240492 459580 240556 459644
rect 241780 459580 241844 459644
rect 243252 459580 243316 459644
rect 244540 459640 244604 459644
rect 244540 459584 244590 459640
rect 244590 459584 244604 459640
rect 244540 459580 244604 459584
rect 246012 459580 246076 459644
rect 247300 459580 247364 459644
rect 248772 459640 248836 459644
rect 248772 459584 248822 459640
rect 248822 459584 248836 459640
rect 248772 459580 248836 459584
rect 251532 459580 251596 459644
rect 252820 459580 252884 459644
rect 342796 459580 342860 459644
rect 344084 459580 344148 459644
rect 345556 459580 345620 459644
rect 346844 459580 346908 459644
rect 348316 459580 348380 459644
rect 280604 320588 280668 320652
rect 251532 320452 251596 320516
rect 299924 320452 299988 320516
rect 309492 320316 309556 320380
rect 280788 320180 280852 320244
rect 338564 320180 338628 320244
rect 512444 320452 512508 320516
rect 512444 320180 512508 320244
rect 551084 320452 551148 320516
rect 551084 320180 551148 320244
rect 299924 320044 299988 320108
rect 309492 320044 309556 320108
rect 338564 319908 338628 319972
rect 385484 319152 385548 319156
rect 385484 319096 385534 319152
rect 385534 319096 385548 319152
rect 385484 319092 385548 319096
rect 385484 318880 385548 318884
rect 385484 318824 385534 318880
rect 385534 318824 385548 318880
rect 385484 318820 385548 318824
rect 252820 304948 252884 305012
rect 341140 290184 341204 290188
rect 341140 290128 341154 290184
rect 341154 290128 341204 290184
rect 341140 290124 341204 290128
rect 341140 289912 341204 289916
rect 341140 289856 341154 289912
rect 341154 289856 341204 289912
rect 341140 289852 341204 289856
rect 319980 282916 320044 282980
rect 319980 278896 320044 278900
rect 319980 278840 320030 278896
rect 320030 278840 320044 278896
rect 319980 278836 320044 278840
rect 248772 258028 248836 258092
rect 319980 251152 320044 251156
rect 319980 251096 320030 251152
rect 320030 251096 320044 251152
rect 319980 251092 320044 251096
rect 235524 244352 235588 244356
rect 235524 244296 235574 244352
rect 235574 244296 235588 244352
rect 235524 244292 235588 244296
rect 319060 242388 319124 242452
rect 377204 242116 377268 242180
rect 247300 241708 247364 241772
rect 319060 241980 319124 242044
rect 299924 241844 299988 241908
rect 300108 241708 300172 241772
rect 235524 241632 235588 241636
rect 235524 241576 235538 241632
rect 235538 241576 235588 241632
rect 235524 241572 235588 241576
rect 319980 241632 320044 241636
rect 377204 241708 377268 241772
rect 319980 241576 320030 241632
rect 320030 241576 320044 241632
rect 319980 241572 320044 241576
rect 551084 241844 551148 241908
rect 551084 241572 551148 241636
rect 319060 227156 319124 227220
rect 319060 226748 319124 226812
rect 244540 226612 244604 226676
rect 261284 226476 261348 226540
rect 288884 226612 288948 226676
rect 288884 226340 288948 226404
rect 551084 226612 551148 226676
rect 551084 226340 551148 226404
rect 261284 226204 261348 226268
rect 276556 221504 276620 221508
rect 276556 221448 276570 221504
rect 276570 221448 276620 221504
rect 276556 221444 276620 221448
rect 319980 216064 320044 216068
rect 319980 216008 320030 216064
rect 320030 216008 320044 216064
rect 319980 216004 320044 216008
rect 246012 211108 246076 211172
rect 276556 208448 276620 208452
rect 276556 208392 276570 208448
rect 276570 208392 276620 208448
rect 276556 208388 276620 208392
rect 319980 206272 320044 206276
rect 319980 206216 320030 206272
rect 320030 206216 320044 206272
rect 319980 206212 320044 206216
rect 553844 183560 553908 183564
rect 553844 183504 553894 183560
rect 553894 183504 553908 183560
rect 553844 183500 553908 183504
rect 242516 182004 242580 182068
rect 288884 179964 288948 180028
rect 241780 179556 241844 179620
rect 269564 179692 269628 179756
rect 288884 179692 288948 179756
rect 327524 179692 327588 179756
rect 299924 179556 299988 179620
rect 269564 179420 269628 179484
rect 308204 179420 308268 179484
rect 327524 179420 327588 179484
rect 356596 179692 356660 179756
rect 396524 179692 396588 179756
rect 396524 179420 396588 179484
rect 551084 179692 551148 179756
rect 551084 179420 551148 179484
rect 356596 179284 356660 179348
rect 299924 179148 299988 179212
rect 308204 179148 308268 179212
rect 285388 177244 285452 177308
rect 553844 174040 553908 174044
rect 553844 173984 553894 174040
rect 553894 173984 553908 174040
rect 553844 173980 553908 173984
rect 91452 173904 91516 173908
rect 91452 173848 91502 173904
rect 91502 173848 91516 173904
rect 91452 173844 91516 173848
rect 225404 173904 225468 173908
rect 225404 173848 225418 173904
rect 225418 173848 225468 173904
rect 225404 173844 225468 173848
rect 357884 173904 357948 173908
rect 357884 173848 357934 173904
rect 357934 173848 357948 173904
rect 357884 173844 357948 173848
rect 560836 164596 560900 164660
rect 357884 164384 357948 164388
rect 357884 164328 357934 164384
rect 357934 164328 357948 164384
rect 357884 164324 357948 164328
rect 91452 164248 91516 164252
rect 91452 164192 91502 164248
rect 91502 164192 91516 164248
rect 91452 164188 91516 164192
rect 225404 164248 225468 164252
rect 225404 164192 225418 164248
rect 225418 164192 225468 164248
rect 225404 164188 225468 164192
rect 243252 164188 243316 164252
rect 560836 164188 560900 164252
rect 285388 164112 285452 164116
rect 285388 164056 285402 164112
rect 285402 164056 285452 164112
rect 285388 164052 285452 164056
rect 242516 163024 242580 163028
rect 242516 162968 242566 163024
rect 242566 162968 242580 163024
rect 242516 162964 242580 162968
rect 242516 157856 242580 157860
rect 242516 157800 242530 157856
rect 242530 157800 242580 157856
rect 242516 157796 242580 157800
rect 309308 151676 309372 151740
rect 242516 144936 242580 144940
rect 242516 144880 242530 144936
rect 242530 144880 242580 144936
rect 242516 144876 242580 144880
rect 309308 142156 309372 142220
rect 239020 133996 239084 134060
rect 357884 133044 357948 133108
rect 366164 133044 366228 133108
rect 308204 132772 308268 132836
rect 317772 132772 317836 132836
rect 327524 132772 327588 132836
rect 308204 132500 308268 132564
rect 317772 132500 317836 132564
rect 327524 132500 327588 132564
rect 357884 132772 357948 132836
rect 366164 132636 366228 132700
rect 551084 132772 551148 132836
rect 551084 132500 551148 132564
rect 342796 126924 342860 126988
rect 240492 117268 240556 117332
rect 377204 101356 377268 101420
rect 237732 101084 237796 101148
rect 316484 100812 316548 100876
rect 377204 101084 377268 101148
rect 396524 101084 396588 101148
rect 396524 100812 396588 100876
rect 551084 101084 551148 101148
rect 551084 100812 551148 100876
rect 316484 100540 316548 100604
rect 344084 92380 344148 92444
rect 345556 75788 345620 75852
rect 236260 70348 236324 70412
rect 346844 42740 346908 42804
rect 327524 39068 327588 39132
rect 232212 38932 232276 38996
rect 317772 38932 317836 38996
rect 346660 39204 346724 39268
rect 346844 38932 346908 38996
rect 356596 38932 356660 38996
rect 317772 38660 317836 38724
rect 327524 38660 327588 38724
rect 346660 38660 346724 38724
rect 346844 38660 346908 38724
rect 551084 38932 551148 38996
rect 551084 38660 551148 38724
rect 356596 38524 356660 38588
rect 233500 23428 233564 23492
rect 177196 10100 177260 10164
rect 177012 9964 177076 10028
rect 348316 9556 348380 9620
rect 250244 7516 250308 7580
rect 501404 7516 501468 7580
rect 393764 7380 393828 7444
rect 250244 7244 250308 7308
rect 308204 7244 308268 7308
rect 292932 7108 292996 7172
rect 293116 7108 293180 7172
rect 299924 7108 299988 7172
rect 375732 7108 375796 7172
rect 537284 7380 537348 7444
rect 443444 7108 443508 7172
rect 346660 6972 346724 7036
rect 346844 6972 346908 7036
rect 300108 6836 300172 6900
rect 308204 6836 308268 6900
rect 393764 6972 393828 7036
rect 346660 6700 346724 6764
rect 346844 6700 346908 6764
rect 375916 6836 375980 6900
rect 382724 6836 382788 6900
rect 443444 6836 443508 6900
rect 501404 7244 501468 7308
rect 537284 7108 537348 7172
rect 382724 6564 382788 6628
rect 222644 6020 222708 6084
rect 347948 3572 348012 3636
rect 348500 3572 348564 3636
rect 145364 3300 145428 3364
rect 145364 3028 145428 3092
rect 222644 2756 222708 2820
<< metal4 >>
rect 0 703278 400 703360
rect 0 703042 82 703278
rect 318 703042 400 703278
rect 0 694934 400 703042
rect 584516 703278 584916 703360
rect 584516 703042 584598 703278
rect 584834 703042 584916 703278
rect 0 694698 82 694934
rect 318 694698 400 694934
rect 0 664298 400 694698
rect 0 664062 82 664298
rect 318 664062 400 664298
rect 0 633662 400 664062
rect 0 633426 82 633662
rect 318 633426 400 633662
rect 0 603026 400 633426
rect 0 602790 82 603026
rect 318 602790 400 603026
rect 0 572390 400 602790
rect 0 572154 82 572390
rect 318 572154 400 572390
rect 0 541754 400 572154
rect 0 541518 82 541754
rect 318 541518 400 541754
rect 0 511118 400 541518
rect 0 510882 82 511118
rect 318 510882 400 511118
rect 0 480482 400 510882
rect 0 480246 82 480482
rect 318 480246 400 480482
rect 0 449846 400 480246
rect 0 449610 82 449846
rect 318 449610 400 449846
rect 0 419210 400 449610
rect 0 418974 82 419210
rect 318 418974 400 419210
rect 0 388574 400 418974
rect 0 388338 82 388574
rect 318 388338 400 388574
rect 0 357938 400 388338
rect 0 357702 82 357938
rect 318 357702 400 357938
rect 0 327302 400 357702
rect 0 327066 82 327302
rect 318 327066 400 327302
rect 0 296666 400 327066
rect 0 296430 82 296666
rect 318 296430 400 296666
rect 0 266030 400 296430
rect 0 265794 82 266030
rect 318 265794 400 266030
rect 0 235394 400 265794
rect 0 235158 82 235394
rect 318 235158 400 235394
rect 0 204758 400 235158
rect 0 204522 82 204758
rect 318 204522 400 204758
rect 0 174122 400 204522
rect 0 173886 82 174122
rect 318 173886 400 174122
rect 0 143486 400 173886
rect 0 143250 82 143486
rect 318 143250 400 143486
rect 0 112850 400 143250
rect 0 112614 82 112850
rect 318 112614 400 112850
rect 0 82214 400 112614
rect 0 81978 82 82214
rect 318 81978 400 82214
rect 0 51578 400 81978
rect 0 51342 82 51578
rect 318 51342 400 51578
rect 0 20942 400 51342
rect 0 20706 82 20942
rect 318 20706 400 20942
rect 0 894 400 20706
rect 800 702478 1200 702560
rect 800 702242 882 702478
rect 1118 702242 1200 702478
rect 800 679616 1200 702242
rect 800 679380 882 679616
rect 1118 679380 1200 679616
rect 800 648980 1200 679380
rect 800 648744 882 648980
rect 1118 648744 1200 648980
rect 800 618344 1200 648744
rect 800 618108 882 618344
rect 1118 618108 1200 618344
rect 583716 702478 584116 702560
rect 583716 702242 583798 702478
rect 584034 702242 584116 702478
rect 583716 679616 584116 702242
rect 583716 679380 583798 679616
rect 584034 679380 584116 679616
rect 583716 648980 584116 679380
rect 583716 648744 583798 648980
rect 584034 648744 584116 648980
rect 583716 618344 584116 648744
rect 443627 618220 443693 618221
rect 443627 618156 443628 618220
rect 443692 618156 443693 618220
rect 443627 618155 443693 618156
rect 800 587708 1200 618108
rect 443630 608701 443690 618155
rect 583716 618108 583798 618344
rect 584034 618108 584116 618344
rect 443627 608700 443693 608701
rect 443627 608636 443628 608700
rect 443692 608636 443693 608700
rect 443627 608635 443693 608636
rect 800 587472 882 587708
rect 1118 587472 1200 587708
rect 800 557072 1200 587472
rect 800 556836 882 557072
rect 1118 556836 1200 557072
rect 800 526436 1200 556836
rect 583716 587708 584116 618108
rect 583716 587472 583798 587708
rect 584034 587472 584116 587708
rect 583716 557072 584116 587472
rect 583716 556836 583798 557072
rect 584034 556836 584116 557072
rect 379043 529820 379109 529821
rect 379043 529756 379044 529820
rect 379108 529756 379109 529820
rect 379043 529755 379109 529756
rect 508763 529820 508829 529821
rect 508763 529756 508764 529820
rect 508828 529756 508829 529820
rect 508763 529755 508829 529756
rect 800 526200 882 526436
rect 1118 526200 1200 526436
rect 800 495800 1200 526200
rect 379046 520301 379106 529755
rect 508766 520301 508826 529755
rect 583716 526436 584116 556836
rect 583716 526200 583798 526436
rect 584034 526200 584116 526436
rect 379043 520300 379109 520301
rect 379043 520236 379044 520300
rect 379108 520236 379109 520300
rect 379043 520235 379109 520236
rect 508763 520300 508829 520301
rect 508763 520236 508764 520300
rect 508828 520236 508829 520300
rect 508763 520235 508829 520236
rect 800 495564 882 495800
rect 1118 495564 1200 495800
rect 800 465164 1200 495564
rect 800 464928 882 465164
rect 1118 464928 1200 465164
rect 800 434528 1200 464928
rect 583716 495800 584116 526200
rect 583716 495564 583798 495800
rect 584034 495564 584116 495800
rect 583716 465164 584116 495564
rect 583716 464928 583798 465164
rect 584034 464928 584116 465164
rect 232211 459644 232277 459645
rect 232211 459580 232212 459644
rect 232276 459580 232277 459644
rect 232211 459579 232277 459580
rect 233499 459644 233565 459645
rect 233499 459580 233500 459644
rect 233564 459580 233565 459644
rect 233499 459579 233565 459580
rect 236259 459644 236325 459645
rect 236259 459580 236260 459644
rect 236324 459580 236325 459644
rect 236259 459579 236325 459580
rect 237731 459644 237797 459645
rect 237731 459580 237732 459644
rect 237796 459580 237797 459644
rect 237731 459579 237797 459580
rect 239019 459644 239085 459645
rect 239019 459580 239020 459644
rect 239084 459580 239085 459644
rect 239019 459579 239085 459580
rect 240491 459644 240557 459645
rect 240491 459580 240492 459644
rect 240556 459580 240557 459644
rect 240491 459579 240557 459580
rect 241779 459644 241845 459645
rect 241779 459580 241780 459644
rect 241844 459580 241845 459644
rect 241779 459579 241845 459580
rect 243251 459644 243317 459645
rect 243251 459580 243252 459644
rect 243316 459580 243317 459644
rect 243251 459579 243317 459580
rect 244539 459644 244605 459645
rect 244539 459580 244540 459644
rect 244604 459580 244605 459644
rect 244539 459579 244605 459580
rect 246011 459644 246077 459645
rect 246011 459580 246012 459644
rect 246076 459580 246077 459644
rect 246011 459579 246077 459580
rect 247299 459644 247365 459645
rect 247299 459580 247300 459644
rect 247364 459580 247365 459644
rect 247299 459579 247365 459580
rect 248771 459644 248837 459645
rect 248771 459580 248772 459644
rect 248836 459580 248837 459644
rect 248771 459579 248837 459580
rect 251531 459644 251597 459645
rect 251531 459580 251532 459644
rect 251596 459580 251597 459644
rect 251531 459579 251597 459580
rect 252819 459644 252885 459645
rect 252819 459580 252820 459644
rect 252884 459580 252885 459644
rect 252819 459579 252885 459580
rect 342795 459644 342861 459645
rect 342795 459580 342796 459644
rect 342860 459580 342861 459644
rect 342795 459579 342861 459580
rect 344083 459644 344149 459645
rect 344083 459580 344084 459644
rect 344148 459580 344149 459644
rect 344083 459579 344149 459580
rect 345555 459644 345621 459645
rect 345555 459580 345556 459644
rect 345620 459580 345621 459644
rect 345555 459579 345621 459580
rect 346843 459644 346909 459645
rect 346843 459580 346844 459644
rect 346908 459580 346909 459644
rect 346843 459579 346909 459580
rect 348315 459644 348381 459645
rect 348315 459580 348316 459644
rect 348380 459580 348381 459644
rect 348315 459579 348381 459580
rect 800 434292 882 434528
rect 1118 434292 1200 434528
rect 800 403892 1200 434292
rect 800 403656 882 403892
rect 1118 403656 1200 403892
rect 800 373256 1200 403656
rect 800 373020 882 373256
rect 1118 373020 1200 373256
rect 800 342620 1200 373020
rect 800 342384 882 342620
rect 1118 342384 1200 342620
rect 800 311984 1200 342384
rect 800 311748 882 311984
rect 1118 311748 1200 311984
rect 800 281348 1200 311748
rect 800 281112 882 281348
rect 1118 281112 1200 281348
rect 800 250712 1200 281112
rect 800 250476 882 250712
rect 1118 250476 1200 250712
rect 800 220076 1200 250476
rect 800 219840 882 220076
rect 1118 219840 1200 220076
rect 800 189440 1200 219840
rect 800 189204 882 189440
rect 1118 189204 1200 189440
rect 800 158804 1200 189204
rect 91451 173908 91517 173909
rect 91451 173844 91452 173908
rect 91516 173844 91517 173908
rect 91451 173843 91517 173844
rect 225403 173908 225469 173909
rect 225403 173844 225404 173908
rect 225468 173844 225469 173908
rect 225403 173843 225469 173844
rect 91454 164253 91514 173843
rect 225406 164253 225466 173843
rect 91451 164252 91517 164253
rect 91451 164188 91452 164252
rect 91516 164188 91517 164252
rect 91451 164187 91517 164188
rect 225403 164252 225469 164253
rect 225403 164188 225404 164252
rect 225468 164188 225469 164252
rect 225403 164187 225469 164188
rect 800 158568 882 158804
rect 1118 158568 1200 158804
rect 800 128168 1200 158568
rect 800 127932 882 128168
rect 1118 127932 1200 128168
rect 800 97532 1200 127932
rect 800 97296 882 97532
rect 1118 97296 1200 97532
rect 800 66896 1200 97296
rect 800 66660 882 66896
rect 1118 66660 1200 66896
rect 800 36260 1200 66660
rect 232214 38997 232274 459579
rect 232211 38996 232277 38997
rect 232211 38932 232212 38996
rect 232276 38932 232277 38996
rect 232211 38931 232277 38932
rect 800 36024 882 36260
rect 1118 36024 1200 36260
rect 800 5624 1200 36024
rect 233502 23493 233562 459579
rect 234598 434528 234918 434570
rect 234598 434292 234640 434528
rect 234876 434292 234918 434528
rect 234598 434250 234918 434292
rect 234598 403892 234918 403934
rect 234598 403656 234640 403892
rect 234876 403656 234918 403892
rect 234598 403614 234918 403656
rect 234598 373256 234918 373298
rect 234598 373020 234640 373256
rect 234876 373020 234918 373256
rect 234598 372978 234918 373020
rect 234598 342620 234918 342662
rect 234598 342384 234640 342620
rect 234876 342384 234918 342620
rect 234598 342342 234918 342384
rect 235523 244356 235589 244357
rect 235523 244292 235524 244356
rect 235588 244292 235589 244356
rect 235523 244291 235589 244292
rect 235526 241637 235586 244291
rect 235523 241636 235589 241637
rect 235523 241572 235524 241636
rect 235588 241572 235589 241636
rect 235523 241571 235589 241572
rect 236262 70413 236322 459579
rect 237734 101149 237794 459579
rect 239022 134061 239082 459579
rect 239019 134060 239085 134061
rect 239019 133996 239020 134060
rect 239084 133996 239085 134060
rect 239019 133995 239085 133996
rect 240494 117333 240554 459579
rect 241782 179621 241842 459579
rect 242515 182068 242581 182069
rect 242515 182004 242516 182068
rect 242580 182004 242581 182068
rect 242515 182003 242581 182004
rect 241779 179620 241845 179621
rect 241779 179556 241780 179620
rect 241844 179556 241845 179620
rect 241779 179555 241845 179556
rect 242518 163029 242578 182003
rect 243254 164253 243314 459579
rect 244542 226677 244602 459579
rect 244539 226676 244605 226677
rect 244539 226612 244540 226676
rect 244604 226612 244605 226676
rect 244539 226611 244605 226612
rect 246014 211173 246074 459579
rect 247302 241773 247362 459579
rect 248774 258093 248834 459579
rect 249958 449846 250278 449888
rect 249958 449610 250000 449846
rect 250236 449610 250278 449846
rect 249958 449568 250278 449610
rect 249958 419210 250278 419252
rect 249958 418974 250000 419210
rect 250236 418974 250278 419210
rect 249958 418932 250278 418974
rect 249958 388574 250278 388616
rect 249958 388338 250000 388574
rect 250236 388338 250278 388574
rect 249958 388296 250278 388338
rect 249958 357938 250278 357980
rect 249958 357702 250000 357938
rect 250236 357702 250278 357938
rect 249958 357660 250278 357702
rect 251534 320517 251594 459579
rect 251531 320516 251597 320517
rect 251531 320452 251532 320516
rect 251596 320452 251597 320516
rect 251531 320451 251597 320452
rect 252822 305013 252882 459579
rect 280603 320652 280669 320653
rect 280603 320588 280604 320652
rect 280668 320650 280669 320652
rect 280668 320590 280850 320650
rect 280668 320588 280669 320590
rect 280603 320587 280669 320588
rect 280790 320245 280850 320590
rect 299923 320516 299989 320517
rect 299923 320452 299924 320516
rect 299988 320452 299989 320516
rect 299923 320451 299989 320452
rect 280787 320244 280853 320245
rect 280787 320180 280788 320244
rect 280852 320180 280853 320244
rect 280787 320179 280853 320180
rect 299926 320109 299986 320451
rect 309491 320380 309557 320381
rect 309491 320316 309492 320380
rect 309556 320316 309557 320380
rect 309491 320315 309557 320316
rect 309494 320109 309554 320315
rect 338563 320244 338629 320245
rect 338563 320180 338564 320244
rect 338628 320180 338629 320244
rect 338563 320179 338629 320180
rect 299923 320108 299989 320109
rect 299923 320044 299924 320108
rect 299988 320044 299989 320108
rect 299923 320043 299989 320044
rect 309491 320108 309557 320109
rect 309491 320044 309492 320108
rect 309556 320044 309557 320108
rect 309491 320043 309557 320044
rect 338566 319973 338626 320179
rect 338563 319972 338629 319973
rect 338563 319908 338564 319972
rect 338628 319908 338629 319972
rect 338563 319907 338629 319908
rect 252819 305012 252885 305013
rect 252819 304948 252820 305012
rect 252884 304948 252885 305012
rect 252819 304947 252885 304948
rect 341139 290188 341205 290189
rect 341139 290124 341140 290188
rect 341204 290124 341205 290188
rect 341139 290123 341205 290124
rect 341142 289917 341202 290123
rect 341139 289916 341205 289917
rect 341139 289852 341140 289916
rect 341204 289852 341205 289916
rect 341139 289851 341205 289852
rect 319979 282980 320045 282981
rect 319979 282916 319980 282980
rect 320044 282916 320045 282980
rect 319979 282915 320045 282916
rect 319982 278901 320042 282915
rect 319979 278900 320045 278901
rect 319979 278836 319980 278900
rect 320044 278836 320045 278900
rect 319979 278835 320045 278836
rect 248771 258092 248837 258093
rect 248771 258028 248772 258092
rect 248836 258028 248837 258092
rect 248771 258027 248837 258028
rect 319979 251156 320045 251157
rect 319979 251092 319980 251156
rect 320044 251092 320045 251156
rect 319979 251091 320045 251092
rect 319059 242452 319125 242453
rect 319059 242388 319060 242452
rect 319124 242388 319125 242452
rect 319059 242387 319125 242388
rect 319062 242045 319122 242387
rect 319059 242044 319125 242045
rect 319059 241980 319060 242044
rect 319124 241980 319125 242044
rect 319059 241979 319125 241980
rect 299923 241908 299989 241909
rect 299923 241844 299924 241908
rect 299988 241844 299989 241908
rect 299923 241843 299989 241844
rect 247299 241772 247365 241773
rect 247299 241708 247300 241772
rect 247364 241708 247365 241772
rect 299926 241770 299986 241843
rect 300107 241772 300173 241773
rect 300107 241770 300108 241772
rect 299926 241710 300108 241770
rect 247299 241707 247365 241708
rect 300107 241708 300108 241710
rect 300172 241708 300173 241772
rect 300107 241707 300173 241708
rect 319982 241637 320042 251091
rect 319979 241636 320045 241637
rect 319979 241572 319980 241636
rect 320044 241572 320045 241636
rect 319979 241571 320045 241572
rect 319059 227220 319125 227221
rect 319059 227156 319060 227220
rect 319124 227156 319125 227220
rect 319059 227155 319125 227156
rect 319062 226813 319122 227155
rect 319059 226812 319125 226813
rect 319059 226748 319060 226812
rect 319124 226748 319125 226812
rect 319059 226747 319125 226748
rect 288883 226676 288949 226677
rect 288883 226612 288884 226676
rect 288948 226612 288949 226676
rect 288883 226611 288949 226612
rect 261283 226540 261349 226541
rect 261283 226476 261284 226540
rect 261348 226476 261349 226540
rect 261283 226475 261349 226476
rect 261286 226269 261346 226475
rect 288886 226405 288946 226611
rect 288883 226404 288949 226405
rect 288883 226340 288884 226404
rect 288948 226340 288949 226404
rect 288883 226339 288949 226340
rect 261283 226268 261349 226269
rect 261283 226204 261284 226268
rect 261348 226204 261349 226268
rect 261283 226203 261349 226204
rect 276555 221508 276621 221509
rect 276555 221444 276556 221508
rect 276620 221444 276621 221508
rect 276555 221443 276621 221444
rect 246011 211172 246077 211173
rect 246011 211108 246012 211172
rect 246076 211108 246077 211172
rect 246011 211107 246077 211108
rect 276558 208453 276618 221443
rect 319979 216068 320045 216069
rect 319979 216004 319980 216068
rect 320044 216004 320045 216068
rect 319979 216003 320045 216004
rect 276555 208452 276621 208453
rect 276555 208388 276556 208452
rect 276620 208388 276621 208452
rect 276555 208387 276621 208388
rect 319982 206277 320042 216003
rect 319979 206276 320045 206277
rect 319979 206212 319980 206276
rect 320044 206212 320045 206276
rect 319979 206211 320045 206212
rect 288883 180028 288949 180029
rect 288883 179964 288884 180028
rect 288948 179964 288949 180028
rect 288883 179963 288949 179964
rect 288886 179757 288946 179963
rect 269563 179756 269629 179757
rect 269563 179692 269564 179756
rect 269628 179692 269629 179756
rect 269563 179691 269629 179692
rect 288883 179756 288949 179757
rect 288883 179692 288884 179756
rect 288948 179692 288949 179756
rect 288883 179691 288949 179692
rect 327523 179756 327589 179757
rect 327523 179692 327524 179756
rect 327588 179692 327589 179756
rect 327523 179691 327589 179692
rect 269566 179485 269626 179691
rect 299923 179620 299989 179621
rect 299923 179556 299924 179620
rect 299988 179556 299989 179620
rect 299923 179555 299989 179556
rect 269563 179484 269629 179485
rect 269563 179420 269564 179484
rect 269628 179420 269629 179484
rect 269563 179419 269629 179420
rect 299926 179213 299986 179555
rect 327526 179485 327586 179691
rect 308203 179484 308269 179485
rect 308203 179420 308204 179484
rect 308268 179420 308269 179484
rect 308203 179419 308269 179420
rect 327523 179484 327589 179485
rect 327523 179420 327524 179484
rect 327588 179420 327589 179484
rect 327523 179419 327589 179420
rect 308206 179213 308266 179419
rect 299923 179212 299989 179213
rect 299923 179148 299924 179212
rect 299988 179148 299989 179212
rect 299923 179147 299989 179148
rect 308203 179212 308269 179213
rect 308203 179148 308204 179212
rect 308268 179148 308269 179212
rect 308203 179147 308269 179148
rect 285387 177308 285453 177309
rect 285387 177244 285388 177308
rect 285452 177244 285453 177308
rect 285387 177243 285453 177244
rect 243251 164252 243317 164253
rect 243251 164188 243252 164252
rect 243316 164188 243317 164252
rect 243251 164187 243317 164188
rect 285390 164117 285450 177243
rect 285387 164116 285453 164117
rect 285387 164052 285388 164116
rect 285452 164052 285453 164116
rect 285387 164051 285453 164052
rect 242515 163028 242581 163029
rect 242515 162964 242516 163028
rect 242580 162964 242581 163028
rect 242515 162963 242581 162964
rect 242515 157860 242581 157861
rect 242515 157796 242516 157860
rect 242580 157796 242581 157860
rect 242515 157795 242581 157796
rect 242518 144941 242578 157795
rect 309307 151740 309373 151741
rect 309307 151676 309308 151740
rect 309372 151676 309373 151740
rect 309307 151675 309373 151676
rect 242515 144940 242581 144941
rect 242515 144876 242516 144940
rect 242580 144876 242581 144940
rect 242515 144875 242581 144876
rect 309310 142221 309370 151675
rect 309307 142220 309373 142221
rect 309307 142156 309308 142220
rect 309372 142156 309373 142220
rect 309307 142155 309373 142156
rect 308203 132836 308269 132837
rect 308203 132772 308204 132836
rect 308268 132772 308269 132836
rect 308203 132771 308269 132772
rect 317771 132836 317837 132837
rect 317771 132772 317772 132836
rect 317836 132772 317837 132836
rect 317771 132771 317837 132772
rect 327523 132836 327589 132837
rect 327523 132772 327524 132836
rect 327588 132772 327589 132836
rect 327523 132771 327589 132772
rect 308206 132565 308266 132771
rect 317774 132565 317834 132771
rect 327526 132565 327586 132771
rect 308203 132564 308269 132565
rect 308203 132500 308204 132564
rect 308268 132500 308269 132564
rect 308203 132499 308269 132500
rect 317771 132564 317837 132565
rect 317771 132500 317772 132564
rect 317836 132500 317837 132564
rect 317771 132499 317837 132500
rect 327523 132564 327589 132565
rect 327523 132500 327524 132564
rect 327588 132500 327589 132564
rect 327523 132499 327589 132500
rect 342798 126989 342858 459579
rect 342795 126988 342861 126989
rect 342795 126924 342796 126988
rect 342860 126924 342861 126988
rect 342795 126923 342861 126924
rect 240491 117332 240557 117333
rect 240491 117268 240492 117332
rect 240556 117268 240557 117332
rect 240491 117267 240557 117268
rect 237731 101148 237797 101149
rect 237731 101084 237732 101148
rect 237796 101084 237797 101148
rect 237731 101083 237797 101084
rect 316483 100876 316549 100877
rect 316483 100812 316484 100876
rect 316548 100812 316549 100876
rect 316483 100811 316549 100812
rect 316486 100605 316546 100811
rect 316483 100604 316549 100605
rect 316483 100540 316484 100604
rect 316548 100540 316549 100604
rect 316483 100539 316549 100540
rect 344086 92445 344146 459579
rect 344083 92444 344149 92445
rect 344083 92380 344084 92444
rect 344148 92380 344149 92444
rect 344083 92379 344149 92380
rect 345558 75853 345618 459579
rect 345555 75852 345621 75853
rect 345555 75788 345556 75852
rect 345620 75788 345621 75852
rect 345555 75787 345621 75788
rect 236259 70412 236325 70413
rect 236259 70348 236260 70412
rect 236324 70348 236325 70412
rect 236259 70347 236325 70348
rect 346846 42805 346906 459579
rect 346843 42804 346909 42805
rect 346843 42740 346844 42804
rect 346908 42740 346909 42804
rect 346843 42739 346909 42740
rect 346659 39268 346725 39269
rect 346659 39204 346660 39268
rect 346724 39204 346725 39268
rect 346659 39203 346725 39204
rect 327523 39132 327589 39133
rect 327523 39068 327524 39132
rect 327588 39068 327589 39132
rect 327523 39067 327589 39068
rect 317771 38996 317837 38997
rect 317771 38932 317772 38996
rect 317836 38932 317837 38996
rect 317771 38931 317837 38932
rect 317774 38725 317834 38931
rect 327526 38725 327586 39067
rect 346662 38725 346722 39203
rect 346843 38996 346909 38997
rect 346843 38932 346844 38996
rect 346908 38932 346909 38996
rect 346843 38931 346909 38932
rect 346846 38725 346906 38931
rect 317771 38724 317837 38725
rect 317771 38660 317772 38724
rect 317836 38660 317837 38724
rect 317771 38659 317837 38660
rect 327523 38724 327589 38725
rect 327523 38660 327524 38724
rect 327588 38660 327589 38724
rect 327523 38659 327589 38660
rect 346659 38724 346725 38725
rect 346659 38660 346660 38724
rect 346724 38660 346725 38724
rect 346659 38659 346725 38660
rect 346843 38724 346909 38725
rect 346843 38660 346844 38724
rect 346908 38660 346909 38724
rect 346843 38659 346909 38660
rect 233499 23492 233565 23493
rect 233499 23428 233500 23492
rect 233564 23428 233565 23492
rect 233499 23427 233565 23428
rect 177195 10164 177261 10165
rect 177195 10100 177196 10164
rect 177260 10100 177261 10164
rect 177195 10099 177261 10100
rect 177011 10028 177077 10029
rect 177011 9964 177012 10028
rect 177076 9964 177077 10028
rect 177011 9963 177077 9964
rect 177014 9890 177074 9963
rect 177198 9890 177258 10099
rect 177014 9830 177258 9890
rect 348318 9621 348378 459579
rect 583716 434528 584116 464928
rect 583716 434292 583798 434528
rect 584034 434292 584116 434528
rect 583716 403892 584116 434292
rect 583716 403656 583798 403892
rect 584034 403656 584116 403892
rect 583716 373256 584116 403656
rect 583716 373020 583798 373256
rect 584034 373020 584116 373256
rect 583716 342620 584116 373020
rect 583716 342384 583798 342620
rect 584034 342384 584116 342620
rect 512443 320516 512509 320517
rect 512443 320452 512444 320516
rect 512508 320452 512509 320516
rect 512443 320451 512509 320452
rect 551083 320516 551149 320517
rect 551083 320452 551084 320516
rect 551148 320452 551149 320516
rect 551083 320451 551149 320452
rect 512446 320245 512506 320451
rect 551086 320245 551146 320451
rect 512443 320244 512509 320245
rect 512443 320180 512444 320244
rect 512508 320180 512509 320244
rect 512443 320179 512509 320180
rect 551083 320244 551149 320245
rect 551083 320180 551084 320244
rect 551148 320180 551149 320244
rect 551083 320179 551149 320180
rect 385483 319156 385549 319157
rect 385483 319092 385484 319156
rect 385548 319092 385549 319156
rect 385483 319091 385549 319092
rect 385486 318885 385546 319091
rect 385483 318884 385549 318885
rect 385483 318820 385484 318884
rect 385548 318820 385549 318884
rect 385483 318819 385549 318820
rect 583716 311984 584116 342384
rect 583716 311748 583798 311984
rect 584034 311748 584116 311984
rect 583716 281348 584116 311748
rect 583716 281112 583798 281348
rect 584034 281112 584116 281348
rect 583716 250712 584116 281112
rect 583716 250476 583798 250712
rect 584034 250476 584116 250712
rect 377203 242180 377269 242181
rect 377203 242116 377204 242180
rect 377268 242116 377269 242180
rect 377203 242115 377269 242116
rect 377206 241773 377266 242115
rect 551083 241908 551149 241909
rect 551083 241844 551084 241908
rect 551148 241844 551149 241908
rect 551083 241843 551149 241844
rect 377203 241772 377269 241773
rect 377203 241708 377204 241772
rect 377268 241708 377269 241772
rect 377203 241707 377269 241708
rect 551086 241637 551146 241843
rect 551083 241636 551149 241637
rect 551083 241572 551084 241636
rect 551148 241572 551149 241636
rect 551083 241571 551149 241572
rect 551083 226676 551149 226677
rect 551083 226612 551084 226676
rect 551148 226612 551149 226676
rect 551083 226611 551149 226612
rect 551086 226405 551146 226611
rect 551083 226404 551149 226405
rect 551083 226340 551084 226404
rect 551148 226340 551149 226404
rect 551083 226339 551149 226340
rect 583716 220076 584116 250476
rect 583716 219840 583798 220076
rect 584034 219840 584116 220076
rect 583716 189440 584116 219840
rect 583716 189204 583798 189440
rect 584034 189204 584116 189440
rect 553843 183564 553909 183565
rect 553843 183500 553844 183564
rect 553908 183500 553909 183564
rect 553843 183499 553909 183500
rect 356595 179756 356661 179757
rect 356595 179692 356596 179756
rect 356660 179692 356661 179756
rect 356595 179691 356661 179692
rect 396523 179756 396589 179757
rect 396523 179692 396524 179756
rect 396588 179692 396589 179756
rect 396523 179691 396589 179692
rect 551083 179756 551149 179757
rect 551083 179692 551084 179756
rect 551148 179692 551149 179756
rect 551083 179691 551149 179692
rect 356598 179349 356658 179691
rect 396526 179485 396586 179691
rect 551086 179485 551146 179691
rect 396523 179484 396589 179485
rect 396523 179420 396524 179484
rect 396588 179420 396589 179484
rect 396523 179419 396589 179420
rect 551083 179484 551149 179485
rect 551083 179420 551084 179484
rect 551148 179420 551149 179484
rect 551083 179419 551149 179420
rect 356595 179348 356661 179349
rect 356595 179284 356596 179348
rect 356660 179284 356661 179348
rect 356595 179283 356661 179284
rect 553846 174045 553906 183499
rect 553843 174044 553909 174045
rect 553843 173980 553844 174044
rect 553908 173980 553909 174044
rect 553843 173979 553909 173980
rect 357883 173908 357949 173909
rect 357883 173844 357884 173908
rect 357948 173844 357949 173908
rect 357883 173843 357949 173844
rect 357886 164389 357946 173843
rect 560835 164660 560901 164661
rect 560835 164596 560836 164660
rect 560900 164596 560901 164660
rect 560835 164595 560901 164596
rect 357883 164388 357949 164389
rect 357883 164324 357884 164388
rect 357948 164324 357949 164388
rect 357883 164323 357949 164324
rect 560838 164253 560898 164595
rect 560835 164252 560901 164253
rect 560835 164188 560836 164252
rect 560900 164188 560901 164252
rect 560835 164187 560901 164188
rect 583716 158804 584116 189204
rect 583716 158568 583798 158804
rect 584034 158568 584116 158804
rect 357883 133108 357949 133109
rect 357883 133044 357884 133108
rect 357948 133044 357949 133108
rect 357883 133043 357949 133044
rect 366163 133108 366229 133109
rect 366163 133044 366164 133108
rect 366228 133044 366229 133108
rect 366163 133043 366229 133044
rect 357886 132837 357946 133043
rect 357883 132836 357949 132837
rect 357883 132772 357884 132836
rect 357948 132772 357949 132836
rect 357883 132771 357949 132772
rect 366166 132701 366226 133043
rect 551083 132836 551149 132837
rect 551083 132772 551084 132836
rect 551148 132772 551149 132836
rect 551083 132771 551149 132772
rect 366163 132700 366229 132701
rect 366163 132636 366164 132700
rect 366228 132636 366229 132700
rect 366163 132635 366229 132636
rect 551086 132565 551146 132771
rect 551083 132564 551149 132565
rect 551083 132500 551084 132564
rect 551148 132500 551149 132564
rect 551083 132499 551149 132500
rect 583716 128168 584116 158568
rect 583716 127932 583798 128168
rect 584034 127932 584116 128168
rect 377203 101420 377269 101421
rect 377203 101356 377204 101420
rect 377268 101356 377269 101420
rect 377203 101355 377269 101356
rect 377206 101149 377266 101355
rect 377203 101148 377269 101149
rect 377203 101084 377204 101148
rect 377268 101084 377269 101148
rect 377203 101083 377269 101084
rect 396523 101148 396589 101149
rect 396523 101084 396524 101148
rect 396588 101084 396589 101148
rect 396523 101083 396589 101084
rect 551083 101148 551149 101149
rect 551083 101084 551084 101148
rect 551148 101084 551149 101148
rect 551083 101083 551149 101084
rect 396526 100877 396586 101083
rect 551086 100877 551146 101083
rect 396523 100876 396589 100877
rect 396523 100812 396524 100876
rect 396588 100812 396589 100876
rect 396523 100811 396589 100812
rect 551083 100876 551149 100877
rect 551083 100812 551084 100876
rect 551148 100812 551149 100876
rect 551083 100811 551149 100812
rect 583716 97532 584116 127932
rect 583716 97296 583798 97532
rect 584034 97296 584116 97532
rect 583716 66896 584116 97296
rect 583716 66660 583798 66896
rect 584034 66660 584116 66896
rect 356595 38996 356661 38997
rect 356595 38932 356596 38996
rect 356660 38932 356661 38996
rect 356595 38931 356661 38932
rect 551083 38996 551149 38997
rect 551083 38932 551084 38996
rect 551148 38932 551149 38996
rect 551083 38931 551149 38932
rect 356598 38589 356658 38931
rect 551086 38725 551146 38931
rect 551083 38724 551149 38725
rect 551083 38660 551084 38724
rect 551148 38660 551149 38724
rect 551083 38659 551149 38660
rect 356595 38588 356661 38589
rect 356595 38524 356596 38588
rect 356660 38524 356661 38588
rect 356595 38523 356661 38524
rect 583716 36260 584116 66660
rect 583716 36024 583798 36260
rect 584034 36024 584116 36260
rect 348315 9620 348381 9621
rect 348315 9556 348316 9620
rect 348380 9556 348381 9620
rect 348315 9555 348381 9556
rect 250243 7580 250309 7581
rect 250243 7516 250244 7580
rect 250308 7516 250309 7580
rect 250243 7515 250309 7516
rect 501403 7580 501469 7581
rect 501403 7516 501404 7580
rect 501468 7516 501469 7580
rect 501403 7515 501469 7516
rect 250246 7309 250306 7515
rect 393763 7444 393829 7445
rect 393763 7380 393764 7444
rect 393828 7380 393829 7444
rect 393763 7379 393829 7380
rect 250243 7308 250309 7309
rect 250243 7244 250244 7308
rect 250308 7244 250309 7308
rect 250243 7243 250309 7244
rect 308203 7308 308269 7309
rect 308203 7244 308204 7308
rect 308268 7244 308269 7308
rect 308203 7243 308269 7244
rect 292931 7172 292997 7173
rect 292931 7108 292932 7172
rect 292996 7170 292997 7172
rect 293115 7172 293181 7173
rect 293115 7170 293116 7172
rect 292996 7110 293116 7170
rect 292996 7108 292997 7110
rect 292931 7107 292997 7108
rect 293115 7108 293116 7110
rect 293180 7108 293181 7172
rect 293115 7107 293181 7108
rect 299923 7172 299989 7173
rect 299923 7108 299924 7172
rect 299988 7170 299989 7172
rect 299988 7110 300170 7170
rect 299988 7108 299989 7110
rect 299923 7107 299989 7108
rect 300110 6901 300170 7110
rect 308206 6901 308266 7243
rect 375731 7172 375797 7173
rect 375731 7108 375732 7172
rect 375796 7170 375797 7172
rect 375796 7110 375978 7170
rect 375796 7108 375797 7110
rect 375731 7107 375797 7108
rect 346659 7036 346725 7037
rect 346659 6972 346660 7036
rect 346724 6972 346725 7036
rect 346659 6971 346725 6972
rect 346843 7036 346909 7037
rect 346843 6972 346844 7036
rect 346908 6972 346909 7036
rect 346843 6971 346909 6972
rect 300107 6900 300173 6901
rect 300107 6836 300108 6900
rect 300172 6836 300173 6900
rect 300107 6835 300173 6836
rect 308203 6900 308269 6901
rect 308203 6836 308204 6900
rect 308268 6836 308269 6900
rect 308203 6835 308269 6836
rect 346662 6765 346722 6971
rect 346846 6765 346906 6971
rect 375918 6901 375978 7110
rect 393766 7037 393826 7379
rect 501406 7309 501466 7515
rect 537283 7444 537349 7445
rect 537283 7380 537284 7444
rect 537348 7380 537349 7444
rect 537283 7379 537349 7380
rect 501403 7308 501469 7309
rect 501403 7244 501404 7308
rect 501468 7244 501469 7308
rect 501403 7243 501469 7244
rect 537286 7173 537346 7379
rect 443443 7172 443509 7173
rect 443443 7108 443444 7172
rect 443508 7108 443509 7172
rect 443443 7107 443509 7108
rect 537283 7172 537349 7173
rect 537283 7108 537284 7172
rect 537348 7108 537349 7172
rect 537283 7107 537349 7108
rect 393763 7036 393829 7037
rect 393763 6972 393764 7036
rect 393828 6972 393829 7036
rect 393763 6971 393829 6972
rect 443446 6901 443506 7107
rect 375915 6900 375981 6901
rect 375915 6836 375916 6900
rect 375980 6836 375981 6900
rect 375915 6835 375981 6836
rect 382723 6900 382789 6901
rect 382723 6836 382724 6900
rect 382788 6836 382789 6900
rect 382723 6835 382789 6836
rect 443443 6900 443509 6901
rect 443443 6836 443444 6900
rect 443508 6836 443509 6900
rect 443443 6835 443509 6836
rect 346659 6764 346725 6765
rect 346659 6700 346660 6764
rect 346724 6700 346725 6764
rect 346659 6699 346725 6700
rect 346843 6764 346909 6765
rect 346843 6700 346844 6764
rect 346908 6700 346909 6764
rect 346843 6699 346909 6700
rect 382726 6629 382786 6835
rect 382723 6628 382789 6629
rect 382723 6564 382724 6628
rect 382788 6564 382789 6628
rect 382723 6563 382789 6564
rect 222643 6084 222709 6085
rect 222643 6020 222644 6084
rect 222708 6020 222709 6084
rect 222643 6019 222709 6020
rect 800 5388 882 5624
rect 1118 5388 1200 5624
rect 800 1694 1200 5388
rect 145363 3364 145429 3365
rect 145363 3300 145364 3364
rect 145428 3300 145429 3364
rect 145363 3299 145429 3300
rect 145366 3093 145426 3299
rect 145363 3092 145429 3093
rect 145363 3028 145364 3092
rect 145428 3028 145429 3092
rect 145363 3027 145429 3028
rect 222646 2821 222706 6019
rect 583716 5624 584116 36024
rect 583716 5388 583798 5624
rect 584034 5388 584116 5624
rect 347950 3710 348562 3770
rect 347950 3637 348010 3710
rect 348502 3637 348562 3710
rect 347947 3636 348013 3637
rect 347947 3572 347948 3636
rect 348012 3572 348013 3636
rect 347947 3571 348013 3572
rect 348499 3636 348565 3637
rect 348499 3572 348500 3636
rect 348564 3572 348565 3636
rect 348499 3571 348565 3572
rect 222643 2820 222709 2821
rect 222643 2756 222644 2820
rect 222708 2756 222709 2820
rect 222643 2755 222709 2756
rect 800 1458 882 1694
rect 1118 1458 1200 1694
rect 800 1376 1200 1458
rect 583716 1694 584116 5388
rect 583716 1458 583798 1694
rect 584034 1458 584116 1694
rect 583716 1376 584116 1458
rect 584516 694934 584916 703042
rect 584516 694698 584598 694934
rect 584834 694698 584916 694934
rect 584516 664298 584916 694698
rect 584516 664062 584598 664298
rect 584834 664062 584916 664298
rect 584516 633662 584916 664062
rect 584516 633426 584598 633662
rect 584834 633426 584916 633662
rect 584516 603026 584916 633426
rect 584516 602790 584598 603026
rect 584834 602790 584916 603026
rect 584516 572390 584916 602790
rect 584516 572154 584598 572390
rect 584834 572154 584916 572390
rect 584516 541754 584916 572154
rect 584516 541518 584598 541754
rect 584834 541518 584916 541754
rect 584516 511118 584916 541518
rect 584516 510882 584598 511118
rect 584834 510882 584916 511118
rect 584516 480482 584916 510882
rect 584516 480246 584598 480482
rect 584834 480246 584916 480482
rect 584516 449846 584916 480246
rect 584516 449610 584598 449846
rect 584834 449610 584916 449846
rect 584516 419210 584916 449610
rect 584516 418974 584598 419210
rect 584834 418974 584916 419210
rect 584516 388574 584916 418974
rect 584516 388338 584598 388574
rect 584834 388338 584916 388574
rect 584516 357938 584916 388338
rect 584516 357702 584598 357938
rect 584834 357702 584916 357938
rect 584516 327302 584916 357702
rect 584516 327066 584598 327302
rect 584834 327066 584916 327302
rect 584516 296666 584916 327066
rect 584516 296430 584598 296666
rect 584834 296430 584916 296666
rect 584516 266030 584916 296430
rect 584516 265794 584598 266030
rect 584834 265794 584916 266030
rect 584516 235394 584916 265794
rect 584516 235158 584598 235394
rect 584834 235158 584916 235394
rect 584516 204758 584916 235158
rect 584516 204522 584598 204758
rect 584834 204522 584916 204758
rect 584516 174122 584916 204522
rect 584516 173886 584598 174122
rect 584834 173886 584916 174122
rect 584516 143486 584916 173886
rect 584516 143250 584598 143486
rect 584834 143250 584916 143486
rect 584516 112850 584916 143250
rect 584516 112614 584598 112850
rect 584834 112614 584916 112850
rect 584516 82214 584916 112614
rect 584516 81978 584598 82214
rect 584834 81978 584916 82214
rect 584516 51578 584916 81978
rect 584516 51342 584598 51578
rect 584834 51342 584916 51578
rect 584516 20942 584916 51342
rect 584516 20706 584598 20942
rect 584834 20706 584916 20942
rect 0 658 82 894
rect 318 658 400 894
rect 0 576 400 658
rect 584516 894 584916 20706
rect 584516 658 584598 894
rect 584834 658 584916 894
rect 584516 576 584916 658
<< via4 >>
rect 82 703042 318 703278
rect 584598 703042 584834 703278
rect 82 694698 318 694934
rect 82 664062 318 664298
rect 82 633426 318 633662
rect 82 602790 318 603026
rect 82 572154 318 572390
rect 82 541518 318 541754
rect 82 510882 318 511118
rect 82 480246 318 480482
rect 82 449610 318 449846
rect 82 418974 318 419210
rect 82 388338 318 388574
rect 82 357702 318 357938
rect 82 327066 318 327302
rect 82 296430 318 296666
rect 82 265794 318 266030
rect 82 235158 318 235394
rect 82 204522 318 204758
rect 82 173886 318 174122
rect 82 143250 318 143486
rect 82 112614 318 112850
rect 82 81978 318 82214
rect 82 51342 318 51578
rect 82 20706 318 20942
rect 882 702242 1118 702478
rect 882 679380 1118 679616
rect 882 648744 1118 648980
rect 882 618108 1118 618344
rect 583798 702242 584034 702478
rect 583798 679380 584034 679616
rect 583798 648744 584034 648980
rect 583798 618108 584034 618344
rect 882 587472 1118 587708
rect 882 556836 1118 557072
rect 583798 587472 584034 587708
rect 583798 556836 584034 557072
rect 882 526200 1118 526436
rect 583798 526200 584034 526436
rect 882 495564 1118 495800
rect 882 464928 1118 465164
rect 583798 495564 584034 495800
rect 583798 464928 584034 465164
rect 882 434292 1118 434528
rect 882 403656 1118 403892
rect 882 373020 1118 373256
rect 882 342384 1118 342620
rect 882 311748 1118 311984
rect 882 281112 1118 281348
rect 882 250476 1118 250712
rect 882 219840 1118 220076
rect 882 189204 1118 189440
rect 882 158568 1118 158804
rect 882 127932 1118 128168
rect 882 97296 1118 97532
rect 882 66660 1118 66896
rect 882 36024 1118 36260
rect 234640 434292 234876 434528
rect 234640 403656 234876 403892
rect 234640 373020 234876 373256
rect 234640 342384 234876 342620
rect 250000 449610 250236 449846
rect 250000 418974 250236 419210
rect 250000 388338 250236 388574
rect 250000 357702 250236 357938
rect 583798 434292 584034 434528
rect 583798 403656 584034 403892
rect 583798 373020 584034 373256
rect 583798 342384 584034 342620
rect 583798 311748 584034 311984
rect 583798 281112 584034 281348
rect 583798 250476 584034 250712
rect 583798 219840 584034 220076
rect 583798 189204 584034 189440
rect 583798 158568 584034 158804
rect 583798 127932 584034 128168
rect 583798 97296 584034 97532
rect 583798 66660 584034 66896
rect 583798 36024 584034 36260
rect 882 5388 1118 5624
rect 583798 5388 584034 5624
rect 882 1458 1118 1694
rect 583798 1458 584034 1694
rect 584598 694698 584834 694934
rect 584598 664062 584834 664298
rect 584598 633426 584834 633662
rect 584598 602790 584834 603026
rect 584598 572154 584834 572390
rect 584598 541518 584834 541754
rect 584598 510882 584834 511118
rect 584598 480246 584834 480482
rect 584598 449610 584834 449846
rect 584598 418974 584834 419210
rect 584598 388338 584834 388574
rect 584598 357702 584834 357938
rect 584598 327066 584834 327302
rect 584598 296430 584834 296666
rect 584598 265794 584834 266030
rect 584598 235158 584834 235394
rect 584598 204522 584834 204758
rect 584598 173886 584834 174122
rect 584598 143250 584834 143486
rect 584598 112614 584834 112850
rect 584598 81978 584834 82214
rect 584598 51342 584834 51578
rect 584598 20706 584834 20942
rect 82 658 318 894
rect 584598 658 584834 894
<< metal5 >>
rect 0 703278 584916 703360
rect 0 703042 82 703278
rect 318 703042 584598 703278
rect 584834 703042 584916 703278
rect 0 702960 584916 703042
rect 800 702478 584116 702560
rect 800 702242 882 702478
rect 1118 702242 583798 702478
rect 584034 702242 584116 702478
rect 800 702160 584116 702242
rect 0 694934 584916 694976
rect 0 694698 82 694934
rect 318 694698 584598 694934
rect 584834 694698 584916 694934
rect 0 694656 584916 694698
rect 0 679616 584916 679658
rect 0 679380 882 679616
rect 1118 679380 583798 679616
rect 584034 679380 584916 679616
rect 0 679338 584916 679380
rect 0 664298 584916 664340
rect 0 664062 82 664298
rect 318 664062 584598 664298
rect 584834 664062 584916 664298
rect 0 664020 584916 664062
rect 0 648980 584916 649022
rect 0 648744 882 648980
rect 1118 648744 583798 648980
rect 584034 648744 584916 648980
rect 0 648702 584916 648744
rect 0 633662 584916 633704
rect 0 633426 82 633662
rect 318 633426 584598 633662
rect 584834 633426 584916 633662
rect 0 633384 584916 633426
rect 0 618344 584916 618386
rect 0 618108 882 618344
rect 1118 618108 583798 618344
rect 584034 618108 584916 618344
rect 0 618066 584916 618108
rect 0 603026 584916 603068
rect 0 602790 82 603026
rect 318 602790 584598 603026
rect 584834 602790 584916 603026
rect 0 602748 584916 602790
rect 0 587708 584916 587750
rect 0 587472 882 587708
rect 1118 587472 583798 587708
rect 584034 587472 584916 587708
rect 0 587430 584916 587472
rect 0 572390 584916 572432
rect 0 572154 82 572390
rect 318 572154 584598 572390
rect 584834 572154 584916 572390
rect 0 572112 584916 572154
rect 0 557072 584916 557114
rect 0 556836 882 557072
rect 1118 556836 583798 557072
rect 584034 556836 584916 557072
rect 0 556794 584916 556836
rect 0 541754 584916 541796
rect 0 541518 82 541754
rect 318 541518 584598 541754
rect 584834 541518 584916 541754
rect 0 541476 584916 541518
rect 0 526436 584916 526478
rect 0 526200 882 526436
rect 1118 526200 583798 526436
rect 584034 526200 584916 526436
rect 0 526158 584916 526200
rect 0 511118 584916 511160
rect 0 510882 82 511118
rect 318 510882 584598 511118
rect 584834 510882 584916 511118
rect 0 510840 584916 510882
rect 0 495800 584916 495842
rect 0 495564 882 495800
rect 1118 495564 583798 495800
rect 584034 495564 584916 495800
rect 0 495522 584916 495564
rect 0 480482 584916 480524
rect 0 480246 82 480482
rect 318 480246 584598 480482
rect 584834 480246 584916 480482
rect 0 480204 584916 480246
rect 0 465164 584916 465206
rect 0 464928 882 465164
rect 1118 464928 583798 465164
rect 584034 464928 584916 465164
rect 0 464886 584916 464928
rect 0 449846 584916 449888
rect 0 449610 82 449846
rect 318 449610 250000 449846
rect 250236 449610 584598 449846
rect 584834 449610 584916 449846
rect 0 449568 584916 449610
rect 0 434528 584916 434570
rect 0 434292 882 434528
rect 1118 434292 234640 434528
rect 234876 434292 583798 434528
rect 584034 434292 584916 434528
rect 0 434250 584916 434292
rect 0 419210 584916 419252
rect 0 418974 82 419210
rect 318 418974 250000 419210
rect 250236 418974 584598 419210
rect 584834 418974 584916 419210
rect 0 418932 584916 418974
rect 0 403892 584916 403934
rect 0 403656 882 403892
rect 1118 403656 234640 403892
rect 234876 403656 583798 403892
rect 584034 403656 584916 403892
rect 0 403614 584916 403656
rect 0 388574 584916 388616
rect 0 388338 82 388574
rect 318 388338 250000 388574
rect 250236 388338 584598 388574
rect 584834 388338 584916 388574
rect 0 388296 584916 388338
rect 0 373256 584916 373298
rect 0 373020 882 373256
rect 1118 373020 234640 373256
rect 234876 373020 583798 373256
rect 584034 373020 584916 373256
rect 0 372978 584916 373020
rect 0 357938 584916 357980
rect 0 357702 82 357938
rect 318 357702 250000 357938
rect 250236 357702 584598 357938
rect 584834 357702 584916 357938
rect 0 357660 584916 357702
rect 0 342620 584916 342662
rect 0 342384 882 342620
rect 1118 342384 234640 342620
rect 234876 342384 583798 342620
rect 584034 342384 584916 342620
rect 0 342342 584916 342384
rect 0 327302 584916 327344
rect 0 327066 82 327302
rect 318 327066 584598 327302
rect 584834 327066 584916 327302
rect 0 327024 584916 327066
rect 0 311984 584916 312026
rect 0 311748 882 311984
rect 1118 311748 583798 311984
rect 584034 311748 584916 311984
rect 0 311706 584916 311748
rect 0 296666 584916 296708
rect 0 296430 82 296666
rect 318 296430 584598 296666
rect 584834 296430 584916 296666
rect 0 296388 584916 296430
rect 0 281348 584916 281390
rect 0 281112 882 281348
rect 1118 281112 583798 281348
rect 584034 281112 584916 281348
rect 0 281070 584916 281112
rect 0 266030 584916 266072
rect 0 265794 82 266030
rect 318 265794 584598 266030
rect 584834 265794 584916 266030
rect 0 265752 584916 265794
rect 0 250712 584916 250754
rect 0 250476 882 250712
rect 1118 250476 583798 250712
rect 584034 250476 584916 250712
rect 0 250434 584916 250476
rect 0 235394 584916 235436
rect 0 235158 82 235394
rect 318 235158 584598 235394
rect 584834 235158 584916 235394
rect 0 235116 584916 235158
rect 0 220076 584916 220118
rect 0 219840 882 220076
rect 1118 219840 583798 220076
rect 584034 219840 584916 220076
rect 0 219798 584916 219840
rect 0 204758 584916 204800
rect 0 204522 82 204758
rect 318 204522 584598 204758
rect 584834 204522 584916 204758
rect 0 204480 584916 204522
rect 0 189440 584916 189482
rect 0 189204 882 189440
rect 1118 189204 583798 189440
rect 584034 189204 584916 189440
rect 0 189162 584916 189204
rect 0 174122 584916 174164
rect 0 173886 82 174122
rect 318 173886 584598 174122
rect 584834 173886 584916 174122
rect 0 173844 584916 173886
rect 0 158804 584916 158846
rect 0 158568 882 158804
rect 1118 158568 583798 158804
rect 584034 158568 584916 158804
rect 0 158526 584916 158568
rect 0 143486 584916 143528
rect 0 143250 82 143486
rect 318 143250 584598 143486
rect 584834 143250 584916 143486
rect 0 143208 584916 143250
rect 0 128168 584916 128210
rect 0 127932 882 128168
rect 1118 127932 583798 128168
rect 584034 127932 584916 128168
rect 0 127890 584916 127932
rect 0 112850 584916 112892
rect 0 112614 82 112850
rect 318 112614 584598 112850
rect 584834 112614 584916 112850
rect 0 112572 584916 112614
rect 0 97532 584916 97574
rect 0 97296 882 97532
rect 1118 97296 583798 97532
rect 584034 97296 584916 97532
rect 0 97254 584916 97296
rect 0 82214 584916 82256
rect 0 81978 82 82214
rect 318 81978 584598 82214
rect 584834 81978 584916 82214
rect 0 81936 584916 81978
rect 0 66896 584916 66938
rect 0 66660 882 66896
rect 1118 66660 583798 66896
rect 584034 66660 584916 66896
rect 0 66618 584916 66660
rect 0 51578 584916 51620
rect 0 51342 82 51578
rect 318 51342 584598 51578
rect 584834 51342 584916 51578
rect 0 51300 584916 51342
rect 0 36260 584916 36302
rect 0 36024 882 36260
rect 1118 36024 583798 36260
rect 584034 36024 584916 36260
rect 0 35982 584916 36024
rect 0 20942 584916 20984
rect 0 20706 82 20942
rect 318 20706 584598 20942
rect 584834 20706 584916 20942
rect 0 20664 584916 20706
rect 0 5624 584916 5666
rect 0 5388 882 5624
rect 1118 5388 583798 5624
rect 584034 5388 584916 5624
rect 0 5346 584916 5388
rect 800 1694 584116 1776
rect 800 1458 882 1694
rect 1118 1458 583798 1694
rect 584034 1458 584116 1694
rect 800 1376 584116 1458
rect 0 894 584916 976
rect 0 658 82 894
rect 318 658 584598 894
rect 584834 658 584916 894
rect 0 576 584916 658
use user_proj_example  mprj
timestamp 1605730173
transform 1 0 230496 0 1 340000
box 0 0 119752 120000
<< labels >>
rlabel metal3 s 584016 7760 584496 7880 4 io_in[0]
port 1 nsew
rlabel metal3 s 584016 476960 584496 477080 4 io_in[10]
port 2 nsew
rlabel metal3 s 584016 523880 584496 524000 4 io_in[11]
port 3 nsew
rlabel metal3 s 584016 570800 584496 570920 4 io_in[12]
port 4 nsew
rlabel metal3 s 584016 617720 584496 617840 4 io_in[13]
port 5 nsew
rlabel metal3 s 584016 664640 584496 664760 4 io_in[14]
port 6 nsew
rlabel metal2 s 573582 703520 573638 704000 4 io_in[15]
port 7 nsew
rlabel metal2 s 508722 703520 508778 704000 4 io_in[16]
port 8 nsew
rlabel metal2 s 443862 703520 443918 704000 4 io_in[17]
port 9 nsew
rlabel metal2 s 378910 703520 378966 704000 4 io_in[18]
port 10 nsew
rlabel metal2 s 314050 703520 314106 704000 4 io_in[19]
port 11 nsew
rlabel metal3 s 584016 54680 584496 54800 4 io_in[1]
port 12 nsew
rlabel metal2 s 249190 703520 249246 704000 4 io_in[20]
port 13 nsew
rlabel metal2 s 184238 703520 184294 704000 4 io_in[21]
port 14 nsew
rlabel metal2 s 119378 703520 119434 704000 4 io_in[22]
port 15 nsew
rlabel metal2 s 54518 703520 54574 704000 4 io_in[23]
port 16 nsew
rlabel metal3 s 496 695376 976 695496 4 io_in[24]
port 17 nsew
rlabel metal3 s 496 645192 976 645312 4 io_in[25]
port 18 nsew
rlabel metal3 s 496 594872 976 594992 4 io_in[26]
port 19 nsew
rlabel metal3 s 496 544552 976 544672 4 io_in[27]
port 20 nsew
rlabel metal3 s 496 494232 976 494352 4 io_in[28]
port 21 nsew
rlabel metal3 s 496 444048 976 444168 4 io_in[29]
port 22 nsew
rlabel metal3 s 584016 101600 584496 101720 4 io_in[2]
port 23 nsew
rlabel metal3 s 496 393728 976 393848 4 io_in[30]
port 24 nsew
rlabel metal3 s 496 343408 976 343528 4 io_in[31]
port 25 nsew
rlabel metal3 s 496 293224 976 293344 4 io_in[32]
port 26 nsew
rlabel metal3 s 496 242904 976 243024 4 io_in[33]
port 27 nsew
rlabel metal3 s 496 192584 976 192704 4 io_in[34]
port 28 nsew
rlabel metal3 s 496 142264 976 142384 4 io_in[35]
port 29 nsew
rlabel metal3 s 496 92080 976 92200 4 io_in[36]
port 30 nsew
rlabel metal3 s 496 41760 976 41880 4 io_in[37]
port 31 nsew
rlabel metal3 s 584016 148520 584496 148640 4 io_in[3]
port 32 nsew
rlabel metal3 s 584016 195440 584496 195560 4 io_in[4]
port 33 nsew
rlabel metal3 s 584016 242360 584496 242480 4 io_in[5]
port 34 nsew
rlabel metal3 s 584016 289280 584496 289400 4 io_in[6]
port 35 nsew
rlabel metal3 s 584016 336200 584496 336320 4 io_in[7]
port 36 nsew
rlabel metal3 s 584016 383120 584496 383240 4 io_in[8]
port 37 nsew
rlabel metal3 s 584016 430040 584496 430160 4 io_in[9]
port 38 nsew
rlabel metal3 s 584016 39040 584496 39160 4 io_oeb[0]
port 39 nsew
rlabel metal3 s 584016 508240 584496 508360 4 io_oeb[10]
port 40 nsew
rlabel metal3 s 584016 555160 584496 555280 4 io_oeb[11]
port 41 nsew
rlabel metal3 s 584016 602080 584496 602200 4 io_oeb[12]
port 42 nsew
rlabel metal3 s 584016 649000 584496 649120 4 io_oeb[13]
port 43 nsew
rlabel metal3 s 584016 695920 584496 696040 4 io_oeb[14]
port 44 nsew
rlabel metal2 s 530342 703520 530398 704000 4 io_oeb[15]
port 45 nsew
rlabel metal2 s 465482 703520 465538 704000 4 io_oeb[16]
port 46 nsew
rlabel metal2 s 400622 703520 400678 704000 4 io_oeb[17]
port 47 nsew
rlabel metal2 s 335670 703520 335726 704000 4 io_oeb[18]
port 48 nsew
rlabel metal2 s 270810 703520 270866 704000 4 io_oeb[19]
port 49 nsew
rlabel metal3 s 584016 85960 584496 86080 4 io_oeb[1]
port 50 nsew
rlabel metal2 s 205950 703520 206006 704000 4 io_oeb[20]
port 51 nsew
rlabel metal2 s 140998 703520 141054 704000 4 io_oeb[21]
port 52 nsew
rlabel metal2 s 76138 703520 76194 704000 4 io_oeb[22]
port 53 nsew
rlabel metal2 s 11278 703520 11334 704000 4 io_oeb[23]
port 54 nsew
rlabel metal3 s 496 661920 976 662040 4 io_oeb[24]
port 55 nsew
rlabel metal3 s 496 611600 976 611720 4 io_oeb[25]
port 56 nsew
rlabel metal3 s 496 561280 976 561400 4 io_oeb[26]
port 57 nsew
rlabel metal3 s 496 511096 976 511216 4 io_oeb[27]
port 58 nsew
rlabel metal3 s 496 460776 976 460896 4 io_oeb[28]
port 59 nsew
rlabel metal3 s 496 410456 976 410576 4 io_oeb[29]
port 60 nsew
rlabel metal3 s 584016 132880 584496 133000 4 io_oeb[2]
port 61 nsew
rlabel metal3 s 496 360272 976 360392 4 io_oeb[30]
port 62 nsew
rlabel metal3 s 496 309952 976 310072 4 io_oeb[31]
port 63 nsew
rlabel metal3 s 496 259632 976 259752 4 io_oeb[32]
port 64 nsew
rlabel metal3 s 496 209312 976 209432 4 io_oeb[33]
port 65 nsew
rlabel metal3 s 496 159128 976 159248 4 io_oeb[34]
port 66 nsew
rlabel metal3 s 496 108808 976 108928 4 io_oeb[35]
port 67 nsew
rlabel metal3 s 496 58488 976 58608 4 io_oeb[36]
port 68 nsew
rlabel metal3 s 496 8304 976 8424 4 io_oeb[37]
port 69 nsew
rlabel metal3 s 584016 179800 584496 179920 4 io_oeb[3]
port 70 nsew
rlabel metal3 s 584016 226720 584496 226840 4 io_oeb[4]
port 71 nsew
rlabel metal3 s 584016 273640 584496 273760 4 io_oeb[5]
port 72 nsew
rlabel metal3 s 584016 320560 584496 320680 4 io_oeb[6]
port 73 nsew
rlabel metal3 s 584016 367480 584496 367600 4 io_oeb[7]
port 74 nsew
rlabel metal3 s 584016 414400 584496 414520 4 io_oeb[8]
port 75 nsew
rlabel metal3 s 584016 461320 584496 461440 4 io_oeb[9]
port 76 nsew
rlabel metal3 s 584016 23400 584496 23520 4 io_out[0]
port 77 nsew
rlabel metal3 s 584016 492600 584496 492720 4 io_out[10]
port 78 nsew
rlabel metal3 s 584016 539520 584496 539640 4 io_out[11]
port 79 nsew
rlabel metal3 s 584016 586440 584496 586560 4 io_out[12]
port 80 nsew
rlabel metal3 s 584016 633360 584496 633480 4 io_out[13]
port 81 nsew
rlabel metal3 s 584016 680280 584496 680400 4 io_out[14]
port 82 nsew
rlabel metal2 s 551962 703520 552018 704000 4 io_out[15]
port 83 nsew
rlabel metal2 s 487102 703520 487158 704000 4 io_out[16]
port 84 nsew
rlabel metal2 s 422242 703520 422298 704000 4 io_out[17]
port 85 nsew
rlabel metal2 s 357290 703520 357346 704000 4 io_out[18]
port 86 nsew
rlabel metal2 s 292430 703520 292486 704000 4 io_out[19]
port 87 nsew
rlabel metal3 s 584016 70320 584496 70440 4 io_out[1]
port 88 nsew
rlabel metal2 s 227570 703520 227626 704000 4 io_out[20]
port 89 nsew
rlabel metal2 s 162618 703520 162674 704000 4 io_out[21]
port 90 nsew
rlabel metal2 s 97758 703520 97814 704000 4 io_out[22]
port 91 nsew
rlabel metal2 s 32898 703520 32954 704000 4 io_out[23]
port 92 nsew
rlabel metal3 s 496 678648 976 678768 4 io_out[24]
port 93 nsew
rlabel metal3 s 496 628328 976 628448 4 io_out[25]
port 94 nsew
rlabel metal3 s 496 578144 976 578264 4 io_out[26]
port 95 nsew
rlabel metal3 s 496 527824 976 527944 4 io_out[27]
port 96 nsew
rlabel metal3 s 496 477504 976 477624 4 io_out[28]
port 97 nsew
rlabel metal3 s 496 427184 976 427304 4 io_out[29]
port 98 nsew
rlabel metal3 s 584016 117240 584496 117360 4 io_out[2]
port 99 nsew
rlabel metal3 s 496 377000 976 377120 4 io_out[30]
port 100 nsew
rlabel metal3 s 496 326680 976 326800 4 io_out[31]
port 101 nsew
rlabel metal3 s 496 276360 976 276480 4 io_out[32]
port 102 nsew
rlabel metal3 s 496 226176 976 226296 4 io_out[33]
port 103 nsew
rlabel metal3 s 496 175856 976 175976 4 io_out[34]
port 104 nsew
rlabel metal3 s 496 125536 976 125656 4 io_out[35]
port 105 nsew
rlabel metal3 s 496 75216 976 75336 4 io_out[36]
port 106 nsew
rlabel metal3 s 496 25032 976 25152 4 io_out[37]
port 107 nsew
rlabel metal3 s 584016 164160 584496 164280 4 io_out[3]
port 108 nsew
rlabel metal3 s 584016 211080 584496 211200 4 io_out[4]
port 109 nsew
rlabel metal3 s 584016 258000 584496 258120 4 io_out[5]
port 110 nsew
rlabel metal3 s 584016 304920 584496 305040 4 io_out[6]
port 111 nsew
rlabel metal3 s 584016 351840 584496 351960 4 io_out[7]
port 112 nsew
rlabel metal3 s 584016 398760 584496 398880 4 io_out[8]
port 113 nsew
rlabel metal3 s 584016 445680 584496 445800 4 io_out[9]
port 114 nsew
rlabel metal2 s 127106 0 127162 480 4 la_data_in[0]
port 115 nsew
rlabel metal2 s 483974 0 484030 480 4 la_data_in[100]
port 116 nsew
rlabel metal2 s 487470 0 487526 480 4 la_data_in[101]
port 117 nsew
rlabel metal2 s 491058 0 491114 480 4 la_data_in[102]
port 118 nsew
rlabel metal2 s 494646 0 494702 480 4 la_data_in[103]
port 119 nsew
rlabel metal2 s 498234 0 498290 480 4 la_data_in[104]
port 120 nsew
rlabel metal2 s 501730 0 501786 480 4 la_data_in[105]
port 121 nsew
rlabel metal2 s 505318 0 505374 480 4 la_data_in[106]
port 122 nsew
rlabel metal2 s 508906 0 508962 480 4 la_data_in[107]
port 123 nsew
rlabel metal2 s 512494 0 512550 480 4 la_data_in[108]
port 124 nsew
rlabel metal2 s 516082 0 516138 480 4 la_data_in[109]
port 125 nsew
rlabel metal2 s 162802 0 162858 480 4 la_data_in[10]
port 126 nsew
rlabel metal2 s 519578 0 519634 480 4 la_data_in[110]
port 127 nsew
rlabel metal2 s 523166 0 523222 480 4 la_data_in[111]
port 128 nsew
rlabel metal2 s 526754 0 526810 480 4 la_data_in[112]
port 129 nsew
rlabel metal2 s 530342 0 530398 480 4 la_data_in[113]
port 130 nsew
rlabel metal2 s 533930 0 533986 480 4 la_data_in[114]
port 131 nsew
rlabel metal2 s 537426 0 537482 480 4 la_data_in[115]
port 132 nsew
rlabel metal2 s 541014 0 541070 480 4 la_data_in[116]
port 133 nsew
rlabel metal2 s 544602 0 544658 480 4 la_data_in[117]
port 134 nsew
rlabel metal2 s 548190 0 548246 480 4 la_data_in[118]
port 135 nsew
rlabel metal2 s 551686 0 551742 480 4 la_data_in[119]
port 136 nsew
rlabel metal2 s 166390 0 166446 480 4 la_data_in[11]
port 137 nsew
rlabel metal2 s 555274 0 555330 480 4 la_data_in[120]
port 138 nsew
rlabel metal2 s 558862 0 558918 480 4 la_data_in[121]
port 139 nsew
rlabel metal2 s 562450 0 562506 480 4 la_data_in[122]
port 140 nsew
rlabel metal2 s 566038 0 566094 480 4 la_data_in[123]
port 141 nsew
rlabel metal2 s 569534 0 569590 480 4 la_data_in[124]
port 142 nsew
rlabel metal2 s 573122 0 573178 480 4 la_data_in[125]
port 143 nsew
rlabel metal2 s 576710 0 576766 480 4 la_data_in[126]
port 144 nsew
rlabel metal2 s 580298 0 580354 480 4 la_data_in[127]
port 145 nsew
rlabel metal2 s 169886 0 169942 480 4 la_data_in[12]
port 146 nsew
rlabel metal2 s 173474 0 173530 480 4 la_data_in[13]
port 147 nsew
rlabel metal2 s 177062 0 177118 480 4 la_data_in[14]
port 148 nsew
rlabel metal2 s 180650 0 180706 480 4 la_data_in[15]
port 149 nsew
rlabel metal2 s 184238 0 184294 480 4 la_data_in[16]
port 150 nsew
rlabel metal2 s 187734 0 187790 480 4 la_data_in[17]
port 151 nsew
rlabel metal2 s 191322 0 191378 480 4 la_data_in[18]
port 152 nsew
rlabel metal2 s 194910 0 194966 480 4 la_data_in[19]
port 153 nsew
rlabel metal2 s 130694 0 130750 480 4 la_data_in[1]
port 154 nsew
rlabel metal2 s 198498 0 198554 480 4 la_data_in[20]
port 155 nsew
rlabel metal2 s 201994 0 202050 480 4 la_data_in[21]
port 156 nsew
rlabel metal2 s 205582 0 205638 480 4 la_data_in[22]
port 157 nsew
rlabel metal2 s 209170 0 209226 480 4 la_data_in[23]
port 158 nsew
rlabel metal2 s 212758 0 212814 480 4 la_data_in[24]
port 159 nsew
rlabel metal2 s 216346 0 216402 480 4 la_data_in[25]
port 160 nsew
rlabel metal2 s 219842 0 219898 480 4 la_data_in[26]
port 161 nsew
rlabel metal2 s 223430 0 223486 480 4 la_data_in[27]
port 162 nsew
rlabel metal2 s 227018 0 227074 480 4 la_data_in[28]
port 163 nsew
rlabel metal2 s 230606 0 230662 480 4 la_data_in[29]
port 164 nsew
rlabel metal2 s 134282 0 134338 480 4 la_data_in[2]
port 165 nsew
rlabel metal2 s 234194 0 234250 480 4 la_data_in[30]
port 166 nsew
rlabel metal2 s 237690 0 237746 480 4 la_data_in[31]
port 167 nsew
rlabel metal2 s 241278 0 241334 480 4 la_data_in[32]
port 168 nsew
rlabel metal2 s 244866 0 244922 480 4 la_data_in[33]
port 169 nsew
rlabel metal2 s 248454 0 248510 480 4 la_data_in[34]
port 170 nsew
rlabel metal2 s 251950 0 252006 480 4 la_data_in[35]
port 171 nsew
rlabel metal2 s 255538 0 255594 480 4 la_data_in[36]
port 172 nsew
rlabel metal2 s 259126 0 259182 480 4 la_data_in[37]
port 173 nsew
rlabel metal2 s 262714 0 262770 480 4 la_data_in[38]
port 174 nsew
rlabel metal2 s 266302 0 266358 480 4 la_data_in[39]
port 175 nsew
rlabel metal2 s 137778 0 137834 480 4 la_data_in[3]
port 176 nsew
rlabel metal2 s 269798 0 269854 480 4 la_data_in[40]
port 177 nsew
rlabel metal2 s 273386 0 273442 480 4 la_data_in[41]
port 178 nsew
rlabel metal2 s 276974 0 277030 480 4 la_data_in[42]
port 179 nsew
rlabel metal2 s 280562 0 280618 480 4 la_data_in[43]
port 180 nsew
rlabel metal2 s 284150 0 284206 480 4 la_data_in[44]
port 181 nsew
rlabel metal2 s 287646 0 287702 480 4 la_data_in[45]
port 182 nsew
rlabel metal2 s 291234 0 291290 480 4 la_data_in[46]
port 183 nsew
rlabel metal2 s 294822 0 294878 480 4 la_data_in[47]
port 184 nsew
rlabel metal2 s 298410 0 298466 480 4 la_data_in[48]
port 185 nsew
rlabel metal2 s 301906 0 301962 480 4 la_data_in[49]
port 186 nsew
rlabel metal2 s 141366 0 141422 480 4 la_data_in[4]
port 187 nsew
rlabel metal2 s 305494 0 305550 480 4 la_data_in[50]
port 188 nsew
rlabel metal2 s 309082 0 309138 480 4 la_data_in[51]
port 189 nsew
rlabel metal2 s 312670 0 312726 480 4 la_data_in[52]
port 190 nsew
rlabel metal2 s 316258 0 316314 480 4 la_data_in[53]
port 191 nsew
rlabel metal2 s 319754 0 319810 480 4 la_data_in[54]
port 192 nsew
rlabel metal2 s 323342 0 323398 480 4 la_data_in[55]
port 193 nsew
rlabel metal2 s 326930 0 326986 480 4 la_data_in[56]
port 194 nsew
rlabel metal2 s 330518 0 330574 480 4 la_data_in[57]
port 195 nsew
rlabel metal2 s 334106 0 334162 480 4 la_data_in[58]
port 196 nsew
rlabel metal2 s 337602 0 337658 480 4 la_data_in[59]
port 197 nsew
rlabel metal2 s 144954 0 145010 480 4 la_data_in[5]
port 198 nsew
rlabel metal2 s 341190 0 341246 480 4 la_data_in[60]
port 199 nsew
rlabel metal2 s 344778 0 344834 480 4 la_data_in[61]
port 200 nsew
rlabel metal2 s 348366 0 348422 480 4 la_data_in[62]
port 201 nsew
rlabel metal2 s 351862 0 351918 480 4 la_data_in[63]
port 202 nsew
rlabel metal2 s 355450 0 355506 480 4 la_data_in[64]
port 203 nsew
rlabel metal2 s 359038 0 359094 480 4 la_data_in[65]
port 204 nsew
rlabel metal2 s 362626 0 362682 480 4 la_data_in[66]
port 205 nsew
rlabel metal2 s 366214 0 366270 480 4 la_data_in[67]
port 206 nsew
rlabel metal2 s 369710 0 369766 480 4 la_data_in[68]
port 207 nsew
rlabel metal2 s 373298 0 373354 480 4 la_data_in[69]
port 208 nsew
rlabel metal2 s 148542 0 148598 480 4 la_data_in[6]
port 209 nsew
rlabel metal2 s 376886 0 376942 480 4 la_data_in[70]
port 210 nsew
rlabel metal2 s 380474 0 380530 480 4 la_data_in[71]
port 211 nsew
rlabel metal2 s 384062 0 384118 480 4 la_data_in[72]
port 212 nsew
rlabel metal2 s 387558 0 387614 480 4 la_data_in[73]
port 213 nsew
rlabel metal2 s 391146 0 391202 480 4 la_data_in[74]
port 214 nsew
rlabel metal2 s 394734 0 394790 480 4 la_data_in[75]
port 215 nsew
rlabel metal2 s 398322 0 398378 480 4 la_data_in[76]
port 216 nsew
rlabel metal2 s 401818 0 401874 480 4 la_data_in[77]
port 217 nsew
rlabel metal2 s 405406 0 405462 480 4 la_data_in[78]
port 218 nsew
rlabel metal2 s 408994 0 409050 480 4 la_data_in[79]
port 219 nsew
rlabel metal2 s 152038 0 152094 480 4 la_data_in[7]
port 220 nsew
rlabel metal2 s 412582 0 412638 480 4 la_data_in[80]
port 221 nsew
rlabel metal2 s 416170 0 416226 480 4 la_data_in[81]
port 222 nsew
rlabel metal2 s 419666 0 419722 480 4 la_data_in[82]
port 223 nsew
rlabel metal2 s 423254 0 423310 480 4 la_data_in[83]
port 224 nsew
rlabel metal2 s 426842 0 426898 480 4 la_data_in[84]
port 225 nsew
rlabel metal2 s 430430 0 430486 480 4 la_data_in[85]
port 226 nsew
rlabel metal2 s 434018 0 434074 480 4 la_data_in[86]
port 227 nsew
rlabel metal2 s 437514 0 437570 480 4 la_data_in[87]
port 228 nsew
rlabel metal2 s 441102 0 441158 480 4 la_data_in[88]
port 229 nsew
rlabel metal2 s 444690 0 444746 480 4 la_data_in[89]
port 230 nsew
rlabel metal2 s 155626 0 155682 480 4 la_data_in[8]
port 231 nsew
rlabel metal2 s 448278 0 448334 480 4 la_data_in[90]
port 232 nsew
rlabel metal2 s 451774 0 451830 480 4 la_data_in[91]
port 233 nsew
rlabel metal2 s 455362 0 455418 480 4 la_data_in[92]
port 234 nsew
rlabel metal2 s 458950 0 459006 480 4 la_data_in[93]
port 235 nsew
rlabel metal2 s 462538 0 462594 480 4 la_data_in[94]
port 236 nsew
rlabel metal2 s 466126 0 466182 480 4 la_data_in[95]
port 237 nsew
rlabel metal2 s 469622 0 469678 480 4 la_data_in[96]
port 238 nsew
rlabel metal2 s 473210 0 473266 480 4 la_data_in[97]
port 239 nsew
rlabel metal2 s 476798 0 476854 480 4 la_data_in[98]
port 240 nsew
rlabel metal2 s 480386 0 480442 480 4 la_data_in[99]
port 241 nsew
rlabel metal2 s 159214 0 159270 480 4 la_data_in[9]
port 242 nsew
rlabel metal2 s 128302 0 128358 480 4 la_data_out[0]
port 243 nsew
rlabel metal2 s 485078 0 485134 480 4 la_data_out[100]
port 244 nsew
rlabel metal2 s 488666 0 488722 480 4 la_data_out[101]
port 245 nsew
rlabel metal2 s 492254 0 492310 480 4 la_data_out[102]
port 246 nsew
rlabel metal2 s 495842 0 495898 480 4 la_data_out[103]
port 247 nsew
rlabel metal2 s 499430 0 499486 480 4 la_data_out[104]
port 248 nsew
rlabel metal2 s 502926 0 502982 480 4 la_data_out[105]
port 249 nsew
rlabel metal2 s 506514 0 506570 480 4 la_data_out[106]
port 250 nsew
rlabel metal2 s 510102 0 510158 480 4 la_data_out[107]
port 251 nsew
rlabel metal2 s 513690 0 513746 480 4 la_data_out[108]
port 252 nsew
rlabel metal2 s 517278 0 517334 480 4 la_data_out[109]
port 253 nsew
rlabel metal2 s 163998 0 164054 480 4 la_data_out[10]
port 254 nsew
rlabel metal2 s 520774 0 520830 480 4 la_data_out[110]
port 255 nsew
rlabel metal2 s 524362 0 524418 480 4 la_data_out[111]
port 256 nsew
rlabel metal2 s 527950 0 528006 480 4 la_data_out[112]
port 257 nsew
rlabel metal2 s 531538 0 531594 480 4 la_data_out[113]
port 258 nsew
rlabel metal2 s 535034 0 535090 480 4 la_data_out[114]
port 259 nsew
rlabel metal2 s 538622 0 538678 480 4 la_data_out[115]
port 260 nsew
rlabel metal2 s 542210 0 542266 480 4 la_data_out[116]
port 261 nsew
rlabel metal2 s 545798 0 545854 480 4 la_data_out[117]
port 262 nsew
rlabel metal2 s 549386 0 549442 480 4 la_data_out[118]
port 263 nsew
rlabel metal2 s 552882 0 552938 480 4 la_data_out[119]
port 264 nsew
rlabel metal2 s 167586 0 167642 480 4 la_data_out[11]
port 265 nsew
rlabel metal2 s 556470 0 556526 480 4 la_data_out[120]
port 266 nsew
rlabel metal2 s 560058 0 560114 480 4 la_data_out[121]
port 267 nsew
rlabel metal2 s 563646 0 563702 480 4 la_data_out[122]
port 268 nsew
rlabel metal2 s 567234 0 567290 480 4 la_data_out[123]
port 269 nsew
rlabel metal2 s 570730 0 570786 480 4 la_data_out[124]
port 270 nsew
rlabel metal2 s 574318 0 574374 480 4 la_data_out[125]
port 271 nsew
rlabel metal2 s 577906 0 577962 480 4 la_data_out[126]
port 272 nsew
rlabel metal2 s 581494 0 581550 480 4 la_data_out[127]
port 273 nsew
rlabel metal2 s 171082 0 171138 480 4 la_data_out[12]
port 274 nsew
rlabel metal2 s 174670 0 174726 480 4 la_data_out[13]
port 275 nsew
rlabel metal2 s 178258 0 178314 480 4 la_data_out[14]
port 276 nsew
rlabel metal2 s 181846 0 181902 480 4 la_data_out[15]
port 277 nsew
rlabel metal2 s 185342 0 185398 480 4 la_data_out[16]
port 278 nsew
rlabel metal2 s 188930 0 188986 480 4 la_data_out[17]
port 279 nsew
rlabel metal2 s 192518 0 192574 480 4 la_data_out[18]
port 280 nsew
rlabel metal2 s 196106 0 196162 480 4 la_data_out[19]
port 281 nsew
rlabel metal2 s 131890 0 131946 480 4 la_data_out[1]
port 282 nsew
rlabel metal2 s 199694 0 199750 480 4 la_data_out[20]
port 283 nsew
rlabel metal2 s 203190 0 203246 480 4 la_data_out[21]
port 284 nsew
rlabel metal2 s 206778 0 206834 480 4 la_data_out[22]
port 285 nsew
rlabel metal2 s 210366 0 210422 480 4 la_data_out[23]
port 286 nsew
rlabel metal2 s 213954 0 214010 480 4 la_data_out[24]
port 287 nsew
rlabel metal2 s 217542 0 217598 480 4 la_data_out[25]
port 288 nsew
rlabel metal2 s 221038 0 221094 480 4 la_data_out[26]
port 289 nsew
rlabel metal2 s 224626 0 224682 480 4 la_data_out[27]
port 290 nsew
rlabel metal2 s 228214 0 228270 480 4 la_data_out[28]
port 291 nsew
rlabel metal2 s 231802 0 231858 480 4 la_data_out[29]
port 292 nsew
rlabel metal2 s 135386 0 135442 480 4 la_data_out[2]
port 293 nsew
rlabel metal2 s 235298 0 235354 480 4 la_data_out[30]
port 294 nsew
rlabel metal2 s 238886 0 238942 480 4 la_data_out[31]
port 295 nsew
rlabel metal2 s 242474 0 242530 480 4 la_data_out[32]
port 296 nsew
rlabel metal2 s 246062 0 246118 480 4 la_data_out[33]
port 297 nsew
rlabel metal2 s 249650 0 249706 480 4 la_data_out[34]
port 298 nsew
rlabel metal2 s 253146 0 253202 480 4 la_data_out[35]
port 299 nsew
rlabel metal2 s 256734 0 256790 480 4 la_data_out[36]
port 300 nsew
rlabel metal2 s 260322 0 260378 480 4 la_data_out[37]
port 301 nsew
rlabel metal2 s 263910 0 263966 480 4 la_data_out[38]
port 302 nsew
rlabel metal2 s 267498 0 267554 480 4 la_data_out[39]
port 303 nsew
rlabel metal2 s 138974 0 139030 480 4 la_data_out[3]
port 304 nsew
rlabel metal2 s 270994 0 271050 480 4 la_data_out[40]
port 305 nsew
rlabel metal2 s 274582 0 274638 480 4 la_data_out[41]
port 306 nsew
rlabel metal2 s 278170 0 278226 480 4 la_data_out[42]
port 307 nsew
rlabel metal2 s 281758 0 281814 480 4 la_data_out[43]
port 308 nsew
rlabel metal2 s 285254 0 285310 480 4 la_data_out[44]
port 309 nsew
rlabel metal2 s 288842 0 288898 480 4 la_data_out[45]
port 310 nsew
rlabel metal2 s 292430 0 292486 480 4 la_data_out[46]
port 311 nsew
rlabel metal2 s 296018 0 296074 480 4 la_data_out[47]
port 312 nsew
rlabel metal2 s 299606 0 299662 480 4 la_data_out[48]
port 313 nsew
rlabel metal2 s 303102 0 303158 480 4 la_data_out[49]
port 314 nsew
rlabel metal2 s 142562 0 142618 480 4 la_data_out[4]
port 315 nsew
rlabel metal2 s 306690 0 306746 480 4 la_data_out[50]
port 316 nsew
rlabel metal2 s 310278 0 310334 480 4 la_data_out[51]
port 317 nsew
rlabel metal2 s 313866 0 313922 480 4 la_data_out[52]
port 318 nsew
rlabel metal2 s 317454 0 317510 480 4 la_data_out[53]
port 319 nsew
rlabel metal2 s 320950 0 321006 480 4 la_data_out[54]
port 320 nsew
rlabel metal2 s 324538 0 324594 480 4 la_data_out[55]
port 321 nsew
rlabel metal2 s 328126 0 328182 480 4 la_data_out[56]
port 322 nsew
rlabel metal2 s 331714 0 331770 480 4 la_data_out[57]
port 323 nsew
rlabel metal2 s 335210 0 335266 480 4 la_data_out[58]
port 324 nsew
rlabel metal2 s 338798 0 338854 480 4 la_data_out[59]
port 325 nsew
rlabel metal2 s 146150 0 146206 480 4 la_data_out[5]
port 326 nsew
rlabel metal2 s 342386 0 342442 480 4 la_data_out[60]
port 327 nsew
rlabel metal2 s 345974 0 346030 480 4 la_data_out[61]
port 328 nsew
rlabel metal2 s 349562 0 349618 480 4 la_data_out[62]
port 329 nsew
rlabel metal2 s 353058 0 353114 480 4 la_data_out[63]
port 330 nsew
rlabel metal2 s 356646 0 356702 480 4 la_data_out[64]
port 331 nsew
rlabel metal2 s 360234 0 360290 480 4 la_data_out[65]
port 332 nsew
rlabel metal2 s 363822 0 363878 480 4 la_data_out[66]
port 333 nsew
rlabel metal2 s 367410 0 367466 480 4 la_data_out[67]
port 334 nsew
rlabel metal2 s 370906 0 370962 480 4 la_data_out[68]
port 335 nsew
rlabel metal2 s 374494 0 374550 480 4 la_data_out[69]
port 336 nsew
rlabel metal2 s 149738 0 149794 480 4 la_data_out[6]
port 337 nsew
rlabel metal2 s 378082 0 378138 480 4 la_data_out[70]
port 338 nsew
rlabel metal2 s 381670 0 381726 480 4 la_data_out[71]
port 339 nsew
rlabel metal2 s 385166 0 385222 480 4 la_data_out[72]
port 340 nsew
rlabel metal2 s 388754 0 388810 480 4 la_data_out[73]
port 341 nsew
rlabel metal2 s 392342 0 392398 480 4 la_data_out[74]
port 342 nsew
rlabel metal2 s 395930 0 395986 480 4 la_data_out[75]
port 343 nsew
rlabel metal2 s 399518 0 399574 480 4 la_data_out[76]
port 344 nsew
rlabel metal2 s 403014 0 403070 480 4 la_data_out[77]
port 345 nsew
rlabel metal2 s 406602 0 406658 480 4 la_data_out[78]
port 346 nsew
rlabel metal2 s 410190 0 410246 480 4 la_data_out[79]
port 347 nsew
rlabel metal2 s 153234 0 153290 480 4 la_data_out[7]
port 348 nsew
rlabel metal2 s 413778 0 413834 480 4 la_data_out[80]
port 349 nsew
rlabel metal2 s 417366 0 417422 480 4 la_data_out[81]
port 350 nsew
rlabel metal2 s 420862 0 420918 480 4 la_data_out[82]
port 351 nsew
rlabel metal2 s 424450 0 424506 480 4 la_data_out[83]
port 352 nsew
rlabel metal2 s 428038 0 428094 480 4 la_data_out[84]
port 353 nsew
rlabel metal2 s 431626 0 431682 480 4 la_data_out[85]
port 354 nsew
rlabel metal2 s 435122 0 435178 480 4 la_data_out[86]
port 355 nsew
rlabel metal2 s 438710 0 438766 480 4 la_data_out[87]
port 356 nsew
rlabel metal2 s 442298 0 442354 480 4 la_data_out[88]
port 357 nsew
rlabel metal2 s 445886 0 445942 480 4 la_data_out[89]
port 358 nsew
rlabel metal2 s 156822 0 156878 480 4 la_data_out[8]
port 359 nsew
rlabel metal2 s 449474 0 449530 480 4 la_data_out[90]
port 360 nsew
rlabel metal2 s 452970 0 453026 480 4 la_data_out[91]
port 361 nsew
rlabel metal2 s 456558 0 456614 480 4 la_data_out[92]
port 362 nsew
rlabel metal2 s 460146 0 460202 480 4 la_data_out[93]
port 363 nsew
rlabel metal2 s 463734 0 463790 480 4 la_data_out[94]
port 364 nsew
rlabel metal2 s 467322 0 467378 480 4 la_data_out[95]
port 365 nsew
rlabel metal2 s 470818 0 470874 480 4 la_data_out[96]
port 366 nsew
rlabel metal2 s 474406 0 474462 480 4 la_data_out[97]
port 367 nsew
rlabel metal2 s 477994 0 478050 480 4 la_data_out[98]
port 368 nsew
rlabel metal2 s 481582 0 481638 480 4 la_data_out[99]
port 369 nsew
rlabel metal2 s 160410 0 160466 480 4 la_data_out[9]
port 370 nsew
rlabel metal2 s 129498 0 129554 480 4 la_oen[0]
port 371 nsew
rlabel metal2 s 486274 0 486330 480 4 la_oen[100]
port 372 nsew
rlabel metal2 s 489862 0 489918 480 4 la_oen[101]
port 373 nsew
rlabel metal2 s 493450 0 493506 480 4 la_oen[102]
port 374 nsew
rlabel metal2 s 497038 0 497094 480 4 la_oen[103]
port 375 nsew
rlabel metal2 s 500626 0 500682 480 4 la_oen[104]
port 376 nsew
rlabel metal2 s 504122 0 504178 480 4 la_oen[105]
port 377 nsew
rlabel metal2 s 507710 0 507766 480 4 la_oen[106]
port 378 nsew
rlabel metal2 s 511298 0 511354 480 4 la_oen[107]
port 379 nsew
rlabel metal2 s 514886 0 514942 480 4 la_oen[108]
port 380 nsew
rlabel metal2 s 518382 0 518438 480 4 la_oen[109]
port 381 nsew
rlabel metal2 s 165194 0 165250 480 4 la_oen[10]
port 382 nsew
rlabel metal2 s 521970 0 522026 480 4 la_oen[110]
port 383 nsew
rlabel metal2 s 525558 0 525614 480 4 la_oen[111]
port 384 nsew
rlabel metal2 s 529146 0 529202 480 4 la_oen[112]
port 385 nsew
rlabel metal2 s 532734 0 532790 480 4 la_oen[113]
port 386 nsew
rlabel metal2 s 536230 0 536286 480 4 la_oen[114]
port 387 nsew
rlabel metal2 s 539818 0 539874 480 4 la_oen[115]
port 388 nsew
rlabel metal2 s 543406 0 543462 480 4 la_oen[116]
port 389 nsew
rlabel metal2 s 546994 0 547050 480 4 la_oen[117]
port 390 nsew
rlabel metal2 s 550582 0 550638 480 4 la_oen[118]
port 391 nsew
rlabel metal2 s 554078 0 554134 480 4 la_oen[119]
port 392 nsew
rlabel metal2 s 168690 0 168746 480 4 la_oen[11]
port 393 nsew
rlabel metal2 s 557666 0 557722 480 4 la_oen[120]
port 394 nsew
rlabel metal2 s 561254 0 561310 480 4 la_oen[121]
port 395 nsew
rlabel metal2 s 564842 0 564898 480 4 la_oen[122]
port 396 nsew
rlabel metal2 s 568338 0 568394 480 4 la_oen[123]
port 397 nsew
rlabel metal2 s 571926 0 571982 480 4 la_oen[124]
port 398 nsew
rlabel metal2 s 575514 0 575570 480 4 la_oen[125]
port 399 nsew
rlabel metal2 s 579102 0 579158 480 4 la_oen[126]
port 400 nsew
rlabel metal2 s 582690 0 582746 480 4 la_oen[127]
port 401 nsew
rlabel metal2 s 172278 0 172334 480 4 la_oen[12]
port 402 nsew
rlabel metal2 s 175866 0 175922 480 4 la_oen[13]
port 403 nsew
rlabel metal2 s 179454 0 179510 480 4 la_oen[14]
port 404 nsew
rlabel metal2 s 183042 0 183098 480 4 la_oen[15]
port 405 nsew
rlabel metal2 s 186538 0 186594 480 4 la_oen[16]
port 406 nsew
rlabel metal2 s 190126 0 190182 480 4 la_oen[17]
port 407 nsew
rlabel metal2 s 193714 0 193770 480 4 la_oen[18]
port 408 nsew
rlabel metal2 s 197302 0 197358 480 4 la_oen[19]
port 409 nsew
rlabel metal2 s 133086 0 133142 480 4 la_oen[1]
port 410 nsew
rlabel metal2 s 200890 0 200946 480 4 la_oen[20]
port 411 nsew
rlabel metal2 s 204386 0 204442 480 4 la_oen[21]
port 412 nsew
rlabel metal2 s 207974 0 208030 480 4 la_oen[22]
port 413 nsew
rlabel metal2 s 211562 0 211618 480 4 la_oen[23]
port 414 nsew
rlabel metal2 s 215150 0 215206 480 4 la_oen[24]
port 415 nsew
rlabel metal2 s 218646 0 218702 480 4 la_oen[25]
port 416 nsew
rlabel metal2 s 222234 0 222290 480 4 la_oen[26]
port 417 nsew
rlabel metal2 s 225822 0 225878 480 4 la_oen[27]
port 418 nsew
rlabel metal2 s 229410 0 229466 480 4 la_oen[28]
port 419 nsew
rlabel metal2 s 232998 0 233054 480 4 la_oen[29]
port 420 nsew
rlabel metal2 s 136582 0 136638 480 4 la_oen[2]
port 421 nsew
rlabel metal2 s 236494 0 236550 480 4 la_oen[30]
port 422 nsew
rlabel metal2 s 240082 0 240138 480 4 la_oen[31]
port 423 nsew
rlabel metal2 s 243670 0 243726 480 4 la_oen[32]
port 424 nsew
rlabel metal2 s 247258 0 247314 480 4 la_oen[33]
port 425 nsew
rlabel metal2 s 250846 0 250902 480 4 la_oen[34]
port 426 nsew
rlabel metal2 s 254342 0 254398 480 4 la_oen[35]
port 427 nsew
rlabel metal2 s 257930 0 257986 480 4 la_oen[36]
port 428 nsew
rlabel metal2 s 261518 0 261574 480 4 la_oen[37]
port 429 nsew
rlabel metal2 s 265106 0 265162 480 4 la_oen[38]
port 430 nsew
rlabel metal2 s 268602 0 268658 480 4 la_oen[39]
port 431 nsew
rlabel metal2 s 140170 0 140226 480 4 la_oen[3]
port 432 nsew
rlabel metal2 s 272190 0 272246 480 4 la_oen[40]
port 433 nsew
rlabel metal2 s 275778 0 275834 480 4 la_oen[41]
port 434 nsew
rlabel metal2 s 279366 0 279422 480 4 la_oen[42]
port 435 nsew
rlabel metal2 s 282954 0 283010 480 4 la_oen[43]
port 436 nsew
rlabel metal2 s 286450 0 286506 480 4 la_oen[44]
port 437 nsew
rlabel metal2 s 290038 0 290094 480 4 la_oen[45]
port 438 nsew
rlabel metal2 s 293626 0 293682 480 4 la_oen[46]
port 439 nsew
rlabel metal2 s 297214 0 297270 480 4 la_oen[47]
port 440 nsew
rlabel metal2 s 300802 0 300858 480 4 la_oen[48]
port 441 nsew
rlabel metal2 s 304298 0 304354 480 4 la_oen[49]
port 442 nsew
rlabel metal2 s 143758 0 143814 480 4 la_oen[4]
port 443 nsew
rlabel metal2 s 307886 0 307942 480 4 la_oen[50]
port 444 nsew
rlabel metal2 s 311474 0 311530 480 4 la_oen[51]
port 445 nsew
rlabel metal2 s 315062 0 315118 480 4 la_oen[52]
port 446 nsew
rlabel metal2 s 318558 0 318614 480 4 la_oen[53]
port 447 nsew
rlabel metal2 s 322146 0 322202 480 4 la_oen[54]
port 448 nsew
rlabel metal2 s 325734 0 325790 480 4 la_oen[55]
port 449 nsew
rlabel metal2 s 329322 0 329378 480 4 la_oen[56]
port 450 nsew
rlabel metal2 s 332910 0 332966 480 4 la_oen[57]
port 451 nsew
rlabel metal2 s 336406 0 336462 480 4 la_oen[58]
port 452 nsew
rlabel metal2 s 339994 0 340050 480 4 la_oen[59]
port 453 nsew
rlabel metal2 s 147346 0 147402 480 4 la_oen[5]
port 454 nsew
rlabel metal2 s 343582 0 343638 480 4 la_oen[60]
port 455 nsew
rlabel metal2 s 347170 0 347226 480 4 la_oen[61]
port 456 nsew
rlabel metal2 s 350758 0 350814 480 4 la_oen[62]
port 457 nsew
rlabel metal2 s 354254 0 354310 480 4 la_oen[63]
port 458 nsew
rlabel metal2 s 357842 0 357898 480 4 la_oen[64]
port 459 nsew
rlabel metal2 s 361430 0 361486 480 4 la_oen[65]
port 460 nsew
rlabel metal2 s 365018 0 365074 480 4 la_oen[66]
port 461 nsew
rlabel metal2 s 368514 0 368570 480 4 la_oen[67]
port 462 nsew
rlabel metal2 s 372102 0 372158 480 4 la_oen[68]
port 463 nsew
rlabel metal2 s 375690 0 375746 480 4 la_oen[69]
port 464 nsew
rlabel metal2 s 150934 0 150990 480 4 la_oen[6]
port 465 nsew
rlabel metal2 s 379278 0 379334 480 4 la_oen[70]
port 466 nsew
rlabel metal2 s 382866 0 382922 480 4 la_oen[71]
port 467 nsew
rlabel metal2 s 386362 0 386418 480 4 la_oen[72]
port 468 nsew
rlabel metal2 s 389950 0 390006 480 4 la_oen[73]
port 469 nsew
rlabel metal2 s 393538 0 393594 480 4 la_oen[74]
port 470 nsew
rlabel metal2 s 397126 0 397182 480 4 la_oen[75]
port 471 nsew
rlabel metal2 s 400714 0 400770 480 4 la_oen[76]
port 472 nsew
rlabel metal2 s 404210 0 404266 480 4 la_oen[77]
port 473 nsew
rlabel metal2 s 407798 0 407854 480 4 la_oen[78]
port 474 nsew
rlabel metal2 s 411386 0 411442 480 4 la_oen[79]
port 475 nsew
rlabel metal2 s 154430 0 154486 480 4 la_oen[7]
port 476 nsew
rlabel metal2 s 414974 0 415030 480 4 la_oen[80]
port 477 nsew
rlabel metal2 s 418470 0 418526 480 4 la_oen[81]
port 478 nsew
rlabel metal2 s 422058 0 422114 480 4 la_oen[82]
port 479 nsew
rlabel metal2 s 425646 0 425702 480 4 la_oen[83]
port 480 nsew
rlabel metal2 s 429234 0 429290 480 4 la_oen[84]
port 481 nsew
rlabel metal2 s 432822 0 432878 480 4 la_oen[85]
port 482 nsew
rlabel metal2 s 436318 0 436374 480 4 la_oen[86]
port 483 nsew
rlabel metal2 s 439906 0 439962 480 4 la_oen[87]
port 484 nsew
rlabel metal2 s 443494 0 443550 480 4 la_oen[88]
port 485 nsew
rlabel metal2 s 447082 0 447138 480 4 la_oen[89]
port 486 nsew
rlabel metal2 s 158018 0 158074 480 4 la_oen[8]
port 487 nsew
rlabel metal2 s 450670 0 450726 480 4 la_oen[90]
port 488 nsew
rlabel metal2 s 454166 0 454222 480 4 la_oen[91]
port 489 nsew
rlabel metal2 s 457754 0 457810 480 4 la_oen[92]
port 490 nsew
rlabel metal2 s 461342 0 461398 480 4 la_oen[93]
port 491 nsew
rlabel metal2 s 464930 0 464986 480 4 la_oen[94]
port 492 nsew
rlabel metal2 s 468426 0 468482 480 4 la_oen[95]
port 493 nsew
rlabel metal2 s 472014 0 472070 480 4 la_oen[96]
port 494 nsew
rlabel metal2 s 475602 0 475658 480 4 la_oen[97]
port 495 nsew
rlabel metal2 s 479190 0 479246 480 4 la_oen[98]
port 496 nsew
rlabel metal2 s 482778 0 482834 480 4 la_oen[99]
port 497 nsew
rlabel metal2 s 161606 0 161662 480 4 la_oen[9]
port 498 nsew
rlabel metal2 s 583886 0 583942 480 4 user_clock2
port 499 nsew
rlabel metal2 s 1066 0 1122 480 4 wb_clk_i
port 500 nsew
rlabel metal2 s 2170 0 2226 480 4 wb_rst_i
port 501 nsew
rlabel metal2 s 3366 0 3422 480 4 wbs_ack_o
port 502 nsew
rlabel metal2 s 8150 0 8206 480 4 wbs_adr_i[0]
port 503 nsew
rlabel metal2 s 48630 0 48686 480 4 wbs_adr_i[10]
port 504 nsew
rlabel metal2 s 52126 0 52182 480 4 wbs_adr_i[11]
port 505 nsew
rlabel metal2 s 55714 0 55770 480 4 wbs_adr_i[12]
port 506 nsew
rlabel metal2 s 59302 0 59358 480 4 wbs_adr_i[13]
port 507 nsew
rlabel metal2 s 62890 0 62946 480 4 wbs_adr_i[14]
port 508 nsew
rlabel metal2 s 66478 0 66534 480 4 wbs_adr_i[15]
port 509 nsew
rlabel metal2 s 69974 0 70030 480 4 wbs_adr_i[16]
port 510 nsew
rlabel metal2 s 73562 0 73618 480 4 wbs_adr_i[17]
port 511 nsew
rlabel metal2 s 77150 0 77206 480 4 wbs_adr_i[18]
port 512 nsew
rlabel metal2 s 80738 0 80794 480 4 wbs_adr_i[19]
port 513 nsew
rlabel metal2 s 12934 0 12990 480 4 wbs_adr_i[1]
port 514 nsew
rlabel metal2 s 84326 0 84382 480 4 wbs_adr_i[20]
port 515 nsew
rlabel metal2 s 87822 0 87878 480 4 wbs_adr_i[21]
port 516 nsew
rlabel metal2 s 91410 0 91466 480 4 wbs_adr_i[22]
port 517 nsew
rlabel metal2 s 94998 0 95054 480 4 wbs_adr_i[23]
port 518 nsew
rlabel metal2 s 98586 0 98642 480 4 wbs_adr_i[24]
port 519 nsew
rlabel metal2 s 102082 0 102138 480 4 wbs_adr_i[25]
port 520 nsew
rlabel metal2 s 105670 0 105726 480 4 wbs_adr_i[26]
port 521 nsew
rlabel metal2 s 109258 0 109314 480 4 wbs_adr_i[27]
port 522 nsew
rlabel metal2 s 112846 0 112902 480 4 wbs_adr_i[28]
port 523 nsew
rlabel metal2 s 116434 0 116490 480 4 wbs_adr_i[29]
port 524 nsew
rlabel metal2 s 17718 0 17774 480 4 wbs_adr_i[2]
port 525 nsew
rlabel metal2 s 119930 0 119986 480 4 wbs_adr_i[30]
port 526 nsew
rlabel metal2 s 123518 0 123574 480 4 wbs_adr_i[31]
port 527 nsew
rlabel metal2 s 22410 0 22466 480 4 wbs_adr_i[3]
port 528 nsew
rlabel metal2 s 27194 0 27250 480 4 wbs_adr_i[4]
port 529 nsew
rlabel metal2 s 30782 0 30838 480 4 wbs_adr_i[5]
port 530 nsew
rlabel metal2 s 34370 0 34426 480 4 wbs_adr_i[6]
port 531 nsew
rlabel metal2 s 37866 0 37922 480 4 wbs_adr_i[7]
port 532 nsew
rlabel metal2 s 41454 0 41510 480 4 wbs_adr_i[8]
port 533 nsew
rlabel metal2 s 45042 0 45098 480 4 wbs_adr_i[9]
port 534 nsew
rlabel metal2 s 4562 0 4618 480 4 wbs_cyc_i
port 535 nsew
rlabel metal2 s 9346 0 9402 480 4 wbs_dat_i[0]
port 536 nsew
rlabel metal2 s 49826 0 49882 480 4 wbs_dat_i[10]
port 537 nsew
rlabel metal2 s 53322 0 53378 480 4 wbs_dat_i[11]
port 538 nsew
rlabel metal2 s 56910 0 56966 480 4 wbs_dat_i[12]
port 539 nsew
rlabel metal2 s 60498 0 60554 480 4 wbs_dat_i[13]
port 540 nsew
rlabel metal2 s 64086 0 64142 480 4 wbs_dat_i[14]
port 541 nsew
rlabel metal2 s 67674 0 67730 480 4 wbs_dat_i[15]
port 542 nsew
rlabel metal2 s 71170 0 71226 480 4 wbs_dat_i[16]
port 543 nsew
rlabel metal2 s 74758 0 74814 480 4 wbs_dat_i[17]
port 544 nsew
rlabel metal2 s 78346 0 78402 480 4 wbs_dat_i[18]
port 545 nsew
rlabel metal2 s 81934 0 81990 480 4 wbs_dat_i[19]
port 546 nsew
rlabel metal2 s 14130 0 14186 480 4 wbs_dat_i[1]
port 547 nsew
rlabel metal2 s 85430 0 85486 480 4 wbs_dat_i[20]
port 548 nsew
rlabel metal2 s 89018 0 89074 480 4 wbs_dat_i[21]
port 549 nsew
rlabel metal2 s 92606 0 92662 480 4 wbs_dat_i[22]
port 550 nsew
rlabel metal2 s 96194 0 96250 480 4 wbs_dat_i[23]
port 551 nsew
rlabel metal2 s 99782 0 99838 480 4 wbs_dat_i[24]
port 552 nsew
rlabel metal2 s 103278 0 103334 480 4 wbs_dat_i[25]
port 553 nsew
rlabel metal2 s 106866 0 106922 480 4 wbs_dat_i[26]
port 554 nsew
rlabel metal2 s 110454 0 110510 480 4 wbs_dat_i[27]
port 555 nsew
rlabel metal2 s 114042 0 114098 480 4 wbs_dat_i[28]
port 556 nsew
rlabel metal2 s 117630 0 117686 480 4 wbs_dat_i[29]
port 557 nsew
rlabel metal2 s 18822 0 18878 480 4 wbs_dat_i[2]
port 558 nsew
rlabel metal2 s 121126 0 121182 480 4 wbs_dat_i[30]
port 559 nsew
rlabel metal2 s 124714 0 124770 480 4 wbs_dat_i[31]
port 560 nsew
rlabel metal2 s 23606 0 23662 480 4 wbs_dat_i[3]
port 561 nsew
rlabel metal2 s 28390 0 28446 480 4 wbs_dat_i[4]
port 562 nsew
rlabel metal2 s 31978 0 32034 480 4 wbs_dat_i[5]
port 563 nsew
rlabel metal2 s 35474 0 35530 480 4 wbs_dat_i[6]
port 564 nsew
rlabel metal2 s 39062 0 39118 480 4 wbs_dat_i[7]
port 565 nsew
rlabel metal2 s 42650 0 42706 480 4 wbs_dat_i[8]
port 566 nsew
rlabel metal2 s 46238 0 46294 480 4 wbs_dat_i[9]
port 567 nsew
rlabel metal2 s 10542 0 10598 480 4 wbs_dat_o[0]
port 568 nsew
rlabel metal2 s 51022 0 51078 480 4 wbs_dat_o[10]
port 569 nsew
rlabel metal2 s 54518 0 54574 480 4 wbs_dat_o[11]
port 570 nsew
rlabel metal2 s 58106 0 58162 480 4 wbs_dat_o[12]
port 571 nsew
rlabel metal2 s 61694 0 61750 480 4 wbs_dat_o[13]
port 572 nsew
rlabel metal2 s 65282 0 65338 480 4 wbs_dat_o[14]
port 573 nsew
rlabel metal2 s 68778 0 68834 480 4 wbs_dat_o[15]
port 574 nsew
rlabel metal2 s 72366 0 72422 480 4 wbs_dat_o[16]
port 575 nsew
rlabel metal2 s 75954 0 76010 480 4 wbs_dat_o[17]
port 576 nsew
rlabel metal2 s 79542 0 79598 480 4 wbs_dat_o[18]
port 577 nsew
rlabel metal2 s 83130 0 83186 480 4 wbs_dat_o[19]
port 578 nsew
rlabel metal2 s 15326 0 15382 480 4 wbs_dat_o[1]
port 579 nsew
rlabel metal2 s 86626 0 86682 480 4 wbs_dat_o[20]
port 580 nsew
rlabel metal2 s 90214 0 90270 480 4 wbs_dat_o[21]
port 581 nsew
rlabel metal2 s 93802 0 93858 480 4 wbs_dat_o[22]
port 582 nsew
rlabel metal2 s 97390 0 97446 480 4 wbs_dat_o[23]
port 583 nsew
rlabel metal2 s 100978 0 101034 480 4 wbs_dat_o[24]
port 584 nsew
rlabel metal2 s 104474 0 104530 480 4 wbs_dat_o[25]
port 585 nsew
rlabel metal2 s 108062 0 108118 480 4 wbs_dat_o[26]
port 586 nsew
rlabel metal2 s 111650 0 111706 480 4 wbs_dat_o[27]
port 587 nsew
rlabel metal2 s 115238 0 115294 480 4 wbs_dat_o[28]
port 588 nsew
rlabel metal2 s 118734 0 118790 480 4 wbs_dat_o[29]
port 589 nsew
rlabel metal2 s 20018 0 20074 480 4 wbs_dat_o[2]
port 590 nsew
rlabel metal2 s 122322 0 122378 480 4 wbs_dat_o[30]
port 591 nsew
rlabel metal2 s 125910 0 125966 480 4 wbs_dat_o[31]
port 592 nsew
rlabel metal2 s 24802 0 24858 480 4 wbs_dat_o[3]
port 593 nsew
rlabel metal2 s 29586 0 29642 480 4 wbs_dat_o[4]
port 594 nsew
rlabel metal2 s 33174 0 33230 480 4 wbs_dat_o[5]
port 595 nsew
rlabel metal2 s 36670 0 36726 480 4 wbs_dat_o[6]
port 596 nsew
rlabel metal2 s 40258 0 40314 480 4 wbs_dat_o[7]
port 597 nsew
rlabel metal2 s 43846 0 43902 480 4 wbs_dat_o[8]
port 598 nsew
rlabel metal2 s 47434 0 47490 480 4 wbs_dat_o[9]
port 599 nsew
rlabel metal2 s 11738 0 11794 480 4 wbs_sel_i[0]
port 600 nsew
rlabel metal2 s 16522 0 16578 480 4 wbs_sel_i[1]
port 601 nsew
rlabel metal2 s 21214 0 21270 480 4 wbs_sel_i[2]
port 602 nsew
rlabel metal2 s 25998 0 26054 480 4 wbs_sel_i[3]
port 603 nsew
rlabel metal2 s 5758 0 5814 480 4 wbs_stb_i
port 604 nsew
rlabel metal2 s 6954 0 7010 480 4 wbs_we_i
port 605 nsew
rlabel metal5 s 800 1376 584116 1776 4 vccd1
port 606 nsew
rlabel metal5 s 0 576 584916 976 4 vssd1
port 607 nsew
<< properties >>
string FIXED_BBOX 0 0 584916 704000
<< end >>
