* NGSPICE file created from caravel.ext - technology: sky130A

* Black-box entry subcircuit for gpio_control_block abstract view
.subckt gpio_control_block mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en
+ pad_gpio_ana_pol pad_gpio_ana_sel pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover
+ pad_gpio_ib_mode_sel pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel
+ pad_gpio_vtrip_sel resetn serial_clock serial_data_in serial_data_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero vccd vssd vccd1 vssd1
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_20um abstract view
.subckt sky130_ef_io__com_bus_slice_20um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_1um abstract view
.subckt sky130_ef_io__com_bus_slice_1um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__gpiov2_pad_wrapped abstract view
.subckt sky130_ef_io__gpiov2_pad_wrapped IN_H PAD_A_NOESD_H PAD_A_ESD_0_H PAD_A_ESD_1_H
+ PAD DM[2] DM[1] DM[0] HLD_H_N IN INP_DIS IB_MODE_SEL ENABLE_H ENABLE_VDDA_H ENABLE_INP_H
+ OE_N TIE_HI_ESD TIE_LO_ESD SLOW VTRIP_SEL HLD_OVR ANALOG_EN ANALOG_SEL ENABLE_VDDIO
+ ENABLE_VSWITCH_H ANALOG_POL OUT AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_5um abstract view
.subckt sky130_ef_io__com_bus_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__com_bus_slice_10um abstract view
.subckt sky130_ef_io__com_bus_slice_10um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__disconnect_vdda_slice_5um abstract view
.subckt sky130_ef_io__disconnect_vdda_slice_5um AMUXBUS_A AMUXBUS_B VSWITCH VDDIO_Q
+ VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__corner_pad abstract view
.subckt sky130_ef_io__corner_pad AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH VDDIO_Q VCCHIB
+ VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vddio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vddio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssio_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssio_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSIO_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um abstract view
.subckt sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um AMUXBUS_A AMUXBUS_B
+ VSSA VDDA VDDIO_Q VDDIO VCCD VSSIO VSSD VSSIO_Q VSWITCH VCCHIB
.ends

* Black-box entry subcircuit for sky130_ef_io__vdda_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vdda_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VDDA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vccd_lvc_clamped2_pad abstract view
.subckt sky130_ef_io__vccd_lvc_clamped2_pad AMUXBUS_A AMUXBUS_B VCCD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssa_hvc_clamped_pad abstract view
.subckt sky130_ef_io__vssa_hvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSA_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__disconnect_vccd_slice_5um abstract view
.subckt sky130_ef_io__disconnect_vccd_slice_5um AMUXBUS_A AMUXBUS_B VSSA VDDA VSWITCH
+ VDDIO_Q VCCHIB VDDIO VSSIO VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_fd_io__top_xres4v2 abstract view
.subckt sky130_fd_io__top_xres4v2 AMUXBUS_A AMUXBUS_B DISABLE_PULLUP_H ENABLE_H ENABLE_VDDIO
+ EN_VDDIO_SIG_H FILT_IN_H INP_SEL_H PAD PAD_A_ESD_H PULLUP_H TIE_HI_ESD TIE_LO_ESD
+ TIE_WEAK_HI_H XRES_H_N VCCD VCCHIB VDDA VDDIO VDDIO_Q VSSA VSSD VSSIO VSSIO_Q VSWITCH
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped2_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped2_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

* Black-box entry subcircuit for sky130_ef_io__vssd_lvc_clamped_pad abstract view
.subckt sky130_ef_io__vssd_lvc_clamped_pad AMUXBUS_A AMUXBUS_B VSSD_PAD VSSA VDDA
+ VSWITCH VDDIO_Q VCCHIB VDDIO VCCD VSSIO VSSD VSSIO_Q
.ends

.subckt chip_io clock clock_core flash_clk flash_clk_core flash_clk_ieb_core flash_clk_oeb_core
+ flash_csb flash_csb_core flash_csb_ieb_core flash_csb_oeb_core flash_io0 flash_io0_di_core
+ flash_io0_do_core flash_io0_ieb_core flash_io0_oeb_core flash_io1 flash_io1_di_core
+ flash_io1_do_core flash_io1_ieb_core flash_io1_oeb_core gpio gpio_in_core gpio_inenb_core
+ gpio_mode0_core gpio_mode1_core gpio_out_core gpio_outenb_core mprj_analog_io[0]
+ mprj_analog_io[10] mprj_analog_io[11] mprj_analog_io[12] mprj_analog_io[13] mprj_analog_io[14]
+ mprj_analog_io[15] mprj_analog_io[16] mprj_analog_io[17] mprj_analog_io[18] mprj_analog_io[19]
+ mprj_analog_io[1] mprj_analog_io[20] mprj_analog_io[21] mprj_analog_io[22] mprj_analog_io[23]
+ mprj_analog_io[24] mprj_analog_io[25] mprj_analog_io[26] mprj_analog_io[27] mprj_analog_io[28]
+ mprj_analog_io[29] mprj_analog_io[2] mprj_analog_io[30] mprj_analog_io[3] mprj_analog_io[4]
+ mprj_analog_io[5] mprj_analog_io[6] mprj_analog_io[7] mprj_analog_io[8] mprj_analog_io[9]
+ mprj_io[0] mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15]
+ mprj_io[16] mprj_io[17] mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21]
+ mprj_io[22] mprj_io[23] mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28]
+ mprj_io[29] mprj_io[2] mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34]
+ mprj_io[35] mprj_io[36] mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6]
+ mprj_io[7] mprj_io[8] mprj_io[9] mprj_io_analog_en[0] mprj_io_analog_en[10] mprj_io_analog_en[11]
+ mprj_io_analog_en[12] mprj_io_analog_en[13] mprj_io_analog_en[14] mprj_io_analog_en[15]
+ mprj_io_analog_en[16] mprj_io_analog_en[17] mprj_io_analog_en[18] mprj_io_analog_en[19]
+ mprj_io_analog_en[1] mprj_io_analog_en[20] mprj_io_analog_en[21] mprj_io_analog_en[22]
+ mprj_io_analog_en[23] mprj_io_analog_en[24] mprj_io_analog_en[25] mprj_io_analog_en[26]
+ mprj_io_analog_en[27] mprj_io_analog_en[28] mprj_io_analog_en[29] mprj_io_analog_en[2]
+ mprj_io_analog_en[30] mprj_io_analog_en[31] mprj_io_analog_en[32] mprj_io_analog_en[33]
+ mprj_io_analog_en[34] mprj_io_analog_en[35] mprj_io_analog_en[36] mprj_io_analog_en[37]
+ mprj_io_analog_en[3] mprj_io_analog_en[4] mprj_io_analog_en[5] mprj_io_analog_en[6]
+ mprj_io_analog_en[7] mprj_io_analog_en[8] mprj_io_analog_en[9] mprj_io_analog_pol[0]
+ mprj_io_analog_pol[10] mprj_io_analog_pol[11] mprj_io_analog_pol[12] mprj_io_analog_pol[13]
+ mprj_io_analog_pol[14] mprj_io_analog_pol[15] mprj_io_analog_pol[16] mprj_io_analog_pol[17]
+ mprj_io_analog_pol[18] mprj_io_analog_pol[19] mprj_io_analog_pol[1] mprj_io_analog_pol[20]
+ mprj_io_analog_pol[21] mprj_io_analog_pol[22] mprj_io_analog_pol[23] mprj_io_analog_pol[24]
+ mprj_io_analog_pol[25] mprj_io_analog_pol[26] mprj_io_analog_pol[27] mprj_io_analog_pol[28]
+ mprj_io_analog_pol[29] mprj_io_analog_pol[2] mprj_io_analog_pol[30] mprj_io_analog_pol[31]
+ mprj_io_analog_pol[32] mprj_io_analog_pol[33] mprj_io_analog_pol[34] mprj_io_analog_pol[35]
+ mprj_io_analog_pol[36] mprj_io_analog_pol[37] mprj_io_analog_pol[3] mprj_io_analog_pol[4]
+ mprj_io_analog_pol[5] mprj_io_analog_pol[6] mprj_io_analog_pol[7] mprj_io_analog_pol[8]
+ mprj_io_analog_pol[9] mprj_io_analog_sel[0] mprj_io_analog_sel[10] mprj_io_analog_sel[11]
+ mprj_io_analog_sel[12] mprj_io_analog_sel[13] mprj_io_analog_sel[14] mprj_io_analog_sel[15]
+ mprj_io_analog_sel[16] mprj_io_analog_sel[17] mprj_io_analog_sel[18] mprj_io_analog_sel[19]
+ mprj_io_analog_sel[1] mprj_io_analog_sel[20] mprj_io_analog_sel[21] mprj_io_analog_sel[22]
+ mprj_io_analog_sel[23] mprj_io_analog_sel[24] mprj_io_analog_sel[25] mprj_io_analog_sel[26]
+ mprj_io_analog_sel[27] mprj_io_analog_sel[28] mprj_io_analog_sel[29] mprj_io_analog_sel[2]
+ mprj_io_analog_sel[30] mprj_io_analog_sel[31] mprj_io_analog_sel[32] mprj_io_analog_sel[33]
+ mprj_io_analog_sel[34] mprj_io_analog_sel[35] mprj_io_analog_sel[36] mprj_io_analog_sel[37]
+ mprj_io_analog_sel[3] mprj_io_analog_sel[4] mprj_io_analog_sel[5] mprj_io_analog_sel[6]
+ mprj_io_analog_sel[7] mprj_io_analog_sel[8] mprj_io_analog_sel[9] mprj_io_dm[0]
+ mprj_io_dm[100] mprj_io_dm[101] mprj_io_dm[102] mprj_io_dm[103] mprj_io_dm[104]
+ mprj_io_dm[105] mprj_io_dm[106] mprj_io_dm[107] mprj_io_dm[108] mprj_io_dm[109]
+ mprj_io_dm[10] mprj_io_dm[110] mprj_io_dm[111] mprj_io_dm[112] mprj_io_dm[113] mprj_io_dm[11]
+ mprj_io_dm[12] mprj_io_dm[13] mprj_io_dm[14] mprj_io_dm[15] mprj_io_dm[16] mprj_io_dm[17]
+ mprj_io_dm[18] mprj_io_dm[19] mprj_io_dm[1] mprj_io_dm[20] mprj_io_dm[21] mprj_io_dm[22]
+ mprj_io_dm[23] mprj_io_dm[24] mprj_io_dm[25] mprj_io_dm[26] mprj_io_dm[27] mprj_io_dm[28]
+ mprj_io_dm[29] mprj_io_dm[2] mprj_io_dm[30] mprj_io_dm[31] mprj_io_dm[32] mprj_io_dm[33]
+ mprj_io_dm[34] mprj_io_dm[35] mprj_io_dm[36] mprj_io_dm[37] mprj_io_dm[38] mprj_io_dm[39]
+ mprj_io_dm[3] mprj_io_dm[40] mprj_io_dm[41] mprj_io_dm[42] mprj_io_dm[43] mprj_io_dm[44]
+ mprj_io_dm[45] mprj_io_dm[46] mprj_io_dm[47] mprj_io_dm[48] mprj_io_dm[49] mprj_io_dm[4]
+ mprj_io_dm[50] mprj_io_dm[51] mprj_io_dm[52] mprj_io_dm[53] mprj_io_dm[54] mprj_io_dm[55]
+ mprj_io_dm[56] mprj_io_dm[57] mprj_io_dm[58] mprj_io_dm[59] mprj_io_dm[5] mprj_io_dm[60]
+ mprj_io_dm[61] mprj_io_dm[62] mprj_io_dm[63] mprj_io_dm[64] mprj_io_dm[65] mprj_io_dm[66]
+ mprj_io_dm[67] mprj_io_dm[68] mprj_io_dm[69] mprj_io_dm[6] mprj_io_dm[70] mprj_io_dm[71]
+ mprj_io_dm[72] mprj_io_dm[73] mprj_io_dm[74] mprj_io_dm[75] mprj_io_dm[76] mprj_io_dm[77]
+ mprj_io_dm[78] mprj_io_dm[79] mprj_io_dm[7] mprj_io_dm[80] mprj_io_dm[81] mprj_io_dm[82]
+ mprj_io_dm[83] mprj_io_dm[84] mprj_io_dm[85] mprj_io_dm[86] mprj_io_dm[87] mprj_io_dm[88]
+ mprj_io_dm[89] mprj_io_dm[8] mprj_io_dm[90] mprj_io_dm[91] mprj_io_dm[92] mprj_io_dm[93]
+ mprj_io_dm[94] mprj_io_dm[95] mprj_io_dm[96] mprj_io_dm[97] mprj_io_dm[98] mprj_io_dm[99]
+ mprj_io_dm[9] mprj_io_enh[0] mprj_io_enh[10] mprj_io_enh[11] mprj_io_enh[12] mprj_io_enh[13]
+ mprj_io_enh[14] mprj_io_enh[15] mprj_io_enh[16] mprj_io_enh[17] mprj_io_enh[18]
+ mprj_io_enh[19] mprj_io_enh[1] mprj_io_enh[20] mprj_io_enh[21] mprj_io_enh[22] mprj_io_enh[23]
+ mprj_io_enh[24] mprj_io_enh[25] mprj_io_enh[26] mprj_io_enh[27] mprj_io_enh[28]
+ mprj_io_enh[29] mprj_io_enh[2] mprj_io_enh[30] mprj_io_enh[31] mprj_io_enh[32] mprj_io_enh[33]
+ mprj_io_enh[34] mprj_io_enh[35] mprj_io_enh[36] mprj_io_enh[37] mprj_io_enh[3] mprj_io_enh[4]
+ mprj_io_enh[5] mprj_io_enh[6] mprj_io_enh[7] mprj_io_enh[8] mprj_io_enh[9] mprj_io_hldh_n[0]
+ mprj_io_hldh_n[10] mprj_io_hldh_n[11] mprj_io_hldh_n[12] mprj_io_hldh_n[13] mprj_io_hldh_n[14]
+ mprj_io_hldh_n[15] mprj_io_hldh_n[16] mprj_io_hldh_n[17] mprj_io_hldh_n[18] mprj_io_hldh_n[19]
+ mprj_io_hldh_n[1] mprj_io_hldh_n[20] mprj_io_hldh_n[21] mprj_io_hldh_n[22] mprj_io_hldh_n[23]
+ mprj_io_hldh_n[24] mprj_io_hldh_n[25] mprj_io_hldh_n[26] mprj_io_hldh_n[27] mprj_io_hldh_n[28]
+ mprj_io_hldh_n[29] mprj_io_hldh_n[2] mprj_io_hldh_n[30] mprj_io_hldh_n[31] mprj_io_hldh_n[32]
+ mprj_io_hldh_n[33] mprj_io_hldh_n[34] mprj_io_hldh_n[35] mprj_io_hldh_n[36] mprj_io_hldh_n[37]
+ mprj_io_hldh_n[3] mprj_io_hldh_n[4] mprj_io_hldh_n[5] mprj_io_hldh_n[6] mprj_io_hldh_n[7]
+ mprj_io_hldh_n[8] mprj_io_hldh_n[9] mprj_io_holdover[0] mprj_io_holdover[10] mprj_io_holdover[11]
+ mprj_io_holdover[12] mprj_io_holdover[13] mprj_io_holdover[14] mprj_io_holdover[15]
+ mprj_io_holdover[16] mprj_io_holdover[17] mprj_io_holdover[18] mprj_io_holdover[19]
+ mprj_io_holdover[1] mprj_io_holdover[20] mprj_io_holdover[21] mprj_io_holdover[22]
+ mprj_io_holdover[23] mprj_io_holdover[24] mprj_io_holdover[25] mprj_io_holdover[26]
+ mprj_io_holdover[27] mprj_io_holdover[28] mprj_io_holdover[29] mprj_io_holdover[2]
+ mprj_io_holdover[30] mprj_io_holdover[31] mprj_io_holdover[32] mprj_io_holdover[33]
+ mprj_io_holdover[34] mprj_io_holdover[35] mprj_io_holdover[36] mprj_io_holdover[37]
+ mprj_io_holdover[3] mprj_io_holdover[4] mprj_io_holdover[5] mprj_io_holdover[6]
+ mprj_io_holdover[7] mprj_io_holdover[8] mprj_io_holdover[9] mprj_io_ib_mode_sel[0]
+ mprj_io_ib_mode_sel[10] mprj_io_ib_mode_sel[11] mprj_io_ib_mode_sel[12] mprj_io_ib_mode_sel[13]
+ mprj_io_ib_mode_sel[14] mprj_io_ib_mode_sel[15] mprj_io_ib_mode_sel[16] mprj_io_ib_mode_sel[17]
+ mprj_io_ib_mode_sel[18] mprj_io_ib_mode_sel[19] mprj_io_ib_mode_sel[1] mprj_io_ib_mode_sel[20]
+ mprj_io_ib_mode_sel[21] mprj_io_ib_mode_sel[22] mprj_io_ib_mode_sel[23] mprj_io_ib_mode_sel[24]
+ mprj_io_ib_mode_sel[25] mprj_io_ib_mode_sel[26] mprj_io_ib_mode_sel[27] mprj_io_ib_mode_sel[28]
+ mprj_io_ib_mode_sel[29] mprj_io_ib_mode_sel[2] mprj_io_ib_mode_sel[30] mprj_io_ib_mode_sel[31]
+ mprj_io_ib_mode_sel[32] mprj_io_ib_mode_sel[33] mprj_io_ib_mode_sel[34] mprj_io_ib_mode_sel[35]
+ mprj_io_ib_mode_sel[36] mprj_io_ib_mode_sel[37] mprj_io_ib_mode_sel[3] mprj_io_ib_mode_sel[4]
+ mprj_io_ib_mode_sel[5] mprj_io_ib_mode_sel[6] mprj_io_ib_mode_sel[7] mprj_io_ib_mode_sel[8]
+ mprj_io_ib_mode_sel[9] mprj_io_in[0] mprj_io_in[10] mprj_io_in[11] mprj_io_in[12]
+ mprj_io_in[13] mprj_io_in[14] mprj_io_in[15] mprj_io_in[16] mprj_io_in[17] mprj_io_in[18]
+ mprj_io_in[19] mprj_io_in[1] mprj_io_in[20] mprj_io_in[21] mprj_io_in[22] mprj_io_in[23]
+ mprj_io_in[24] mprj_io_in[25] mprj_io_in[26] mprj_io_in[27] mprj_io_in[28] mprj_io_in[29]
+ mprj_io_in[2] mprj_io_in[30] mprj_io_in[31] mprj_io_in[32] mprj_io_in[33] mprj_io_in[34]
+ mprj_io_in[35] mprj_io_in[36] mprj_io_in[37] mprj_io_in[3] mprj_io_in[4] mprj_io_in[5]
+ mprj_io_in[6] mprj_io_in[7] mprj_io_in[8] mprj_io_in[9] mprj_io_inp_dis[0] mprj_io_inp_dis[10]
+ mprj_io_inp_dis[11] mprj_io_inp_dis[12] mprj_io_inp_dis[13] mprj_io_inp_dis[14]
+ mprj_io_inp_dis[15] mprj_io_inp_dis[16] mprj_io_inp_dis[17] mprj_io_inp_dis[18]
+ mprj_io_inp_dis[19] mprj_io_inp_dis[1] mprj_io_inp_dis[20] mprj_io_inp_dis[21] mprj_io_inp_dis[22]
+ mprj_io_inp_dis[23] mprj_io_inp_dis[24] mprj_io_inp_dis[25] mprj_io_inp_dis[26]
+ mprj_io_inp_dis[27] mprj_io_inp_dis[28] mprj_io_inp_dis[29] mprj_io_inp_dis[2] mprj_io_inp_dis[30]
+ mprj_io_inp_dis[31] mprj_io_inp_dis[32] mprj_io_inp_dis[33] mprj_io_inp_dis[34]
+ mprj_io_inp_dis[35] mprj_io_inp_dis[36] mprj_io_inp_dis[37] mprj_io_inp_dis[3] mprj_io_inp_dis[4]
+ mprj_io_inp_dis[5] mprj_io_inp_dis[6] mprj_io_inp_dis[7] mprj_io_inp_dis[8] mprj_io_inp_dis[9]
+ mprj_io_oeb[0] mprj_io_oeb[10] mprj_io_oeb[11] mprj_io_oeb[12] mprj_io_oeb[13] mprj_io_oeb[14]
+ mprj_io_oeb[15] mprj_io_oeb[16] mprj_io_oeb[17] mprj_io_oeb[18] mprj_io_oeb[19]
+ mprj_io_oeb[1] mprj_io_oeb[20] mprj_io_oeb[21] mprj_io_oeb[22] mprj_io_oeb[23] mprj_io_oeb[24]
+ mprj_io_oeb[25] mprj_io_oeb[26] mprj_io_oeb[27] mprj_io_oeb[28] mprj_io_oeb[29]
+ mprj_io_oeb[2] mprj_io_oeb[30] mprj_io_oeb[31] mprj_io_oeb[32] mprj_io_oeb[33] mprj_io_oeb[34]
+ mprj_io_oeb[35] mprj_io_oeb[36] mprj_io_oeb[37] mprj_io_oeb[3] mprj_io_oeb[4] mprj_io_oeb[5]
+ mprj_io_oeb[6] mprj_io_oeb[7] mprj_io_oeb[8] mprj_io_oeb[9] mprj_io_out[0] mprj_io_out[10]
+ mprj_io_out[11] mprj_io_out[12] mprj_io_out[13] mprj_io_out[14] mprj_io_out[15]
+ mprj_io_out[16] mprj_io_out[17] mprj_io_out[18] mprj_io_out[19] mprj_io_out[1] mprj_io_out[20]
+ mprj_io_out[21] mprj_io_out[22] mprj_io_out[23] mprj_io_out[24] mprj_io_out[25]
+ mprj_io_out[26] mprj_io_out[27] mprj_io_out[28] mprj_io_out[29] mprj_io_out[2] mprj_io_out[30]
+ mprj_io_out[31] mprj_io_out[32] mprj_io_out[33] mprj_io_out[34] mprj_io_out[35]
+ mprj_io_out[36] mprj_io_out[37] mprj_io_out[3] mprj_io_out[4] mprj_io_out[5] mprj_io_out[6]
+ mprj_io_out[7] mprj_io_out[8] mprj_io_out[9] mprj_io_slow_sel[0] mprj_io_slow_sel[10]
+ mprj_io_slow_sel[11] mprj_io_slow_sel[12] mprj_io_slow_sel[13] mprj_io_slow_sel[14]
+ mprj_io_slow_sel[15] mprj_io_slow_sel[16] mprj_io_slow_sel[17] mprj_io_slow_sel[18]
+ mprj_io_slow_sel[19] mprj_io_slow_sel[1] mprj_io_slow_sel[20] mprj_io_slow_sel[21]
+ mprj_io_slow_sel[22] mprj_io_slow_sel[23] mprj_io_slow_sel[24] mprj_io_slow_sel[25]
+ mprj_io_slow_sel[26] mprj_io_slow_sel[27] mprj_io_slow_sel[28] mprj_io_slow_sel[29]
+ mprj_io_slow_sel[2] mprj_io_slow_sel[30] mprj_io_slow_sel[31] mprj_io_slow_sel[32]
+ mprj_io_slow_sel[33] mprj_io_slow_sel[34] mprj_io_slow_sel[35] mprj_io_slow_sel[36]
+ mprj_io_slow_sel[37] mprj_io_slow_sel[3] mprj_io_slow_sel[4] mprj_io_slow_sel[5]
+ mprj_io_slow_sel[6] mprj_io_slow_sel[7] mprj_io_slow_sel[8] mprj_io_slow_sel[9]
+ mprj_io_vtrip_sel[0] mprj_io_vtrip_sel[10] mprj_io_vtrip_sel[11] mprj_io_vtrip_sel[12]
+ mprj_io_vtrip_sel[13] mprj_io_vtrip_sel[14] mprj_io_vtrip_sel[15] mprj_io_vtrip_sel[16]
+ mprj_io_vtrip_sel[17] mprj_io_vtrip_sel[18] mprj_io_vtrip_sel[19] mprj_io_vtrip_sel[1]
+ mprj_io_vtrip_sel[20] mprj_io_vtrip_sel[21] mprj_io_vtrip_sel[22] mprj_io_vtrip_sel[23]
+ mprj_io_vtrip_sel[24] mprj_io_vtrip_sel[25] mprj_io_vtrip_sel[26] mprj_io_vtrip_sel[27]
+ mprj_io_vtrip_sel[28] mprj_io_vtrip_sel[29] mprj_io_vtrip_sel[2] mprj_io_vtrip_sel[30]
+ mprj_io_vtrip_sel[31] mprj_io_vtrip_sel[32] mprj_io_vtrip_sel[33] mprj_io_vtrip_sel[34]
+ mprj_io_vtrip_sel[35] mprj_io_vtrip_sel[36] mprj_io_vtrip_sel[37] mprj_io_vtrip_sel[3]
+ mprj_io_vtrip_sel[4] mprj_io_vtrip_sel[5] mprj_io_vtrip_sel[6] mprj_io_vtrip_sel[7]
+ mprj_io_vtrip_sel[8] mprj_io_vtrip_sel[9] por porb_h resetb resetb_core_h vccd vccd1
+ vccd1_pad vccd2 vccd2_pad vccd_pad vdda vdda1 vdda1_pad vdda2 vdda2_pad vdda_pad
+ vddio vddio_pad vssa vssa1 vssa1_pad vssa2 vssa2_pad vssa_pad vssd vssd1 vssd1_pad
+ vssd2 vssd2_pad vssd_pad vssio vssio_pad vssio_pad2 vddio_pad2 vssa1_pad2 vdda1_pad2
+ VSUBS
XFILLER_592 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_570 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xclock_pad clock_pad/IN_H clock_pad/PAD_A_NOESD_H clock_pad/PAD_A_ESD_0_H clock_pad/PAD_A_ESD_1_H
+ clock vssd vssd vccd vddio clock_core por vssd porb_h porb_h clock_pad/TIE_LO_ESD
+ vccd clock_pad/TIE_HI_ESD clock_pad/TIE_LO_ESD vssd vssd vssd vssd vssd vccd vssa
+ vssd vssd gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[17\] mprj_pads.area2_io_pad\[17\]/IN_H mprj_pads.area2_io_pad\[17\]/PAD_A_NOESD_H
+ mprj_analog_io[28] mprj_pads.area2_io_pad\[17\]/PAD_A_ESD_1_H mprj_io[35] mprj_io_dm[107]
+ mprj_io_dm[106] mprj_io_dm[105] mprj_io_hldh_n[35] mprj_io_in[35] mprj_io_inp_dis[35]
+ mprj_io_ib_mode_sel[35] mprj_io_enh[35] porb_h mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD
+ mprj_io_oeb[35] mprj_pads.area2_io_pad\[17\]/TIE_HI_ESD mprj_pads.area2_io_pad\[17\]/TIE_LO_ESD
+ mprj_io_slow_sel[35] mprj_io_vtrip_sel[35] mprj_io_holdover[35] mprj_io_analog_en[35]
+ mprj_io_analog_sel[35] vccd vssio mprj_io_analog_pol[35] mprj_io_out[35] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_25 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_14 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_69 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_58 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_47 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_36 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vccd_lvc_clamped_pad
Xmprj_pads.area2_io_pad\[7\] mprj_pads.area2_io_pad\[7\]/IN_H mprj_pads.area2_io_pad\[7\]/PAD_A_NOESD_H
+ mprj_analog_io[18] mprj_pads.area2_io_pad\[7\]/PAD_A_ESD_1_H mprj_io[25] mprj_io_dm[77]
+ mprj_io_dm[76] mprj_io_dm[75] mprj_io_hldh_n[25] mprj_io_in[25] mprj_io_inp_dis[25]
+ mprj_io_ib_mode_sel[25] mprj_io_enh[25] porb_h mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD
+ mprj_io_oeb[25] mprj_pads.area2_io_pad\[7\]/TIE_HI_ESD mprj_pads.area2_io_pad\[7\]/TIE_LO_ESD
+ mprj_io_slow_sel[25] mprj_io_vtrip_sel[25] mprj_io_holdover[25] mprj_io_analog_en[25]
+ mprj_io_analog_sel[25] vccd vssio mprj_io_analog_pol[25] mprj_io_out[25] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_229 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_207 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_796 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_785 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_774 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_763 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_752 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_741 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_730 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_593 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_582 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_560 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[7\] mprj_pads.area1_io_pad\[7\]/IN_H mprj_pads.area1_io_pad\[7\]/PAD_A_NOESD_H
+ mprj_analog_io[0] mprj_pads.area1_io_pad\[7\]/PAD_A_ESD_1_H mprj_io[7] mprj_io_dm[23]
+ mprj_io_dm[22] mprj_io_dm[21] mprj_io_hldh_n[7] mprj_io_in[7] mprj_io_inp_dis[7]
+ mprj_io_ib_mode_sel[7] mprj_io_enh[7] porb_h mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD
+ mprj_io_oeb[7] mprj_pads.area1_io_pad\[7\]/TIE_HI_ESD mprj_pads.area1_io_pad\[7\]/TIE_LO_ESD
+ mprj_io_slow_sel[7] mprj_io_vtrip_sel[7] mprj_io_holdover[7] mprj_io_analog_en[7]
+ mprj_io_analog_sel[7] vccd vssio mprj_io_analog_pol[7] mprj_io_out[7] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_59 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_48 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_37 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_26 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_15 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_208 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_797 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_786 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_775 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_764 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_742 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_731 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_720 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_594 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_583 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_572 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_550 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_380 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_391 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[11\] mprj_pads.area1_io_pad\[11\]/IN_H mprj_pads.area1_io_pad\[11\]/PAD_A_NOESD_H
+ mprj_analog_io[4] mprj_pads.area1_io_pad\[11\]/PAD_A_ESD_1_H mprj_io[11] mprj_io_dm[35]
+ mprj_io_dm[34] mprj_io_dm[33] mprj_io_hldh_n[11] mprj_io_in[11] mprj_io_inp_dis[11]
+ mprj_io_ib_mode_sel[11] mprj_io_enh[11] porb_h mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD
+ mprj_io_oeb[11] mprj_pads.area1_io_pad\[11\]/TIE_HI_ESD mprj_pads.area1_io_pad\[11\]/TIE_LO_ESD
+ mprj_io_slow_sel[11] mprj_io_vtrip_sel[11] mprj_io_holdover[11] mprj_io_analog_en[11]
+ mprj_io_analog_sel[11] vccd vssio mprj_io_analog_pol[11] mprj_io_out[11] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_49 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_38 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_27 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_16 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_209 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_798 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_787 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_776 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_765 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_754 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_732 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_721 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_710 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_595 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_584 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_573 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_562 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_540 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_381 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_392 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[15\] mprj_pads.area2_io_pad\[15\]/IN_H mprj_pads.area2_io_pad\[15\]/PAD_A_NOESD_H
+ mprj_analog_io[26] mprj_pads.area2_io_pad\[15\]/PAD_A_ESD_1_H mprj_io[33] mprj_io_dm[101]
+ mprj_io_dm[100] mprj_io_dm[99] mprj_io_hldh_n[33] mprj_io_in[33] mprj_io_inp_dis[33]
+ mprj_io_ib_mode_sel[33] mprj_io_enh[33] porb_h mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD
+ mprj_io_oeb[33] mprj_pads.area2_io_pad\[15\]/TIE_HI_ESD mprj_pads.area2_io_pad\[15\]/TIE_LO_ESD
+ mprj_io_slow_sel[33] mprj_io_vtrip_sel[33] mprj_io_holdover[33] mprj_io_analog_en[33]
+ mprj_io_analog_sel[33] vccd vssio mprj_io_analog_pol[33] mprj_io_out[33] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_39 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_28 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[5\] mprj_pads.area2_io_pad\[5\]/IN_H mprj_pads.area2_io_pad\[5\]/PAD_A_NOESD_H
+ mprj_analog_io[16] mprj_pads.area2_io_pad\[5\]/PAD_A_ESD_1_H mprj_io[23] mprj_io_dm[71]
+ mprj_io_dm[70] mprj_io_dm[69] mprj_io_hldh_n[23] mprj_io_in[23] mprj_io_inp_dis[23]
+ mprj_io_ib_mode_sel[23] mprj_io_enh[23] porb_h mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD
+ mprj_io_oeb[23] mprj_pads.area2_io_pad\[5\]/TIE_HI_ESD mprj_pads.area2_io_pad\[5\]/TIE_LO_ESD
+ mprj_io_slow_sel[23] mprj_io_vtrip_sel[23] mprj_io_holdover[23] mprj_io_analog_en[23]
+ mprj_io_analog_sel[23] vccd vssio mprj_io_analog_pol[23] mprj_io_out[23] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_799 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_788 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_777 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_766 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_755 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_744 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_733 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_722 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_711 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_700 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_596 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_585 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_574 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_563 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_552 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_530 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_360 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_382 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_393 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_190 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_29 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_18 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[5\] mprj_pads.area1_io_pad\[5\]/IN_H mprj_pads.area1_io_pad\[5\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[5\]/PAD_A_ESD_1_H
+ mprj_io[5] mprj_io_dm[17] mprj_io_dm[16] mprj_io_dm[15] mprj_io_hldh_n[5] mprj_io_in[5]
+ mprj_io_inp_dis[5] mprj_io_ib_mode_sel[5] mprj_io_enh[5] porb_h mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD
+ mprj_io_oeb[5] mprj_pads.area1_io_pad\[5\]/TIE_HI_ESD mprj_pads.area1_io_pad\[5\]/TIE_LO_ESD
+ mprj_io_slow_sel[5] mprj_io_vtrip_sel[5] mprj_io_holdover[5] mprj_io_analog_en[5]
+ mprj_io_analog_sel[5] vccd vssio mprj_io_analog_pol[5] mprj_io_out[5] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xdisconnect_vdda_0 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
XFILLER_723 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_712 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_701 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_789 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_778 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_767 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_756 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_745 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_597 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_586 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_575 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_564 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_553 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_542 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_520 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_350 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_361 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_383 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_394 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_19 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_191 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_180 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xdisconnect_vdda_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
XFILLER_779 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_768 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_757 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_746 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_735 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_713 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_702 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_598 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_587 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_576 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_565 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_554 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_543 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_532 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_510 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser2_corner gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xmgmt_vddio_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio_pad vssa
+ vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vddio_hvc_clamped_pad
XFILLER_351 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_362 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_384 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_395 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_170 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_192 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_181 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[13\] mprj_pads.area2_io_pad\[13\]/IN_H mprj_pads.area2_io_pad\[13\]/PAD_A_NOESD_H
+ mprj_analog_io[24] mprj_pads.area2_io_pad\[13\]/PAD_A_ESD_1_H mprj_io[31] mprj_io_dm[95]
+ mprj_io_dm[94] mprj_io_dm[93] mprj_io_hldh_n[31] mprj_io_in[31] mprj_io_inp_dis[31]
+ mprj_io_ib_mode_sel[31] mprj_io_enh[31] porb_h mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD
+ mprj_io_oeb[31] mprj_pads.area2_io_pad\[13\]/TIE_HI_ESD mprj_pads.area2_io_pad\[13\]/TIE_LO_ESD
+ mprj_io_slow_sel[31] mprj_io_vtrip_sel[31] mprj_io_holdover[31] mprj_io_analog_en[31]
+ mprj_io_analog_sel[31] vccd vssio mprj_io_analog_pol[31] mprj_io_out[31] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xdisconnect_vdda_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio gpio_pad/VDDIO_Q vccd
+ vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vdda_slice_5um
Xmgmt_vssio_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio_pad vssa
+ vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssio_hvc_clamped_pad
XFILLER_769 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_758 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_747 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_736 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_725 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_714 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_703 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[3\] mprj_pads.area2_io_pad\[3\]/IN_H mprj_pads.area2_io_pad\[3\]/PAD_A_NOESD_H
+ mprj_analog_io[14] mprj_pads.area2_io_pad\[3\]/PAD_A_ESD_1_H mprj_io[21] mprj_io_dm[65]
+ mprj_io_dm[64] mprj_io_dm[63] mprj_io_hldh_n[21] mprj_io_in[21] mprj_io_inp_dis[21]
+ mprj_io_ib_mode_sel[21] mprj_io_enh[21] porb_h mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD
+ mprj_io_oeb[21] mprj_pads.area2_io_pad\[3\]/TIE_HI_ESD mprj_pads.area2_io_pad\[3\]/TIE_LO_ESD
+ mprj_io_slow_sel[21] mprj_io_vtrip_sel[21] mprj_io_holdover[21] mprj_io_analog_en[21]
+ mprj_io_analog_sel[21] vccd vssio mprj_io_analog_pol[21] mprj_io_out[21] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_500 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_599 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_588 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_577 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_566 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_555 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_544 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_533 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_522 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_330 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_341 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_385 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_396 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_171 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_160 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xbus_tie_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area1_io_pad\[3\] mprj_pads.area1_io_pad\[3\]/IN_H mprj_pads.area1_io_pad\[3\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[3\]/PAD_A_ESD_1_H
+ mprj_io[3] mprj_io_dm[11] mprj_io_dm[10] mprj_io_dm[9] mprj_io_hldh_n[3] mprj_io_in[3]
+ mprj_io_inp_dis[3] mprj_io_ib_mode_sel[3] mprj_io_enh[3] porb_h mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD
+ mprj_io_oeb[3] mprj_pads.area1_io_pad\[3\]/TIE_HI_ESD mprj_pads.area1_io_pad\[3\]/TIE_LO_ESD
+ mprj_io_slow_sel[3] mprj_io_vtrip_sel[3] mprj_io_holdover[3] mprj_io_analog_en[3]
+ mprj_io_analog_sel[3] vccd vssio mprj_io_analog_pol[3] mprj_io_out[3] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_759 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_748 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_737 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_726 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_704 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_589 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_578 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_567 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_556 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_545 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_534 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_523 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_512 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_331 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_342 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_364 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_375 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_386 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_397 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_172 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_161 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_194 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_749 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_738 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_727 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_716 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_705 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser2_vdda_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
XFILLER_579 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_568 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_557 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_546 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_535 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_524 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_513 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_502 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_310 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_332 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_343 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_365 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_376 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_387 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_398 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_173 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_162 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_151 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_140 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_195 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xbus_tie_70 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[11\] mprj_pads.area2_io_pad\[11\]/IN_H mprj_pads.area2_io_pad\[11\]/PAD_A_NOESD_H
+ mprj_analog_io[22] mprj_pads.area2_io_pad\[11\]/PAD_A_ESD_1_H mprj_io[29] mprj_io_dm[89]
+ mprj_io_dm[88] mprj_io_dm[87] mprj_io_hldh_n[29] mprj_io_in[29] mprj_io_inp_dis[29]
+ mprj_io_ib_mode_sel[29] mprj_io_enh[29] porb_h mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD
+ mprj_io_oeb[29] mprj_pads.area2_io_pad\[11\]/TIE_HI_ESD mprj_pads.area2_io_pad\[11\]/TIE_LO_ESD
+ mprj_io_slow_sel[29] mprj_io_vtrip_sel[29] mprj_io_holdover[29] mprj_io_analog_en[29]
+ mprj_io_analog_sel[29] vccd vssio mprj_io_analog_pol[29] mprj_io_out[29] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_3 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_739 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_728 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_717 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_569 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_558 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_547 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_536 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_525 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_514 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_503 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[1\] mprj_pads.area2_io_pad\[1\]/IN_H mprj_pads.area2_io_pad\[1\]/PAD_A_NOESD_H
+ mprj_analog_io[12] mprj_pads.area2_io_pad\[1\]/PAD_A_ESD_1_H mprj_io[19] mprj_io_dm[59]
+ mprj_io_dm[58] mprj_io_dm[57] mprj_io_hldh_n[19] mprj_io_in[19] mprj_io_inp_dis[19]
+ mprj_io_ib_mode_sel[19] mprj_io_enh[19] porb_h mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD
+ mprj_io_oeb[19] mprj_pads.area2_io_pad\[1\]/TIE_HI_ESD mprj_pads.area2_io_pad\[1\]/TIE_LO_ESD
+ mprj_io_slow_sel[19] mprj_io_vtrip_sel[19] mprj_io_holdover[19] mprj_io_analog_en[19]
+ mprj_io_analog_sel[19] vccd vssio mprj_io_analog_pol[19] mprj_io_out[19] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_300 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_311 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_333 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_344 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_366 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_377 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_388 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_399 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_141 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_130 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_174 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_152 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_196 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xbus_tie_4 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_60 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_71 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_729 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_718 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_707 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[1\] mprj_pads.area1_io_pad\[1\]/IN_H mprj_pads.area1_io_pad\[1\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[1\]/PAD_A_ESD_1_H
+ mprj_io[1] mprj_io_dm[5] mprj_io_dm[4] mprj_io_dm[3] mprj_io_hldh_n[1] mprj_io_in[1]
+ mprj_io_inp_dis[1] mprj_io_ib_mode_sel[1] mprj_io_enh[1] porb_h mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD
+ mprj_io_oeb[1] mprj_pads.area1_io_pad\[1\]/TIE_HI_ESD mprj_pads.area1_io_pad\[1\]/TIE_LO_ESD
+ mprj_io_slow_sel[1] mprj_io_vtrip_sel[1] mprj_io_holdover[1] mprj_io_analog_en[1]
+ mprj_io_analog_sel[1] vccd vssio mprj_io_analog_pol[1] mprj_io_out[1] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_559 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_548 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_537 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_526 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_515 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_504 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_334 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_345 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_367 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_378 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_389 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_175 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_164 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_153 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_142 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_131 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_120 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_197 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xgpio_pad gpio_pad/IN_H gpio_pad/PAD_A_NOESD_H gpio_pad/PAD_A_ESD_0_H gpio_pad/PAD_A_ESD_1_H
+ gpio gpio_mode1_core gpio_mode1_core gpio_mode0_core vddio gpio_in_core gpio_inenb_core
+ vssd porb_h porb_h gpio_pad/TIE_LO_ESD gpio_outenb_core gpio_pad/TIE_HI_ESD gpio_pad/TIE_LO_ESD
+ vssd vssd vssd vssd vssd vccd vssa vssd gpio_out_core gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_5 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_50 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_61 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_72 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_719 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_708 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_516 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_505 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_549 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_538 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_527 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_313 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_324 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_368 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_379 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_176 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_165 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_154 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_143 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[16\] mprj_pads.area1_io_pad\[16\]/IN_H mprj_pads.area1_io_pad\[16\]/PAD_A_NOESD_H
+ mprj_analog_io[9] mprj_pads.area1_io_pad\[16\]/PAD_A_ESD_1_H mprj_io[16] mprj_io_dm[50]
+ mprj_io_dm[49] mprj_io_dm[48] mprj_io_hldh_n[16] mprj_io_in[16] mprj_io_inp_dis[16]
+ mprj_io_ib_mode_sel[16] mprj_io_enh[16] porb_h mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD
+ mprj_io_oeb[16] mprj_pads.area1_io_pad\[16\]/TIE_HI_ESD mprj_pads.area1_io_pad\[16\]/TIE_LO_ESD
+ mprj_io_slow_sel[16] mprj_io_vtrip_sel[16] mprj_io_holdover[16] mprj_io_analog_en[16]
+ mprj_io_analog_sel[16] vccd vssio mprj_io_analog_pol[16] mprj_io_out[16] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_132 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_121 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_198 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser1_vdda_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda1_pad vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xbus_tie_6 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_40 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_51 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_62 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_709 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_539 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_528 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_517 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_506 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_314 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_325 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_347 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_358 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_166 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_155 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_144 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_133 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_122 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_111 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_100 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_188 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_177 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__vccd_lvc_clamped2_pad
Xbus_tie_30 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_41 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_52 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_63 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_7 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_529 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_518 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_507 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_315 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_326 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_348 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_359 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xmgmt_vssa_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
XFILLER_167 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_156 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_145 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_134 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_123 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_112 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_101 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_189 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_178 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xmgmt_corner\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
XFILLER_690 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vssa_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1_pad2 vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xbus_tie_31 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_20 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_42 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_53 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_64 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_8 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_519 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_508 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_316 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_327 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_349 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_157 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_146 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_135 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_113 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_102 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_168 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_179 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_680 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_691 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[14\] mprj_pads.area1_io_pad\[14\]/IN_H mprj_pads.area1_io_pad\[14\]/PAD_A_NOESD_H
+ mprj_analog_io[7] mprj_pads.area1_io_pad\[14\]/PAD_A_ESD_1_H mprj_io[14] mprj_io_dm[44]
+ mprj_io_dm[43] mprj_io_dm[42] mprj_io_hldh_n[14] mprj_io_in[14] mprj_io_inp_dis[14]
+ mprj_io_ib_mode_sel[14] mprj_io_enh[14] porb_h mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD
+ mprj_io_oeb[14] mprj_pads.area1_io_pad\[14\]/TIE_HI_ESD mprj_pads.area1_io_pad\[14\]/TIE_LO_ESD
+ mprj_io_slow_sel[14] mprj_io_vtrip_sel[14] mprj_io_holdover[14] mprj_io_analog_en[14]
+ mprj_io_analog_sel[14] vccd vssio mprj_io_analog_pol[14] mprj_io_out[14] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xbus_tie_32 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_21 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_10 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_9 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_43 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_54 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_65 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_509 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_317 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_328 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_169 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_158 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_147 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_136 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_125 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_114 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_103 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_670 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_681 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_692 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[18\] mprj_pads.area2_io_pad\[18\]/IN_H mprj_pads.area2_io_pad\[18\]/PAD_A_NOESD_H
+ mprj_analog_io[29] mprj_pads.area2_io_pad\[18\]/PAD_A_ESD_1_H mprj_io[36] mprj_io_dm[110]
+ mprj_io_dm[109] mprj_io_dm[108] mprj_io_hldh_n[36] mprj_io_in[36] mprj_io_inp_dis[36]
+ mprj_io_ib_mode_sel[36] mprj_io_enh[36] porb_h mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD
+ mprj_io_oeb[36] mprj_pads.area2_io_pad\[18\]/TIE_HI_ESD mprj_pads.area2_io_pad\[18\]/TIE_LO_ESD
+ mprj_io_slow_sel[36] mprj_io_vtrip_sel[36] mprj_io_holdover[36] mprj_io_analog_en[36]
+ mprj_io_analog_sel[36] vccd vssio mprj_io_analog_pol[36] mprj_io_out[36] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xdisconnect_vccd_0 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vssio gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vccd_slice_5um
Xbus_tie_33 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_22 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_11 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_44 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_55 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_66 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmprj_pads.area2_io_pad\[8\] mprj_pads.area2_io_pad\[8\]/IN_H mprj_pads.area2_io_pad\[8\]/PAD_A_NOESD_H
+ mprj_analog_io[19] mprj_pads.area2_io_pad\[8\]/PAD_A_ESD_1_H mprj_io[26] mprj_io_dm[80]
+ mprj_io_dm[79] mprj_io_dm[78] mprj_io_hldh_n[26] mprj_io_in[26] mprj_io_inp_dis[26]
+ mprj_io_ib_mode_sel[26] mprj_io_enh[26] porb_h mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD
+ mprj_io_oeb[26] mprj_pads.area2_io_pad\[8\]/TIE_HI_ESD mprj_pads.area2_io_pad\[8\]/TIE_LO_ESD
+ mprj_io_slow_sel[26] mprj_io_vtrip_sel[26] mprj_io_holdover[26] mprj_io_analog_en[26]
+ mprj_io_analog_sel[26] vccd vssio mprj_io_analog_pol[26] mprj_io_out[26] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_307 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_159 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_148 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_126 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_115 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_104 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_660 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_671 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_682 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_693 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_490 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_34 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_23 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_12 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_45 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_56 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_67 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xdisconnect_vccd_1 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vssio gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vccd_slice_5um
Xmprj_pads.area1_io_pad\[8\] mprj_pads.area1_io_pad\[8\]/IN_H mprj_pads.area1_io_pad\[8\]/PAD_A_NOESD_H
+ mprj_analog_io[1] mprj_pads.area1_io_pad\[8\]/PAD_A_ESD_1_H mprj_io[8] mprj_io_dm[26]
+ mprj_io_dm[25] mprj_io_dm[24] mprj_io_hldh_n[8] mprj_io_in[8] mprj_io_inp_dis[8]
+ mprj_io_ib_mode_sel[8] mprj_io_enh[8] porb_h mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD
+ mprj_io_oeb[8] mprj_pads.area1_io_pad\[8\]/TIE_HI_ESD mprj_pads.area1_io_pad\[8\]/TIE_LO_ESD
+ mprj_io_slow_sel[8] mprj_io_vtrip_sel[8] mprj_io_holdover[8] mprj_io_analog_en[8]
+ mprj_io_analog_sel[8] vccd vssio mprj_io_analog_pol[8] mprj_io_out[8] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xresetb_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio porb_h vccd vssio vssio vssio
+ resetb resetb_pad/PAD_A_ESD_H vssio resetb_pad/TIE_HI_ESD resetb_pad/TIE_LO_ESD
+ resetb_pad/PAD_A_ESD_H resetb_core_h vccd vccd vdda vddio gpio_pad/VDDIO_Q vssa
+ vssd vssio gpio_pad/VSSIO_Q vddio sky130_fd_io__top_xres4v2
XFILLER_308 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_149 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_138 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_127 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_116 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_105 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_650 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_661 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_672 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_683 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_694 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_480 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_24 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_13 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_35 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_46 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_57 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_68 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xdisconnect_vccd_2 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vssio gpio_pad/VSSIO_Q sky130_ef_io__disconnect_vccd_slice_5um
Xmprj_pads.area1_io_pad\[12\] mprj_pads.area1_io_pad\[12\]/IN_H mprj_pads.area1_io_pad\[12\]/PAD_A_NOESD_H
+ mprj_analog_io[5] mprj_pads.area1_io_pad\[12\]/PAD_A_ESD_1_H mprj_io[12] mprj_io_dm[38]
+ mprj_io_dm[37] mprj_io_dm[36] mprj_io_hldh_n[12] mprj_io_in[12] mprj_io_inp_dis[12]
+ mprj_io_ib_mode_sel[12] mprj_io_enh[12] porb_h mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD
+ mprj_io_oeb[12] mprj_pads.area1_io_pad\[12\]/TIE_HI_ESD mprj_pads.area1_io_pad\[12\]/TIE_LO_ESD
+ mprj_io_slow_sel[12] mprj_io_vtrip_sel[12] mprj_io_holdover[12] mprj_io_analog_en[12]
+ mprj_io_analog_sel[12] vccd vssio mprj_io_analog_pol[12] mprj_io_out[12] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_810 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_309 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_139 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_128 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_117 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_106 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_651 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_662 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_673 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_684 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_695 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_492 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_25 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_14 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_36 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_47 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_58 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_69 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_470 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[16\] mprj_pads.area2_io_pad\[16\]/IN_H mprj_pads.area2_io_pad\[16\]/PAD_A_NOESD_H
+ mprj_analog_io[27] mprj_pads.area2_io_pad\[16\]/PAD_A_ESD_1_H mprj_io[34] mprj_io_dm[104]
+ mprj_io_dm[103] mprj_io_dm[102] mprj_io_hldh_n[34] mprj_io_in[34] mprj_io_inp_dis[34]
+ mprj_io_ib_mode_sel[34] mprj_io_enh[34] porb_h mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD
+ mprj_io_oeb[34] mprj_pads.area2_io_pad\[16\]/TIE_HI_ESD mprj_pads.area2_io_pad\[16\]/TIE_LO_ESD
+ mprj_io_slow_sel[34] mprj_io_vtrip_sel[34] mprj_io_holdover[34] mprj_io_analog_en[34]
+ mprj_io_analog_sel[34] vccd vssio mprj_io_analog_pol[34] mprj_io_out[34] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[6\] mprj_pads.area2_io_pad\[6\]/IN_H mprj_pads.area2_io_pad\[6\]/PAD_A_NOESD_H
+ mprj_analog_io[17] mprj_pads.area2_io_pad\[6\]/PAD_A_ESD_1_H mprj_io[24] mprj_io_dm[74]
+ mprj_io_dm[73] mprj_io_dm[72] mprj_io_hldh_n[24] mprj_io_in[24] mprj_io_inp_dis[24]
+ mprj_io_ib_mode_sel[24] mprj_io_enh[24] porb_h mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD
+ mprj_io_oeb[24] mprj_pads.area2_io_pad\[6\]/TIE_HI_ESD mprj_pads.area2_io_pad\[6\]/TIE_LO_ESD
+ mprj_io_slow_sel[24] mprj_io_vtrip_sel[24] mprj_io_holdover[24] mprj_io_analog_en[24]
+ mprj_io_analog_sel[24] vccd vssio mprj_io_analog_pol[24] mprj_io_out[24] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_811 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xflash_csb_pad flash_csb_pad/IN_H flash_csb_pad/PAD_A_NOESD_H flash_csb_pad/PAD_A_ESD_0_H
+ flash_csb_pad/PAD_A_ESD_1_H flash_csb vccd vccd vssd vddio flash_csb_pad/IN flash_csb_ieb_core
+ vssd porb_h porb_h flash_csb_pad/TIE_LO_ESD flash_csb_oeb_core flash_csb_pad/TIE_HI_ESD
+ flash_csb_pad/TIE_LO_ESD vssd vssd vssd vssd vssd vccd vssa vssd flash_csb_core
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_129 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_118 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_107 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_641 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_652 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_663 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_674 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_685 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_493 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_482 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_460 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xbus_tie_26 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_15 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_37 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_48 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_59 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_290 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area1_io_pad\[6\] mprj_pads.area1_io_pad\[6\]/IN_H mprj_pads.area1_io_pad\[6\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[6\]/PAD_A_ESD_1_H
+ mprj_io[6] mprj_io_dm[20] mprj_io_dm[19] mprj_io_dm[18] mprj_io_hldh_n[6] mprj_io_in[6]
+ mprj_io_inp_dis[6] mprj_io_ib_mode_sel[6] mprj_io_enh[6] porb_h mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD
+ mprj_io_oeb[6] mprj_pads.area1_io_pad\[6\]/TIE_HI_ESD mprj_pads.area1_io_pad\[6\]/TIE_LO_ESD
+ mprj_io_slow_sel[6] mprj_io_vtrip_sel[6] mprj_io_holdover[6] mprj_io_analog_en[6]
+ mprj_io_analog_sel[6] vccd vssio mprj_io_analog_pol[6] mprj_io_out[6] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_812 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_801 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vssd_lvclmap_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd1_pad vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__vssd_lvc_clamped2_pad
XFILLER_119 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_108 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_697 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_631 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_642 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_653 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_664 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_675 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_686 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_494 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_483 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_450 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_472 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_27 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_16 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_38 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_49 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_280 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_291 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xmprj_pads.area1_io_pad\[10\] mprj_pads.area1_io_pad\[10\]/IN_H mprj_pads.area1_io_pad\[10\]/PAD_A_NOESD_H
+ mprj_analog_io[3] mprj_pads.area1_io_pad\[10\]/PAD_A_ESD_1_H mprj_io[10] mprj_io_dm[32]
+ mprj_io_dm[31] mprj_io_dm[30] mprj_io_hldh_n[10] mprj_io_in[10] mprj_io_inp_dis[10]
+ mprj_io_ib_mode_sel[10] mprj_io_enh[10] porb_h mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD
+ mprj_io_oeb[10] mprj_pads.area1_io_pad\[10\]/TIE_HI_ESD mprj_pads.area1_io_pad\[10\]/TIE_LO_ESD
+ mprj_io_slow_sel[10] mprj_io_vtrip_sel[10] mprj_io_holdover[10] mprj_io_analog_en[10]
+ mprj_io_analog_sel[10] vccd vssio mprj_io_analog_pol[10] mprj_io_out[10] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_813 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_802 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xflash_io1_pad flash_io1_pad/IN_H flash_io1_pad/PAD_A_NOESD_H flash_io1_pad/PAD_A_ESD_0_H
+ flash_io1_pad/PAD_A_ESD_1_H flash_io1 flash_io1_ieb_core flash_io1_ieb_core flash_io1_oeb_core
+ vddio flash_io1_di_core flash_io1_ieb_core vssd porb_h porb_h flash_io1_pad/TIE_LO_ESD
+ flash_io1_oeb_core flash_io1_pad/TIE_HI_ESD flash_io1_pad/TIE_LO_ESD vssd vssd vssd
+ vssd vssd vccd vssa vssd flash_io1_do_core gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_610 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_698 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_632 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_643 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_654 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_665 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_676 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmgmt_vddio_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vddio_pad2 vssa2
+ vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__vddio_hvc_clamped_pad
XFILLER_495 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_484 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_440 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_462 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_473 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_28 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_17 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_39 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xmgmt_vssd_lvclmap_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vssd_lvc_clamped_pad
XFILLER_281 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_292 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area2_io_pad\[14\] mprj_pads.area2_io_pad\[14\]/IN_H mprj_pads.area2_io_pad\[14\]/PAD_A_NOESD_H
+ mprj_analog_io[25] mprj_pads.area2_io_pad\[14\]/PAD_A_ESD_1_H mprj_io[32] mprj_io_dm[98]
+ mprj_io_dm[97] mprj_io_dm[96] mprj_io_hldh_n[32] mprj_io_in[32] mprj_io_inp_dis[32]
+ mprj_io_ib_mode_sel[32] mprj_io_enh[32] porb_h mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD
+ mprj_io_oeb[32] mprj_pads.area2_io_pad\[14\]/TIE_HI_ESD mprj_pads.area2_io_pad\[14\]/TIE_LO_ESD
+ mprj_io_slow_sel[32] mprj_io_vtrip_sel[32] mprj_io_holdover[32] mprj_io_analog_en[32]
+ mprj_io_analog_sel[32] vccd vssio mprj_io_analog_pol[32] mprj_io_out[32] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_814 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_803 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[4\] mprj_pads.area2_io_pad\[4\]/IN_H mprj_pads.area2_io_pad\[4\]/PAD_A_NOESD_H
+ mprj_analog_io[15] mprj_pads.area2_io_pad\[4\]/PAD_A_ESD_1_H mprj_io[22] mprj_io_dm[68]
+ mprj_io_dm[67] mprj_io_dm[66] mprj_io_hldh_n[22] mprj_io_in[22] mprj_io_inp_dis[22]
+ mprj_io_ib_mode_sel[22] mprj_io_enh[22] porb_h mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD
+ mprj_io_oeb[22] mprj_pads.area2_io_pad\[4\]/TIE_HI_ESD mprj_pads.area2_io_pad\[4\]/TIE_LO_ESD
+ mprj_io_slow_sel[22] mprj_io_vtrip_sel[22] mprj_io_holdover[22] mprj_io_analog_en[22]
+ mprj_io_analog_sel[22] vccd vssio mprj_io_analog_pol[22] mprj_io_out[22] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_611 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_600 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_699 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_622 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_633 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_644 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_655 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_666 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_688 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_496 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_485 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_29 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
Xbus_tie_18 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_430 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_452 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_463 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_474 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_260 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_282 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_293 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[4\] mprj_pads.area1_io_pad\[4\]/IN_H mprj_pads.area1_io_pad\[4\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[4\]/PAD_A_ESD_1_H
+ mprj_io[4] mprj_io_dm[14] mprj_io_dm[13] mprj_io_dm[12] mprj_io_hldh_n[4] mprj_io_in[4]
+ mprj_io_inp_dis[4] mprj_io_ib_mode_sel[4] mprj_io_enh[4] porb_h mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD
+ mprj_io_oeb[4] mprj_pads.area1_io_pad\[4\]/TIE_HI_ESD mprj_pads.area1_io_pad\[4\]/TIE_LO_ESD
+ mprj_io_slow_sel[4] mprj_io_vtrip_sel[4] mprj_io_holdover[4] mprj_io_analog_en[4]
+ mprj_io_analog_sel[4] vccd vssio mprj_io_analog_pol[4] mprj_io_out[4] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_815 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_804 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_612 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_623 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_634 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_645 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_656 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_667 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_678 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_689 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_90 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_497 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_486 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_475 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xbus_tie_19 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda gpio_pad/VDDIO_Q vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q vddio vccd sky130_ef_io__connect_vcchib_vccd_and_vswitch_vddio_slice_20um
XFILLER_420 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_442 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_453 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_464 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_283 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_294 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_816 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_805 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_602 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_613 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_624 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_635 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_646 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_657 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_679 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_91 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_80 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_498 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_487 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_476 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_432 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_443 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_454 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_465 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_262 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_240 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_273 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmprj_pads.area2_io_pad\[12\] mprj_pads.area2_io_pad\[12\]/IN_H mprj_pads.area2_io_pad\[12\]/PAD_A_NOESD_H
+ mprj_analog_io[23] mprj_pads.area2_io_pad\[12\]/PAD_A_ESD_1_H mprj_io[30] mprj_io_dm[92]
+ mprj_io_dm[91] mprj_io_dm[90] mprj_io_hldh_n[30] mprj_io_in[30] mprj_io_inp_dis[30]
+ mprj_io_ib_mode_sel[30] mprj_io_enh[30] porb_h mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD
+ mprj_io_oeb[30] mprj_pads.area2_io_pad\[12\]/TIE_HI_ESD mprj_pads.area2_io_pad\[12\]/TIE_LO_ESD
+ mprj_io_slow_sel[30] mprj_io_vtrip_sel[30] mprj_io_holdover[30] mprj_io_analog_en[30]
+ mprj_io_analog_sel[30] vccd vssio mprj_io_analog_pol[30] mprj_io_out[30] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_817 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_806 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xmgmt_vssio_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssio_pad2 vssa2
+ vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__vssio_hvc_clamped_pad
XFILLER_603 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_614 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_625 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_636 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_647 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_658 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_669 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_92 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_81 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area2_io_pad\[2\] mprj_pads.area2_io_pad\[2\]/IN_H mprj_pads.area2_io_pad\[2\]/PAD_A_NOESD_H
+ mprj_analog_io[13] mprj_pads.area2_io_pad\[2\]/PAD_A_ESD_1_H mprj_io[20] mprj_io_dm[62]
+ mprj_io_dm[61] mprj_io_dm[60] mprj_io_hldh_n[20] mprj_io_in[20] mprj_io_inp_dis[20]
+ mprj_io_ib_mode_sel[20] mprj_io_enh[20] porb_h mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD
+ mprj_io_oeb[20] mprj_pads.area2_io_pad\[2\]/TIE_HI_ESD mprj_pads.area2_io_pad\[2\]/TIE_LO_ESD
+ mprj_io_slow_sel[20] mprj_io_vtrip_sel[20] mprj_io_holdover[20] mprj_io_analog_en[20]
+ mprj_io_analog_sel[20] vccd vssio mprj_io_analog_pol[20] mprj_io_out[20] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_499 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_488 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_477 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_422 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_433 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_444 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_455 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_466 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_263 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_241 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_230 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_274 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_296 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_818 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_807 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser2_vssa_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[2\] mprj_pads.area1_io_pad\[2\]/IN_H mprj_pads.area1_io_pad\[2\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[2\]/PAD_A_ESD_1_H
+ mprj_io[2] mprj_io_dm[8] mprj_io_dm[7] mprj_io_dm[6] mprj_io_hldh_n[2] mprj_io_in[2]
+ mprj_io_inp_dis[2] mprj_io_ib_mode_sel[2] mprj_io_enh[2] porb_h mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD
+ mprj_io_oeb[2] mprj_pads.area1_io_pad\[2\]/TIE_HI_ESD mprj_pads.area1_io_pad\[2\]/TIE_LO_ESD
+ mprj_io_slow_sel[2] mprj_io_vtrip_sel[2] mprj_io_holdover[2] mprj_io_analog_en[2]
+ mprj_io_analog_sel[2] vccd vssio mprj_io_analog_pol[2] mprj_io_out[2] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_5 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_604 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_615 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_626 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_637 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_648 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_93 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_82 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_71 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_60 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_489 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_478 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_401 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_412 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_423 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_434 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_445 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_456 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_467 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_264 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_242 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_231 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_275 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_297 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_808 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_6 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_605 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_616 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_627 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_638 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_94 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_72 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_61 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_50 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_479 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_402 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_413 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_424 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_435 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_446 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_457 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_468 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_265 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_243 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_232 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_276 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_298 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area1_io_pad\[17\] mprj_pads.area1_io_pad\[17\]/IN_H mprj_pads.area1_io_pad\[17\]/PAD_A_NOESD_H
+ mprj_analog_io[10] mprj_pads.area1_io_pad\[17\]/PAD_A_ESD_1_H mprj_io[17] mprj_io_dm[53]
+ mprj_io_dm[52] mprj_io_dm[51] mprj_io_hldh_n[17] mprj_io_in[17] mprj_io_inp_dis[17]
+ mprj_io_ib_mode_sel[17] mprj_io_enh[17] porb_h mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD
+ mprj_io_oeb[17] mprj_pads.area1_io_pad\[17\]/TIE_HI_ESD mprj_pads.area1_io_pad\[17\]/TIE_LO_ESD
+ mprj_io_slow_sel[17] mprj_io_vtrip_sel[17] mprj_io_holdover[17] mprj_io_analog_en[17]
+ mprj_io_analog_sel[17] vccd vssio mprj_io_analog_pol[17] mprj_io_out[17] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xuser1_vdda_hvclamp_pad\[1\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda1_pad2 vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xmprj_pads.area2_io_pad\[10\] mprj_pads.area2_io_pad\[10\]/IN_H mprj_pads.area2_io_pad\[10\]/PAD_A_NOESD_H
+ mprj_analog_io[21] mprj_pads.area2_io_pad\[10\]/PAD_A_ESD_1_H mprj_io[28] mprj_io_dm[86]
+ mprj_io_dm[85] mprj_io_dm[84] mprj_io_hldh_n[28] mprj_io_in[28] mprj_io_inp_dis[28]
+ mprj_io_ib_mode_sel[28] mprj_io_enh[28] porb_h mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD
+ mprj_io_oeb[28] mprj_pads.area2_io_pad\[10\]/TIE_HI_ESD mprj_pads.area2_io_pad\[10\]/TIE_LO_ESD
+ mprj_io_slow_sel[28] mprj_io_vtrip_sel[28] mprj_io_holdover[28] mprj_io_analog_en[28]
+ mprj_io_analog_sel[28] vccd vssio mprj_io_analog_pol[28] mprj_io_out[28] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_7 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_606 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_617 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_628 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_639 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_95 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_84 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_73 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_62 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_51 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_40 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_403 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_414 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_425 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_436 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_447 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_458 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_469 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area2_io_pad\[0\] mprj_pads.area2_io_pad\[0\]/IN_H mprj_pads.area2_io_pad\[0\]/PAD_A_NOESD_H
+ mprj_analog_io[11] mprj_pads.area2_io_pad\[0\]/PAD_A_ESD_1_H mprj_io[18] mprj_io_dm[56]
+ mprj_io_dm[55] mprj_io_dm[54] mprj_io_hldh_n[18] mprj_io_in[18] mprj_io_inp_dis[18]
+ mprj_io_ib_mode_sel[18] mprj_io_enh[18] porb_h mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD
+ mprj_io_oeb[18] mprj_pads.area2_io_pad\[0\]/TIE_HI_ESD mprj_pads.area2_io_pad\[0\]/TIE_LO_ESD
+ mprj_io_slow_sel[18] mprj_io_vtrip_sel[18] mprj_io_holdover[18] mprj_io_analog_en[18]
+ mprj_io_analog_sel[18] vccd vssio mprj_io_analog_pol[18] mprj_io_out[18] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_266 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_222 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_211 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_277 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_299 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_8 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_607 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_618 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_629 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_85 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_74 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_63 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_52 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_41 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[0\] mprj_pads.area1_io_pad\[0\]/IN_H mprj_pads.area1_io_pad\[0\]/PAD_A_NOESD_H
+ mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_0_H mprj_pads.area1_io_pad\[0\]/PAD_A_ESD_1_H
+ mprj_io[0] mprj_io_dm[2] mprj_io_dm[1] mprj_io_dm[0] mprj_io_hldh_n[0] mprj_io_in[0]
+ mprj_io_inp_dis[0] mprj_io_ib_mode_sel[0] mprj_io_enh[0] porb_h mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD
+ mprj_io_oeb[0] mprj_pads.area1_io_pad\[0\]/TIE_HI_ESD mprj_pads.area1_io_pad\[0\]/TIE_LO_ESD
+ mprj_io_slow_sel[0] mprj_io_vtrip_sel[0] mprj_io_holdover[0] mprj_io_analog_en[0]
+ mprj_io_analog_sel[0] vccd vssio mprj_io_analog_pol[0] mprj_io_out[0] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_404 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_415 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_426 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_437 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_448 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_459 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_256 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_245 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_223 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_212 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_9 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_608 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_619 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_97 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_86 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_75 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_64 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_53 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_42 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_31 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_20 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_405 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_416 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_427 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_438 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_449 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_257 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_246 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_224 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_213 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_279 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_791 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_780 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmgmt_vdda_hvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vdda_pad vssa vdda vddio
+ gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__vdda_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[15\] mprj_pads.area1_io_pad\[15\]/IN_H mprj_pads.area1_io_pad\[15\]/PAD_A_NOESD_H
+ mprj_analog_io[8] mprj_pads.area1_io_pad\[15\]/PAD_A_ESD_1_H mprj_io[15] mprj_io_dm[47]
+ mprj_io_dm[46] mprj_io_dm[45] mprj_io_hldh_n[15] mprj_io_in[15] mprj_io_inp_dis[15]
+ mprj_io_ib_mode_sel[15] mprj_io_enh[15] porb_h mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD
+ mprj_io_oeb[15] mprj_pads.area1_io_pad\[15\]/TIE_HI_ESD mprj_pads.area1_io_pad\[15\]/TIE_LO_ESD
+ mprj_io_slow_sel[15] mprj_io_vtrip_sel[15] mprj_io_holdover[15] mprj_io_analog_en[15]
+ mprj_io_analog_sel[15] vccd vssio mprj_io_analog_pol[15] mprj_io_out[15] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_609 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_98 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_87 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_76 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_65 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_54 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_32 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_21 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_10 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_406 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_417 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_428 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_439 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_258 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_247 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_225 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_214 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_792 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_770 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
Xmprj_pads.area2_io_pad\[19\] mprj_pads.area2_io_pad\[19\]/IN_H mprj_pads.area2_io_pad\[19\]/PAD_A_NOESD_H
+ mprj_analog_io[30] mprj_pads.area2_io_pad\[19\]/PAD_A_ESD_1_H mprj_io[37] mprj_io_dm[113]
+ mprj_io_dm[112] mprj_io_dm[111] mprj_io_hldh_n[37] mprj_io_in[37] mprj_io_inp_dis[37]
+ mprj_io_ib_mode_sel[37] mprj_io_enh[37] porb_h mprj_pads.area2_io_pad\[19\]/TIE_LO_ESD
+ mprj_io_oeb[37] mprj_pads.area2_io_pad\[19\]/TIE_HI_ESD mprj_pads.area2_io_pad\[19\]/TIE_LO_ESD
+ mprj_io_slow_sel[37] mprj_io_vtrip_sel[37] mprj_io_holdover[37] mprj_io_analog_en[37]
+ mprj_io_analog_sel[37] vccd vssio mprj_io_analog_pol[37] mprj_io_out[37] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xmprj_pads.area2_io_pad\[9\] mprj_pads.area2_io_pad\[9\]/IN_H mprj_pads.area2_io_pad\[9\]/PAD_A_NOESD_H
+ mprj_analog_io[20] mprj_pads.area2_io_pad\[9\]/PAD_A_ESD_1_H mprj_io[27] mprj_io_dm[83]
+ mprj_io_dm[82] mprj_io_dm[81] mprj_io_hldh_n[27] mprj_io_in[27] mprj_io_inp_dis[27]
+ mprj_io_ib_mode_sel[27] mprj_io_enh[27] porb_h mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD
+ mprj_io_oeb[27] mprj_pads.area2_io_pad\[9\]/TIE_HI_ESD mprj_pads.area2_io_pad\[9\]/TIE_LO_ESD
+ mprj_io_slow_sel[27] mprj_io_vtrip_sel[27] mprj_io_holdover[27] mprj_io_analog_en[27]
+ mprj_io_analog_sel[27] vccd vssio mprj_io_analog_pol[27] mprj_io_out[27] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
Xflash_io0_pad flash_io0_pad/IN_H flash_io0_pad/PAD_A_NOESD_H flash_io0_pad/PAD_A_ESD_0_H
+ flash_io0_pad/PAD_A_ESD_1_H flash_io0 flash_io0_ieb_core flash_io0_ieb_core flash_io0_oeb_core
+ vddio flash_io0_di_core flash_io0_ieb_core vssd porb_h porb_h flash_io0_pad/TIE_LO_ESD
+ flash_io0_oeb_core flash_io0_pad/TIE_HI_ESD flash_io0_pad/TIE_LO_ESD vssd vssd vssd
+ vssd vssd vccd vssa vssd flash_io0_do_core gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B
+ vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_99 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_88 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_77 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_66 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_55 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_44 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_33 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_22 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_11 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_407 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_418 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_429 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_259 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_248 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_226 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_215 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_793 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_782 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_760 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_590 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmgmt_corner\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
Xuser1_vssa_hvclamp_pad\[0\] gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1_pad vssa1
+ vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__vssa_hvc_clamped_pad
Xmprj_pads.area1_io_pad\[9\] mprj_pads.area1_io_pad\[9\]/IN_H mprj_pads.area1_io_pad\[9\]/PAD_A_NOESD_H
+ mprj_analog_io[2] mprj_pads.area1_io_pad\[9\]/PAD_A_ESD_1_H mprj_io[9] mprj_io_dm[29]
+ mprj_io_dm[28] mprj_io_dm[27] mprj_io_hldh_n[9] mprj_io_in[9] mprj_io_inp_dis[9]
+ mprj_io_ib_mode_sel[9] mprj_io_enh[9] porb_h mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD
+ mprj_io_oeb[9] mprj_pads.area1_io_pad\[9\]/TIE_HI_ESD mprj_pads.area1_io_pad\[9\]/TIE_LO_ESD
+ mprj_io_slow_sel[9] mprj_io_vtrip_sel[9] mprj_io_holdover[9] mprj_io_analog_en[9]
+ mprj_io_analog_sel[9] vccd vssio mprj_io_analog_pol[9] mprj_io_out[9] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_89 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_78 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_67 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_45 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_34 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_23 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_12 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xflash_clk_pad flash_clk_pad/IN_H flash_clk_pad/PAD_A_NOESD_H flash_clk_pad/PAD_A_ESD_0_H
+ flash_clk_pad/PAD_A_ESD_1_H flash_clk vccd vccd vssd vddio flash_clk_pad/IN flash_clk_ieb_core
+ vssd porb_h porb_h flash_clk_pad/TIE_LO_ESD flash_clk_oeb_core flash_clk_pad/TIE_HI_ESD
+ flash_clk_pad/TIE_LO_ESD vssd vssd vssd vssd vssd vccd vssa vssd flash_clk_core
+ gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q vccd vddio
+ vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_408 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_419 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_249 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_205 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_794 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_783 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_772 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_761 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_750 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
Xuser1_vccd_lvclamp_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vccd1_pad vssa1 vdda1
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__vccd_lvc_clamped2_pad
XFILLER_580 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xmprj_pads.area1_io_pad\[13\] mprj_pads.area1_io_pad\[13\]/IN_H mprj_pads.area1_io_pad\[13\]/PAD_A_NOESD_H
+ mprj_analog_io[6] mprj_pads.area1_io_pad\[13\]/PAD_A_ESD_1_H mprj_io[13] mprj_io_dm[41]
+ mprj_io_dm[40] mprj_io_dm[39] mprj_io_hldh_n[13] mprj_io_in[13] mprj_io_inp_dis[13]
+ mprj_io_ib_mode_sel[13] mprj_io_enh[13] porb_h mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD
+ mprj_io_oeb[13] mprj_pads.area1_io_pad\[13\]/TIE_HI_ESD mprj_pads.area1_io_pad\[13\]/TIE_LO_ESD
+ mprj_io_slow_sel[13] mprj_io_vtrip_sel[13] mprj_io_holdover[13] mprj_io_analog_en[13]
+ mprj_io_analog_sel[13] vccd vssio mprj_io_analog_pol[13] mprj_io_out[13] gpio_pad/AMUXBUS_A
+ gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q vccd vddio vccd1 vssio vssd1
+ gpio_pad/VSSIO_Q sky130_ef_io__gpiov2_pad_wrapped
XFILLER_79 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_68 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
XFILLER_57 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_46 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_35 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_24 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_13 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa2 vdda2 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
Xuser1_corner gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__corner_pad
XFILLER_409 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_1um
Xuser2_vssd_lvclmap_pad gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssd2_pad vssa2 vdda2
+ vddio gpio_pad/VDDIO_Q vccd vddio vccd2 vssio vssd2 gpio_pad/VSSIO_Q sky130_ef_io__vssd_lvc_clamped2_pad
XFILLER_239 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_228 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_206 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa vdda vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd vssio vssd gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_10um
XFILLER_795 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_784 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_773 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
XFILLER_751 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_5um
XFILLER_740 gpio_pad/AMUXBUS_A gpio_pad/AMUXBUS_B vssa1 vdda1 vddio gpio_pad/VDDIO_Q
+ vccd vddio vccd1 vssio vssd1 gpio_pad/VSSIO_Q sky130_ef_io__com_bus_slice_20um
.ends

* Black-box entry subcircuit for mgmt_core abstract view
.subckt mgmt_core clock core_clk core_rstn flash_clk flash_clk_ieb flash_clk_oeb flash_csb
+ flash_csb_ieb flash_csb_oeb flash_io0_di flash_io0_do flash_io0_ieb flash_io0_oeb
+ flash_io1_di flash_io1_do flash_io1_ieb flash_io1_oeb gpio_in_pad gpio_inenb_pad
+ gpio_mode0_pad gpio_mode1_pad gpio_out_pad gpio_outenb_pad jtag_out jtag_outenb
+ la_input[0] la_input[100] la_input[101] la_input[102] la_input[103] la_input[104]
+ la_input[105] la_input[106] la_input[107] la_input[108] la_input[109] la_input[10]
+ la_input[110] la_input[111] la_input[112] la_input[113] la_input[114] la_input[115]
+ la_input[116] la_input[117] la_input[118] la_input[119] la_input[11] la_input[120]
+ la_input[121] la_input[122] la_input[123] la_input[124] la_input[125] la_input[126]
+ la_input[127] la_input[12] la_input[13] la_input[14] la_input[15] la_input[16] la_input[17]
+ la_input[18] la_input[19] la_input[1] la_input[20] la_input[21] la_input[22] la_input[23]
+ la_input[24] la_input[25] la_input[26] la_input[27] la_input[28] la_input[29] la_input[2]
+ la_input[30] la_input[31] la_input[32] la_input[33] la_input[34] la_input[35] la_input[36]
+ la_input[37] la_input[38] la_input[39] la_input[3] la_input[40] la_input[41] la_input[42]
+ la_input[43] la_input[44] la_input[45] la_input[46] la_input[47] la_input[48] la_input[49]
+ la_input[4] la_input[50] la_input[51] la_input[52] la_input[53] la_input[54] la_input[55]
+ la_input[56] la_input[57] la_input[58] la_input[59] la_input[5] la_input[60] la_input[61]
+ la_input[62] la_input[63] la_input[64] la_input[65] la_input[66] la_input[67] la_input[68]
+ la_input[69] la_input[6] la_input[70] la_input[71] la_input[72] la_input[73] la_input[74]
+ la_input[75] la_input[76] la_input[77] la_input[78] la_input[79] la_input[7] la_input[80]
+ la_input[81] la_input[82] la_input[83] la_input[84] la_input[85] la_input[86] la_input[87]
+ la_input[88] la_input[89] la_input[8] la_input[90] la_input[91] la_input[92] la_input[93]
+ la_input[94] la_input[95] la_input[96] la_input[97] la_input[98] la_input[99] la_input[9]
+ la_oen[0] la_oen[100] la_oen[101] la_oen[102] la_oen[103] la_oen[104] la_oen[105]
+ la_oen[106] la_oen[107] la_oen[108] la_oen[109] la_oen[10] la_oen[110] la_oen[111]
+ la_oen[112] la_oen[113] la_oen[114] la_oen[115] la_oen[116] la_oen[117] la_oen[118]
+ la_oen[119] la_oen[11] la_oen[120] la_oen[121] la_oen[122] la_oen[123] la_oen[124]
+ la_oen[125] la_oen[126] la_oen[127] la_oen[12] la_oen[13] la_oen[14] la_oen[15]
+ la_oen[16] la_oen[17] la_oen[18] la_oen[19] la_oen[1] la_oen[20] la_oen[21] la_oen[22]
+ la_oen[23] la_oen[24] la_oen[25] la_oen[26] la_oen[27] la_oen[28] la_oen[29] la_oen[2]
+ la_oen[30] la_oen[31] la_oen[32] la_oen[33] la_oen[34] la_oen[35] la_oen[36] la_oen[37]
+ la_oen[38] la_oen[39] la_oen[3] la_oen[40] la_oen[41] la_oen[42] la_oen[43] la_oen[44]
+ la_oen[45] la_oen[46] la_oen[47] la_oen[48] la_oen[49] la_oen[4] la_oen[50] la_oen[51]
+ la_oen[52] la_oen[53] la_oen[54] la_oen[55] la_oen[56] la_oen[57] la_oen[58] la_oen[59]
+ la_oen[5] la_oen[60] la_oen[61] la_oen[62] la_oen[63] la_oen[64] la_oen[65] la_oen[66]
+ la_oen[67] la_oen[68] la_oen[69] la_oen[6] la_oen[70] la_oen[71] la_oen[72] la_oen[73]
+ la_oen[74] la_oen[75] la_oen[76] la_oen[77] la_oen[78] la_oen[79] la_oen[7] la_oen[80]
+ la_oen[81] la_oen[82] la_oen[83] la_oen[84] la_oen[85] la_oen[86] la_oen[87] la_oen[88]
+ la_oen[89] la_oen[8] la_oen[90] la_oen[91] la_oen[92] la_oen[93] la_oen[94] la_oen[95]
+ la_oen[96] la_oen[97] la_oen[98] la_oen[99] la_oen[9] la_output[0] la_output[100]
+ la_output[101] la_output[102] la_output[103] la_output[104] la_output[105] la_output[106]
+ la_output[107] la_output[108] la_output[109] la_output[10] la_output[110] la_output[111]
+ la_output[112] la_output[113] la_output[114] la_output[115] la_output[116] la_output[117]
+ la_output[118] la_output[119] la_output[11] la_output[120] la_output[121] la_output[122]
+ la_output[123] la_output[124] la_output[125] la_output[126] la_output[127] la_output[12]
+ la_output[13] la_output[14] la_output[15] la_output[16] la_output[17] la_output[18]
+ la_output[19] la_output[1] la_output[20] la_output[21] la_output[22] la_output[23]
+ la_output[24] la_output[25] la_output[26] la_output[27] la_output[28] la_output[29]
+ la_output[2] la_output[30] la_output[31] la_output[32] la_output[33] la_output[34]
+ la_output[35] la_output[36] la_output[37] la_output[38] la_output[39] la_output[3]
+ la_output[40] la_output[41] la_output[42] la_output[43] la_output[44] la_output[45]
+ la_output[46] la_output[47] la_output[48] la_output[49] la_output[4] la_output[50]
+ la_output[51] la_output[52] la_output[53] la_output[54] la_output[55] la_output[56]
+ la_output[57] la_output[58] la_output[59] la_output[5] la_output[60] la_output[61]
+ la_output[62] la_output[63] la_output[64] la_output[65] la_output[66] la_output[67]
+ la_output[68] la_output[69] la_output[6] la_output[70] la_output[71] la_output[72]
+ la_output[73] la_output[74] la_output[75] la_output[76] la_output[77] la_output[78]
+ la_output[79] la_output[7] la_output[80] la_output[81] la_output[82] la_output[83]
+ la_output[84] la_output[85] la_output[86] la_output[87] la_output[88] la_output[89]
+ la_output[8] la_output[90] la_output[91] la_output[92] la_output[93] la_output[94]
+ la_output[95] la_output[96] la_output[97] la_output[98] la_output[99] la_output[9]
+ mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13] mask_rev[14] mask_rev[15]
+ mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1] mask_rev[20] mask_rev[21]
+ mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26] mask_rev[27] mask_rev[28]
+ mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3] mask_rev[4] mask_rev[5]
+ mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] mgmt_addr[0] mgmt_addr[1] mgmt_addr[2]
+ mgmt_addr[3] mgmt_addr[4] mgmt_addr[5] mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0]
+ mgmt_addr_ro[1] mgmt_addr_ro[2] mgmt_addr_ro[3] mgmt_addr_ro[4] mgmt_addr_ro[5]
+ mgmt_addr_ro[6] mgmt_addr_ro[7] mgmt_ena[0] mgmt_ena[1] mgmt_ena_ro mgmt_in_data[0]
+ mgmt_in_data[10] mgmt_in_data[11] mgmt_in_data[12] mgmt_in_data[13] mgmt_in_data[14]
+ mgmt_in_data[15] mgmt_in_data[16] mgmt_in_data[17] mgmt_in_data[18] mgmt_in_data[19]
+ mgmt_in_data[1] mgmt_in_data[20] mgmt_in_data[21] mgmt_in_data[22] mgmt_in_data[23]
+ mgmt_in_data[24] mgmt_in_data[25] mgmt_in_data[26] mgmt_in_data[27] mgmt_in_data[28]
+ mgmt_in_data[29] mgmt_in_data[2] mgmt_in_data[30] mgmt_in_data[31] mgmt_in_data[32]
+ mgmt_in_data[33] mgmt_in_data[34] mgmt_in_data[35] mgmt_in_data[36] mgmt_in_data[37]
+ mgmt_in_data[3] mgmt_in_data[4] mgmt_in_data[5] mgmt_in_data[6] mgmt_in_data[7]
+ mgmt_in_data[8] mgmt_in_data[9] mgmt_out_data[0] mgmt_out_data[10] mgmt_out_data[11]
+ mgmt_out_data[12] mgmt_out_data[13] mgmt_out_data[14] mgmt_out_data[15] mgmt_out_data[16]
+ mgmt_out_data[17] mgmt_out_data[18] mgmt_out_data[19] mgmt_out_data[1] mgmt_out_data[20]
+ mgmt_out_data[21] mgmt_out_data[22] mgmt_out_data[23] mgmt_out_data[24] mgmt_out_data[25]
+ mgmt_out_data[26] mgmt_out_data[27] mgmt_out_data[28] mgmt_out_data[29] mgmt_out_data[2]
+ mgmt_out_data[30] mgmt_out_data[31] mgmt_out_data[32] mgmt_out_data[33] mgmt_out_data[34]
+ mgmt_out_data[35] mgmt_out_data[36] mgmt_out_data[37] mgmt_out_data[3] mgmt_out_data[4]
+ mgmt_out_data[5] mgmt_out_data[6] mgmt_out_data[7] mgmt_out_data[8] mgmt_out_data[9]
+ mgmt_rdata[0] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12] mgmt_rdata[13] mgmt_rdata[14]
+ mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18] mgmt_rdata[19] mgmt_rdata[1]
+ mgmt_rdata[20] mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23] mgmt_rdata[24] mgmt_rdata[25]
+ mgmt_rdata[26] mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29] mgmt_rdata[2] mgmt_rdata[30]
+ mgmt_rdata[31] mgmt_rdata[32] mgmt_rdata[33] mgmt_rdata[34] mgmt_rdata[35] mgmt_rdata[36]
+ mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39] mgmt_rdata[3] mgmt_rdata[40] mgmt_rdata[41]
+ mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45] mgmt_rdata[46] mgmt_rdata[47]
+ mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[4] mgmt_rdata[50] mgmt_rdata[51] mgmt_rdata[52]
+ mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56] mgmt_rdata[57] mgmt_rdata[58]
+ mgmt_rdata[59] mgmt_rdata[5] mgmt_rdata[60] mgmt_rdata[61] mgmt_rdata[62] mgmt_rdata[63]
+ mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8] mgmt_rdata[9] mgmt_rdata_ro[0] mgmt_rdata_ro[10]
+ mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13] mgmt_rdata_ro[14] mgmt_rdata_ro[15]
+ mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18] mgmt_rdata_ro[19] mgmt_rdata_ro[1]
+ mgmt_rdata_ro[20] mgmt_rdata_ro[21] mgmt_rdata_ro[22] mgmt_rdata_ro[23] mgmt_rdata_ro[24]
+ mgmt_rdata_ro[25] mgmt_rdata_ro[26] mgmt_rdata_ro[27] mgmt_rdata_ro[28] mgmt_rdata_ro[29]
+ mgmt_rdata_ro[2] mgmt_rdata_ro[30] mgmt_rdata_ro[31] mgmt_rdata_ro[3] mgmt_rdata_ro[4]
+ mgmt_rdata_ro[5] mgmt_rdata_ro[6] mgmt_rdata_ro[7] mgmt_rdata_ro[8] mgmt_rdata_ro[9]
+ mgmt_wdata[0] mgmt_wdata[10] mgmt_wdata[11] mgmt_wdata[12] mgmt_wdata[13] mgmt_wdata[14]
+ mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17] mgmt_wdata[18] mgmt_wdata[19] mgmt_wdata[1]
+ mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23] mgmt_wdata[24] mgmt_wdata[25]
+ mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29] mgmt_wdata[2] mgmt_wdata[30]
+ mgmt_wdata[31] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5] mgmt_wdata[6] mgmt_wdata[7]
+ mgmt_wdata[8] mgmt_wdata[9] mgmt_wen[0] mgmt_wen[1] mgmt_wen_mask[0] mgmt_wen_mask[1]
+ mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_wen_mask[4] mgmt_wen_mask[5] mgmt_wen_mask[6]
+ mgmt_wen_mask[7] mprj2_vcc_pwrgood mprj2_vdd_pwrgood mprj_ack_i mprj_adr_o[0] mprj_adr_o[10]
+ mprj_adr_o[11] mprj_adr_o[12] mprj_adr_o[13] mprj_adr_o[14] mprj_adr_o[15] mprj_adr_o[16]
+ mprj_adr_o[17] mprj_adr_o[18] mprj_adr_o[19] mprj_adr_o[1] mprj_adr_o[20] mprj_adr_o[21]
+ mprj_adr_o[22] mprj_adr_o[23] mprj_adr_o[24] mprj_adr_o[25] mprj_adr_o[26] mprj_adr_o[27]
+ mprj_adr_o[28] mprj_adr_o[29] mprj_adr_o[2] mprj_adr_o[30] mprj_adr_o[31] mprj_adr_o[3]
+ mprj_adr_o[4] mprj_adr_o[5] mprj_adr_o[6] mprj_adr_o[7] mprj_adr_o[8] mprj_adr_o[9]
+ mprj_cyc_o mprj_dat_i[0] mprj_dat_i[10] mprj_dat_i[11] mprj_dat_i[12] mprj_dat_i[13]
+ mprj_dat_i[14] mprj_dat_i[15] mprj_dat_i[16] mprj_dat_i[17] mprj_dat_i[18] mprj_dat_i[19]
+ mprj_dat_i[1] mprj_dat_i[20] mprj_dat_i[21] mprj_dat_i[22] mprj_dat_i[23] mprj_dat_i[24]
+ mprj_dat_i[25] mprj_dat_i[26] mprj_dat_i[27] mprj_dat_i[28] mprj_dat_i[29] mprj_dat_i[2]
+ mprj_dat_i[30] mprj_dat_i[31] mprj_dat_i[3] mprj_dat_i[4] mprj_dat_i[5] mprj_dat_i[6]
+ mprj_dat_i[7] mprj_dat_i[8] mprj_dat_i[9] mprj_dat_o[0] mprj_dat_o[10] mprj_dat_o[11]
+ mprj_dat_o[12] mprj_dat_o[13] mprj_dat_o[14] mprj_dat_o[15] mprj_dat_o[16] mprj_dat_o[17]
+ mprj_dat_o[18] mprj_dat_o[19] mprj_dat_o[1] mprj_dat_o[20] mprj_dat_o[21] mprj_dat_o[22]
+ mprj_dat_o[23] mprj_dat_o[24] mprj_dat_o[25] mprj_dat_o[26] mprj_dat_o[27] mprj_dat_o[28]
+ mprj_dat_o[29] mprj_dat_o[2] mprj_dat_o[30] mprj_dat_o[31] mprj_dat_o[3] mprj_dat_o[4]
+ mprj_dat_o[5] mprj_dat_o[6] mprj_dat_o[7] mprj_dat_o[8] mprj_dat_o[9] mprj_io_loader_clock
+ mprj_io_loader_data mprj_io_loader_resetn mprj_sel_o[0] mprj_sel_o[1] mprj_sel_o[2]
+ mprj_sel_o[3] mprj_stb_o mprj_vcc_pwrgood mprj_vdd_pwrgood mprj_we_o porb pwr_ctrl_out[0]
+ pwr_ctrl_out[1] pwr_ctrl_out[2] pwr_ctrl_out[3] resetb sdo_out sdo_outenb user_clk
+ VPWR VGND
.ends

* Black-box entry subcircuit for simple_por abstract view
.subckt simple_por vdd3v3 vdd1v8 vss porb_h por_l porb_l
.ends

* Black-box entry subcircuit for user_id_programming abstract view
.subckt user_id_programming mask_rev[0] mask_rev[10] mask_rev[11] mask_rev[12] mask_rev[13]
+ mask_rev[14] mask_rev[15] mask_rev[16] mask_rev[17] mask_rev[18] mask_rev[19] mask_rev[1]
+ mask_rev[20] mask_rev[21] mask_rev[22] mask_rev[23] mask_rev[24] mask_rev[25] mask_rev[26]
+ mask_rev[27] mask_rev[28] mask_rev[29] mask_rev[2] mask_rev[30] mask_rev[31] mask_rev[3]
+ mask_rev[4] mask_rev[5] mask_rev[6] mask_rev[7] mask_rev[8] mask_rev[9] VPWR VGND
.ends

* Black-box entry subcircuit for mgmt_protect abstract view
.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_oen_core[0] la_oen_core[100] la_oen_core[101] la_oen_core[102]
+ la_oen_core[103] la_oen_core[104] la_oen_core[105] la_oen_core[106] la_oen_core[107]
+ la_oen_core[108] la_oen_core[109] la_oen_core[10] la_oen_core[110] la_oen_core[111]
+ la_oen_core[112] la_oen_core[113] la_oen_core[114] la_oen_core[115] la_oen_core[116]
+ la_oen_core[117] la_oen_core[118] la_oen_core[119] la_oen_core[11] la_oen_core[120]
+ la_oen_core[121] la_oen_core[122] la_oen_core[123] la_oen_core[124] la_oen_core[125]
+ la_oen_core[126] la_oen_core[127] la_oen_core[12] la_oen_core[13] la_oen_core[14]
+ la_oen_core[15] la_oen_core[16] la_oen_core[17] la_oen_core[18] la_oen_core[19]
+ la_oen_core[1] la_oen_core[20] la_oen_core[21] la_oen_core[22] la_oen_core[23] la_oen_core[24]
+ la_oen_core[25] la_oen_core[26] la_oen_core[27] la_oen_core[28] la_oen_core[29]
+ la_oen_core[2] la_oen_core[30] la_oen_core[31] la_oen_core[32] la_oen_core[33] la_oen_core[34]
+ la_oen_core[35] la_oen_core[36] la_oen_core[37] la_oen_core[38] la_oen_core[39]
+ la_oen_core[3] la_oen_core[40] la_oen_core[41] la_oen_core[42] la_oen_core[43] la_oen_core[44]
+ la_oen_core[45] la_oen_core[46] la_oen_core[47] la_oen_core[48] la_oen_core[49]
+ la_oen_core[4] la_oen_core[50] la_oen_core[51] la_oen_core[52] la_oen_core[53] la_oen_core[54]
+ la_oen_core[55] la_oen_core[56] la_oen_core[57] la_oen_core[58] la_oen_core[59]
+ la_oen_core[5] la_oen_core[60] la_oen_core[61] la_oen_core[62] la_oen_core[63] la_oen_core[64]
+ la_oen_core[65] la_oen_core[66] la_oen_core[67] la_oen_core[68] la_oen_core[69]
+ la_oen_core[6] la_oen_core[70] la_oen_core[71] la_oen_core[72] la_oen_core[73] la_oen_core[74]
+ la_oen_core[75] la_oen_core[76] la_oen_core[77] la_oen_core[78] la_oen_core[79]
+ la_oen_core[7] la_oen_core[80] la_oen_core[81] la_oen_core[82] la_oen_core[83] la_oen_core[84]
+ la_oen_core[85] la_oen_core[86] la_oen_core[87] la_oen_core[88] la_oen_core[89]
+ la_oen_core[8] la_oen_core[90] la_oen_core[91] la_oen_core[92] la_oen_core[93] la_oen_core[94]
+ la_oen_core[95] la_oen_core[96] la_oen_core[97] la_oen_core[98] la_oen_core[99]
+ la_oen_core[9] la_oen_mprj[0] la_oen_mprj[100] la_oen_mprj[101] la_oen_mprj[102]
+ la_oen_mprj[103] la_oen_mprj[104] la_oen_mprj[105] la_oen_mprj[106] la_oen_mprj[107]
+ la_oen_mprj[108] la_oen_mprj[109] la_oen_mprj[10] la_oen_mprj[110] la_oen_mprj[111]
+ la_oen_mprj[112] la_oen_mprj[113] la_oen_mprj[114] la_oen_mprj[115] la_oen_mprj[116]
+ la_oen_mprj[117] la_oen_mprj[118] la_oen_mprj[119] la_oen_mprj[11] la_oen_mprj[120]
+ la_oen_mprj[121] la_oen_mprj[122] la_oen_mprj[123] la_oen_mprj[124] la_oen_mprj[125]
+ la_oen_mprj[126] la_oen_mprj[127] la_oen_mprj[12] la_oen_mprj[13] la_oen_mprj[14]
+ la_oen_mprj[15] la_oen_mprj[16] la_oen_mprj[17] la_oen_mprj[18] la_oen_mprj[19]
+ la_oen_mprj[1] la_oen_mprj[20] la_oen_mprj[21] la_oen_mprj[22] la_oen_mprj[23] la_oen_mprj[24]
+ la_oen_mprj[25] la_oen_mprj[26] la_oen_mprj[27] la_oen_mprj[28] la_oen_mprj[29]
+ la_oen_mprj[2] la_oen_mprj[30] la_oen_mprj[31] la_oen_mprj[32] la_oen_mprj[33] la_oen_mprj[34]
+ la_oen_mprj[35] la_oen_mprj[36] la_oen_mprj[37] la_oen_mprj[38] la_oen_mprj[39]
+ la_oen_mprj[3] la_oen_mprj[40] la_oen_mprj[41] la_oen_mprj[42] la_oen_mprj[43] la_oen_mprj[44]
+ la_oen_mprj[45] la_oen_mprj[46] la_oen_mprj[47] la_oen_mprj[48] la_oen_mprj[49]
+ la_oen_mprj[4] la_oen_mprj[50] la_oen_mprj[51] la_oen_mprj[52] la_oen_mprj[53] la_oen_mprj[54]
+ la_oen_mprj[55] la_oen_mprj[56] la_oen_mprj[57] la_oen_mprj[58] la_oen_mprj[59]
+ la_oen_mprj[5] la_oen_mprj[60] la_oen_mprj[61] la_oen_mprj[62] la_oen_mprj[63] la_oen_mprj[64]
+ la_oen_mprj[65] la_oen_mprj[66] la_oen_mprj[67] la_oen_mprj[68] la_oen_mprj[69]
+ la_oen_mprj[6] la_oen_mprj[70] la_oen_mprj[71] la_oen_mprj[72] la_oen_mprj[73] la_oen_mprj[74]
+ la_oen_mprj[75] la_oen_mprj[76] la_oen_mprj[77] la_oen_mprj[78] la_oen_mprj[79]
+ la_oen_mprj[7] la_oen_mprj[80] la_oen_mprj[81] la_oen_mprj[82] la_oen_mprj[83] la_oen_mprj[84]
+ la_oen_mprj[85] la_oen_mprj[86] la_oen_mprj[87] la_oen_mprj[88] la_oen_mprj[89]
+ la_oen_mprj[8] la_oen_mprj[90] la_oen_mprj[91] la_oen_mprj[92] la_oen_mprj[93] la_oen_mprj[94]
+ la_oen_mprj[95] la_oen_mprj[96] la_oen_mprj[97] la_oen_mprj[98] la_oen_mprj[99]
+ la_oen_mprj[9] mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12]
+ mprj_adr_o_core[13] mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16]
+ mprj_adr_o_core[17] mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20]
+ mprj_adr_o_core[21] mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24]
+ mprj_adr_o_core[25] mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28]
+ mprj_adr_o_core[29] mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3]
+ mprj_adr_o_core[4] mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8]
+ mprj_adr_o_core[9] mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12]
+ mprj_adr_o_user[13] mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16]
+ mprj_adr_o_user[17] mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20]
+ mprj_adr_o_user[21] mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24]
+ mprj_adr_o_user[25] mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28]
+ mprj_adr_o_user[29] mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3]
+ mprj_adr_o_user[4] mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8]
+ mprj_adr_o_user[9] mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10]
+ mprj_dat_o_core[11] mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14]
+ mprj_dat_o_core[15] mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18]
+ mprj_dat_o_core[19] mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22]
+ mprj_dat_o_core[23] mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26]
+ mprj_dat_o_core[27] mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30]
+ mprj_dat_o_core[31] mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6]
+ mprj_dat_o_core[7] mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10]
+ mprj_dat_o_user[11] mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14]
+ mprj_dat_o_user[15] mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18]
+ mprj_dat_o_user[19] mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22]
+ mprj_dat_o_user[23] mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26]
+ mprj_dat_o_user[27] mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30]
+ mprj_dat_o_user[31] mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6]
+ mprj_dat_o_user[7] mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1]
+ mprj_sel_o_core[2] mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2]
+ mprj_sel_o_user[3] mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user
+ user1_vcc_powergood user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood
+ user_clock user_clock2 user_reset user_resetn vccd vssd vccd1 vssd1 vccd2 vssd2
+ vdda1 vssa1 vdda2 vssa2
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_4 abstract view
.subckt sky130_fd_sc_hvl__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__decap_8 abstract view
.subckt sky130_fd_sc_hvl__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_2 abstract view
.subckt sky130_fd_sc_hvl__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__fill_1 abstract view
.subckt sky130_fd_sc_hvl__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__diode_2 abstract view
.subckt sky130_fd_sc_hvl__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hvl__lsbufhv2lv_1 abstract view
.subckt sky130_fd_sc_hvl__lsbufhv2lv_1 A LVPWR VGND VNB VPB VPWR X
.ends

.subckt sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped A X VPWR VGND LVPWR LVGND VSUBS
XFILLER_0_24 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_28 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_2
XFILLER_0_16 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_1_30 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XFILLER_1_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_4
XFILLER_1_12 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XANTENNA_lvlshiftdown_A A VGND VGND VPWR VPWR sky130_fd_sc_hvl__diode_2
XFILLER_2_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_30 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XFILLER_2_10 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
XFILLER_0_0 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_2_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_2
Xlvlshiftdown A LVPWR VGND VGND VPWR VPWR X sky130_fd_sc_hvl__lsbufhv2lv_1
XFILLER_0_8 VGND VGND VPWR VPWR sky130_fd_sc_hvl__decap_8
XFILLER_0_30 VGND VGND VPWR VPWR sky130_fd_sc_hvl__fill_1
.ends

* Black-box entry subcircuit for user_project_wrapper abstract view
.subckt user_project_wrapper analog_io[0] analog_io[10] analog_io[11] analog_io[12]
+ analog_io[13] analog_io[14] analog_io[15] analog_io[16] analog_io[17] analog_io[18]
+ analog_io[19] analog_io[1] analog_io[20] analog_io[21] analog_io[22] analog_io[23]
+ analog_io[24] analog_io[25] analog_io[26] analog_io[27] analog_io[28] analog_io[29]
+ analog_io[2] analog_io[30] analog_io[3] analog_io[4] analog_io[5] analog_io[6] analog_io[7]
+ analog_io[8] analog_io[9] io_in[0] io_in[10] io_in[11] io_in[12] io_in[13] io_in[14]
+ io_in[15] io_in[16] io_in[17] io_in[18] io_in[19] io_in[1] io_in[20] io_in[21] io_in[22]
+ io_in[23] io_in[24] io_in[25] io_in[26] io_in[27] io_in[28] io_in[29] io_in[2] io_in[30]
+ io_in[31] io_in[32] io_in[33] io_in[34] io_in[35] io_in[36] io_in[37] io_in[3] io_in[4]
+ io_in[5] io_in[6] io_in[7] io_in[8] io_in[9] io_oeb[0] io_oeb[10] io_oeb[11] io_oeb[12]
+ io_oeb[13] io_oeb[14] io_oeb[15] io_oeb[16] io_oeb[17] io_oeb[18] io_oeb[19] io_oeb[1]
+ io_oeb[20] io_oeb[21] io_oeb[22] io_oeb[23] io_oeb[24] io_oeb[25] io_oeb[26] io_oeb[27]
+ io_oeb[28] io_oeb[29] io_oeb[2] io_oeb[30] io_oeb[31] io_oeb[32] io_oeb[33] io_oeb[34]
+ io_oeb[35] io_oeb[36] io_oeb[37] io_oeb[3] io_oeb[4] io_oeb[5] io_oeb[6] io_oeb[7]
+ io_oeb[8] io_oeb[9] io_out[0] io_out[10] io_out[11] io_out[12] io_out[13] io_out[14]
+ io_out[15] io_out[16] io_out[17] io_out[18] io_out[19] io_out[1] io_out[20] io_out[21]
+ io_out[22] io_out[23] io_out[24] io_out[25] io_out[26] io_out[27] io_out[28] io_out[29]
+ io_out[2] io_out[30] io_out[31] io_out[32] io_out[33] io_out[34] io_out[35] io_out[36]
+ io_out[37] io_out[3] io_out[4] io_out[5] io_out[6] io_out[7] io_out[8] io_out[9]
+ la_data_in[0] la_data_in[100] la_data_in[101] la_data_in[102] la_data_in[103] la_data_in[104]
+ la_data_in[105] la_data_in[106] la_data_in[107] la_data_in[108] la_data_in[109]
+ la_data_in[10] la_data_in[110] la_data_in[111] la_data_in[112] la_data_in[113] la_data_in[114]
+ la_data_in[115] la_data_in[116] la_data_in[117] la_data_in[118] la_data_in[119]
+ la_data_in[11] la_data_in[120] la_data_in[121] la_data_in[122] la_data_in[123] la_data_in[124]
+ la_data_in[125] la_data_in[126] la_data_in[127] la_data_in[12] la_data_in[13] la_data_in[14]
+ la_data_in[15] la_data_in[16] la_data_in[17] la_data_in[18] la_data_in[19] la_data_in[1]
+ la_data_in[20] la_data_in[21] la_data_in[22] la_data_in[23] la_data_in[24] la_data_in[25]
+ la_data_in[26] la_data_in[27] la_data_in[28] la_data_in[29] la_data_in[2] la_data_in[30]
+ la_data_in[31] la_data_in[32] la_data_in[33] la_data_in[34] la_data_in[35] la_data_in[36]
+ la_data_in[37] la_data_in[38] la_data_in[39] la_data_in[3] la_data_in[40] la_data_in[41]
+ la_data_in[42] la_data_in[43] la_data_in[44] la_data_in[45] la_data_in[46] la_data_in[47]
+ la_data_in[48] la_data_in[49] la_data_in[4] la_data_in[50] la_data_in[51] la_data_in[52]
+ la_data_in[53] la_data_in[54] la_data_in[55] la_data_in[56] la_data_in[57] la_data_in[58]
+ la_data_in[59] la_data_in[5] la_data_in[60] la_data_in[61] la_data_in[62] la_data_in[63]
+ la_data_in[64] la_data_in[65] la_data_in[66] la_data_in[67] la_data_in[68] la_data_in[69]
+ la_data_in[6] la_data_in[70] la_data_in[71] la_data_in[72] la_data_in[73] la_data_in[74]
+ la_data_in[75] la_data_in[76] la_data_in[77] la_data_in[78] la_data_in[79] la_data_in[7]
+ la_data_in[80] la_data_in[81] la_data_in[82] la_data_in[83] la_data_in[84] la_data_in[85]
+ la_data_in[86] la_data_in[87] la_data_in[88] la_data_in[89] la_data_in[8] la_data_in[90]
+ la_data_in[91] la_data_in[92] la_data_in[93] la_data_in[94] la_data_in[95] la_data_in[96]
+ la_data_in[97] la_data_in[98] la_data_in[99] la_data_in[9] la_data_out[0] la_data_out[100]
+ la_data_out[101] la_data_out[102] la_data_out[103] la_data_out[104] la_data_out[105]
+ la_data_out[106] la_data_out[107] la_data_out[108] la_data_out[109] la_data_out[10]
+ la_data_out[110] la_data_out[111] la_data_out[112] la_data_out[113] la_data_out[114]
+ la_data_out[115] la_data_out[116] la_data_out[117] la_data_out[118] la_data_out[119]
+ la_data_out[11] la_data_out[120] la_data_out[121] la_data_out[122] la_data_out[123]
+ la_data_out[124] la_data_out[125] la_data_out[126] la_data_out[127] la_data_out[12]
+ la_data_out[13] la_data_out[14] la_data_out[15] la_data_out[16] la_data_out[17]
+ la_data_out[18] la_data_out[19] la_data_out[1] la_data_out[20] la_data_out[21] la_data_out[22]
+ la_data_out[23] la_data_out[24] la_data_out[25] la_data_out[26] la_data_out[27]
+ la_data_out[28] la_data_out[29] la_data_out[2] la_data_out[30] la_data_out[31] la_data_out[32]
+ la_data_out[33] la_data_out[34] la_data_out[35] la_data_out[36] la_data_out[37]
+ la_data_out[38] la_data_out[39] la_data_out[3] la_data_out[40] la_data_out[41] la_data_out[42]
+ la_data_out[43] la_data_out[44] la_data_out[45] la_data_out[46] la_data_out[47]
+ la_data_out[48] la_data_out[49] la_data_out[4] la_data_out[50] la_data_out[51] la_data_out[52]
+ la_data_out[53] la_data_out[54] la_data_out[55] la_data_out[56] la_data_out[57]
+ la_data_out[58] la_data_out[59] la_data_out[5] la_data_out[60] la_data_out[61] la_data_out[62]
+ la_data_out[63] la_data_out[64] la_data_out[65] la_data_out[66] la_data_out[67]
+ la_data_out[68] la_data_out[69] la_data_out[6] la_data_out[70] la_data_out[71] la_data_out[72]
+ la_data_out[73] la_data_out[74] la_data_out[75] la_data_out[76] la_data_out[77]
+ la_data_out[78] la_data_out[79] la_data_out[7] la_data_out[80] la_data_out[81] la_data_out[82]
+ la_data_out[83] la_data_out[84] la_data_out[85] la_data_out[86] la_data_out[87]
+ la_data_out[88] la_data_out[89] la_data_out[8] la_data_out[90] la_data_out[91] la_data_out[92]
+ la_data_out[93] la_data_out[94] la_data_out[95] la_data_out[96] la_data_out[97]
+ la_data_out[98] la_data_out[99] la_data_out[9] la_oen[0] la_oen[100] la_oen[101]
+ la_oen[102] la_oen[103] la_oen[104] la_oen[105] la_oen[106] la_oen[107] la_oen[108]
+ la_oen[109] la_oen[10] la_oen[110] la_oen[111] la_oen[112] la_oen[113] la_oen[114]
+ la_oen[115] la_oen[116] la_oen[117] la_oen[118] la_oen[119] la_oen[11] la_oen[120]
+ la_oen[121] la_oen[122] la_oen[123] la_oen[124] la_oen[125] la_oen[126] la_oen[127]
+ la_oen[12] la_oen[13] la_oen[14] la_oen[15] la_oen[16] la_oen[17] la_oen[18] la_oen[19]
+ la_oen[1] la_oen[20] la_oen[21] la_oen[22] la_oen[23] la_oen[24] la_oen[25] la_oen[26]
+ la_oen[27] la_oen[28] la_oen[29] la_oen[2] la_oen[30] la_oen[31] la_oen[32] la_oen[33]
+ la_oen[34] la_oen[35] la_oen[36] la_oen[37] la_oen[38] la_oen[39] la_oen[3] la_oen[40]
+ la_oen[41] la_oen[42] la_oen[43] la_oen[44] la_oen[45] la_oen[46] la_oen[47] la_oen[48]
+ la_oen[49] la_oen[4] la_oen[50] la_oen[51] la_oen[52] la_oen[53] la_oen[54] la_oen[55]
+ la_oen[56] la_oen[57] la_oen[58] la_oen[59] la_oen[5] la_oen[60] la_oen[61] la_oen[62]
+ la_oen[63] la_oen[64] la_oen[65] la_oen[66] la_oen[67] la_oen[68] la_oen[69] la_oen[6]
+ la_oen[70] la_oen[71] la_oen[72] la_oen[73] la_oen[74] la_oen[75] la_oen[76] la_oen[77]
+ la_oen[78] la_oen[79] la_oen[7] la_oen[80] la_oen[81] la_oen[82] la_oen[83] la_oen[84]
+ la_oen[85] la_oen[86] la_oen[87] la_oen[88] la_oen[89] la_oen[8] la_oen[90] la_oen[91]
+ la_oen[92] la_oen[93] la_oen[94] la_oen[95] la_oen[96] la_oen[97] la_oen[98] la_oen[99]
+ la_oen[9] user_clock2 wb_clk_i wb_rst_i wbs_ack_o wbs_adr_i[0] wbs_adr_i[10] wbs_adr_i[11]
+ wbs_adr_i[12] wbs_adr_i[13] wbs_adr_i[14] wbs_adr_i[15] wbs_adr_i[16] wbs_adr_i[17]
+ wbs_adr_i[18] wbs_adr_i[19] wbs_adr_i[1] wbs_adr_i[20] wbs_adr_i[21] wbs_adr_i[22]
+ wbs_adr_i[23] wbs_adr_i[24] wbs_adr_i[25] wbs_adr_i[26] wbs_adr_i[27] wbs_adr_i[28]
+ wbs_adr_i[29] wbs_adr_i[2] wbs_adr_i[30] wbs_adr_i[31] wbs_adr_i[3] wbs_adr_i[4]
+ wbs_adr_i[5] wbs_adr_i[6] wbs_adr_i[7] wbs_adr_i[8] wbs_adr_i[9] wbs_cyc_i wbs_dat_i[0]
+ wbs_dat_i[10] wbs_dat_i[11] wbs_dat_i[12] wbs_dat_i[13] wbs_dat_i[14] wbs_dat_i[15]
+ wbs_dat_i[16] wbs_dat_i[17] wbs_dat_i[18] wbs_dat_i[19] wbs_dat_i[1] wbs_dat_i[20]
+ wbs_dat_i[21] wbs_dat_i[22] wbs_dat_i[23] wbs_dat_i[24] wbs_dat_i[25] wbs_dat_i[26]
+ wbs_dat_i[27] wbs_dat_i[28] wbs_dat_i[29] wbs_dat_i[2] wbs_dat_i[30] wbs_dat_i[31]
+ wbs_dat_i[3] wbs_dat_i[4] wbs_dat_i[5] wbs_dat_i[6] wbs_dat_i[7] wbs_dat_i[8] wbs_dat_i[9]
+ wbs_dat_o[0] wbs_dat_o[10] wbs_dat_o[11] wbs_dat_o[12] wbs_dat_o[13] wbs_dat_o[14]
+ wbs_dat_o[15] wbs_dat_o[16] wbs_dat_o[17] wbs_dat_o[18] wbs_dat_o[19] wbs_dat_o[1]
+ wbs_dat_o[20] wbs_dat_o[21] wbs_dat_o[22] wbs_dat_o[23] wbs_dat_o[24] wbs_dat_o[25]
+ wbs_dat_o[26] wbs_dat_o[27] wbs_dat_o[28] wbs_dat_o[29] wbs_dat_o[2] wbs_dat_o[30]
+ wbs_dat_o[31] wbs_dat_o[3] wbs_dat_o[4] wbs_dat_o[5] wbs_dat_o[6] wbs_dat_o[7] wbs_dat_o[8]
+ wbs_dat_o[9] wbs_sel_i[0] wbs_sel_i[1] wbs_sel_i[2] wbs_sel_i[3] wbs_stb_i wbs_we_i
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
.ends

* Black-box entry subcircuit for storage abstract view
.subckt storage mgmt_addr[0] mgmt_addr[1] mgmt_addr[2] mgmt_addr[3] mgmt_addr[4] mgmt_addr[5]
+ mgmt_addr[6] mgmt_addr[7] mgmt_addr_ro[0] mgmt_addr_ro[1] mgmt_addr_ro[2] mgmt_addr_ro[3]
+ mgmt_addr_ro[4] mgmt_addr_ro[5] mgmt_addr_ro[6] mgmt_addr_ro[7] mgmt_clk mgmt_ena[0]
+ mgmt_ena[1] mgmt_ena_ro mgmt_rdata[0] mgmt_rdata[10] mgmt_rdata[11] mgmt_rdata[12]
+ mgmt_rdata[13] mgmt_rdata[14] mgmt_rdata[15] mgmt_rdata[16] mgmt_rdata[17] mgmt_rdata[18]
+ mgmt_rdata[19] mgmt_rdata[1] mgmt_rdata[20] mgmt_rdata[21] mgmt_rdata[22] mgmt_rdata[23]
+ mgmt_rdata[24] mgmt_rdata[25] mgmt_rdata[26] mgmt_rdata[27] mgmt_rdata[28] mgmt_rdata[29]
+ mgmt_rdata[2] mgmt_rdata[30] mgmt_rdata[31] mgmt_rdata[32] mgmt_rdata[33] mgmt_rdata[34]
+ mgmt_rdata[35] mgmt_rdata[36] mgmt_rdata[37] mgmt_rdata[38] mgmt_rdata[39] mgmt_rdata[3]
+ mgmt_rdata[40] mgmt_rdata[41] mgmt_rdata[42] mgmt_rdata[43] mgmt_rdata[44] mgmt_rdata[45]
+ mgmt_rdata[46] mgmt_rdata[47] mgmt_rdata[48] mgmt_rdata[49] mgmt_rdata[4] mgmt_rdata[50]
+ mgmt_rdata[51] mgmt_rdata[52] mgmt_rdata[53] mgmt_rdata[54] mgmt_rdata[55] mgmt_rdata[56]
+ mgmt_rdata[57] mgmt_rdata[58] mgmt_rdata[59] mgmt_rdata[5] mgmt_rdata[60] mgmt_rdata[61]
+ mgmt_rdata[62] mgmt_rdata[63] mgmt_rdata[6] mgmt_rdata[7] mgmt_rdata[8] mgmt_rdata[9]
+ mgmt_rdata_ro[0] mgmt_rdata_ro[10] mgmt_rdata_ro[11] mgmt_rdata_ro[12] mgmt_rdata_ro[13]
+ mgmt_rdata_ro[14] mgmt_rdata_ro[15] mgmt_rdata_ro[16] mgmt_rdata_ro[17] mgmt_rdata_ro[18]
+ mgmt_rdata_ro[19] mgmt_rdata_ro[1] mgmt_rdata_ro[20] mgmt_rdata_ro[21] mgmt_rdata_ro[22]
+ mgmt_rdata_ro[23] mgmt_rdata_ro[24] mgmt_rdata_ro[25] mgmt_rdata_ro[26] mgmt_rdata_ro[27]
+ mgmt_rdata_ro[28] mgmt_rdata_ro[29] mgmt_rdata_ro[2] mgmt_rdata_ro[30] mgmt_rdata_ro[31]
+ mgmt_rdata_ro[3] mgmt_rdata_ro[4] mgmt_rdata_ro[5] mgmt_rdata_ro[6] mgmt_rdata_ro[7]
+ mgmt_rdata_ro[8] mgmt_rdata_ro[9] mgmt_wdata[0] mgmt_wdata[10] mgmt_wdata[11] mgmt_wdata[12]
+ mgmt_wdata[13] mgmt_wdata[14] mgmt_wdata[15] mgmt_wdata[16] mgmt_wdata[17] mgmt_wdata[18]
+ mgmt_wdata[19] mgmt_wdata[1] mgmt_wdata[20] mgmt_wdata[21] mgmt_wdata[22] mgmt_wdata[23]
+ mgmt_wdata[24] mgmt_wdata[25] mgmt_wdata[26] mgmt_wdata[27] mgmt_wdata[28] mgmt_wdata[29]
+ mgmt_wdata[2] mgmt_wdata[30] mgmt_wdata[31] mgmt_wdata[3] mgmt_wdata[4] mgmt_wdata[5]
+ mgmt_wdata[6] mgmt_wdata[7] mgmt_wdata[8] mgmt_wdata[9] mgmt_wen[0] mgmt_wen[1]
+ mgmt_wen_mask[0] mgmt_wen_mask[1] mgmt_wen_mask[2] mgmt_wen_mask[3] mgmt_wen_mask[4]
+ mgmt_wen_mask[5] mgmt_wen_mask[6] mgmt_wen_mask[7] VPWR VGND
.ends

.subckt caravel clock flash_clk flash_csb flash_io0 flash_io1 gpio mprj_io[0] mprj_io[10]
+ mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15] mprj_io[16] mprj_io[17]
+ mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21] mprj_io[22] mprj_io[23]
+ mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28] mprj_io[29] mprj_io[2]
+ mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34] mprj_io[35] mprj_io[36]
+ mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] mprj_io[7] mprj_io[8] mprj_io[9]
+ resetb pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2] pwr_ctrl_out[3] vssa_pad
+ vssd_pad vssio_pad vdda_pad vssd1_pad vdda1_pad vccd1_pad vssa1_pad vccd2_pad vssa2_pad
+ vdda2_pad vssd2_pad vddio_pad vccd_pad vssio_pad2 vddio_pad2 vssa1_pad2 vdda1_pad2
Xgpio_control_in\[28\] soc/mgmt_in_data[28] gpio_control_in\[28\]/one soc/mgmt_in_data[28]
+ gpio_control_in\[28\]/one padframe/mprj_io_analog_en[28] padframe/mprj_io_analog_pol[28]
+ padframe/mprj_io_analog_sel[28] padframe/mprj_io_dm[84] padframe/mprj_io_dm[85]
+ padframe/mprj_io_dm[86] padframe/mprj_io_holdover[28] padframe/mprj_io_ib_mode_sel[28]
+ padframe/mprj_io_in[28] padframe/mprj_io_inp_dis[28] padframe/mprj_io_out[28] padframe/mprj_io_oeb[28]
+ padframe/mprj_io_slow_sel[28] padframe/mprj_io_vtrip_sel[28] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[28\]/serial_data_in gpio_control_in\[29\]/serial_data_in
+ mprj/io_in[28] mprj/io_oeb[28] mprj/io_out[28] gpio_control_in\[28\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[10\] soc/mgmt_in_data[10] gpio_control_in\[10\]/one soc/mgmt_in_data[10]
+ gpio_control_in\[10\]/one padframe/mprj_io_analog_en[10] padframe/mprj_io_analog_pol[10]
+ padframe/mprj_io_analog_sel[10] padframe/mprj_io_dm[30] padframe/mprj_io_dm[31]
+ padframe/mprj_io_dm[32] padframe/mprj_io_holdover[10] padframe/mprj_io_ib_mode_sel[10]
+ padframe/mprj_io_in[10] padframe/mprj_io_inp_dis[10] padframe/mprj_io_out[10] padframe/mprj_io_oeb[10]
+ padframe/mprj_io_slow_sel[10] padframe/mprj_io_vtrip_sel[10] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[9\]/serial_data_out gpio_control_in\[11\]/serial_data_in
+ mprj/io_in[10] mprj/io_oeb[10] mprj/io_out[10] gpio_control_in\[10\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xpadframe clock soc/clock flash_clk soc/flash_clk soc/flash_clk_ieb soc/flash_clk_oeb
+ flash_csb soc/flash_csb soc/flash_csb_ieb soc/flash_csb_oeb flash_io0 soc/flash_io0_di
+ soc/flash_io0_do soc/flash_io0_ieb soc/flash_io0_oeb flash_io1 soc/flash_io1_di
+ soc/flash_io1_do soc/flash_io1_ieb soc/flash_io1_oeb gpio soc/gpio_in_pad soc/gpio_inenb_pad
+ soc/gpio_mode0_pad soc/gpio_mode1_pad soc/gpio_out_pad soc/gpio_outenb_pad mprj/analog_io[0]
+ mprj/analog_io[10] mprj/analog_io[11] mprj/analog_io[12] mprj/analog_io[13] mprj/analog_io[14]
+ mprj/analog_io[15] mprj/analog_io[16] mprj/analog_io[17] mprj/analog_io[18] mprj/analog_io[19]
+ mprj/analog_io[1] mprj/analog_io[20] mprj/analog_io[21] mprj/analog_io[22] mprj/analog_io[23]
+ mprj/analog_io[24] mprj/analog_io[25] mprj/analog_io[26] mprj/analog_io[27] mprj/analog_io[28]
+ mprj/analog_io[29] mprj/analog_io[2] mprj/analog_io[30] mprj/analog_io[3] mprj/analog_io[4]
+ mprj/analog_io[5] mprj/analog_io[6] mprj/analog_io[7] mprj/analog_io[8] mprj/analog_io[9]
+ mprj_io[0] mprj_io[10] mprj_io[11] mprj_io[12] mprj_io[13] mprj_io[14] mprj_io[15]
+ mprj_io[16] mprj_io[17] mprj_io[18] mprj_io[19] mprj_io[1] mprj_io[20] mprj_io[21]
+ mprj_io[22] mprj_io[23] mprj_io[24] mprj_io[25] mprj_io[26] mprj_io[27] mprj_io[28]
+ mprj_io[29] mprj_io[2] mprj_io[30] mprj_io[31] mprj_io[32] mprj_io[33] mprj_io[34]
+ mprj_io[35] mprj_io[36] mprj_io[37] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6]
+ mprj_io[7] mprj_io[8] mprj_io[9] padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_en[10]
+ padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_en[12] padframe/mprj_io_analog_en[13]
+ padframe/mprj_io_analog_en[14] padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_en[16]
+ padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_en[18] padframe/mprj_io_analog_en[19]
+ padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_en[20] padframe/mprj_io_analog_en[21]
+ padframe/mprj_io_analog_en[22] padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_en[24]
+ padframe/mprj_io_analog_en[25] padframe/mprj_io_analog_en[26] padframe/mprj_io_analog_en[27]
+ padframe/mprj_io_analog_en[28] padframe/mprj_io_analog_en[29] padframe/mprj_io_analog_en[2]
+ padframe/mprj_io_analog_en[30] padframe/mprj_io_analog_en[31] padframe/mprj_io_analog_en[32]
+ padframe/mprj_io_analog_en[33] padframe/mprj_io_analog_en[34] padframe/mprj_io_analog_en[35]
+ padframe/mprj_io_analog_en[36] padframe/mprj_io_analog_en[37] padframe/mprj_io_analog_en[3]
+ padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_en[6]
+ padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_en[9]
+ padframe/mprj_io_analog_pol[0] padframe/mprj_io_analog_pol[10] padframe/mprj_io_analog_pol[11]
+ padframe/mprj_io_analog_pol[12] padframe/mprj_io_analog_pol[13] padframe/mprj_io_analog_pol[14]
+ padframe/mprj_io_analog_pol[15] padframe/mprj_io_analog_pol[16] padframe/mprj_io_analog_pol[17]
+ padframe/mprj_io_analog_pol[18] padframe/mprj_io_analog_pol[19] padframe/mprj_io_analog_pol[1]
+ padframe/mprj_io_analog_pol[20] padframe/mprj_io_analog_pol[21] padframe/mprj_io_analog_pol[22]
+ padframe/mprj_io_analog_pol[23] padframe/mprj_io_analog_pol[24] padframe/mprj_io_analog_pol[25]
+ padframe/mprj_io_analog_pol[26] padframe/mprj_io_analog_pol[27] padframe/mprj_io_analog_pol[28]
+ padframe/mprj_io_analog_pol[29] padframe/mprj_io_analog_pol[2] padframe/mprj_io_analog_pol[30]
+ padframe/mprj_io_analog_pol[31] padframe/mprj_io_analog_pol[32] padframe/mprj_io_analog_pol[33]
+ padframe/mprj_io_analog_pol[34] padframe/mprj_io_analog_pol[35] padframe/mprj_io_analog_pol[36]
+ padframe/mprj_io_analog_pol[37] padframe/mprj_io_analog_pol[3] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_pol[5] padframe/mprj_io_analog_pol[6] padframe/mprj_io_analog_pol[7]
+ padframe/mprj_io_analog_pol[8] padframe/mprj_io_analog_pol[9] padframe/mprj_io_analog_sel[0]
+ padframe/mprj_io_analog_sel[10] padframe/mprj_io_analog_sel[11] padframe/mprj_io_analog_sel[12]
+ padframe/mprj_io_analog_sel[13] padframe/mprj_io_analog_sel[14] padframe/mprj_io_analog_sel[15]
+ padframe/mprj_io_analog_sel[16] padframe/mprj_io_analog_sel[17] padframe/mprj_io_analog_sel[18]
+ padframe/mprj_io_analog_sel[19] padframe/mprj_io_analog_sel[1] padframe/mprj_io_analog_sel[20]
+ padframe/mprj_io_analog_sel[21] padframe/mprj_io_analog_sel[22] padframe/mprj_io_analog_sel[23]
+ padframe/mprj_io_analog_sel[24] padframe/mprj_io_analog_sel[25] padframe/mprj_io_analog_sel[26]
+ padframe/mprj_io_analog_sel[27] padframe/mprj_io_analog_sel[28] padframe/mprj_io_analog_sel[29]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_analog_sel[30] padframe/mprj_io_analog_sel[31]
+ padframe/mprj_io_analog_sel[32] padframe/mprj_io_analog_sel[33] padframe/mprj_io_analog_sel[34]
+ padframe/mprj_io_analog_sel[35] padframe/mprj_io_analog_sel[36] padframe/mprj_io_analog_sel[37]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_analog_sel[4] padframe/mprj_io_analog_sel[5]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_analog_sel[7] padframe/mprj_io_analog_sel[8]
+ padframe/mprj_io_analog_sel[9] padframe/mprj_io_dm[0] padframe/mprj_io_dm[100] padframe/mprj_io_dm[101]
+ padframe/mprj_io_dm[102] padframe/mprj_io_dm[103] padframe/mprj_io_dm[104] padframe/mprj_io_dm[105]
+ padframe/mprj_io_dm[106] padframe/mprj_io_dm[107] padframe/mprj_io_dm[108] padframe/mprj_io_dm[109]
+ padframe/mprj_io_dm[10] padframe/mprj_io_dm[110] padframe/mprj_io_dm[111] padframe/mprj_io_dm[112]
+ padframe/mprj_io_dm[113] padframe/mprj_io_dm[11] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13]
+ padframe/mprj_io_dm[14] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[1] padframe/mprj_io_dm[20]
+ padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23] padframe/mprj_io_dm[24]
+ padframe/mprj_io_dm[25] padframe/mprj_io_dm[26] padframe/mprj_io_dm[27] padframe/mprj_io_dm[28]
+ padframe/mprj_io_dm[29] padframe/mprj_io_dm[2] padframe/mprj_io_dm[30] padframe/mprj_io_dm[31]
+ padframe/mprj_io_dm[32] padframe/mprj_io_dm[33] padframe/mprj_io_dm[34] padframe/mprj_io_dm[35]
+ padframe/mprj_io_dm[36] padframe/mprj_io_dm[37] padframe/mprj_io_dm[38] padframe/mprj_io_dm[39]
+ padframe/mprj_io_dm[3] padframe/mprj_io_dm[40] padframe/mprj_io_dm[41] padframe/mprj_io_dm[42]
+ padframe/mprj_io_dm[43] padframe/mprj_io_dm[44] padframe/mprj_io_dm[45] padframe/mprj_io_dm[46]
+ padframe/mprj_io_dm[47] padframe/mprj_io_dm[48] padframe/mprj_io_dm[49] padframe/mprj_io_dm[4]
+ padframe/mprj_io_dm[50] padframe/mprj_io_dm[51] padframe/mprj_io_dm[52] padframe/mprj_io_dm[53]
+ padframe/mprj_io_dm[54] padframe/mprj_io_dm[55] padframe/mprj_io_dm[56] padframe/mprj_io_dm[57]
+ padframe/mprj_io_dm[58] padframe/mprj_io_dm[59] padframe/mprj_io_dm[5] padframe/mprj_io_dm[60]
+ padframe/mprj_io_dm[61] padframe/mprj_io_dm[62] padframe/mprj_io_dm[63] padframe/mprj_io_dm[64]
+ padframe/mprj_io_dm[65] padframe/mprj_io_dm[66] padframe/mprj_io_dm[67] padframe/mprj_io_dm[68]
+ padframe/mprj_io_dm[69] padframe/mprj_io_dm[6] padframe/mprj_io_dm[70] padframe/mprj_io_dm[71]
+ padframe/mprj_io_dm[72] padframe/mprj_io_dm[73] padframe/mprj_io_dm[74] padframe/mprj_io_dm[75]
+ padframe/mprj_io_dm[76] padframe/mprj_io_dm[77] padframe/mprj_io_dm[78] padframe/mprj_io_dm[79]
+ padframe/mprj_io_dm[7] padframe/mprj_io_dm[80] padframe/mprj_io_dm[81] padframe/mprj_io_dm[82]
+ padframe/mprj_io_dm[83] padframe/mprj_io_dm[84] padframe/mprj_io_dm[85] padframe/mprj_io_dm[86]
+ padframe/mprj_io_dm[87] padframe/mprj_io_dm[88] padframe/mprj_io_dm[89] padframe/mprj_io_dm[8]
+ padframe/mprj_io_dm[90] padframe/mprj_io_dm[91] padframe/mprj_io_dm[92] padframe/mprj_io_dm[93]
+ padframe/mprj_io_dm[94] padframe/mprj_io_dm[95] padframe/mprj_io_dm[96] padframe/mprj_io_dm[97]
+ padframe/mprj_io_dm[98] padframe/mprj_io_dm[99] padframe/mprj_io_dm[9] por/porb_h
+ por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h
+ por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h
+ por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h
+ por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h
+ por/porb_h por/porb_h por/porb_h por/porb_h por/porb_h vddio vddio vddio vddio vddio
+ vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio
+ vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio vddio
+ vddio vddio vddio vddio vddio padframe/mprj_io_holdover[0] padframe/mprj_io_holdover[10]
+ padframe/mprj_io_holdover[11] padframe/mprj_io_holdover[12] padframe/mprj_io_holdover[13]
+ padframe/mprj_io_holdover[14] padframe/mprj_io_holdover[15] padframe/mprj_io_holdover[16]
+ padframe/mprj_io_holdover[17] padframe/mprj_io_holdover[18] padframe/mprj_io_holdover[19]
+ padframe/mprj_io_holdover[1] padframe/mprj_io_holdover[20] padframe/mprj_io_holdover[21]
+ padframe/mprj_io_holdover[22] padframe/mprj_io_holdover[23] padframe/mprj_io_holdover[24]
+ padframe/mprj_io_holdover[25] padframe/mprj_io_holdover[26] padframe/mprj_io_holdover[27]
+ padframe/mprj_io_holdover[28] padframe/mprj_io_holdover[29] padframe/mprj_io_holdover[2]
+ padframe/mprj_io_holdover[30] padframe/mprj_io_holdover[31] padframe/mprj_io_holdover[32]
+ padframe/mprj_io_holdover[33] padframe/mprj_io_holdover[34] padframe/mprj_io_holdover[35]
+ padframe/mprj_io_holdover[36] padframe/mprj_io_holdover[37] padframe/mprj_io_holdover[3]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_holdover[5] padframe/mprj_io_holdover[6]
+ padframe/mprj_io_holdover[7] padframe/mprj_io_holdover[8] padframe/mprj_io_holdover[9]
+ padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_ib_mode_sel[10] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_ib_mode_sel[12] padframe/mprj_io_ib_mode_sel[13] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_ib_mode_sel[15] padframe/mprj_io_ib_mode_sel[16] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_ib_mode_sel[18] padframe/mprj_io_ib_mode_sel[19] padframe/mprj_io_ib_mode_sel[1]
+ padframe/mprj_io_ib_mode_sel[20] padframe/mprj_io_ib_mode_sel[21] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_ib_mode_sel[23] padframe/mprj_io_ib_mode_sel[24] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_ib_mode_sel[26] padframe/mprj_io_ib_mode_sel[27] padframe/mprj_io_ib_mode_sel[28]
+ padframe/mprj_io_ib_mode_sel[29] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_ib_mode_sel[30]
+ padframe/mprj_io_ib_mode_sel[31] padframe/mprj_io_ib_mode_sel[32] padframe/mprj_io_ib_mode_sel[33]
+ padframe/mprj_io_ib_mode_sel[34] padframe/mprj_io_ib_mode_sel[35] padframe/mprj_io_ib_mode_sel[36]
+ padframe/mprj_io_ib_mode_sel[37] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_ib_mode_sel[4]
+ padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_ib_mode_sel[7]
+ padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[0]
+ padframe/mprj_io_in[10] padframe/mprj_io_in[11] padframe/mprj_io_in[12] padframe/mprj_io_in[13]
+ padframe/mprj_io_in[14] padframe/mprj_io_in[15] padframe/mprj_io_in[16] padframe/mprj_io_in[17]
+ padframe/mprj_io_in[18] padframe/mprj_io_in[19] padframe/mprj_io_in[1] padframe/mprj_io_in[20]
+ padframe/mprj_io_in[21] padframe/mprj_io_in[22] padframe/mprj_io_in[23] padframe/mprj_io_in[24]
+ padframe/mprj_io_in[25] padframe/mprj_io_in[26] padframe/mprj_io_in[27] padframe/mprj_io_in[28]
+ padframe/mprj_io_in[29] padframe/mprj_io_in[2] padframe/mprj_io_in[30] padframe/mprj_io_in[31]
+ padframe/mprj_io_in[32] padframe/mprj_io_in[33] padframe/mprj_io_in[34] padframe/mprj_io_in[35]
+ padframe/mprj_io_in[36] padframe/mprj_io_in[37] padframe/mprj_io_in[3] padframe/mprj_io_in[4]
+ padframe/mprj_io_in[5] padframe/mprj_io_in[6] padframe/mprj_io_in[7] padframe/mprj_io_in[8]
+ padframe/mprj_io_in[9] padframe/mprj_io_inp_dis[0] padframe/mprj_io_inp_dis[10]
+ padframe/mprj_io_inp_dis[11] padframe/mprj_io_inp_dis[12] padframe/mprj_io_inp_dis[13]
+ padframe/mprj_io_inp_dis[14] padframe/mprj_io_inp_dis[15] padframe/mprj_io_inp_dis[16]
+ padframe/mprj_io_inp_dis[17] padframe/mprj_io_inp_dis[18] padframe/mprj_io_inp_dis[19]
+ padframe/mprj_io_inp_dis[1] padframe/mprj_io_inp_dis[20] padframe/mprj_io_inp_dis[21]
+ padframe/mprj_io_inp_dis[22] padframe/mprj_io_inp_dis[23] padframe/mprj_io_inp_dis[24]
+ padframe/mprj_io_inp_dis[25] padframe/mprj_io_inp_dis[26] padframe/mprj_io_inp_dis[27]
+ padframe/mprj_io_inp_dis[28] padframe/mprj_io_inp_dis[29] padframe/mprj_io_inp_dis[2]
+ padframe/mprj_io_inp_dis[30] padframe/mprj_io_inp_dis[31] padframe/mprj_io_inp_dis[32]
+ padframe/mprj_io_inp_dis[33] padframe/mprj_io_inp_dis[34] padframe/mprj_io_inp_dis[35]
+ padframe/mprj_io_inp_dis[36] padframe/mprj_io_inp_dis[37] padframe/mprj_io_inp_dis[3]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_inp_dis[5] padframe/mprj_io_inp_dis[6]
+ padframe/mprj_io_inp_dis[7] padframe/mprj_io_inp_dis[8] padframe/mprj_io_inp_dis[9]
+ padframe/mprj_io_oeb[0] padframe/mprj_io_oeb[10] padframe/mprj_io_oeb[11] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_oeb[13] padframe/mprj_io_oeb[14] padframe/mprj_io_oeb[15] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_oeb[17] padframe/mprj_io_oeb[18] padframe/mprj_io_oeb[19] padframe/mprj_io_oeb[1]
+ padframe/mprj_io_oeb[20] padframe/mprj_io_oeb[21] padframe/mprj_io_oeb[22] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_oeb[24] padframe/mprj_io_oeb[25] padframe/mprj_io_oeb[26] padframe/mprj_io_oeb[27]
+ padframe/mprj_io_oeb[28] padframe/mprj_io_oeb[29] padframe/mprj_io_oeb[2] padframe/mprj_io_oeb[30]
+ padframe/mprj_io_oeb[31] padframe/mprj_io_oeb[32] padframe/mprj_io_oeb[33] padframe/mprj_io_oeb[34]
+ padframe/mprj_io_oeb[35] padframe/mprj_io_oeb[36] padframe/mprj_io_oeb[37] padframe/mprj_io_oeb[3]
+ padframe/mprj_io_oeb[4] padframe/mprj_io_oeb[5] padframe/mprj_io_oeb[6] padframe/mprj_io_oeb[7]
+ padframe/mprj_io_oeb[8] padframe/mprj_io_oeb[9] padframe/mprj_io_out[0] padframe/mprj_io_out[10]
+ padframe/mprj_io_out[11] padframe/mprj_io_out[12] padframe/mprj_io_out[13] padframe/mprj_io_out[14]
+ padframe/mprj_io_out[15] padframe/mprj_io_out[16] padframe/mprj_io_out[17] padframe/mprj_io_out[18]
+ padframe/mprj_io_out[19] padframe/mprj_io_out[1] padframe/mprj_io_out[20] padframe/mprj_io_out[21]
+ padframe/mprj_io_out[22] padframe/mprj_io_out[23] padframe/mprj_io_out[24] padframe/mprj_io_out[25]
+ padframe/mprj_io_out[26] padframe/mprj_io_out[27] padframe/mprj_io_out[28] padframe/mprj_io_out[29]
+ padframe/mprj_io_out[2] padframe/mprj_io_out[30] padframe/mprj_io_out[31] padframe/mprj_io_out[32]
+ padframe/mprj_io_out[33] padframe/mprj_io_out[34] padframe/mprj_io_out[35] padframe/mprj_io_out[36]
+ padframe/mprj_io_out[37] padframe/mprj_io_out[3] padframe/mprj_io_out[4] padframe/mprj_io_out[5]
+ padframe/mprj_io_out[6] padframe/mprj_io_out[7] padframe/mprj_io_out[8] padframe/mprj_io_out[9]
+ padframe/mprj_io_slow_sel[0] padframe/mprj_io_slow_sel[10] padframe/mprj_io_slow_sel[11]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_slow_sel[13] padframe/mprj_io_slow_sel[14]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_slow_sel[16] padframe/mprj_io_slow_sel[17]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_slow_sel[19] padframe/mprj_io_slow_sel[1]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_slow_sel[21] padframe/mprj_io_slow_sel[22]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_slow_sel[24] padframe/mprj_io_slow_sel[25]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_slow_sel[27] padframe/mprj_io_slow_sel[28]
+ padframe/mprj_io_slow_sel[29] padframe/mprj_io_slow_sel[2] padframe/mprj_io_slow_sel[30]
+ padframe/mprj_io_slow_sel[31] padframe/mprj_io_slow_sel[32] padframe/mprj_io_slow_sel[33]
+ padframe/mprj_io_slow_sel[34] padframe/mprj_io_slow_sel[35] padframe/mprj_io_slow_sel[36]
+ padframe/mprj_io_slow_sel[37] padframe/mprj_io_slow_sel[3] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_slow_sel[5] padframe/mprj_io_slow_sel[6] padframe/mprj_io_slow_sel[7]
+ padframe/mprj_io_slow_sel[8] padframe/mprj_io_slow_sel[9] padframe/mprj_io_vtrip_sel[0]
+ padframe/mprj_io_vtrip_sel[10] padframe/mprj_io_vtrip_sel[11] padframe/mprj_io_vtrip_sel[12]
+ padframe/mprj_io_vtrip_sel[13] padframe/mprj_io_vtrip_sel[14] padframe/mprj_io_vtrip_sel[15]
+ padframe/mprj_io_vtrip_sel[16] padframe/mprj_io_vtrip_sel[17] padframe/mprj_io_vtrip_sel[18]
+ padframe/mprj_io_vtrip_sel[19] padframe/mprj_io_vtrip_sel[1] padframe/mprj_io_vtrip_sel[20]
+ padframe/mprj_io_vtrip_sel[21] padframe/mprj_io_vtrip_sel[22] padframe/mprj_io_vtrip_sel[23]
+ padframe/mprj_io_vtrip_sel[24] padframe/mprj_io_vtrip_sel[25] padframe/mprj_io_vtrip_sel[26]
+ padframe/mprj_io_vtrip_sel[27] padframe/mprj_io_vtrip_sel[28] padframe/mprj_io_vtrip_sel[29]
+ padframe/mprj_io_vtrip_sel[2] padframe/mprj_io_vtrip_sel[30] padframe/mprj_io_vtrip_sel[31]
+ padframe/mprj_io_vtrip_sel[32] padframe/mprj_io_vtrip_sel[33] padframe/mprj_io_vtrip_sel[34]
+ padframe/mprj_io_vtrip_sel[35] padframe/mprj_io_vtrip_sel[36] padframe/mprj_io_vtrip_sel[37]
+ padframe/mprj_io_vtrip_sel[3] padframe/mprj_io_vtrip_sel[4] padframe/mprj_io_vtrip_sel[5]
+ padframe/mprj_io_vtrip_sel[6] padframe/mprj_io_vtrip_sel[7] padframe/mprj_io_vtrip_sel[8]
+ padframe/mprj_io_vtrip_sel[9] por/por_l por/porb_h resetb rstb_level/A vccd vccd1
+ vccd1_pad vccd2 vccd2_pad vccd_pad padframe/vdda vdda1 vdda1_pad vdda2 vdda2_pad
+ vdda_pad vddio vddio_pad padframe/vssa vssa1 vssa1_pad vssa2 vssa2_pad vssa_pad
+ vssd vssd1 vssd1_pad vssd2 vssd2_pad vssd_pad vssio vssio_pad vssio_pad2 vddio_pad2
+ vssa1_pad2 vdda1_pad2 VSUBS chip_io
Xgpio_control_in\[26\] soc/mgmt_in_data[26] gpio_control_in\[26\]/one soc/mgmt_in_data[26]
+ gpio_control_in\[26\]/one padframe/mprj_io_analog_en[26] padframe/mprj_io_analog_pol[26]
+ padframe/mprj_io_analog_sel[26] padframe/mprj_io_dm[78] padframe/mprj_io_dm[79]
+ padframe/mprj_io_dm[80] padframe/mprj_io_holdover[26] padframe/mprj_io_ib_mode_sel[26]
+ padframe/mprj_io_in[26] padframe/mprj_io_inp_dis[26] padframe/mprj_io_out[26] padframe/mprj_io_oeb[26]
+ padframe/mprj_io_slow_sel[26] padframe/mprj_io_vtrip_sel[26] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[26\]/serial_data_in gpio_control_in\[27\]/serial_data_in
+ mprj/io_in[26] mprj/io_oeb[26] mprj/io_out[26] gpio_control_in\[26\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[33\] soc/mgmt_in_data[33] gpio_control_in\[33\]/one soc/mgmt_in_data[33]
+ gpio_control_in\[33\]/one padframe/mprj_io_analog_en[33] padframe/mprj_io_analog_pol[33]
+ padframe/mprj_io_analog_sel[33] padframe/mprj_io_dm[99] padframe/mprj_io_dm[100]
+ padframe/mprj_io_dm[101] padframe/mprj_io_holdover[33] padframe/mprj_io_ib_mode_sel[33]
+ padframe/mprj_io_in[33] padframe/mprj_io_inp_dis[33] padframe/mprj_io_out[33] padframe/mprj_io_oeb[33]
+ padframe/mprj_io_slow_sel[33] padframe/mprj_io_vtrip_sel[33] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[33\]/serial_data_in gpio_control_in\[34\]/serial_data_in
+ mprj/io_in[33] mprj/io_oeb[33] mprj/io_out[33] gpio_control_in\[33\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xsoc soc/clock soc/core_clk soc/resetb soc/flash_clk soc/flash_clk_ieb soc/flash_clk_oeb
+ soc/flash_csb soc/flash_csb_ieb soc/flash_csb_oeb soc/flash_io0_di soc/flash_io0_do
+ soc/flash_io0_ieb soc/flash_io0_oeb soc/flash_io1_di soc/flash_io1_do soc/flash_io1_ieb
+ soc/flash_io1_oeb soc/gpio_in_pad soc/gpio_inenb_pad soc/gpio_mode0_pad soc/gpio_mode1_pad
+ soc/gpio_out_pad soc/gpio_outenb_pad soc/jtag_out soc/jtag_outenb soc/la_input[0]
+ soc/la_input[100] soc/la_input[101] soc/la_input[102] soc/la_input[103] soc/la_input[104]
+ soc/la_input[105] soc/la_input[106] soc/la_input[107] soc/la_input[108] soc/la_input[109]
+ soc/la_input[10] soc/la_input[110] soc/la_input[111] soc/la_input[112] soc/la_input[113]
+ soc/la_input[114] soc/la_input[115] soc/la_input[116] soc/la_input[117] soc/la_input[118]
+ soc/la_input[119] soc/la_input[11] soc/la_input[120] soc/la_input[121] soc/la_input[122]
+ soc/la_input[123] soc/la_input[124] soc/la_input[125] soc/la_input[126] soc/la_input[127]
+ soc/la_input[12] soc/la_input[13] soc/la_input[14] soc/la_input[15] soc/la_input[16]
+ soc/la_input[17] soc/la_input[18] soc/la_input[19] soc/la_input[1] soc/la_input[20]
+ soc/la_input[21] soc/la_input[22] soc/la_input[23] soc/la_input[24] soc/la_input[25]
+ soc/la_input[26] soc/la_input[27] soc/la_input[28] soc/la_input[29] soc/la_input[2]
+ soc/la_input[30] soc/la_input[31] soc/la_input[32] soc/la_input[33] soc/la_input[34]
+ soc/la_input[35] soc/la_input[36] soc/la_input[37] soc/la_input[38] soc/la_input[39]
+ soc/la_input[3] soc/la_input[40] soc/la_input[41] soc/la_input[42] soc/la_input[43]
+ soc/la_input[44] soc/la_input[45] soc/la_input[46] soc/la_input[47] soc/la_input[48]
+ soc/la_input[49] soc/la_input[4] soc/la_input[50] soc/la_input[51] soc/la_input[52]
+ soc/la_input[53] soc/la_input[54] soc/la_input[55] soc/la_input[56] soc/la_input[57]
+ soc/la_input[58] soc/la_input[59] soc/la_input[5] soc/la_input[60] soc/la_input[61]
+ soc/la_input[62] soc/la_input[63] soc/la_input[64] soc/la_input[65] soc/la_input[66]
+ soc/la_input[67] soc/la_input[68] soc/la_input[69] soc/la_input[6] soc/la_input[70]
+ soc/la_input[71] soc/la_input[72] soc/la_input[73] soc/la_input[74] soc/la_input[75]
+ soc/la_input[76] soc/la_input[77] soc/la_input[78] soc/la_input[79] soc/la_input[7]
+ soc/la_input[80] soc/la_input[81] soc/la_input[82] soc/la_input[83] soc/la_input[84]
+ soc/la_input[85] soc/la_input[86] soc/la_input[87] soc/la_input[88] soc/la_input[89]
+ soc/la_input[8] soc/la_input[90] soc/la_input[91] soc/la_input[92] soc/la_input[93]
+ soc/la_input[94] soc/la_input[95] soc/la_input[96] soc/la_input[97] soc/la_input[98]
+ soc/la_input[99] soc/la_input[9] soc/la_oen[0] soc/la_oen[100] soc/la_oen[101] soc/la_oen[102]
+ soc/la_oen[103] soc/la_oen[104] soc/la_oen[105] soc/la_oen[106] soc/la_oen[107]
+ soc/la_oen[108] soc/la_oen[109] soc/la_oen[10] soc/la_oen[110] soc/la_oen[111] soc/la_oen[112]
+ soc/la_oen[113] soc/la_oen[114] soc/la_oen[115] soc/la_oen[116] soc/la_oen[117]
+ soc/la_oen[118] soc/la_oen[119] soc/la_oen[11] soc/la_oen[120] soc/la_oen[121] soc/la_oen[122]
+ soc/la_oen[123] soc/la_oen[124] soc/la_oen[125] soc/la_oen[126] soc/la_oen[127]
+ soc/la_oen[12] soc/la_oen[13] soc/la_oen[14] soc/la_oen[15] soc/la_oen[16] soc/la_oen[17]
+ soc/la_oen[18] soc/la_oen[19] soc/la_oen[1] soc/la_oen[20] soc/la_oen[21] soc/la_oen[22]
+ soc/la_oen[23] soc/la_oen[24] soc/la_oen[25] soc/la_oen[26] soc/la_oen[27] soc/la_oen[28]
+ soc/la_oen[29] soc/la_oen[2] soc/la_oen[30] soc/la_oen[31] soc/la_oen[32] soc/la_oen[33]
+ soc/la_oen[34] soc/la_oen[35] soc/la_oen[36] soc/la_oen[37] soc/la_oen[38] soc/la_oen[39]
+ soc/la_oen[3] soc/la_oen[40] soc/la_oen[41] soc/la_oen[42] soc/la_oen[43] soc/la_oen[44]
+ soc/la_oen[45] soc/la_oen[46] soc/la_oen[47] soc/la_oen[48] soc/la_oen[49] soc/la_oen[4]
+ soc/la_oen[50] soc/la_oen[51] soc/la_oen[52] soc/la_oen[53] soc/la_oen[54] soc/la_oen[55]
+ soc/la_oen[56] soc/la_oen[57] soc/la_oen[58] soc/la_oen[59] soc/la_oen[5] soc/la_oen[60]
+ soc/la_oen[61] soc/la_oen[62] soc/la_oen[63] soc/la_oen[64] soc/la_oen[65] soc/la_oen[66]
+ soc/la_oen[67] soc/la_oen[68] soc/la_oen[69] soc/la_oen[6] soc/la_oen[70] soc/la_oen[71]
+ soc/la_oen[72] soc/la_oen[73] soc/la_oen[74] soc/la_oen[75] soc/la_oen[76] soc/la_oen[77]
+ soc/la_oen[78] soc/la_oen[79] soc/la_oen[7] soc/la_oen[80] soc/la_oen[81] soc/la_oen[82]
+ soc/la_oen[83] soc/la_oen[84] soc/la_oen[85] soc/la_oen[86] soc/la_oen[87] soc/la_oen[88]
+ soc/la_oen[89] soc/la_oen[8] soc/la_oen[90] soc/la_oen[91] soc/la_oen[92] soc/la_oen[93]
+ soc/la_oen[94] soc/la_oen[95] soc/la_oen[96] soc/la_oen[97] soc/la_oen[98] soc/la_oen[99]
+ soc/la_oen[9] soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102]
+ soc/la_output[103] soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107]
+ soc/la_output[108] soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111]
+ soc/la_output[112] soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116]
+ soc/la_output[117] soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120]
+ soc/la_output[121] soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125]
+ soc/la_output[126] soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14]
+ soc/la_output[15] soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19]
+ soc/la_output[1] soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23]
+ soc/la_output[24] soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28]
+ soc/la_output[29] soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32]
+ soc/la_output[33] soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37]
+ soc/la_output[38] soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41]
+ soc/la_output[42] soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46]
+ soc/la_output[47] soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50]
+ soc/la_output[51] soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55]
+ soc/la_output[56] soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5]
+ soc/la_output[60] soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64]
+ soc/la_output[65] soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69]
+ soc/la_output[6] soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73]
+ soc/la_output[74] soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78]
+ soc/la_output[79] soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82]
+ soc/la_output[83] soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87]
+ soc/la_output[88] soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91]
+ soc/la_output[92] soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96]
+ soc/la_output[97] soc/la_output[98] soc/la_output[99] soc/la_output[9] soc/mask_rev[0]
+ soc/mask_rev[10] soc/mask_rev[11] soc/mask_rev[12] soc/mask_rev[13] soc/mask_rev[14]
+ soc/mask_rev[15] soc/mask_rev[16] soc/mask_rev[17] soc/mask_rev[18] soc/mask_rev[19]
+ soc/mask_rev[1] soc/mask_rev[20] soc/mask_rev[21] soc/mask_rev[22] soc/mask_rev[23]
+ soc/mask_rev[24] soc/mask_rev[25] soc/mask_rev[26] soc/mask_rev[27] soc/mask_rev[28]
+ soc/mask_rev[29] soc/mask_rev[2] soc/mask_rev[30] soc/mask_rev[31] soc/mask_rev[3]
+ soc/mask_rev[4] soc/mask_rev[5] soc/mask_rev[6] soc/mask_rev[7] soc/mask_rev[8]
+ soc/mask_rev[9] soc/mgmt_addr[0] soc/mgmt_addr[1] soc/mgmt_addr[2] soc/mgmt_addr[3]
+ soc/mgmt_addr[4] soc/mgmt_addr[5] soc/mgmt_addr[6] soc/mgmt_addr[7] soc/mgmt_addr_ro[0]
+ soc/mgmt_addr_ro[1] soc/mgmt_addr_ro[2] soc/mgmt_addr_ro[3] soc/mgmt_addr_ro[4]
+ soc/mgmt_addr_ro[5] soc/mgmt_addr_ro[6] soc/mgmt_addr_ro[7] soc/mgmt_ena[0] soc/mgmt_ena[1]
+ soc/mgmt_ena_ro soc/mgmt_in_data[0] soc/mgmt_in_data[10] soc/mgmt_in_data[11] soc/mgmt_in_data[12]
+ soc/mgmt_in_data[13] soc/mgmt_in_data[14] soc/mgmt_in_data[15] soc/mgmt_in_data[16]
+ soc/mgmt_in_data[17] soc/mgmt_in_data[18] soc/mgmt_in_data[19] soc/mgmt_in_data[1]
+ soc/mgmt_in_data[20] soc/mgmt_in_data[21] soc/mgmt_in_data[22] soc/mgmt_in_data[23]
+ soc/mgmt_in_data[24] soc/mgmt_in_data[25] soc/mgmt_in_data[26] soc/mgmt_in_data[27]
+ soc/mgmt_in_data[28] soc/mgmt_in_data[29] soc/mgmt_in_data[2] soc/mgmt_in_data[30]
+ soc/mgmt_in_data[31] soc/mgmt_in_data[32] soc/mgmt_in_data[33] soc/mgmt_in_data[34]
+ soc/mgmt_in_data[35] soc/mgmt_in_data[36] soc/mgmt_in_data[37] soc/mgmt_in_data[3]
+ soc/mgmt_in_data[4] soc/mgmt_in_data[5] soc/mgmt_in_data[6] soc/mgmt_in_data[7]
+ soc/mgmt_in_data[8] soc/mgmt_in_data[9] soc/mgmt_out_data[0] soc/mgmt_in_data[10]
+ soc/mgmt_in_data[11] soc/mgmt_in_data[12] soc/mgmt_in_data[13] soc/mgmt_in_data[14]
+ soc/mgmt_in_data[15] soc/mgmt_in_data[16] soc/mgmt_in_data[17] soc/mgmt_in_data[18]
+ soc/mgmt_in_data[19] soc/mgmt_out_data[1] soc/mgmt_in_data[20] soc/mgmt_in_data[21]
+ soc/mgmt_in_data[22] soc/mgmt_in_data[23] soc/mgmt_in_data[24] soc/mgmt_in_data[25]
+ soc/mgmt_in_data[26] soc/mgmt_in_data[27] soc/mgmt_in_data[28] soc/mgmt_in_data[29]
+ soc/mgmt_in_data[2] soc/mgmt_in_data[30] soc/mgmt_in_data[31] soc/mgmt_in_data[32]
+ soc/mgmt_in_data[33] soc/mgmt_in_data[34] soc/mgmt_in_data[35] soc/mgmt_in_data[36]
+ soc/mgmt_in_data[37] soc/mgmt_in_data[3] soc/mgmt_in_data[4] soc/mgmt_in_data[5]
+ soc/mgmt_in_data[6] soc/mgmt_in_data[7] soc/mgmt_in_data[8] soc/mgmt_in_data[9]
+ soc/mgmt_rdata[0] soc/mgmt_rdata[10] soc/mgmt_rdata[11] soc/mgmt_rdata[12] soc/mgmt_rdata[13]
+ soc/mgmt_rdata[14] soc/mgmt_rdata[15] soc/mgmt_rdata[16] soc/mgmt_rdata[17] soc/mgmt_rdata[18]
+ soc/mgmt_rdata[19] soc/mgmt_rdata[1] soc/mgmt_rdata[20] soc/mgmt_rdata[21] soc/mgmt_rdata[22]
+ soc/mgmt_rdata[23] soc/mgmt_rdata[24] soc/mgmt_rdata[25] soc/mgmt_rdata[26] soc/mgmt_rdata[27]
+ soc/mgmt_rdata[28] soc/mgmt_rdata[29] soc/mgmt_rdata[2] soc/mgmt_rdata[30] soc/mgmt_rdata[31]
+ soc/mgmt_rdata[32] soc/mgmt_rdata[33] soc/mgmt_rdata[34] soc/mgmt_rdata[35] soc/mgmt_rdata[36]
+ soc/mgmt_rdata[37] soc/mgmt_rdata[38] soc/mgmt_rdata[39] soc/mgmt_rdata[3] soc/mgmt_rdata[40]
+ soc/mgmt_rdata[41] soc/mgmt_rdata[42] soc/mgmt_rdata[43] soc/mgmt_rdata[44] soc/mgmt_rdata[45]
+ soc/mgmt_rdata[46] soc/mgmt_rdata[47] soc/mgmt_rdata[48] soc/mgmt_rdata[49] soc/mgmt_rdata[4]
+ soc/mgmt_rdata[50] soc/mgmt_rdata[51] soc/mgmt_rdata[52] soc/mgmt_rdata[53] soc/mgmt_rdata[54]
+ soc/mgmt_rdata[55] soc/mgmt_rdata[56] soc/mgmt_rdata[57] soc/mgmt_rdata[58] soc/mgmt_rdata[59]
+ soc/mgmt_rdata[5] soc/mgmt_rdata[60] soc/mgmt_rdata[61] soc/mgmt_rdata[62] soc/mgmt_rdata[63]
+ soc/mgmt_rdata[6] soc/mgmt_rdata[7] soc/mgmt_rdata[8] soc/mgmt_rdata[9] soc/mgmt_rdata_ro[0]
+ soc/mgmt_rdata_ro[10] soc/mgmt_rdata_ro[11] soc/mgmt_rdata_ro[12] soc/mgmt_rdata_ro[13]
+ soc/mgmt_rdata_ro[14] soc/mgmt_rdata_ro[15] soc/mgmt_rdata_ro[16] soc/mgmt_rdata_ro[17]
+ soc/mgmt_rdata_ro[18] soc/mgmt_rdata_ro[19] soc/mgmt_rdata_ro[1] soc/mgmt_rdata_ro[20]
+ soc/mgmt_rdata_ro[21] soc/mgmt_rdata_ro[22] soc/mgmt_rdata_ro[23] soc/mgmt_rdata_ro[24]
+ soc/mgmt_rdata_ro[25] soc/mgmt_rdata_ro[26] soc/mgmt_rdata_ro[27] soc/mgmt_rdata_ro[28]
+ soc/mgmt_rdata_ro[29] soc/mgmt_rdata_ro[2] soc/mgmt_rdata_ro[30] soc/mgmt_rdata_ro[31]
+ soc/mgmt_rdata_ro[3] soc/mgmt_rdata_ro[4] soc/mgmt_rdata_ro[5] soc/mgmt_rdata_ro[6]
+ soc/mgmt_rdata_ro[7] soc/mgmt_rdata_ro[8] soc/mgmt_rdata_ro[9] soc/mgmt_wdata[0]
+ soc/mgmt_wdata[10] soc/mgmt_wdata[11] soc/mgmt_wdata[12] soc/mgmt_wdata[13] soc/mgmt_wdata[14]
+ soc/mgmt_wdata[15] soc/mgmt_wdata[16] soc/mgmt_wdata[17] soc/mgmt_wdata[18] soc/mgmt_wdata[19]
+ soc/mgmt_wdata[1] soc/mgmt_wdata[20] soc/mgmt_wdata[21] soc/mgmt_wdata[22] soc/mgmt_wdata[23]
+ soc/mgmt_wdata[24] soc/mgmt_wdata[25] soc/mgmt_wdata[26] soc/mgmt_wdata[27] soc/mgmt_wdata[28]
+ soc/mgmt_wdata[29] soc/mgmt_wdata[2] soc/mgmt_wdata[30] soc/mgmt_wdata[31] soc/mgmt_wdata[3]
+ soc/mgmt_wdata[4] soc/mgmt_wdata[5] soc/mgmt_wdata[6] soc/mgmt_wdata[7] soc/mgmt_wdata[8]
+ soc/mgmt_wdata[9] soc/mgmt_wen[0] soc/mgmt_wen[1] soc/mgmt_wen_mask[0] soc/mgmt_wen_mask[1]
+ soc/mgmt_wen_mask[2] soc/mgmt_wen_mask[3] soc/mgmt_wen_mask[4] soc/mgmt_wen_mask[5]
+ soc/mgmt_wen_mask[6] soc/mgmt_wen_mask[7] soc/mprj2_vcc_pwrgood soc/mprj2_vdd_pwrgood
+ soc/mprj_ack_i soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11] soc/mprj_adr_o[12]
+ soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16] soc/mprj_adr_o[17]
+ soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20] soc/mprj_adr_o[21]
+ soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25] soc/mprj_adr_o[26]
+ soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2] soc/mprj_adr_o[30]
+ soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5] soc/mprj_adr_o[6]
+ soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] soc/mprj_cyc_o soc/mprj_dat_i[0]
+ soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12] soc/mprj_dat_i[13] soc/mprj_dat_i[14]
+ soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17] soc/mprj_dat_i[18] soc/mprj_dat_i[19]
+ soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21] soc/mprj_dat_i[22] soc/mprj_dat_i[23]
+ soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26] soc/mprj_dat_i[27] soc/mprj_dat_i[28]
+ soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30] soc/mprj_dat_i[31] soc/mprj_dat_i[3]
+ soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6] soc/mprj_dat_i[7] soc/mprj_dat_i[8]
+ soc/mprj_dat_i[9] soc/mprj_dat_o[0] soc/mprj_dat_o[10] soc/mprj_dat_o[11] soc/mprj_dat_o[12]
+ soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15] soc/mprj_dat_o[16] soc/mprj_dat_o[17]
+ soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1] soc/mprj_dat_o[20] soc/mprj_dat_o[21]
+ soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24] soc/mprj_dat_o[25] soc/mprj_dat_o[26]
+ soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29] soc/mprj_dat_o[2] soc/mprj_dat_o[30]
+ soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4] soc/mprj_dat_o[5] soc/mprj_dat_o[6]
+ soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9] soc/mprj_io_loader_clock soc/mprj_io_loader_data
+ soc/mprj_io_loader_resetn soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2]
+ soc/mprj_sel_o[3] soc/mprj_stb_o soc/mprj_vcc_pwrgood soc/mprj_vdd_pwrgood soc/mprj_we_o
+ soc/porb pwr_ctrl_out[0] pwr_ctrl_out[1] pwr_ctrl_out[2] pwr_ctrl_out[3] soc/resetb
+ soc/sdo_out soc/sdo_outenb soc/user_clk vccd vssd mgmt_core
Xgpio_control_in\[19\] soc/mgmt_in_data[19] gpio_control_in\[19\]/one soc/mgmt_in_data[19]
+ gpio_control_in\[19\]/one padframe/mprj_io_analog_en[19] padframe/mprj_io_analog_pol[19]
+ padframe/mprj_io_analog_sel[19] padframe/mprj_io_dm[57] padframe/mprj_io_dm[58]
+ padframe/mprj_io_dm[59] padframe/mprj_io_holdover[19] padframe/mprj_io_ib_mode_sel[19]
+ padframe/mprj_io_in[19] padframe/mprj_io_inp_dis[19] padframe/mprj_io_out[19] padframe/mprj_io_oeb[19]
+ padframe/mprj_io_slow_sel[19] padframe/mprj_io_vtrip_sel[19] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[19\]/serial_data_in gpio_control_in\[20\]/serial_data_in
+ mprj/io_in[19] mprj/io_oeb[19] mprj/io_out[19] gpio_control_in\[19\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[31\] soc/mgmt_in_data[31] gpio_control_in\[31\]/one soc/mgmt_in_data[31]
+ gpio_control_in\[31\]/one padframe/mprj_io_analog_en[31] padframe/mprj_io_analog_pol[31]
+ padframe/mprj_io_analog_sel[31] padframe/mprj_io_dm[93] padframe/mprj_io_dm[94]
+ padframe/mprj_io_dm[95] padframe/mprj_io_holdover[31] padframe/mprj_io_ib_mode_sel[31]
+ padframe/mprj_io_in[31] padframe/mprj_io_inp_dis[31] padframe/mprj_io_out[31] padframe/mprj_io_oeb[31]
+ padframe/mprj_io_slow_sel[31] padframe/mprj_io_vtrip_sel[31] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[31\]/serial_data_in gpio_control_in\[32\]/serial_data_in
+ mprj/io_in[31] mprj/io_oeb[31] mprj/io_out[31] gpio_control_in\[31\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xpor vddio vccd vssio por/porb_h por/por_l soc/porb simple_por
Xgpio_control_in\[24\] soc/mgmt_in_data[24] gpio_control_in\[24\]/one soc/mgmt_in_data[24]
+ gpio_control_in\[24\]/one padframe/mprj_io_analog_en[24] padframe/mprj_io_analog_pol[24]
+ padframe/mprj_io_analog_sel[24] padframe/mprj_io_dm[72] padframe/mprj_io_dm[73]
+ padframe/mprj_io_dm[74] padframe/mprj_io_holdover[24] padframe/mprj_io_ib_mode_sel[24]
+ padframe/mprj_io_in[24] padframe/mprj_io_inp_dis[24] padframe/mprj_io_out[24] padframe/mprj_io_oeb[24]
+ padframe/mprj_io_slow_sel[24] padframe/mprj_io_vtrip_sel[24] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[24\]/serial_data_in gpio_control_in\[25\]/serial_data_in
+ mprj/io_in[24] mprj/io_oeb[24] mprj/io_out[24] gpio_control_in\[24\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_bidir\[1\] soc/mgmt_in_data[1] soc/sdo_outenb soc/sdo_out gpio_control_bidir\[1\]/one
+ padframe/mprj_io_analog_en[1] padframe/mprj_io_analog_pol[1] padframe/mprj_io_analog_sel[1]
+ padframe/mprj_io_dm[3] padframe/mprj_io_dm[4] padframe/mprj_io_dm[5] padframe/mprj_io_holdover[1]
+ padframe/mprj_io_ib_mode_sel[1] padframe/mprj_io_in[1] padframe/mprj_io_inp_dis[1]
+ padframe/mprj_io_out[1] padframe/mprj_io_oeb[1] padframe/mprj_io_slow_sel[1] padframe/mprj_io_vtrip_sel[1]
+ soc/mprj_io_loader_resetn soc/mprj_io_loader_clock gpio_control_bidir\[1\]/serial_data_in
+ gpio_control_in\[2\]/serial_data_in mprj/io_in[1] mprj/io_oeb[1] mprj/io_out[1]
+ gpio_control_bidir\[1\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[17\] soc/mgmt_in_data[17] gpio_control_in\[17\]/one soc/mgmt_in_data[17]
+ gpio_control_in\[17\]/one padframe/mprj_io_analog_en[17] padframe/mprj_io_analog_pol[17]
+ padframe/mprj_io_analog_sel[17] padframe/mprj_io_dm[51] padframe/mprj_io_dm[52]
+ padframe/mprj_io_dm[53] padframe/mprj_io_holdover[17] padframe/mprj_io_ib_mode_sel[17]
+ padframe/mprj_io_in[17] padframe/mprj_io_inp_dis[17] padframe/mprj_io_out[17] padframe/mprj_io_oeb[17]
+ padframe/mprj_io_slow_sel[17] padframe/mprj_io_vtrip_sel[17] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[17\]/serial_data_in gpio_control_in\[18\]/serial_data_in
+ mprj/io_in[17] mprj/io_oeb[17] mprj/io_out[17] gpio_control_in\[17\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[22\] soc/mgmt_in_data[22] gpio_control_in\[22\]/one soc/mgmt_in_data[22]
+ gpio_control_in\[22\]/one padframe/mprj_io_analog_en[22] padframe/mprj_io_analog_pol[22]
+ padframe/mprj_io_analog_sel[22] padframe/mprj_io_dm[66] padframe/mprj_io_dm[67]
+ padframe/mprj_io_dm[68] padframe/mprj_io_holdover[22] padframe/mprj_io_ib_mode_sel[22]
+ padframe/mprj_io_in[22] padframe/mprj_io_inp_dis[22] padframe/mprj_io_out[22] padframe/mprj_io_oeb[22]
+ padframe/mprj_io_slow_sel[22] padframe/mprj_io_vtrip_sel[22] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[22\]/serial_data_in gpio_control_in\[23\]/serial_data_in
+ mprj/io_in[22] mprj/io_oeb[22] mprj/io_out[22] gpio_control_in\[22\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[8\] soc/mgmt_in_data[8] gpio_control_in\[8\]/one soc/mgmt_in_data[8]
+ gpio_control_in\[8\]/one padframe/mprj_io_analog_en[8] padframe/mprj_io_analog_pol[8]
+ padframe/mprj_io_analog_sel[8] padframe/mprj_io_dm[24] padframe/mprj_io_dm[25] padframe/mprj_io_dm[26]
+ padframe/mprj_io_holdover[8] padframe/mprj_io_ib_mode_sel[8] padframe/mprj_io_in[8]
+ padframe/mprj_io_inp_dis[8] padframe/mprj_io_out[8] padframe/mprj_io_oeb[8] padframe/mprj_io_slow_sel[8]
+ padframe/mprj_io_vtrip_sel[8] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[8\]/serial_data_in gpio_control_in\[9\]/serial_data_in mprj/io_in[8]
+ mprj/io_oeb[8] mprj/io_out[8] gpio_control_in\[8\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[15\] soc/mgmt_in_data[15] gpio_control_in\[15\]/one soc/mgmt_in_data[15]
+ gpio_control_in\[15\]/one padframe/mprj_io_analog_en[15] padframe/mprj_io_analog_pol[15]
+ padframe/mprj_io_analog_sel[15] padframe/mprj_io_dm[45] padframe/mprj_io_dm[46]
+ padframe/mprj_io_dm[47] padframe/mprj_io_holdover[15] padframe/mprj_io_ib_mode_sel[15]
+ padframe/mprj_io_in[15] padframe/mprj_io_inp_dis[15] padframe/mprj_io_out[15] padframe/mprj_io_oeb[15]
+ padframe/mprj_io_slow_sel[15] padframe/mprj_io_vtrip_sel[15] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[15\]/serial_data_in gpio_control_in\[16\]/serial_data_in
+ mprj/io_in[15] mprj/io_oeb[15] mprj/io_out[15] gpio_control_in\[15\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xuser_id_value soc/mask_rev[0] soc/mask_rev[10] soc/mask_rev[11] soc/mask_rev[12]
+ soc/mask_rev[13] soc/mask_rev[14] soc/mask_rev[15] soc/mask_rev[16] soc/mask_rev[17]
+ soc/mask_rev[18] soc/mask_rev[19] soc/mask_rev[1] soc/mask_rev[20] soc/mask_rev[21]
+ soc/mask_rev[22] soc/mask_rev[23] soc/mask_rev[24] soc/mask_rev[25] soc/mask_rev[26]
+ soc/mask_rev[27] soc/mask_rev[28] soc/mask_rev[29] soc/mask_rev[2] soc/mask_rev[30]
+ soc/mask_rev[31] soc/mask_rev[3] soc/mask_rev[4] soc/mask_rev[5] soc/mask_rev[6]
+ soc/mask_rev[7] soc/mask_rev[8] soc/mask_rev[9] vccd vssd user_id_programming
Xgpio_control_in\[20\] soc/mgmt_in_data[20] gpio_control_in\[20\]/one soc/mgmt_in_data[20]
+ gpio_control_in\[20\]/one padframe/mprj_io_analog_en[20] padframe/mprj_io_analog_pol[20]
+ padframe/mprj_io_analog_sel[20] padframe/mprj_io_dm[60] padframe/mprj_io_dm[61]
+ padframe/mprj_io_dm[62] padframe/mprj_io_holdover[20] padframe/mprj_io_ib_mode_sel[20]
+ padframe/mprj_io_in[20] padframe/mprj_io_inp_dis[20] padframe/mprj_io_out[20] padframe/mprj_io_oeb[20]
+ padframe/mprj_io_slow_sel[20] padframe/mprj_io_vtrip_sel[20] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[20\]/serial_data_in gpio_control_in\[21\]/serial_data_in
+ mprj/io_in[20] mprj/io_oeb[20] mprj/io_out[20] gpio_control_in\[20\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[6\] soc/mgmt_in_data[6] gpio_control_in\[6\]/one soc/mgmt_in_data[6]
+ gpio_control_in\[6\]/one padframe/mprj_io_analog_en[6] padframe/mprj_io_analog_pol[6]
+ padframe/mprj_io_analog_sel[6] padframe/mprj_io_dm[18] padframe/mprj_io_dm[19] padframe/mprj_io_dm[20]
+ padframe/mprj_io_holdover[6] padframe/mprj_io_ib_mode_sel[6] padframe/mprj_io_in[6]
+ padframe/mprj_io_inp_dis[6] padframe/mprj_io_out[6] padframe/mprj_io_oeb[6] padframe/mprj_io_slow_sel[6]
+ padframe/mprj_io_vtrip_sel[6] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[6\]/serial_data_in gpio_control_in\[7\]/serial_data_in mprj/io_in[6]
+ mprj/io_oeb[6] mprj/io_out[6] gpio_control_in\[6\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[13\] soc/mgmt_in_data[13] gpio_control_in\[13\]/one soc/mgmt_in_data[13]
+ gpio_control_in\[13\]/one padframe/mprj_io_analog_en[13] padframe/mprj_io_analog_pol[13]
+ padframe/mprj_io_analog_sel[13] padframe/mprj_io_dm[39] padframe/mprj_io_dm[40]
+ padframe/mprj_io_dm[41] padframe/mprj_io_holdover[13] padframe/mprj_io_ib_mode_sel[13]
+ padframe/mprj_io_in[13] padframe/mprj_io_inp_dis[13] padframe/mprj_io_out[13] padframe/mprj_io_oeb[13]
+ padframe/mprj_io_slow_sel[13] padframe/mprj_io_vtrip_sel[13] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[13\]/serial_data_in gpio_control_in\[14\]/serial_data_in
+ mprj/io_in[13] mprj/io_oeb[13] mprj/io_out[13] gpio_control_in\[13\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[36\] soc/mgmt_in_data[36] gpio_control_in\[36\]/one soc/mgmt_in_data[36]
+ gpio_control_in\[36\]/one padframe/mprj_io_analog_en[36] padframe/mprj_io_analog_pol[36]
+ padframe/mprj_io_analog_sel[36] padframe/mprj_io_dm[108] padframe/mprj_io_dm[109]
+ padframe/mprj_io_dm[110] padframe/mprj_io_holdover[36] padframe/mprj_io_ib_mode_sel[36]
+ padframe/mprj_io_in[36] padframe/mprj_io_inp_dis[36] padframe/mprj_io_out[36] padframe/mprj_io_oeb[36]
+ padframe/mprj_io_slow_sel[36] padframe/mprj_io_vtrip_sel[36] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[36\]/serial_data_in gpio_control_in\[37\]/serial_data_in
+ mprj/io_in[36] mprj/io_oeb[36] mprj/io_out[36] gpio_control_in\[36\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[29\] soc/mgmt_in_data[29] gpio_control_in\[29\]/one soc/mgmt_in_data[29]
+ gpio_control_in\[29\]/one padframe/mprj_io_analog_en[29] padframe/mprj_io_analog_pol[29]
+ padframe/mprj_io_analog_sel[29] padframe/mprj_io_dm[87] padframe/mprj_io_dm[88]
+ padframe/mprj_io_dm[89] padframe/mprj_io_holdover[29] padframe/mprj_io_ib_mode_sel[29]
+ padframe/mprj_io_in[29] padframe/mprj_io_inp_dis[29] padframe/mprj_io_out[29] padframe/mprj_io_oeb[29]
+ padframe/mprj_io_slow_sel[29] padframe/mprj_io_vtrip_sel[29] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[29\]/serial_data_in gpio_control_in\[30\]/serial_data_in
+ mprj/io_in[29] mprj/io_oeb[29] mprj/io_out[29] gpio_control_in\[29\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[4\] soc/mgmt_in_data[4] gpio_control_in\[4\]/one soc/mgmt_in_data[4]
+ gpio_control_in\[4\]/one padframe/mprj_io_analog_en[4] padframe/mprj_io_analog_pol[4]
+ padframe/mprj_io_analog_sel[4] padframe/mprj_io_dm[12] padframe/mprj_io_dm[13] padframe/mprj_io_dm[14]
+ padframe/mprj_io_holdover[4] padframe/mprj_io_ib_mode_sel[4] padframe/mprj_io_in[4]
+ padframe/mprj_io_inp_dis[4] padframe/mprj_io_out[4] padframe/mprj_io_oeb[4] padframe/mprj_io_slow_sel[4]
+ padframe/mprj_io_vtrip_sel[4] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[4\]/serial_data_in gpio_control_in\[5\]/serial_data_in mprj/io_in[4]
+ mprj/io_oeb[4] mprj/io_out[4] gpio_control_in\[4\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[11\] soc/mgmt_in_data[11] gpio_control_in\[11\]/one soc/mgmt_in_data[11]
+ gpio_control_in\[11\]/one padframe/mprj_io_analog_en[11] padframe/mprj_io_analog_pol[11]
+ padframe/mprj_io_analog_sel[11] padframe/mprj_io_dm[33] padframe/mprj_io_dm[34]
+ padframe/mprj_io_dm[35] padframe/mprj_io_holdover[11] padframe/mprj_io_ib_mode_sel[11]
+ padframe/mprj_io_in[11] padframe/mprj_io_inp_dis[11] padframe/mprj_io_out[11] padframe/mprj_io_oeb[11]
+ padframe/mprj_io_slow_sel[11] padframe/mprj_io_vtrip_sel[11] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[11\]/serial_data_in gpio_control_in\[12\]/serial_data_in
+ mprj/io_in[11] mprj/io_oeb[11] mprj/io_out[11] gpio_control_in\[11\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[34\] soc/mgmt_in_data[34] gpio_control_in\[34\]/one soc/mgmt_in_data[34]
+ gpio_control_in\[34\]/one padframe/mprj_io_analog_en[34] padframe/mprj_io_analog_pol[34]
+ padframe/mprj_io_analog_sel[34] padframe/mprj_io_dm[102] padframe/mprj_io_dm[103]
+ padframe/mprj_io_dm[104] padframe/mprj_io_holdover[34] padframe/mprj_io_ib_mode_sel[34]
+ padframe/mprj_io_in[34] padframe/mprj_io_inp_dis[34] padframe/mprj_io_out[34] padframe/mprj_io_oeb[34]
+ padframe/mprj_io_slow_sel[34] padframe/mprj_io_vtrip_sel[34] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[34\]/serial_data_in gpio_control_in\[35\]/serial_data_in
+ mprj/io_in[34] mprj/io_oeb[34] mprj/io_out[34] gpio_control_in\[34\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xmgmt_buffers soc/core_clk soc/user_clk soc/resetb mprj/la_data_in[0] mprj/la_data_in[100]
+ mprj/la_data_in[101] mprj/la_data_in[102] mprj/la_data_in[103] mprj/la_data_in[104]
+ mprj/la_data_in[105] mprj/la_data_in[106] mprj/la_data_in[107] mprj/la_data_in[108]
+ mprj/la_data_in[109] mprj/la_data_in[10] mprj/la_data_in[110] mprj/la_data_in[111]
+ mprj/la_data_in[112] mprj/la_data_in[113] mprj/la_data_in[114] mprj/la_data_in[115]
+ mprj/la_data_in[116] mprj/la_data_in[117] mprj/la_data_in[118] mprj/la_data_in[119]
+ mprj/la_data_in[11] mprj/la_data_in[120] mprj/la_data_in[121] mprj/la_data_in[122]
+ mprj/la_data_in[123] mprj/la_data_in[124] mprj/la_data_in[125] mprj/la_data_in[126]
+ mprj/la_data_in[127] mprj/la_data_in[12] mprj/la_data_in[13] mprj/la_data_in[14]
+ mprj/la_data_in[15] mprj/la_data_in[16] mprj/la_data_in[17] mprj/la_data_in[18]
+ mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20] mprj/la_data_in[21] mprj/la_data_in[22]
+ mprj/la_data_in[23] mprj/la_data_in[24] mprj/la_data_in[25] mprj/la_data_in[26]
+ mprj/la_data_in[27] mprj/la_data_in[28] mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30]
+ mprj/la_data_in[31] mprj/la_data_in[32] mprj/la_data_in[33] mprj/la_data_in[34]
+ mprj/la_data_in[35] mprj/la_data_in[36] mprj/la_data_in[37] mprj/la_data_in[38]
+ mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40] mprj/la_data_in[41] mprj/la_data_in[42]
+ mprj/la_data_in[43] mprj/la_data_in[44] mprj/la_data_in[45] mprj/la_data_in[46]
+ mprj/la_data_in[47] mprj/la_data_in[48] mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50]
+ mprj/la_data_in[51] mprj/la_data_in[52] mprj/la_data_in[53] mprj/la_data_in[54]
+ mprj/la_data_in[55] mprj/la_data_in[56] mprj/la_data_in[57] mprj/la_data_in[58]
+ mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60] mprj/la_data_in[61] mprj/la_data_in[62]
+ mprj/la_data_in[63] mprj/la_data_in[64] mprj/la_data_in[65] mprj/la_data_in[66]
+ mprj/la_data_in[67] mprj/la_data_in[68] mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70]
+ mprj/la_data_in[71] mprj/la_data_in[72] mprj/la_data_in[73] mprj/la_data_in[74]
+ mprj/la_data_in[75] mprj/la_data_in[76] mprj/la_data_in[77] mprj/la_data_in[78]
+ mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80] mprj/la_data_in[81] mprj/la_data_in[82]
+ mprj/la_data_in[83] mprj/la_data_in[84] mprj/la_data_in[85] mprj/la_data_in[86]
+ mprj/la_data_in[87] mprj/la_data_in[88] mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90]
+ mprj/la_data_in[91] mprj/la_data_in[92] mprj/la_data_in[93] mprj/la_data_in[94]
+ mprj/la_data_in[95] mprj/la_data_in[96] mprj/la_data_in[97] mprj/la_data_in[98]
+ mprj/la_data_in[99] mprj/la_data_in[9] soc/la_input[0] soc/la_input[100] soc/la_input[101]
+ soc/la_input[102] soc/la_input[103] soc/la_input[104] soc/la_input[105] soc/la_input[106]
+ soc/la_input[107] soc/la_input[108] soc/la_input[109] soc/la_input[10] soc/la_input[110]
+ soc/la_input[111] soc/la_input[112] soc/la_input[113] soc/la_input[114] soc/la_input[115]
+ soc/la_input[116] soc/la_input[117] soc/la_input[118] soc/la_input[119] soc/la_input[11]
+ soc/la_input[120] soc/la_input[121] soc/la_input[122] soc/la_input[123] soc/la_input[124]
+ soc/la_input[125] soc/la_input[126] soc/la_input[127] soc/la_input[12] soc/la_input[13]
+ soc/la_input[14] soc/la_input[15] soc/la_input[16] soc/la_input[17] soc/la_input[18]
+ soc/la_input[19] soc/la_input[1] soc/la_input[20] soc/la_input[21] soc/la_input[22]
+ soc/la_input[23] soc/la_input[24] soc/la_input[25] soc/la_input[26] soc/la_input[27]
+ soc/la_input[28] soc/la_input[29] soc/la_input[2] soc/la_input[30] soc/la_input[31]
+ soc/la_input[32] soc/la_input[33] soc/la_input[34] soc/la_input[35] soc/la_input[36]
+ soc/la_input[37] soc/la_input[38] soc/la_input[39] soc/la_input[3] soc/la_input[40]
+ soc/la_input[41] soc/la_input[42] soc/la_input[43] soc/la_input[44] soc/la_input[45]
+ soc/la_input[46] soc/la_input[47] soc/la_input[48] soc/la_input[49] soc/la_input[4]
+ soc/la_input[50] soc/la_input[51] soc/la_input[52] soc/la_input[53] soc/la_input[54]
+ soc/la_input[55] soc/la_input[56] soc/la_input[57] soc/la_input[58] soc/la_input[59]
+ soc/la_input[5] soc/la_input[60] soc/la_input[61] soc/la_input[62] soc/la_input[63]
+ soc/la_input[64] soc/la_input[65] soc/la_input[66] soc/la_input[67] soc/la_input[68]
+ soc/la_input[69] soc/la_input[6] soc/la_input[70] soc/la_input[71] soc/la_input[72]
+ soc/la_input[73] soc/la_input[74] soc/la_input[75] soc/la_input[76] soc/la_input[77]
+ soc/la_input[78] soc/la_input[79] soc/la_input[7] soc/la_input[80] soc/la_input[81]
+ soc/la_input[82] soc/la_input[83] soc/la_input[84] soc/la_input[85] soc/la_input[86]
+ soc/la_input[87] soc/la_input[88] soc/la_input[89] soc/la_input[8] soc/la_input[90]
+ soc/la_input[91] soc/la_input[92] soc/la_input[93] soc/la_input[94] soc/la_input[95]
+ soc/la_input[96] soc/la_input[97] soc/la_input[98] soc/la_input[99] soc/la_input[9]
+ mprj/la_data_out[0] mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102]
+ mprj/la_data_out[103] mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106]
+ mprj/la_data_out[107] mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10]
+ mprj/la_data_out[110] mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113]
+ mprj/la_data_out[114] mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117]
+ mprj/la_data_out[118] mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120]
+ mprj/la_data_out[121] mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124]
+ mprj/la_data_out[125] mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12]
+ mprj/la_data_out[13] mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16]
+ mprj/la_data_out[17] mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1]
+ mprj/la_data_out[20] mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23]
+ mprj/la_data_out[24] mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27]
+ mprj/la_data_out[28] mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30]
+ mprj/la_data_out[31] mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34]
+ mprj/la_data_out[35] mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38]
+ mprj/la_data_out[39] mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41]
+ mprj/la_data_out[42] mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45]
+ mprj/la_data_out[46] mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49]
+ mprj/la_data_out[4] mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52]
+ mprj/la_data_out[53] mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56]
+ mprj/la_data_out[57] mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5]
+ mprj/la_data_out[60] mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63]
+ mprj/la_data_out[64] mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67]
+ mprj/la_data_out[68] mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70]
+ mprj/la_data_out[71] mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74]
+ mprj/la_data_out[75] mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78]
+ mprj/la_data_out[79] mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81]
+ mprj/la_data_out[82] mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85]
+ mprj/la_data_out[86] mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89]
+ mprj/la_data_out[8] mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92]
+ mprj/la_data_out[93] mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96]
+ mprj/la_data_out[97] mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9]
+ soc/la_output[0] soc/la_output[100] soc/la_output[101] soc/la_output[102] soc/la_output[103]
+ soc/la_output[104] soc/la_output[105] soc/la_output[106] soc/la_output[107] soc/la_output[108]
+ soc/la_output[109] soc/la_output[10] soc/la_output[110] soc/la_output[111] soc/la_output[112]
+ soc/la_output[113] soc/la_output[114] soc/la_output[115] soc/la_output[116] soc/la_output[117]
+ soc/la_output[118] soc/la_output[119] soc/la_output[11] soc/la_output[120] soc/la_output[121]
+ soc/la_output[122] soc/la_output[123] soc/la_output[124] soc/la_output[125] soc/la_output[126]
+ soc/la_output[127] soc/la_output[12] soc/la_output[13] soc/la_output[14] soc/la_output[15]
+ soc/la_output[16] soc/la_output[17] soc/la_output[18] soc/la_output[19] soc/la_output[1]
+ soc/la_output[20] soc/la_output[21] soc/la_output[22] soc/la_output[23] soc/la_output[24]
+ soc/la_output[25] soc/la_output[26] soc/la_output[27] soc/la_output[28] soc/la_output[29]
+ soc/la_output[2] soc/la_output[30] soc/la_output[31] soc/la_output[32] soc/la_output[33]
+ soc/la_output[34] soc/la_output[35] soc/la_output[36] soc/la_output[37] soc/la_output[38]
+ soc/la_output[39] soc/la_output[3] soc/la_output[40] soc/la_output[41] soc/la_output[42]
+ soc/la_output[43] soc/la_output[44] soc/la_output[45] soc/la_output[46] soc/la_output[47]
+ soc/la_output[48] soc/la_output[49] soc/la_output[4] soc/la_output[50] soc/la_output[51]
+ soc/la_output[52] soc/la_output[53] soc/la_output[54] soc/la_output[55] soc/la_output[56]
+ soc/la_output[57] soc/la_output[58] soc/la_output[59] soc/la_output[5] soc/la_output[60]
+ soc/la_output[61] soc/la_output[62] soc/la_output[63] soc/la_output[64] soc/la_output[65]
+ soc/la_output[66] soc/la_output[67] soc/la_output[68] soc/la_output[69] soc/la_output[6]
+ soc/la_output[70] soc/la_output[71] soc/la_output[72] soc/la_output[73] soc/la_output[74]
+ soc/la_output[75] soc/la_output[76] soc/la_output[77] soc/la_output[78] soc/la_output[79]
+ soc/la_output[7] soc/la_output[80] soc/la_output[81] soc/la_output[82] soc/la_output[83]
+ soc/la_output[84] soc/la_output[85] soc/la_output[86] soc/la_output[87] soc/la_output[88]
+ soc/la_output[89] soc/la_output[8] soc/la_output[90] soc/la_output[91] soc/la_output[92]
+ soc/la_output[93] soc/la_output[94] soc/la_output[95] soc/la_output[96] soc/la_output[97]
+ soc/la_output[98] soc/la_output[99] soc/la_output[9] mprj/la_oen[0] mprj/la_oen[100]
+ mprj/la_oen[101] mprj/la_oen[102] mprj/la_oen[103] mprj/la_oen[104] mprj/la_oen[105]
+ mprj/la_oen[106] mprj/la_oen[107] mprj/la_oen[108] mprj/la_oen[109] mprj/la_oen[10]
+ mprj/la_oen[110] mprj/la_oen[111] mprj/la_oen[112] mprj/la_oen[113] mprj/la_oen[114]
+ mprj/la_oen[115] mprj/la_oen[116] mprj/la_oen[117] mprj/la_oen[118] mprj/la_oen[119]
+ mprj/la_oen[11] mprj/la_oen[120] mprj/la_oen[121] mprj/la_oen[122] mprj/la_oen[123]
+ mprj/la_oen[124] mprj/la_oen[125] mprj/la_oen[126] mprj/la_oen[127] mprj/la_oen[12]
+ mprj/la_oen[13] mprj/la_oen[14] mprj/la_oen[15] mprj/la_oen[16] mprj/la_oen[17]
+ mprj/la_oen[18] mprj/la_oen[19] mprj/la_oen[1] mprj/la_oen[20] mprj/la_oen[21] mprj/la_oen[22]
+ mprj/la_oen[23] mprj/la_oen[24] mprj/la_oen[25] mprj/la_oen[26] mprj/la_oen[27]
+ mprj/la_oen[28] mprj/la_oen[29] mprj/la_oen[2] mprj/la_oen[30] mprj/la_oen[31] mprj/la_oen[32]
+ mprj/la_oen[33] mprj/la_oen[34] mprj/la_oen[35] mprj/la_oen[36] mprj/la_oen[37]
+ mprj/la_oen[38] mprj/la_oen[39] mprj/la_oen[3] mprj/la_oen[40] mprj/la_oen[41] mprj/la_oen[42]
+ mprj/la_oen[43] mprj/la_oen[44] mprj/la_oen[45] mprj/la_oen[46] mprj/la_oen[47]
+ mprj/la_oen[48] mprj/la_oen[49] mprj/la_oen[4] mprj/la_oen[50] mprj/la_oen[51] mprj/la_oen[52]
+ mprj/la_oen[53] mprj/la_oen[54] mprj/la_oen[55] mprj/la_oen[56] mprj/la_oen[57]
+ mprj/la_oen[58] mprj/la_oen[59] mprj/la_oen[5] mprj/la_oen[60] mprj/la_oen[61] mprj/la_oen[62]
+ mprj/la_oen[63] mprj/la_oen[64] mprj/la_oen[65] mprj/la_oen[66] mprj/la_oen[67]
+ mprj/la_oen[68] mprj/la_oen[69] mprj/la_oen[6] mprj/la_oen[70] mprj/la_oen[71] mprj/la_oen[72]
+ mprj/la_oen[73] mprj/la_oen[74] mprj/la_oen[75] mprj/la_oen[76] mprj/la_oen[77]
+ mprj/la_oen[78] mprj/la_oen[79] mprj/la_oen[7] mprj/la_oen[80] mprj/la_oen[81] mprj/la_oen[82]
+ mprj/la_oen[83] mprj/la_oen[84] mprj/la_oen[85] mprj/la_oen[86] mprj/la_oen[87]
+ mprj/la_oen[88] mprj/la_oen[89] mprj/la_oen[8] mprj/la_oen[90] mprj/la_oen[91] mprj/la_oen[92]
+ mprj/la_oen[93] mprj/la_oen[94] mprj/la_oen[95] mprj/la_oen[96] mprj/la_oen[97]
+ mprj/la_oen[98] mprj/la_oen[99] mprj/la_oen[9] soc/la_oen[0] soc/la_oen[100] soc/la_oen[101]
+ soc/la_oen[102] soc/la_oen[103] soc/la_oen[104] soc/la_oen[105] soc/la_oen[106]
+ soc/la_oen[107] soc/la_oen[108] soc/la_oen[109] soc/la_oen[10] soc/la_oen[110] soc/la_oen[111]
+ soc/la_oen[112] soc/la_oen[113] soc/la_oen[114] soc/la_oen[115] soc/la_oen[116]
+ soc/la_oen[117] soc/la_oen[118] soc/la_oen[119] soc/la_oen[11] soc/la_oen[120] soc/la_oen[121]
+ soc/la_oen[122] soc/la_oen[123] soc/la_oen[124] soc/la_oen[125] soc/la_oen[126]
+ soc/la_oen[127] soc/la_oen[12] soc/la_oen[13] soc/la_oen[14] soc/la_oen[15] soc/la_oen[16]
+ soc/la_oen[17] soc/la_oen[18] soc/la_oen[19] soc/la_oen[1] soc/la_oen[20] soc/la_oen[21]
+ soc/la_oen[22] soc/la_oen[23] soc/la_oen[24] soc/la_oen[25] soc/la_oen[26] soc/la_oen[27]
+ soc/la_oen[28] soc/la_oen[29] soc/la_oen[2] soc/la_oen[30] soc/la_oen[31] soc/la_oen[32]
+ soc/la_oen[33] soc/la_oen[34] soc/la_oen[35] soc/la_oen[36] soc/la_oen[37] soc/la_oen[38]
+ soc/la_oen[39] soc/la_oen[3] soc/la_oen[40] soc/la_oen[41] soc/la_oen[42] soc/la_oen[43]
+ soc/la_oen[44] soc/la_oen[45] soc/la_oen[46] soc/la_oen[47] soc/la_oen[48] soc/la_oen[49]
+ soc/la_oen[4] soc/la_oen[50] soc/la_oen[51] soc/la_oen[52] soc/la_oen[53] soc/la_oen[54]
+ soc/la_oen[55] soc/la_oen[56] soc/la_oen[57] soc/la_oen[58] soc/la_oen[59] soc/la_oen[5]
+ soc/la_oen[60] soc/la_oen[61] soc/la_oen[62] soc/la_oen[63] soc/la_oen[64] soc/la_oen[65]
+ soc/la_oen[66] soc/la_oen[67] soc/la_oen[68] soc/la_oen[69] soc/la_oen[6] soc/la_oen[70]
+ soc/la_oen[71] soc/la_oen[72] soc/la_oen[73] soc/la_oen[74] soc/la_oen[75] soc/la_oen[76]
+ soc/la_oen[77] soc/la_oen[78] soc/la_oen[79] soc/la_oen[7] soc/la_oen[80] soc/la_oen[81]
+ soc/la_oen[82] soc/la_oen[83] soc/la_oen[84] soc/la_oen[85] soc/la_oen[86] soc/la_oen[87]
+ soc/la_oen[88] soc/la_oen[89] soc/la_oen[8] soc/la_oen[90] soc/la_oen[91] soc/la_oen[92]
+ soc/la_oen[93] soc/la_oen[94] soc/la_oen[95] soc/la_oen[96] soc/la_oen[97] soc/la_oen[98]
+ soc/la_oen[99] soc/la_oen[9] soc/mprj_adr_o[0] soc/mprj_adr_o[10] soc/mprj_adr_o[11]
+ soc/mprj_adr_o[12] soc/mprj_adr_o[13] soc/mprj_adr_o[14] soc/mprj_adr_o[15] soc/mprj_adr_o[16]
+ soc/mprj_adr_o[17] soc/mprj_adr_o[18] soc/mprj_adr_o[19] soc/mprj_adr_o[1] soc/mprj_adr_o[20]
+ soc/mprj_adr_o[21] soc/mprj_adr_o[22] soc/mprj_adr_o[23] soc/mprj_adr_o[24] soc/mprj_adr_o[25]
+ soc/mprj_adr_o[26] soc/mprj_adr_o[27] soc/mprj_adr_o[28] soc/mprj_adr_o[29] soc/mprj_adr_o[2]
+ soc/mprj_adr_o[30] soc/mprj_adr_o[31] soc/mprj_adr_o[3] soc/mprj_adr_o[4] soc/mprj_adr_o[5]
+ soc/mprj_adr_o[6] soc/mprj_adr_o[7] soc/mprj_adr_o[8] soc/mprj_adr_o[9] mprj/wbs_adr_i[0]
+ mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12] mprj/wbs_adr_i[13] mprj/wbs_adr_i[14]
+ mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17] mprj/wbs_adr_i[18] mprj/wbs_adr_i[19]
+ mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21] mprj/wbs_adr_i[22] mprj/wbs_adr_i[23]
+ mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26] mprj/wbs_adr_i[27] mprj/wbs_adr_i[28]
+ mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30] mprj/wbs_adr_i[31] mprj/wbs_adr_i[3]
+ mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6] mprj/wbs_adr_i[7] mprj/wbs_adr_i[8]
+ mprj/wbs_adr_i[9] soc/mprj_cyc_o mprj/wbs_cyc_i soc/mprj_dat_o[0] soc/mprj_dat_o[10]
+ soc/mprj_dat_o[11] soc/mprj_dat_o[12] soc/mprj_dat_o[13] soc/mprj_dat_o[14] soc/mprj_dat_o[15]
+ soc/mprj_dat_o[16] soc/mprj_dat_o[17] soc/mprj_dat_o[18] soc/mprj_dat_o[19] soc/mprj_dat_o[1]
+ soc/mprj_dat_o[20] soc/mprj_dat_o[21] soc/mprj_dat_o[22] soc/mprj_dat_o[23] soc/mprj_dat_o[24]
+ soc/mprj_dat_o[25] soc/mprj_dat_o[26] soc/mprj_dat_o[27] soc/mprj_dat_o[28] soc/mprj_dat_o[29]
+ soc/mprj_dat_o[2] soc/mprj_dat_o[30] soc/mprj_dat_o[31] soc/mprj_dat_o[3] soc/mprj_dat_o[4]
+ soc/mprj_dat_o[5] soc/mprj_dat_o[6] soc/mprj_dat_o[7] soc/mprj_dat_o[8] soc/mprj_dat_o[9]
+ mprj/wbs_dat_i[0] mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13]
+ mprj/wbs_dat_i[14] mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18]
+ mprj/wbs_dat_i[19] mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22]
+ mprj/wbs_dat_i[23] mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27]
+ mprj/wbs_dat_i[28] mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31]
+ mprj/wbs_dat_i[3] mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7]
+ mprj/wbs_dat_i[8] mprj/wbs_dat_i[9] soc/mprj_sel_o[0] soc/mprj_sel_o[1] soc/mprj_sel_o[2]
+ soc/mprj_sel_o[3] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1] mprj/wbs_sel_i[2] mprj/wbs_sel_i[3]
+ soc/mprj_stb_o mprj/wbs_stb_i soc/mprj_we_o mprj/wbs_we_i soc/mprj_vcc_pwrgood soc/mprj_vdd_pwrgood
+ soc/mprj2_vcc_pwrgood soc/mprj2_vdd_pwrgood mprj/wb_clk_i mprj/user_clock2 mprj/wb_rst_i
+ mgmt_buffers/user_resetn vccd vssd vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
+ mgmt_protect
Xrstb_level rstb_level/A soc/resetb vddio vssio vccd rstb_level/LVGND VSUBS sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped
Xgpio_control_in\[27\] soc/mgmt_in_data[27] gpio_control_in\[27\]/one soc/mgmt_in_data[27]
+ gpio_control_in\[27\]/one padframe/mprj_io_analog_en[27] padframe/mprj_io_analog_pol[27]
+ padframe/mprj_io_analog_sel[27] padframe/mprj_io_dm[81] padframe/mprj_io_dm[82]
+ padframe/mprj_io_dm[83] padframe/mprj_io_holdover[27] padframe/mprj_io_ib_mode_sel[27]
+ padframe/mprj_io_in[27] padframe/mprj_io_inp_dis[27] padframe/mprj_io_out[27] padframe/mprj_io_oeb[27]
+ padframe/mprj_io_slow_sel[27] padframe/mprj_io_vtrip_sel[27] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[27\]/serial_data_in gpio_control_in\[28\]/serial_data_in
+ mprj/io_in[27] mprj/io_oeb[27] mprj/io_out[27] gpio_control_in\[27\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[2\] soc/mgmt_in_data[2] gpio_control_in\[2\]/one soc/mgmt_in_data[2]
+ gpio_control_in\[2\]/one padframe/mprj_io_analog_en[2] padframe/mprj_io_analog_pol[2]
+ padframe/mprj_io_analog_sel[2] padframe/mprj_io_dm[6] padframe/mprj_io_dm[7] padframe/mprj_io_dm[8]
+ padframe/mprj_io_holdover[2] padframe/mprj_io_ib_mode_sel[2] padframe/mprj_io_in[2]
+ padframe/mprj_io_inp_dis[2] padframe/mprj_io_out[2] padframe/mprj_io_oeb[2] padframe/mprj_io_slow_sel[2]
+ padframe/mprj_io_vtrip_sel[2] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[2\]/serial_data_in gpio_control_in\[3\]/serial_data_in mprj/io_in[2]
+ mprj/io_oeb[2] mprj/io_out[2] gpio_control_in\[2\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[32\] soc/mgmt_in_data[32] gpio_control_in\[32\]/one soc/mgmt_in_data[32]
+ gpio_control_in\[32\]/one padframe/mprj_io_analog_en[32] padframe/mprj_io_analog_pol[32]
+ padframe/mprj_io_analog_sel[32] padframe/mprj_io_dm[96] padframe/mprj_io_dm[97]
+ padframe/mprj_io_dm[98] padframe/mprj_io_holdover[32] padframe/mprj_io_ib_mode_sel[32]
+ padframe/mprj_io_in[32] padframe/mprj_io_inp_dis[32] padframe/mprj_io_out[32] padframe/mprj_io_oeb[32]
+ padframe/mprj_io_slow_sel[32] padframe/mprj_io_vtrip_sel[32] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[32\]/serial_data_in gpio_control_in\[33\]/serial_data_in
+ mprj/io_in[32] mprj/io_oeb[32] mprj/io_out[32] gpio_control_in\[32\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[25\] soc/mgmt_in_data[25] gpio_control_in\[25\]/one soc/mgmt_in_data[25]
+ gpio_control_in\[25\]/one padframe/mprj_io_analog_en[25] padframe/mprj_io_analog_pol[25]
+ padframe/mprj_io_analog_sel[25] padframe/mprj_io_dm[75] padframe/mprj_io_dm[76]
+ padframe/mprj_io_dm[77] padframe/mprj_io_holdover[25] padframe/mprj_io_ib_mode_sel[25]
+ padframe/mprj_io_in[25] padframe/mprj_io_inp_dis[25] padframe/mprj_io_out[25] padframe/mprj_io_oeb[25]
+ padframe/mprj_io_slow_sel[25] padframe/mprj_io_vtrip_sel[25] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[25\]/serial_data_in gpio_control_in\[26\]/serial_data_in
+ mprj/io_in[25] mprj/io_oeb[25] mprj/io_out[25] gpio_control_in\[25\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[18\] soc/mgmt_in_data[18] gpio_control_in\[18\]/one soc/mgmt_in_data[18]
+ gpio_control_in\[18\]/one padframe/mprj_io_analog_en[18] padframe/mprj_io_analog_pol[18]
+ padframe/mprj_io_analog_sel[18] padframe/mprj_io_dm[54] padframe/mprj_io_dm[55]
+ padframe/mprj_io_dm[56] padframe/mprj_io_holdover[18] padframe/mprj_io_ib_mode_sel[18]
+ padframe/mprj_io_in[18] padframe/mprj_io_inp_dis[18] padframe/mprj_io_out[18] padframe/mprj_io_oeb[18]
+ padframe/mprj_io_slow_sel[18] padframe/mprj_io_vtrip_sel[18] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[18\]/serial_data_in gpio_control_in\[19\]/serial_data_in
+ mprj/io_in[18] mprj/io_oeb[18] mprj/io_out[18] gpio_control_in\[18\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[30\] soc/mgmt_in_data[30] gpio_control_in\[30\]/one soc/mgmt_in_data[30]
+ gpio_control_in\[30\]/one padframe/mprj_io_analog_en[30] padframe/mprj_io_analog_pol[30]
+ padframe/mprj_io_analog_sel[30] padframe/mprj_io_dm[90] padframe/mprj_io_dm[91]
+ padframe/mprj_io_dm[92] padframe/mprj_io_holdover[30] padframe/mprj_io_ib_mode_sel[30]
+ padframe/mprj_io_in[30] padframe/mprj_io_inp_dis[30] padframe/mprj_io_out[30] padframe/mprj_io_oeb[30]
+ padframe/mprj_io_slow_sel[30] padframe/mprj_io_vtrip_sel[30] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[30\]/serial_data_in gpio_control_in\[31\]/serial_data_in
+ mprj/io_in[30] mprj/io_oeb[30] mprj/io_out[30] gpio_control_in\[30\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[23\] soc/mgmt_in_data[23] gpio_control_in\[23\]/one soc/mgmt_in_data[23]
+ gpio_control_in\[23\]/one padframe/mprj_io_analog_en[23] padframe/mprj_io_analog_pol[23]
+ padframe/mprj_io_analog_sel[23] padframe/mprj_io_dm[69] padframe/mprj_io_dm[70]
+ padframe/mprj_io_dm[71] padframe/mprj_io_holdover[23] padframe/mprj_io_ib_mode_sel[23]
+ padframe/mprj_io_in[23] padframe/mprj_io_inp_dis[23] padframe/mprj_io_out[23] padframe/mprj_io_oeb[23]
+ padframe/mprj_io_slow_sel[23] padframe/mprj_io_vtrip_sel[23] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[23\]/serial_data_in gpio_control_in\[24\]/serial_data_in
+ mprj/io_in[23] mprj/io_oeb[23] mprj/io_out[23] gpio_control_in\[23\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[9\] soc/mgmt_in_data[9] gpio_control_in\[9\]/one soc/mgmt_in_data[9]
+ gpio_control_in\[9\]/one padframe/mprj_io_analog_en[9] padframe/mprj_io_analog_pol[9]
+ padframe/mprj_io_analog_sel[9] padframe/mprj_io_dm[27] padframe/mprj_io_dm[28] padframe/mprj_io_dm[29]
+ padframe/mprj_io_holdover[9] padframe/mprj_io_ib_mode_sel[9] padframe/mprj_io_in[9]
+ padframe/mprj_io_inp_dis[9] padframe/mprj_io_out[9] padframe/mprj_io_oeb[9] padframe/mprj_io_slow_sel[9]
+ padframe/mprj_io_vtrip_sel[9] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[9\]/serial_data_in gpio_control_in\[9\]/serial_data_out mprj/io_in[9]
+ mprj/io_oeb[9] mprj/io_out[9] gpio_control_in\[9\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_bidir\[0\] soc/mgmt_in_data[0] soc/jtag_outenb soc/jtag_out gpio_control_bidir\[0\]/one
+ padframe/mprj_io_analog_en[0] padframe/mprj_io_analog_pol[0] padframe/mprj_io_analog_sel[0]
+ padframe/mprj_io_dm[0] padframe/mprj_io_dm[1] padframe/mprj_io_dm[2] padframe/mprj_io_holdover[0]
+ padframe/mprj_io_ib_mode_sel[0] padframe/mprj_io_in[0] padframe/mprj_io_inp_dis[0]
+ padframe/mprj_io_out[0] padframe/mprj_io_oeb[0] padframe/mprj_io_slow_sel[0] padframe/mprj_io_vtrip_sel[0]
+ soc/mprj_io_loader_resetn soc/mprj_io_loader_clock soc/mprj_io_loader_data gpio_control_bidir\[1\]/serial_data_in
+ mprj/io_in[0] mprj/io_oeb[0] mprj/io_out[0] gpio_control_bidir\[0\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[16\] soc/mgmt_in_data[16] gpio_control_in\[16\]/one soc/mgmt_in_data[16]
+ gpio_control_in\[16\]/one padframe/mprj_io_analog_en[16] padframe/mprj_io_analog_pol[16]
+ padframe/mprj_io_analog_sel[16] padframe/mprj_io_dm[48] padframe/mprj_io_dm[49]
+ padframe/mprj_io_dm[50] padframe/mprj_io_holdover[16] padframe/mprj_io_ib_mode_sel[16]
+ padframe/mprj_io_in[16] padframe/mprj_io_inp_dis[16] padframe/mprj_io_out[16] padframe/mprj_io_oeb[16]
+ padframe/mprj_io_slow_sel[16] padframe/mprj_io_vtrip_sel[16] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[16\]/serial_data_in gpio_control_in\[17\]/serial_data_in
+ mprj/io_in[16] mprj/io_oeb[16] mprj/io_out[16] gpio_control_in\[16\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[21\] soc/mgmt_in_data[21] gpio_control_in\[21\]/one soc/mgmt_in_data[21]
+ gpio_control_in\[21\]/one padframe/mprj_io_analog_en[21] padframe/mprj_io_analog_pol[21]
+ padframe/mprj_io_analog_sel[21] padframe/mprj_io_dm[63] padframe/mprj_io_dm[64]
+ padframe/mprj_io_dm[65] padframe/mprj_io_holdover[21] padframe/mprj_io_ib_mode_sel[21]
+ padframe/mprj_io_in[21] padframe/mprj_io_inp_dis[21] padframe/mprj_io_out[21] padframe/mprj_io_oeb[21]
+ padframe/mprj_io_slow_sel[21] padframe/mprj_io_vtrip_sel[21] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[21\]/serial_data_in gpio_control_in\[22\]/serial_data_in
+ mprj/io_in[21] mprj/io_oeb[21] mprj/io_out[21] gpio_control_in\[21\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xmprj mprj/analog_io[0] mprj/analog_io[10] mprj/analog_io[11] mprj/analog_io[12] mprj/analog_io[13]
+ mprj/analog_io[14] mprj/analog_io[15] mprj/analog_io[16] mprj/analog_io[17] mprj/analog_io[18]
+ mprj/analog_io[19] mprj/analog_io[1] mprj/analog_io[20] mprj/analog_io[21] mprj/analog_io[22]
+ mprj/analog_io[23] mprj/analog_io[24] mprj/analog_io[25] mprj/analog_io[26] mprj/analog_io[27]
+ mprj/analog_io[28] mprj/analog_io[29] mprj/analog_io[2] mprj/analog_io[30] mprj/analog_io[3]
+ mprj/analog_io[4] mprj/analog_io[5] mprj/analog_io[6] mprj/analog_io[7] mprj/analog_io[8]
+ mprj/analog_io[9] mprj/io_in[0] mprj/io_in[10] mprj/io_in[11] mprj/io_in[12] mprj/io_in[13]
+ mprj/io_in[14] mprj/io_in[15] mprj/io_in[16] mprj/io_in[17] mprj/io_in[18] mprj/io_in[19]
+ mprj/io_in[1] mprj/io_in[20] mprj/io_in[21] mprj/io_in[22] mprj/io_in[23] mprj/io_in[24]
+ mprj/io_in[25] mprj/io_in[26] mprj/io_in[27] mprj/io_in[28] mprj/io_in[29] mprj/io_in[2]
+ mprj/io_in[30] mprj/io_in[31] mprj/io_in[32] mprj/io_in[33] mprj/io_in[34] mprj/io_in[35]
+ mprj/io_in[36] mprj/io_in[37] mprj/io_in[3] mprj/io_in[4] mprj/io_in[5] mprj/io_in[6]
+ mprj/io_in[7] mprj/io_in[8] mprj/io_in[9] mprj/io_oeb[0] mprj/io_oeb[10] mprj/io_oeb[11]
+ mprj/io_oeb[12] mprj/io_oeb[13] mprj/io_oeb[14] mprj/io_oeb[15] mprj/io_oeb[16]
+ mprj/io_oeb[17] mprj/io_oeb[18] mprj/io_oeb[19] mprj/io_oeb[1] mprj/io_oeb[20] mprj/io_oeb[21]
+ mprj/io_oeb[22] mprj/io_oeb[23] mprj/io_oeb[24] mprj/io_oeb[25] mprj/io_oeb[26]
+ mprj/io_oeb[27] mprj/io_oeb[28] mprj/io_oeb[29] mprj/io_oeb[2] mprj/io_oeb[30] mprj/io_oeb[31]
+ mprj/io_oeb[32] mprj/io_oeb[33] mprj/io_oeb[34] mprj/io_oeb[35] mprj/io_oeb[36]
+ mprj/io_oeb[37] mprj/io_oeb[3] mprj/io_oeb[4] mprj/io_oeb[5] mprj/io_oeb[6] mprj/io_oeb[7]
+ mprj/io_oeb[8] mprj/io_oeb[9] mprj/io_out[0] mprj/io_out[10] mprj/io_out[11] mprj/io_out[12]
+ mprj/io_out[13] mprj/io_out[14] mprj/io_out[15] mprj/io_out[16] mprj/io_out[17]
+ mprj/io_out[18] mprj/io_out[19] mprj/io_out[1] mprj/io_out[20] mprj/io_out[21] mprj/io_out[22]
+ mprj/io_out[23] mprj/io_out[24] mprj/io_out[25] mprj/io_out[26] mprj/io_out[27]
+ mprj/io_out[28] mprj/io_out[29] mprj/io_out[2] mprj/io_out[30] mprj/io_out[31] mprj/io_out[32]
+ mprj/io_out[33] mprj/io_out[34] mprj/io_out[35] mprj/io_out[36] mprj/io_out[37]
+ mprj/io_out[3] mprj/io_out[4] mprj/io_out[5] mprj/io_out[6] mprj/io_out[7] mprj/io_out[8]
+ mprj/io_out[9] mprj/la_data_in[0] mprj/la_data_in[100] mprj/la_data_in[101] mprj/la_data_in[102]
+ mprj/la_data_in[103] mprj/la_data_in[104] mprj/la_data_in[105] mprj/la_data_in[106]
+ mprj/la_data_in[107] mprj/la_data_in[108] mprj/la_data_in[109] mprj/la_data_in[10]
+ mprj/la_data_in[110] mprj/la_data_in[111] mprj/la_data_in[112] mprj/la_data_in[113]
+ mprj/la_data_in[114] mprj/la_data_in[115] mprj/la_data_in[116] mprj/la_data_in[117]
+ mprj/la_data_in[118] mprj/la_data_in[119] mprj/la_data_in[11] mprj/la_data_in[120]
+ mprj/la_data_in[121] mprj/la_data_in[122] mprj/la_data_in[123] mprj/la_data_in[124]
+ mprj/la_data_in[125] mprj/la_data_in[126] mprj/la_data_in[127] mprj/la_data_in[12]
+ mprj/la_data_in[13] mprj/la_data_in[14] mprj/la_data_in[15] mprj/la_data_in[16]
+ mprj/la_data_in[17] mprj/la_data_in[18] mprj/la_data_in[19] mprj/la_data_in[1] mprj/la_data_in[20]
+ mprj/la_data_in[21] mprj/la_data_in[22] mprj/la_data_in[23] mprj/la_data_in[24]
+ mprj/la_data_in[25] mprj/la_data_in[26] mprj/la_data_in[27] mprj/la_data_in[28]
+ mprj/la_data_in[29] mprj/la_data_in[2] mprj/la_data_in[30] mprj/la_data_in[31] mprj/la_data_in[32]
+ mprj/la_data_in[33] mprj/la_data_in[34] mprj/la_data_in[35] mprj/la_data_in[36]
+ mprj/la_data_in[37] mprj/la_data_in[38] mprj/la_data_in[39] mprj/la_data_in[3] mprj/la_data_in[40]
+ mprj/la_data_in[41] mprj/la_data_in[42] mprj/la_data_in[43] mprj/la_data_in[44]
+ mprj/la_data_in[45] mprj/la_data_in[46] mprj/la_data_in[47] mprj/la_data_in[48]
+ mprj/la_data_in[49] mprj/la_data_in[4] mprj/la_data_in[50] mprj/la_data_in[51] mprj/la_data_in[52]
+ mprj/la_data_in[53] mprj/la_data_in[54] mprj/la_data_in[55] mprj/la_data_in[56]
+ mprj/la_data_in[57] mprj/la_data_in[58] mprj/la_data_in[59] mprj/la_data_in[5] mprj/la_data_in[60]
+ mprj/la_data_in[61] mprj/la_data_in[62] mprj/la_data_in[63] mprj/la_data_in[64]
+ mprj/la_data_in[65] mprj/la_data_in[66] mprj/la_data_in[67] mprj/la_data_in[68]
+ mprj/la_data_in[69] mprj/la_data_in[6] mprj/la_data_in[70] mprj/la_data_in[71] mprj/la_data_in[72]
+ mprj/la_data_in[73] mprj/la_data_in[74] mprj/la_data_in[75] mprj/la_data_in[76]
+ mprj/la_data_in[77] mprj/la_data_in[78] mprj/la_data_in[79] mprj/la_data_in[7] mprj/la_data_in[80]
+ mprj/la_data_in[81] mprj/la_data_in[82] mprj/la_data_in[83] mprj/la_data_in[84]
+ mprj/la_data_in[85] mprj/la_data_in[86] mprj/la_data_in[87] mprj/la_data_in[88]
+ mprj/la_data_in[89] mprj/la_data_in[8] mprj/la_data_in[90] mprj/la_data_in[91] mprj/la_data_in[92]
+ mprj/la_data_in[93] mprj/la_data_in[94] mprj/la_data_in[95] mprj/la_data_in[96]
+ mprj/la_data_in[97] mprj/la_data_in[98] mprj/la_data_in[99] mprj/la_data_in[9] mprj/la_data_out[0]
+ mprj/la_data_out[100] mprj/la_data_out[101] mprj/la_data_out[102] mprj/la_data_out[103]
+ mprj/la_data_out[104] mprj/la_data_out[105] mprj/la_data_out[106] mprj/la_data_out[107]
+ mprj/la_data_out[108] mprj/la_data_out[109] mprj/la_data_out[10] mprj/la_data_out[110]
+ mprj/la_data_out[111] mprj/la_data_out[112] mprj/la_data_out[113] mprj/la_data_out[114]
+ mprj/la_data_out[115] mprj/la_data_out[116] mprj/la_data_out[117] mprj/la_data_out[118]
+ mprj/la_data_out[119] mprj/la_data_out[11] mprj/la_data_out[120] mprj/la_data_out[121]
+ mprj/la_data_out[122] mprj/la_data_out[123] mprj/la_data_out[124] mprj/la_data_out[125]
+ mprj/la_data_out[126] mprj/la_data_out[127] mprj/la_data_out[12] mprj/la_data_out[13]
+ mprj/la_data_out[14] mprj/la_data_out[15] mprj/la_data_out[16] mprj/la_data_out[17]
+ mprj/la_data_out[18] mprj/la_data_out[19] mprj/la_data_out[1] mprj/la_data_out[20]
+ mprj/la_data_out[21] mprj/la_data_out[22] mprj/la_data_out[23] mprj/la_data_out[24]
+ mprj/la_data_out[25] mprj/la_data_out[26] mprj/la_data_out[27] mprj/la_data_out[28]
+ mprj/la_data_out[29] mprj/la_data_out[2] mprj/la_data_out[30] mprj/la_data_out[31]
+ mprj/la_data_out[32] mprj/la_data_out[33] mprj/la_data_out[34] mprj/la_data_out[35]
+ mprj/la_data_out[36] mprj/la_data_out[37] mprj/la_data_out[38] mprj/la_data_out[39]
+ mprj/la_data_out[3] mprj/la_data_out[40] mprj/la_data_out[41] mprj/la_data_out[42]
+ mprj/la_data_out[43] mprj/la_data_out[44] mprj/la_data_out[45] mprj/la_data_out[46]
+ mprj/la_data_out[47] mprj/la_data_out[48] mprj/la_data_out[49] mprj/la_data_out[4]
+ mprj/la_data_out[50] mprj/la_data_out[51] mprj/la_data_out[52] mprj/la_data_out[53]
+ mprj/la_data_out[54] mprj/la_data_out[55] mprj/la_data_out[56] mprj/la_data_out[57]
+ mprj/la_data_out[58] mprj/la_data_out[59] mprj/la_data_out[5] mprj/la_data_out[60]
+ mprj/la_data_out[61] mprj/la_data_out[62] mprj/la_data_out[63] mprj/la_data_out[64]
+ mprj/la_data_out[65] mprj/la_data_out[66] mprj/la_data_out[67] mprj/la_data_out[68]
+ mprj/la_data_out[69] mprj/la_data_out[6] mprj/la_data_out[70] mprj/la_data_out[71]
+ mprj/la_data_out[72] mprj/la_data_out[73] mprj/la_data_out[74] mprj/la_data_out[75]
+ mprj/la_data_out[76] mprj/la_data_out[77] mprj/la_data_out[78] mprj/la_data_out[79]
+ mprj/la_data_out[7] mprj/la_data_out[80] mprj/la_data_out[81] mprj/la_data_out[82]
+ mprj/la_data_out[83] mprj/la_data_out[84] mprj/la_data_out[85] mprj/la_data_out[86]
+ mprj/la_data_out[87] mprj/la_data_out[88] mprj/la_data_out[89] mprj/la_data_out[8]
+ mprj/la_data_out[90] mprj/la_data_out[91] mprj/la_data_out[92] mprj/la_data_out[93]
+ mprj/la_data_out[94] mprj/la_data_out[95] mprj/la_data_out[96] mprj/la_data_out[97]
+ mprj/la_data_out[98] mprj/la_data_out[99] mprj/la_data_out[9] mprj/la_oen[0] mprj/la_oen[100]
+ mprj/la_oen[101] mprj/la_oen[102] mprj/la_oen[103] mprj/la_oen[104] mprj/la_oen[105]
+ mprj/la_oen[106] mprj/la_oen[107] mprj/la_oen[108] mprj/la_oen[109] mprj/la_oen[10]
+ mprj/la_oen[110] mprj/la_oen[111] mprj/la_oen[112] mprj/la_oen[113] mprj/la_oen[114]
+ mprj/la_oen[115] mprj/la_oen[116] mprj/la_oen[117] mprj/la_oen[118] mprj/la_oen[119]
+ mprj/la_oen[11] mprj/la_oen[120] mprj/la_oen[121] mprj/la_oen[122] mprj/la_oen[123]
+ mprj/la_oen[124] mprj/la_oen[125] mprj/la_oen[126] mprj/la_oen[127] mprj/la_oen[12]
+ mprj/la_oen[13] mprj/la_oen[14] mprj/la_oen[15] mprj/la_oen[16] mprj/la_oen[17]
+ mprj/la_oen[18] mprj/la_oen[19] mprj/la_oen[1] mprj/la_oen[20] mprj/la_oen[21] mprj/la_oen[22]
+ mprj/la_oen[23] mprj/la_oen[24] mprj/la_oen[25] mprj/la_oen[26] mprj/la_oen[27]
+ mprj/la_oen[28] mprj/la_oen[29] mprj/la_oen[2] mprj/la_oen[30] mprj/la_oen[31] mprj/la_oen[32]
+ mprj/la_oen[33] mprj/la_oen[34] mprj/la_oen[35] mprj/la_oen[36] mprj/la_oen[37]
+ mprj/la_oen[38] mprj/la_oen[39] mprj/la_oen[3] mprj/la_oen[40] mprj/la_oen[41] mprj/la_oen[42]
+ mprj/la_oen[43] mprj/la_oen[44] mprj/la_oen[45] mprj/la_oen[46] mprj/la_oen[47]
+ mprj/la_oen[48] mprj/la_oen[49] mprj/la_oen[4] mprj/la_oen[50] mprj/la_oen[51] mprj/la_oen[52]
+ mprj/la_oen[53] mprj/la_oen[54] mprj/la_oen[55] mprj/la_oen[56] mprj/la_oen[57]
+ mprj/la_oen[58] mprj/la_oen[59] mprj/la_oen[5] mprj/la_oen[60] mprj/la_oen[61] mprj/la_oen[62]
+ mprj/la_oen[63] mprj/la_oen[64] mprj/la_oen[65] mprj/la_oen[66] mprj/la_oen[67]
+ mprj/la_oen[68] mprj/la_oen[69] mprj/la_oen[6] mprj/la_oen[70] mprj/la_oen[71] mprj/la_oen[72]
+ mprj/la_oen[73] mprj/la_oen[74] mprj/la_oen[75] mprj/la_oen[76] mprj/la_oen[77]
+ mprj/la_oen[78] mprj/la_oen[79] mprj/la_oen[7] mprj/la_oen[80] mprj/la_oen[81] mprj/la_oen[82]
+ mprj/la_oen[83] mprj/la_oen[84] mprj/la_oen[85] mprj/la_oen[86] mprj/la_oen[87]
+ mprj/la_oen[88] mprj/la_oen[89] mprj/la_oen[8] mprj/la_oen[90] mprj/la_oen[91] mprj/la_oen[92]
+ mprj/la_oen[93] mprj/la_oen[94] mprj/la_oen[95] mprj/la_oen[96] mprj/la_oen[97]
+ mprj/la_oen[98] mprj/la_oen[99] mprj/la_oen[9] mprj/user_clock2 mprj/wb_clk_i mprj/wb_rst_i
+ soc/mprj_ack_i mprj/wbs_adr_i[0] mprj/wbs_adr_i[10] mprj/wbs_adr_i[11] mprj/wbs_adr_i[12]
+ mprj/wbs_adr_i[13] mprj/wbs_adr_i[14] mprj/wbs_adr_i[15] mprj/wbs_adr_i[16] mprj/wbs_adr_i[17]
+ mprj/wbs_adr_i[18] mprj/wbs_adr_i[19] mprj/wbs_adr_i[1] mprj/wbs_adr_i[20] mprj/wbs_adr_i[21]
+ mprj/wbs_adr_i[22] mprj/wbs_adr_i[23] mprj/wbs_adr_i[24] mprj/wbs_adr_i[25] mprj/wbs_adr_i[26]
+ mprj/wbs_adr_i[27] mprj/wbs_adr_i[28] mprj/wbs_adr_i[29] mprj/wbs_adr_i[2] mprj/wbs_adr_i[30]
+ mprj/wbs_adr_i[31] mprj/wbs_adr_i[3] mprj/wbs_adr_i[4] mprj/wbs_adr_i[5] mprj/wbs_adr_i[6]
+ mprj/wbs_adr_i[7] mprj/wbs_adr_i[8] mprj/wbs_adr_i[9] mprj/wbs_cyc_i mprj/wbs_dat_i[0]
+ mprj/wbs_dat_i[10] mprj/wbs_dat_i[11] mprj/wbs_dat_i[12] mprj/wbs_dat_i[13] mprj/wbs_dat_i[14]
+ mprj/wbs_dat_i[15] mprj/wbs_dat_i[16] mprj/wbs_dat_i[17] mprj/wbs_dat_i[18] mprj/wbs_dat_i[19]
+ mprj/wbs_dat_i[1] mprj/wbs_dat_i[20] mprj/wbs_dat_i[21] mprj/wbs_dat_i[22] mprj/wbs_dat_i[23]
+ mprj/wbs_dat_i[24] mprj/wbs_dat_i[25] mprj/wbs_dat_i[26] mprj/wbs_dat_i[27] mprj/wbs_dat_i[28]
+ mprj/wbs_dat_i[29] mprj/wbs_dat_i[2] mprj/wbs_dat_i[30] mprj/wbs_dat_i[31] mprj/wbs_dat_i[3]
+ mprj/wbs_dat_i[4] mprj/wbs_dat_i[5] mprj/wbs_dat_i[6] mprj/wbs_dat_i[7] mprj/wbs_dat_i[8]
+ mprj/wbs_dat_i[9] soc/mprj_dat_i[0] soc/mprj_dat_i[10] soc/mprj_dat_i[11] soc/mprj_dat_i[12]
+ soc/mprj_dat_i[13] soc/mprj_dat_i[14] soc/mprj_dat_i[15] soc/mprj_dat_i[16] soc/mprj_dat_i[17]
+ soc/mprj_dat_i[18] soc/mprj_dat_i[19] soc/mprj_dat_i[1] soc/mprj_dat_i[20] soc/mprj_dat_i[21]
+ soc/mprj_dat_i[22] soc/mprj_dat_i[23] soc/mprj_dat_i[24] soc/mprj_dat_i[25] soc/mprj_dat_i[26]
+ soc/mprj_dat_i[27] soc/mprj_dat_i[28] soc/mprj_dat_i[29] soc/mprj_dat_i[2] soc/mprj_dat_i[30]
+ soc/mprj_dat_i[31] soc/mprj_dat_i[3] soc/mprj_dat_i[4] soc/mprj_dat_i[5] soc/mprj_dat_i[6]
+ soc/mprj_dat_i[7] soc/mprj_dat_i[8] soc/mprj_dat_i[9] mprj/wbs_sel_i[0] mprj/wbs_sel_i[1]
+ mprj/wbs_sel_i[2] mprj/wbs_sel_i[3] mprj/wbs_stb_i mprj/wbs_we_i vccd1 vssd1 vccd2
+ vssd2 vdda1 vssa1 vdda2 vssa2 user_project_wrapper
Xgpio_control_in\[14\] soc/mgmt_in_data[14] gpio_control_in\[14\]/one soc/mgmt_in_data[14]
+ gpio_control_in\[14\]/one padframe/mprj_io_analog_en[14] padframe/mprj_io_analog_pol[14]
+ padframe/mprj_io_analog_sel[14] padframe/mprj_io_dm[42] padframe/mprj_io_dm[43]
+ padframe/mprj_io_dm[44] padframe/mprj_io_holdover[14] padframe/mprj_io_ib_mode_sel[14]
+ padframe/mprj_io_in[14] padframe/mprj_io_inp_dis[14] padframe/mprj_io_out[14] padframe/mprj_io_oeb[14]
+ padframe/mprj_io_slow_sel[14] padframe/mprj_io_vtrip_sel[14] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[14\]/serial_data_in gpio_control_in\[15\]/serial_data_in
+ mprj/io_in[14] mprj/io_oeb[14] mprj/io_out[14] gpio_control_in\[14\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[7\] soc/mgmt_in_data[7] gpio_control_in\[7\]/one soc/mgmt_in_data[7]
+ gpio_control_in\[7\]/one padframe/mprj_io_analog_en[7] padframe/mprj_io_analog_pol[7]
+ padframe/mprj_io_analog_sel[7] padframe/mprj_io_dm[21] padframe/mprj_io_dm[22] padframe/mprj_io_dm[23]
+ padframe/mprj_io_holdover[7] padframe/mprj_io_ib_mode_sel[7] padframe/mprj_io_in[7]
+ padframe/mprj_io_inp_dis[7] padframe/mprj_io_out[7] padframe/mprj_io_oeb[7] padframe/mprj_io_slow_sel[7]
+ padframe/mprj_io_vtrip_sel[7] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[7\]/serial_data_in gpio_control_in\[8\]/serial_data_in mprj/io_in[7]
+ mprj/io_oeb[7] mprj/io_out[7] gpio_control_in\[7\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[5\] soc/mgmt_in_data[5] gpio_control_in\[5\]/one soc/mgmt_in_data[5]
+ gpio_control_in\[5\]/one padframe/mprj_io_analog_en[5] padframe/mprj_io_analog_pol[5]
+ padframe/mprj_io_analog_sel[5] padframe/mprj_io_dm[15] padframe/mprj_io_dm[16] padframe/mprj_io_dm[17]
+ padframe/mprj_io_holdover[5] padframe/mprj_io_ib_mode_sel[5] padframe/mprj_io_in[5]
+ padframe/mprj_io_inp_dis[5] padframe/mprj_io_out[5] padframe/mprj_io_oeb[5] padframe/mprj_io_slow_sel[5]
+ padframe/mprj_io_vtrip_sel[5] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[5\]/serial_data_in gpio_control_in\[6\]/serial_data_in mprj/io_in[5]
+ mprj/io_oeb[5] mprj/io_out[5] gpio_control_in\[5\]/zero vccd vssd vccd1 vssd1 gpio_control_block
Xgpio_control_in\[37\] soc/mgmt_in_data[37] gpio_control_in\[37\]/one soc/mgmt_in_data[37]
+ gpio_control_in\[37\]/one padframe/mprj_io_analog_en[37] padframe/mprj_io_analog_pol[37]
+ padframe/mprj_io_analog_sel[37] padframe/mprj_io_dm[111] padframe/mprj_io_dm[112]
+ padframe/mprj_io_dm[113] padframe/mprj_io_holdover[37] padframe/mprj_io_ib_mode_sel[37]
+ padframe/mprj_io_in[37] padframe/mprj_io_inp_dis[37] padframe/mprj_io_out[37] padframe/mprj_io_oeb[37]
+ padframe/mprj_io_slow_sel[37] padframe/mprj_io_vtrip_sel[37] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[37\]/serial_data_in gpio_control_in\[37\]/serial_data_out
+ mprj/io_in[37] mprj/io_oeb[37] mprj/io_out[37] gpio_control_in\[37\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[12\] soc/mgmt_in_data[12] gpio_control_in\[12\]/one soc/mgmt_in_data[12]
+ gpio_control_in\[12\]/one padframe/mprj_io_analog_en[12] padframe/mprj_io_analog_pol[12]
+ padframe/mprj_io_analog_sel[12] padframe/mprj_io_dm[36] padframe/mprj_io_dm[37]
+ padframe/mprj_io_dm[38] padframe/mprj_io_holdover[12] padframe/mprj_io_ib_mode_sel[12]
+ padframe/mprj_io_in[12] padframe/mprj_io_inp_dis[12] padframe/mprj_io_out[12] padframe/mprj_io_oeb[12]
+ padframe/mprj_io_slow_sel[12] padframe/mprj_io_vtrip_sel[12] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[12\]/serial_data_in gpio_control_in\[13\]/serial_data_in
+ mprj/io_in[12] mprj/io_oeb[12] mprj/io_out[12] gpio_control_in\[12\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xstorage soc/mgmt_addr[0] soc/mgmt_addr[1] soc/mgmt_addr[2] soc/mgmt_addr[3] soc/mgmt_addr[4]
+ soc/mgmt_addr[5] soc/mgmt_addr[6] soc/mgmt_addr[7] soc/mgmt_addr_ro[0] soc/mgmt_addr_ro[1]
+ soc/mgmt_addr_ro[2] soc/mgmt_addr_ro[3] soc/mgmt_addr_ro[4] soc/mgmt_addr_ro[5]
+ soc/mgmt_addr_ro[6] soc/mgmt_addr_ro[7] soc/core_clk soc/mgmt_ena[0] soc/mgmt_ena[1]
+ soc/mgmt_ena_ro soc/mgmt_rdata[0] soc/mgmt_rdata[10] soc/mgmt_rdata[11] soc/mgmt_rdata[12]
+ soc/mgmt_rdata[13] soc/mgmt_rdata[14] soc/mgmt_rdata[15] soc/mgmt_rdata[16] soc/mgmt_rdata[17]
+ soc/mgmt_rdata[18] soc/mgmt_rdata[19] soc/mgmt_rdata[1] soc/mgmt_rdata[20] soc/mgmt_rdata[21]
+ soc/mgmt_rdata[22] soc/mgmt_rdata[23] soc/mgmt_rdata[24] soc/mgmt_rdata[25] soc/mgmt_rdata[26]
+ soc/mgmt_rdata[27] soc/mgmt_rdata[28] soc/mgmt_rdata[29] soc/mgmt_rdata[2] soc/mgmt_rdata[30]
+ soc/mgmt_rdata[31] soc/mgmt_rdata[32] soc/mgmt_rdata[33] soc/mgmt_rdata[34] soc/mgmt_rdata[35]
+ soc/mgmt_rdata[36] soc/mgmt_rdata[37] soc/mgmt_rdata[38] soc/mgmt_rdata[39] soc/mgmt_rdata[3]
+ soc/mgmt_rdata[40] soc/mgmt_rdata[41] soc/mgmt_rdata[42] soc/mgmt_rdata[43] soc/mgmt_rdata[44]
+ soc/mgmt_rdata[45] soc/mgmt_rdata[46] soc/mgmt_rdata[47] soc/mgmt_rdata[48] soc/mgmt_rdata[49]
+ soc/mgmt_rdata[4] soc/mgmt_rdata[50] soc/mgmt_rdata[51] soc/mgmt_rdata[52] soc/mgmt_rdata[53]
+ soc/mgmt_rdata[54] soc/mgmt_rdata[55] soc/mgmt_rdata[56] soc/mgmt_rdata[57] soc/mgmt_rdata[58]
+ soc/mgmt_rdata[59] soc/mgmt_rdata[5] soc/mgmt_rdata[60] soc/mgmt_rdata[61] soc/mgmt_rdata[62]
+ soc/mgmt_rdata[63] soc/mgmt_rdata[6] soc/mgmt_rdata[7] soc/mgmt_rdata[8] soc/mgmt_rdata[9]
+ soc/mgmt_rdata_ro[0] soc/mgmt_rdata_ro[10] soc/mgmt_rdata_ro[11] soc/mgmt_rdata_ro[12]
+ soc/mgmt_rdata_ro[13] soc/mgmt_rdata_ro[14] soc/mgmt_rdata_ro[15] soc/mgmt_rdata_ro[16]
+ soc/mgmt_rdata_ro[17] soc/mgmt_rdata_ro[18] soc/mgmt_rdata_ro[19] soc/mgmt_rdata_ro[1]
+ soc/mgmt_rdata_ro[20] soc/mgmt_rdata_ro[21] soc/mgmt_rdata_ro[22] soc/mgmt_rdata_ro[23]
+ soc/mgmt_rdata_ro[24] soc/mgmt_rdata_ro[25] soc/mgmt_rdata_ro[26] soc/mgmt_rdata_ro[27]
+ soc/mgmt_rdata_ro[28] soc/mgmt_rdata_ro[29] soc/mgmt_rdata_ro[2] soc/mgmt_rdata_ro[30]
+ soc/mgmt_rdata_ro[31] soc/mgmt_rdata_ro[3] soc/mgmt_rdata_ro[4] soc/mgmt_rdata_ro[5]
+ soc/mgmt_rdata_ro[6] soc/mgmt_rdata_ro[7] soc/mgmt_rdata_ro[8] soc/mgmt_rdata_ro[9]
+ soc/mgmt_wdata[0] soc/mgmt_wdata[10] soc/mgmt_wdata[11] soc/mgmt_wdata[12] soc/mgmt_wdata[13]
+ soc/mgmt_wdata[14] soc/mgmt_wdata[15] soc/mgmt_wdata[16] soc/mgmt_wdata[17] soc/mgmt_wdata[18]
+ soc/mgmt_wdata[19] soc/mgmt_wdata[1] soc/mgmt_wdata[20] soc/mgmt_wdata[21] soc/mgmt_wdata[22]
+ soc/mgmt_wdata[23] soc/mgmt_wdata[24] soc/mgmt_wdata[25] soc/mgmt_wdata[26] soc/mgmt_wdata[27]
+ soc/mgmt_wdata[28] soc/mgmt_wdata[29] soc/mgmt_wdata[2] soc/mgmt_wdata[30] soc/mgmt_wdata[31]
+ soc/mgmt_wdata[3] soc/mgmt_wdata[4] soc/mgmt_wdata[5] soc/mgmt_wdata[6] soc/mgmt_wdata[7]
+ soc/mgmt_wdata[8] soc/mgmt_wdata[9] soc/mgmt_wen[0] soc/mgmt_wen[1] soc/mgmt_wen_mask[0]
+ soc/mgmt_wen_mask[1] soc/mgmt_wen_mask[2] soc/mgmt_wen_mask[3] soc/mgmt_wen_mask[4]
+ soc/mgmt_wen_mask[5] soc/mgmt_wen_mask[6] soc/mgmt_wen_mask[7] vccd vssd storage
Xgpio_control_in\[35\] soc/mgmt_in_data[35] gpio_control_in\[35\]/one soc/mgmt_in_data[35]
+ gpio_control_in\[35\]/one padframe/mprj_io_analog_en[35] padframe/mprj_io_analog_pol[35]
+ padframe/mprj_io_analog_sel[35] padframe/mprj_io_dm[105] padframe/mprj_io_dm[106]
+ padframe/mprj_io_dm[107] padframe/mprj_io_holdover[35] padframe/mprj_io_ib_mode_sel[35]
+ padframe/mprj_io_in[35] padframe/mprj_io_inp_dis[35] padframe/mprj_io_out[35] padframe/mprj_io_oeb[35]
+ padframe/mprj_io_slow_sel[35] padframe/mprj_io_vtrip_sel[35] soc/mprj_io_loader_resetn
+ soc/mprj_io_loader_clock gpio_control_in\[35\]/serial_data_in gpio_control_in\[36\]/serial_data_in
+ mprj/io_in[35] mprj/io_oeb[35] mprj/io_out[35] gpio_control_in\[35\]/zero vccd vssd
+ vccd1 vssd1 gpio_control_block
Xgpio_control_in\[3\] soc/mgmt_in_data[3] gpio_control_in\[3\]/one soc/mgmt_in_data[3]
+ gpio_control_in\[3\]/one padframe/mprj_io_analog_en[3] padframe/mprj_io_analog_pol[3]
+ padframe/mprj_io_analog_sel[3] padframe/mprj_io_dm[9] padframe/mprj_io_dm[10] padframe/mprj_io_dm[11]
+ padframe/mprj_io_holdover[3] padframe/mprj_io_ib_mode_sel[3] padframe/mprj_io_in[3]
+ padframe/mprj_io_inp_dis[3] padframe/mprj_io_out[3] padframe/mprj_io_oeb[3] padframe/mprj_io_slow_sel[3]
+ padframe/mprj_io_vtrip_sel[3] soc/mprj_io_loader_resetn soc/mprj_io_loader_clock
+ gpio_control_in\[3\]/serial_data_in gpio_control_in\[4\]/serial_data_in mprj/io_in[3]
+ mprj/io_oeb[3] mprj/io_out[3] gpio_control_in\[3\]/zero vccd vssd vccd1 vssd1 gpio_control_block
.ends

