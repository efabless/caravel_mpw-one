.SUBCKT icecap c0
*.PININFO c0:B
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch_levelshifter fbk fbk_n hold reset 
+ switch_lv switch_lv_n vgnd vpwr_hv vpwr_lv
*.PININFO hold:I reset:I switch_lv:I switch_lv_n:I fbk:O fbk_n:O vgnd:B 
*.PININFO vpwr_hv:B vpwr_lv:B
XICEnet97 net97 / icecap
XICEhold hold / icecap
XICEnet105 net105 / icecap
XICEfbk fbk / icecap
XICEfbk_n fbk_n / icecap
XICEreset reset / icecap
XICEnet109 net109 / icecap
XICEnet117 net117 / icecap
XICEswitch_lv_n switch_lv_n / icecap
XICEswitch_lv switch_lv / icecap
mI184 fbk reset vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI183 net97 vpwr_lv net109 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 fbk hold net105 vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI182 net105 vpwr_lv net117 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 net109 switch_lv vgnd vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 fbk_n hold net97 vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 net117 switch_lv_n vgnd vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI185 fbk_n fbk vpwr_hv vpwr_hv phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 fbk fbk_n vpwr_hv vpwr_hv phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch_s0 hold in_lv out_h reset vccd vdda vssa 
+ vssd
*.PININFO hold:I in_lv:I reset:I out_h:O vccd:B vdda:B vssa:B vssd:B
XICEnet17 net17 / icecap
XICEout_h out_h / icecap
XICEreset reset / icecap
XICEin_lv_n in_lv_n / icecap
XICEin_lv_i in_lv_i / icecap
XICEnet13 net13 / icecap
XICEhold hold / icecap
XICEin_lv in_lv / icecap
XI0 net17 net13 hold reset in_lv_i in_lv_n vssa vdda vccd / 
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
mI22 in_lv_n in_lv vssd vssd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 in_lv_i in_lv_n vssd vssd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 out_h net13 vssa vssa nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 in_lv_n in_lv vccd vccd phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 in_lv_i in_lv_n vccd vccd phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 out_h net13 vdda vdda phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch_sl hold in_lv out_h out_h_n reset vccd 
+ vdda vssa vssd vswitch
*.PININFO hold:I in_lv:I reset:I out_h:O out_h_n:O vccd:B vdda:B vssa:B vssd:B 
*.PININFO vswitch:B
XICEin_lv_i in_lv_i / icecap
XICEin_lv_n in_lv_n / icecap
XICEnet39 net39 / icecap
XICEhold hold / icecap
XICEout_h_n out_h_n / icecap
XICEout_h out_h / icecap
XICEnet48 net48 / icecap
XICEnet44 net44 / icecap
XICEin_lv in_lv / icecap
XICEnet35 net35 / icecap
XICEreset reset / icecap
mI14 out_h net44 vswitch vswitch phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 out_h_n net39 vdda vdda phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 in_lv_i in_lv_n vccd vccd phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 in_lv_n in_lv vccd vccd phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h net44 vssa vssa nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 out_h_n net39 vssa vssa nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 in_lv_i in_lv_n vssd vssd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI22 in_lv_n in_lv vssd vssd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI0 net39 net35 hold reset in_lv_i in_lv_n vssa vdda vccd / 
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
XI1 net48 net44 hold reset in_lv_i in_lv_n vssa vswitch vccd / 
+ sky130_fd_io__amuxsplitv2_switch_levelshifter
.ENDS
.SUBCKT s8_esd_res75only_small pad rout
*.PININFO pad:B rout:B
rI175 pad rout mrp1 m=1 w=2 l=3.15
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_switch amuxbus_l amuxbus_r ngate_sl_h ngate_sr_h 
+ nmid_h pgate_sl_h_n pgate_sr_h_n vdda vssa
*.PININFO ngate_sl_h:I ngate_sr_h:I nmid_h:I pgate_sl_h_n:I pgate_sr_h_n:I 
*.PININFO amuxbus_l:B amuxbus_r:B vdda:B vssa:B
XICEpgate_sl_h_n pgate_sl_h_n / icecap
XICEpgate_sr_h_n pgate_sr_h_n / icecap
XICEnmid_h nmid_h / icecap
XICEngate_sl_h ngate_sl_h / icecap
XICEamuxbus_l amuxbus_l / icecap
XICEngate_sr_h ngate_sr_h / icecap
XICEnmid_h_s nmid_h_s / icecap
XICEamuxbus_r amuxbus_r / icecap
XICEmid mid / icecap
xI20 mid vdda condiode
xI19 vssa vdda condiode
XI18 vssa nmid_h_s / s8_esd_res75only_small
mI1 amuxbus_l ngate_sl_h mid mid nhv m=30 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 mid ngate_sr_h amuxbus_r mid nhv m=30 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI4 mid nmid_h nmid_h_s vssa nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI0 mid pgate_sl_h_n amuxbus_l vdda phv m=14 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI3 amuxbus_r pgate_sr_h_n mid vdda phv m=14 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__hvsbt_nand2 in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 out in0 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out in1 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net25 vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net25 in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__amuxsplitv2_delay enable_vdda_h hld_vdda_h_n hold reset 
+ vcc_io vgnd
*.PININFO enable_vdda_h:I hld_vdda_h_n:I hold:O reset:O vcc_io:B vgnd:B
XICEhold hold / icecap
XICEhld_vdda_h hld_vdda_h / icecap
XICEreset reset / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEhld_vdda_h_n_switch hld_vdda_h_n_switch / icecap
XICEhld_vdda_h_n hld_vdda_h_n / icecap
XICEenable_vdda_switch enable_vdda_switch / icecap
XI33 enable_vdda_switch hld_vdda_h_n_switch reset vgnd vcc_io / 
+ sky130_fd_io__hvsbt_nand2
mI29 hld_vdda_h_n_switch hld_vdda_h vcc_io vcc_io phv m=2 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI28 hld_vdda_h hld_vdda_h_n vcc_io vcc_io phv m=1 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 enable_vdda_switch enable_vdda_h_n vcc_io vcc_io phv m=2 w=3.00 l=0.60 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 enable_vdda_h_n enable_vdda_h vcc_io vcc_io phv m=1 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 hold reset vcc_io vcc_io phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 hld_vdda_h_n_switch hld_vdda_h vgnd vgnd nhv m=2 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 hld_vdda_h hld_vdda_h_n vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 enable_vdda_switch enable_vdda_h_n vgnd vgnd nhv m=2 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 enable_vdda_h_n enable_vdda_h vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI37 hold reset vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__top_amuxsplitv2 amuxbus_a_l amuxbus_a_r amuxbus_b_l 
+ amuxbus_b_r enable_vdda_h hld_vdda_h_n switch_aa_s0 switch_aa_sl 
+ switch_aa_sr switch_bb_s0 switch_bb_sl switch_bb_sr vccd vcchib vdda vddio 
+ vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO enable_vdda_h:I hld_vdda_h_n:I switch_aa_s0:I switch_aa_sl:I 
*.PININFO switch_aa_sr:I switch_bb_s0:I switch_bb_sl:I switch_bb_sr:I 
*.PININFO amuxbus_a_l:B amuxbus_a_r:B amuxbus_b_l:B amuxbus_b_r:B vccd:B 
*.PININFO vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B 
*.PININFO vswitch:B
xI22 vssa vdda condiode
XI18 hold switch_aa_s0 ng_vdda_aa_s0_h reset vccd vdda vssa vssd / 
+ sky130_fd_io__amuxsplitv2_switch_s0
XI348 hold switch_bb_s0 ng_vdda_bb_s0_h reset vccd vdda vssa vssd / 
+ sky130_fd_io__amuxsplitv2_switch_s0
XI347 hold switch_aa_sl ng_vswitch_aa_sl_h pg_vdda_aa_sl_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI24 hold switch_aa_sr ng_vswitch_aa_sr_h pg_vdda_aa_sr_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI349 hold switch_bb_sr ng_vswitch_bb_sr_h pg_vdda_bb_sr_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI350 hold switch_bb_sl ng_vswitch_bb_sl_h pg_vdda_bb_sl_h_n reset vccd vdda 
+ vssa vssd vswitch / sky130_fd_io__amuxsplitv2_switch_sl
XI6 amuxbus_a_l amuxbus_a_r ng_vswitch_aa_sl_h ng_vswitch_aa_sr_h 
+ ng_vdda_aa_s0_h pg_vdda_aa_sl_h_n pg_vdda_aa_sr_h_n vdda vssa / 
+ sky130_fd_io__amuxsplitv2_switch
XI8 amuxbus_b_l amuxbus_b_r ng_vswitch_bb_sl_h ng_vswitch_bb_sr_h 
+ ng_vdda_bb_s0_h pg_vdda_bb_sl_h_n pg_vdda_bb_sr_h_n vdda vssa / 
+ sky130_fd_io__amuxsplitv2_switch
XI342 enable_vdda_h hld_vdda_h_n hold reset vdda vssa / 
+ sky130_fd_io__amuxsplitv2_delay
XICEnet27 enable_vdda_h / icecap
XICEamuxbus_b_r amuxbus_b_r / icecap
XICEswitch_aa_sl_h ng_vswitch_aa_sl_h / icecap
XICEamuxbus_a_l amuxbus_a_l / icecap
XICEswitch_bb_sl_h_n pg_vdda_bb_sl_h_n / icecap
XICEswitch_bb_sr_h ng_vswitch_bb_sr_h / icecap
XICEswitch_aa_s0_h ng_vdda_aa_s0_h / icecap
XICEswitch_aa_s0 hold / icecap
XICEswitch_aa_sr_h ng_vswitch_aa_sr_h / icecap
XICEswitch_aa_sl_h_n pg_vdda_aa_sl_h_n / icecap
XICEswitch_bb_sl_h ng_vswitch_bb_sl_h / icecap
XICEswitch_bb_s0_h ng_vdda_bb_s0_h / icecap
XICEswitch_bb_sr_h_n pg_vdda_bb_sr_h_n / icecap
XICEswitch_aa_sr_h_n pg_vdda_aa_sr_h_n / icecap
XI355 hold / icecap
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix p1g p1gb p2g padlo 
+ vgnd vpwr
*.PININFO padlo:I vgnd:I vpwr:I p1g:O p1gb:O p2g:O
XICEpadlo_bar padlo_bar / icecap
XICEp2gb p2gb / icecap
XICEp1gb p1gb / icecap
XICEp2g p2g / icecap
XICEp1g_new p1g_new / icecap
XICEp1g p1g / icecap
XICEpadlo padlo / icecap
XICEp2g_new p2g_new / icecap
mI76 p1g p1gb vpwr vpwr phv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI64 p1g_new padlo vpwr vpwr phv m=2 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI53 padlo_bar padlo vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI50 p2g_new p1g_new vpwr vpwr phv m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI49 p2g_new padlo_bar vpwr vpwr phv m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI65 p1g_new p2g_new vpwr vpwr phv m=2 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI77 p2g p2gb vpwr vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI70 p2gb p2g_new vpwr vpwr phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI72 p1gb p1g_new vpwr vpwr phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI54 padlo_bar padlo vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI69 p1g_new padlo net140 vgnd nhv m=1 w=1.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI78 p2g p2gb vgnd vgnd nhv m=2 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI67 net140 p2g_new vgnd vgnd nhv m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI71 p2gb p2g_new vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI79 p1g p1gb vgnd vgnd nhv m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI51 p2g_new padlo_bar net124 vgnd nhv m=1 w=1.00 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI73 p1gb p1g_new vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI52 net124 p1g_new vgnd vgnd nhv m=1 w=1.00 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix padlo pug4_h pug7_h tie_hi 
+ vpb_drvr
*.PININFO padlo:I tie_hi:I vpb_drvr:I pug4_h:O pug7_h:O
mI52 pug4_h padlo tie_hi vpb_drvr phv m=1 w=15.0 l=0.50 mult=1 sa=1.825 
+ sb=1.825 sd=280e-3 topography=normal area=0.063 perim=1.14
mI53 pug7_h padlo tie_hi vpb_drvr phv m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_nand2 in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpb phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out in1 vpwr vpb phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net25 vnb nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net25 in0 vgnd vnb nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_inv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vnb nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI1 out in vpwr vpb phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_nor in0 in1 out vgnd vnb vpb vpwr
*.PININFO in0:I in1:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEin0 in0 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
mI3 net17 in0 vpwr vpb phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out in1 net17 vpb phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in0 vgnd vnb nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out in1 vgnd vnb nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__tk_em1o a b
*.PININFO a:B b:B
rI1 a net11 short
rI2 b net7 short
.ENDS
.SUBCKT sky130_fd_io__tk_em1s a b
*.PININFO a:B b:B
rI1 a net8 short
rI2 b net8 short
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_dly in out out_n vcc_io vgnd
*.PININFO in:I vcc_io:I vgnd:I out:O out_n:O
XICEa5 a5 / icecap
XICEa3 a3 / icecap
XICEout out / icecap
XICEa2 a2 / icecap
XICEa7 a7 / icecap
XICEout_n out_n / icecap
XICEa4 a4 / icecap
XICEa6 a6 / icecap
XICEa1 a1 / icecap
XICEin in / icecap
XI228 out_n a5 / sky130_fd_io__tk_em1o
XI229 out_n a7 / sky130_fd_io__tk_em1o
XI227 a6 out / sky130_fd_io__tk_em1o
XI214 out_n a1 / sky130_fd_io__tk_em1o
XI215 a2 out / sky130_fd_io__tk_em1o
XEdly0 in out / sky130_fd_io__tk_em1o
XI217 out_n a3 / sky130_fd_io__tk_em1s
XEdly2 a4 out / sky130_fd_io__tk_em1s
mI196 a1 in vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI204 a4 a3 vgnd vgnd nhv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI199 a2 a1 vgnd vgnd nhv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI198 a3 a2 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI232 a5 a4 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI231 a6 a5 vgnd vgnd nhv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI230 a7 a6 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI197 a1 in vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI202 a4 a3 vcc_io vcc_io phv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI201 a2 a1 vcc_io vcc_io phv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI200 a3 a2 vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI235 a5 a4 vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI234 a6 a5 vcc_io vcc_io phv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI233 a7 a6 vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_log_i2c_fix dishs_h dishs_h_n en_h enhs_h 
+ enhs_h_n enhs_lat_h_n exiths_h forcehi_h<1> od_i_h_n vcc_io vgnd
*.PININFO en_h:I enhs_lat_h_n:I forcehi_h<1>:I od_i_h_n:I vcc_io:I vgnd:I 
*.PININFO dishs_h:O dishs_h_n:O enhs_h:O enhs_h_n:O exiths_h:O
XICEdishs_h_n dishs_h_n / icecap
XICEnet39 net39 / icecap
XICEdishs_h dishs_h / icecap
XICEnet74 net74 / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEen_h en_h / icecap
XICEenhs_dly_h_n enhs_dly_h_n / icecap
XICEenhs_h_n enhs_h_n / icecap
XICEnet46 net46 / icecap
XICEnet80 net80 / icecap
XICEforcehi_h<1> forcehi_h<1> / icecap
XICEenhs_dly_h enhs_dly_h / icecap
XICEexiths_h exiths_h / icecap
XICEenhs_lat_h_n enhs_lat_h_n / icecap
XICEenhs_h enhs_h / icecap
XI664 net39 net46 dishs_h vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_nand2
XI663 net80 forcehi_h<1> net46 vgnd vgnd vcc_io vcc_io / 
+ sky130_fd_io__sio_hvsbt_nand2
XI662 od_i_h_n en_h net39 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_nand2
XI658 od_i_h_n net80 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI666 enhs_lat_h_n net74 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI565 net74 enhs_h_n vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI667 dishs_h dishs_h_n vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI637 enhs_h_n enhs_h vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI553 net74 enhs_dly_h_n exiths_h vgnd vgnd vcc_io vcc_io / 
+ sky130_fd_io__sio_hvsbt_nor
XI521 net74 enhs_dly_h enhs_dly_h_n vcc_io vgnd / sky130_fd_io__sio_hotswap_dly
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_hys in out vcc_io vgnd
*.PININFO in:I vcc_io:I vgnd:I out:O
XICEvcc_io_buf vcc_io_buf / icecap
XICEout out / icecap
XICEvgnd_buf vgnd_buf / icecap
XICEin in / icecap
XICEint_p int_p / icecap
XICEint_n int_n / icecap
mI650 vcc_io_buf out int_n vgnd nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI649 int_n in vgnd vgnd nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI648 out in int_n vgnd nhv m=2 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI655 vgnd_buf vcc_io vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI647 vgnd_buf out int_p vcc_io phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI656 vcc_io_buf vgnd vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI646 out in int_p vcc_io phv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI645 int_p in vcc_io vcc_io phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_pghspd in1 in2 out vgnd
*.PININFO in1:I in2:I vgnd:I out:O
XICEin2 in2 / icecap
XICEnet25 net25 / icecap
XICEnet34 net34 / icecap
XICEnet27 net27 / icecap
XICEnet30 net30 / icecap
XICEnet42 net42 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
XICEnet38 net38 / icecap
XEin2b vgnd net25 / sky130_fd_io__tk_em1o
XEoutb net38 out / sky130_fd_io__tk_em1o
XEin1b vgnd net27 / sky130_fd_io__tk_em1o
XEin1a in1 net27 / sky130_fd_io__tk_em1s
XEouta net42 out / sky130_fd_io__tk_em1s
XEin2a in2 net25 / sky130_fd_io__tk_em1s
mI481 net50 in2 vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI507 out in1 net50 vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI651 net42 net27 net34 vgnd nhv m=6 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI654 net38 net27 net30 vgnd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI652 net34 net25 vgnd vgnd nhv m=6 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI653 net30 net25 vgnd vgnd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_hotswap_wpd en out vgnd
*.PININFO en:I vgnd:I out:O
XICEout out / icecap
XICEnpd<17> npd<17> / icecap
XICEen en / icecap
XICEnpd<14> npd<14> / icecap
XICEnpd<15> npd<15> / icecap
XICEnpd<18> npd<18> / icecap
XICEnpd<16> npd<16> / icecap
XI198 npd<15> npd<16> / sky130_fd_io__tk_em1o
XI209 vgnd npd<14> / sky130_fd_io__tk_em1o
XI196 npd<17> npd<18> / sky130_fd_io__tk_em1o
XI197 npd<16> npd<17> / sky130_fd_io__tk_em1o
XE20 npd<18> out / sky130_fd_io__tk_em1o
XI208 npd<14> npd<15> / sky130_fd_io__tk_em1o
mnen17 npd<17> en npd<16> vgnd nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnen15 npd<15> en npd<14> vgnd nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnen14 npd<14> en vgnd vgnd nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mnen16 npd<16> en npd<15> vgnd nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnen19 out en npd<18> vgnd nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mnen18 npd<18> en npd<17> vgnd nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_latch dishs_h dishs_h_n enhs_h enhs_h_n 
+ enhs_lat_h_n enhs_lathys_h_n exiths_h p3out pad_esd pghs_h vcc_io vgnd 
+ vpb_drvr vpwr_ka
*.PININFO dishs_h:I dishs_h_n:I enhs_h:I enhs_h_n:I exiths_h:I pad_esd:I 
*.PININFO vcc_io:I vgnd:I vpb_drvr:I vpwr_ka:I enhs_lat_h_n:O 
*.PININFO enhs_lathys_h_n:O p3out:O pghs_h:B
XI660 vgnd net102 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XI528 n6 net96 vgnd vgnd vcc_io vcc_io / sky130_fd_io__sio_hvsbt_inv_x1
XEhys2 enhs_lathys_h_n enhs_lat_h_n / sky130_fd_io__tk_em1o
XI658 net96 enhs_lat_h_n / sky130_fd_io__tk_em1s
XEhys1 net117 enhs_lathys_h_n / sky130_fd_io__tk_em1s
Xhys n6 net117 vcc_io vgnd / sky130_fd_io__sio_hotswap_hys
Xpghspd enhs_h n2 pghs_h vgnd / sky130_fd_io__sio_hotswap_pghspd
Xwpdenhs vpwr_ka net127 vgnd / sky130_fd_io__sio_hotswap_wpd
Xwpdexhs vpwr_ka net124 vgnd / sky130_fd_io__sio_hotswap_wpd
mI502 net186 pghs_h vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI484 net161 enhs_h pghs_h vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI491 n5 n6 vgnd vgnd nhv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI498 n2 n6 net124 vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI500 net170 enhs_h_n n2 vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mnexiths pghs_h exiths_h vgnd vgnd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI485 n3 n2 net161 vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI499 n4 pghs_h net170 vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI497 n6 n5 vgnd vgnd nhv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mndishs pghs_h dishs_h vgnd vgnd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI508 n2 enhs_h_n net186 vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI696 vgnd exiths_h vgnd vgnd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI487 pghs_h n5 net127 vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI697 vgnd dishs_h vgnd vgnd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI492 n5 n6 vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI503 n4 vgnd vcc_io vcc_io phv m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI488 n3 vgnd vcc_io vcc_io phv m=1 w=0.42 l=2.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI505 n6 n5 vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI493 n5 n3 vcc_io vcc_io phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI323 n2 dishs_h_n vcc_io vcc_io phv m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI279 n2 pad_esd vcc_io vcc_io phv m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI504 n6 n4 vcc_io vcc_io phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI689 p3out pad_esd vcc_io vpb_drvr phv m=12 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix en_h enhs_lat_h_n forcehi_h<1> 
+ od_i_h_n p3out pad_esd pghs_h vddio vpb_drvr vpwr_ka vssd
*.PININFO en_h:I forcehi_h<1>:I od_i_h_n:I pad_esd:I vddio:I vpb_drvr:I 
*.PININFO vpwr_ka:I vssd:I enhs_lat_h_n:O p3out:O pghs_h:B
XICEvpb_drvr vpb_drvr / icecap
XICEpghs_h pghs_h / icecap
XICEforcehi_h<1> forcehi_h<1> / icecap
XICEdishs_h dishs_h / icecap
XICEdishs_h_n dishs_h_n / icecap
XICEpad_esd pad_esd / icecap
XICEenhs_lathys_h_n enhs_lathys_h_n / icecap
XICEp3out p3out / icecap
XICEen_h en_h / icecap
XICEenhs_h_n enhs_h_n / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEenhs_h enhs_h / icecap
XICEenhs_lat_h_n enhs_lat_h_n / icecap
XICEexiths_h exiths_h / icecap
Xhslog dishs_h dishs_h_n en_h enhs_h enhs_h_n enhs_lathys_h_n exiths_h 
+ forcehi_h<1> od_i_h_n vddio vssd / sky130_fd_io__sio_hotswap_log_i2c_fix
Xhslatch dishs_h dishs_h_n enhs_h enhs_h_n enhs_lat_h_n enhs_lathys_h_n 
+ exiths_h p3out pad_esd pghs_h vddio vssd vpb_drvr vpwr_ka / 
+ sky130_fd_io__gpio_ovtv2_hotswap_latch
.ENDS
.SUBCKT sky130_fd_io__sio_tk_em1s a b
*.PININFO a:B b:B
rI1 a net8 short
rI2 b net8 short
.ENDS
.SUBCKT sky130_fd_io__sio_tk_em1o a b
*.PININFO a:B b:B
rI1 a net11 short
rI2 b net7 short
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_inv_x4 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vnb nhv m=4 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI1 out in vpwr vpb phv m=4 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghspu pad pghs_h pghs_h_latch tie_hi 
+ vcc_io_soft vpb_drvr
*.PININFO pad:I tie_hi:I vcc_io_soft:I vpb_drvr:I pghs_h:O pghs_h_latch:O
XEg9 tie_hi pg8 / sky130_fd_io__sio_tk_em1o
XEg2 pg2 vcc_io_soft / sky130_fd_io__sio_tk_em1s
XEg5 pg6 pg4 / sky130_fd_io__sio_tk_em1s
XEg4 pg4 pg3 / sky130_fd_io__sio_tk_em1s
XEpghs3 padhi3 pghs_h_latch / sky130_fd_io__sio_tk_em1s
XEg3 pg3 pg2 / sky130_fd_io__sio_tk_em1s
XEpghs7 padhi7 net36 / sky130_fd_io__sio_tk_em1s
XEg7 pg7 pg6 / sky130_fd_io__sio_tk_em1s
XEg8 pg8 pg7 / sky130_fd_io__sio_tk_em1s
XEpghs2 padhi2 padhi3 / sky130_fd_io__sio_tk_em1s
XEpghs8 pghs_h padhi7 / sky130_fd_io__sio_tk_em1s
XICEpg2 pg2 / icecap
XICEpadhi7 padhi7 / icecap
XICEpg3 pg3 / icecap
XICEpadhi6 net36 / icecap
XICEpg7 pg7 / icecap
XICEpadhi4 pghs_h_latch / icecap
XICEpg8 pg8 / icecap
XICEpg4 pg4 / icecap
XICEpadhi3 padhi3 / icecap
XICEpadhi2 padhi2 / icecap
XICEpadhi8 pghs_h / icecap
XICEpg5 pg6 / icecap
XICEtie_hi tie_hi / icecap
mpghs8 pghs_h pg8 pad vpb_drvr phv m=1 w=20.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpghs2 padhi2 pg2 pad vpb_drvr phv m=1 w=20.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpghs3 padhi3 pg3 pad vpb_drvr phv m=1 w=20.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpghs6 net36 pg6 pad vpb_drvr phv m=1 w=15.0 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mpghs4 pghs_h_latch pg4 pad vpb_drvr phv m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpghs7 padhi7 pg7 pad vpb_drvr phv m=1 w=20.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT s8_esd_signal_5_sym_hv_local_5term gate in nbody nwellRing vgnd
*.PININFO gate:I in:B nbody:B nwellRing:B vgnd:B
mI1 in gate vgnd nbody nhvesd m=1 w=5.40 l=0.60 mult=1 sa=0.0 sb=0.0 sd=0.0 
+ topography=normal area=0.048 perim=0.94
rI9 net18 nbody short
rI8 net16 nwellRing short
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix en_h force_h<1> od_i_h_n 
+ p3out pad padlo pghs_h tie_hi vcc_io_soft vddio vpb_drvr vpwr_ka vssd
*.PININFO en_h:I force_h<1>:I od_i_h_n:I pad:I tie_hi:I vcc_io_soft:I vddio:I 
*.PININFO vpb_drvr:I vpwr_ka:I vssd:I p3out:O padlo:O pghs_h:O
XICEtie_hi tie_hi / icecap
XICEen_h en_h / icecap
XICEenhs_latbuf_h_n enhs_latbuf_h_n / icecap
XICEpad pad / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEp3out p3out / icecap
XICEenhs_lat_h enhs_lat_h / icecap
XICEnet54 net54 / icecap
XICEforce_h<1> force_h<1> / icecap
XICEvcc_io_soft vcc_io_soft / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEenhs_lat_h_n enhs_lat_h_n / icecap
XICEnet50 net50 / icecap
XICEpadlo padlo / icecap
XICEpghs_h pghs_h / icecap
Xhsctl en_h enhs_lat_h_n force_h<1> od_i_h_n p3out pad net50 vddio vpb_drvr 
+ vpwr_ka vssd / sky130_fd_io__gpio_ovtv2_hotswap_ctl_i2c_fix
XI3 enhs_latbuf_h_n padlo / sky130_fd_io__sio_tk_em1s
XEpghs12 pghs_h net54 / sky130_fd_io__sio_tk_em1o
XI2 enhs_lat_h enhs_latbuf_h_n vssd vssd vddio vddio / 
+ sky130_fd_io__sio_hvsbt_inv_x4
XI1 enhs_lat_h_n enhs_lat_h vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x1
Xpghspu pad pghs_h net50 tie_hi vcc_io_soft vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pghspu
Xclamp vssd vddio vssd vddio pad / s8_esd_signal_5_sym_hv_local_5term
mpghs12 net54 padlo vpb_drvr vpb_drvr phv m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__sio_tk_tie_r_out_esd a b
*.PININFO a:B b:B
resd_r a b mrp1 m=1 w=0.5 l=10.2
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_pug pad padlo pug_h tie_hi vpb_drvr
*.PININFO pad:I padlo:I tie_hi:I vpb_drvr:I pug_h:O
XEg1 padlo net22 / sky130_fd_io__sio_tk_em1s
XI65 net24 tie_hi / sky130_fd_io__sio_tk_em1s
XEs2 net26 tie_hi / sky130_fd_io__sio_tk_em1s
XEs1 pad net26 / sky130_fd_io__sio_tk_em1o
XEg2 net22 net24 / sky130_fd_io__sio_tk_em1o
mI52 pug_h net22 net26 vpb_drvr phv m=1 w=15.0 l=0.50 mult=1 sa=1.825 sb=1.825 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI53 pug_h net24 net26 vpb_drvr phv m=1 w=15.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_bias pswg_h vcc_io vpb_drvr
*.PININFO pswg_h:I vcc_io:I vpb_drvr:O
XICEvpb_drvr vpb_drvr / icecap
XICEpswg_h pswg_h / icecap
mpsw_vccio vpb_drvr pswg_h vcc_io vpb_drvr phv m=22 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 vpb_drvr pswg_h vcc_io vpb_drvr phv m=9 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit pb pd pgin ps
*.PININFO pb:I pgin:I pd:B ps:B
XICEpd pd / icecap
XICEnet15 pgin / icecap
XICEpgin pgin / icecap
mpdrv pd pgin ps pb phvesd m=2 w=15.50 l=0.55 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias p2g pad soft_vcc_io tie_hi 
+ vpb_drvr
*.PININFO p2g:I pad:I soft_vcc_io:I tie_hi:I vpb_drvr:B
XICEsoft_vcc_io soft_vcc_io / icecap
XICEp2g p2g / icecap
XICEtie_hi tie_hi / icecap
Xpsw_pad4 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad0 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad3 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad2 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad5 vpb_drvr vpb_drvr soft_vcc_io pad / 
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
Xpsw_pad1 vpb_drvr vpb_drvr p2g pad / sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias_unit
XI5 tie_hi soft_vcc_io / sky130_fd_io__tk_em1o
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix force_h<1> nghs_h 
+ od_i_h_n oe_hs_h p2g pad pad_esd pghs_h pug_h<7> pug_h<6> pug_h<5> pug_h<4> 
+ pug_h<3> pug_h<2> pug_h<1> pug_h<0> vcc_io_soft vddio vpb_drvr vpwr_ka vssd
*.PININFO force_h<1>:I od_i_h_n:I oe_hs_h:I pad:I pad_esd:I vddio:I vpwr_ka:I 
*.PININFO vssd:I nghs_h:O p2g:O pghs_h:O vcc_io_soft:O vpb_drvr:O pug_h<7>:B 
*.PININFO pug_h<6>:B pug_h<5>:B pug_h<4>:B pug_h<3>:B pug_h<2>:B pug_h<1>:B 
*.PININFO pug_h<0>:B
Xnon_overlap p1g nghs_h p2g padlo vssd vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_nonoverlap_leak_fix
Xpug47 padlo pug_h<4> pug_h<7> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug_ovtfix
Xpghs oe_hs_h force_h<1> od_i_h_n net74 pad_esd padlo p1g tie_hi vcc_io_soft 
+ vddio vpb_drvr vpwr_ka vssd / sky130_fd_io__gpio_ovtv2_hotswap_pghs_i2c_fix
Xresd_tiehi vpb_drvr tie_hi / sky130_fd_io__sio_tk_tie_r_out_esd
Xresd_vccio vddio vcc_io_soft / sky130_fd_io__sio_tk_tie_r_out_esd
Xpug<3> pad_esd padlo pug_h<3> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<2> pad_esd padlo pug_h<2> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<1> pad_esd padlo pug_h<1> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<0> pad_esd padlo pug_h<0> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<6> pad_esd padlo pug_h<6> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xpug<5> pad_esd padlo pug_h<5> tie_hi vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_pug
Xp1_bias p1g vddio vpb_drvr / sky130_fd_io__gpio_ovtv2_hotswap_bias
Xp2p4_bias p2g pad vcc_io_soft vcc_io_soft vpb_drvr / 
+ sky130_fd_io__gpio_ovtv2_hotswap_vpb_bias
XICEnet84 vpb_drvr / icecap
XICEnet135 vpb_drvr / icecap
XICEod_h od_i_h_n / icecap
XICEp1g p1g / icecap
XICEnet89 vpb_drvr / icecap
XICEp2g p2g / icecap
XICEoe_hs_h oe_hs_h / icecap
XICEnet136 vpb_drvr / icecap
XICEnet148 tie_hi / icecap
XICEnet152 padlo / icecap
XICEforce_h<1> force_h<1> / icecap
XICEpadlo padlo / icecap
XICEnet149 p1g / icecap
XICEvcc_io_soft vcc_io_soft / icecap
XICEnet142 vpb_drvr / icecap
XICEtie_hi tie_hi / icecap
XICEvpb_drvr vpb_drvr / icecap
rI26 p2g net137 short
rI39 p2g net74 short
rI49 pghs_h p1g short
.ENDS
.SUBCKT sky130_fd_io__com_pad pad vgnd_io
*.PININFO pad:B vgnd_io:B
XICEpad pad / icecap
.ENDS
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_slow pad pd_h vcc_io vgnd_io
*.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
XICEpd_h pd_h / icecap
XICEpad pad / icecap
XICEvcc_io vcc_io / icecap
mndrv pad pd_h vgnd_io vgnd_io nhv m=4 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_pddrvr_weak pad pd_h vcc_io vgnd_io
*.PININFO pd_h:I vcc_io:I vgnd_io:I pad:O
XICEvcc_io vcc_io / icecap
XICEpd_h pd_h / icecap
XICEpad pad / icecap
mndrv1 pad pd_h vgnd_io vgnd_io nhv m=6 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_res_strong_slow ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
XICErb rb / icecap
XICEnet30 net30 / icecap
XICEra ra / icecap
XICEnet34 net34 / icecap
XI28 net34 net30 / sky130_fd_io__tk_em1s
rI32 rb net30 mrp1 m=1 w=2 l=2
rI29 net30 net34 mrp1 m=1 w=2 l=3
rr1 net34 ra mrp1 m=1 w=2 l=5
.ENDS
.SUBCKT sky130_fd_io__com_res_weak ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
XICEn<3> n<3> / icecap
XICEn<2> n<2> / icecap
XICErb rb / icecap
XICEn<0> n<0> / icecap
XICEn<4> n<4> / icecap
XICEra ra / icecap
XICEnet64 net64 / icecap
XICEn<1> n<1> / icecap
XICEn<5> n<5> / icecap
Xe9 n<0> n<1> / sky130_fd_io__tk_em1s
Xe11 n<2> n<3> / sky130_fd_io__tk_em1s
Xe10 n<1> n<2> / sky130_fd_io__tk_em1s
Xe12 n<3> rb / sky130_fd_io__tk_em1s
Xe13 n<4> n<0> / sky130_fd_io__tk_em1s
Xe14 n<5> n<4> / sky130_fd_io__tk_em1o
rI84 n<0> n<1> mrp1 m=1 w=0.8 l=1.5
rI62 n<3> rb mrp1 m=1 w=0.8 l=1.5
rI82 n<2> n<3> mrp1 m=1 w=0.8 l=1.5
rI85 ra net64 mrp1 m=1 w=0.8 l=50
rI83 n<1> n<2> mrp1 m=1 w=0.8 l=1.5
rI116 net64 n<5> mrp1 m=1 w=0.8 l=12
rI104 n<4> n<0> mrp1 m=1 w=0.8 l=6
rI134 n<5> n<4> mrp1 m=1 w=0.8 l=6
.ENDS
.SUBCKT sky130_fd_io__tk_tie_r_out_esd a b
*.PININFO a:B b:B
resd_r a b mrp1 m=1 w=0.5 l=10.2
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr_unit nd ngin ns
*.PININFO ngin:I nd:B ns:B
XICEngin ngin / icecap
XICEnet13 ngin / icecap
XICEnd nd / icecap
mndrv nd ngin ns ns nhvesd m=1 w=40.31 l=0.55 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pddrvr pad pd_csd pd_h<3> pd_h<2> tie_lo_esd vddio 
+ vssio vssio_q
*.PININFO pd_csd:I pd_h<3>:I pd_h<2>:I tie_lo_esd:O pad:B vddio:B vssio:B 
*.PININFO vssio_q:B
XICEpd_csd pd_csd / icecap
XICEpd_h<2> pd_h<2> / icecap
XICEpd_h<3> pd_h<3> / icecap
XICEpad pad / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XICEvssio_q vssio_q / icecap
XI26 vssio tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
Xn1 pad pd_h<2> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn2 pad pd_h<2> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn3 pad pd_h<2> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn8 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn7 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn6 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn5 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn9 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn10 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
Xn11 pad pd_h<3> vssio / sky130_fd_io__gpio_ovtv2_pddrvr_unit
rI8 vddio net96 short
mn14 pad pd_csd vssio_q vssio_q nhvesd m=1 w=40.31 l=0.55 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mn13 pad pd_csd vssio_q vssio_q nhvesd m=1 w=40.31 l=0.55 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
xI9 vssio vddio condiode
xI62 vssio_q vddio condiode
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_weak nghs_h pad pghs_h pu_h_n pug_h vddio 
+ vpb_drvr vssd vssio
*.PININFO nghs_h:I pghs_h:I pu_h_n:I vddio:I vpb_drvr:I vssd:I vssio:I pad:B 
*.PININFO pug_h:B
XICEnet26 net26 / icecap
XICEpghs_h pghs_h / icecap
XICEnghs_h nghs_h / icecap
XICEpad pad / icecap
XICEpug_h pug_h / icecap
XICEpu_h_n pu_h_n / icecap
XI36 pad net26 / sky130_fd_io__tk_em1o
mI51 pug_h nghs_h pu_h_n vssio nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI50 pu_h_n pghs_h pug_h vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpdrv pad pug_h vddio vpb_drvr phv m=3 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI35 net26 pug_h vddio vpb_drvr phv m=1 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 pad pug_h vddio vpb_drvr phv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow nghs_h pad pghs_h pu_h_n pug_h 
+ vddio vpb_drvr vssd vssio
*.PININFO nghs_h:I pghs_h:I pu_h_n:I vddio:I vpb_drvr:I vssd:I vssio:I pad:B 
*.PININFO pug_h:B
XICEvssio vssio / icecap
XICEpghs_h pghs_h / icecap
XICEnghs_h nghs_h / icecap
XICEpug_h pug_h / icecap
XICEpu_h_n pu_h_n / icecap
XICEpad pad / icecap
mI20 pug_h nghs_h pu_h_n vssio nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 pu_h_n pghs_h pug_h vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpdrv pad pug_h vddio vpb_drvr phv m=12 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__tk_em2o a b
*.PININFO a:B b:B
rI1 a net11 short
rI2 b net7 short
.ENDS
.SUBCKT sky130_fd_io__tk_em2s a b
*.PININFO a:B b:B
rI1 a net8 short
rI2 b net8 short
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5 pb pd pgin ps
*.PININFO pgin:I pb:B pd:B ps:B
XICEnet15 pgin / icecap
XICEpgin pgin / icecap
XICEpd pd / icecap
mpdrv pd pgin ps pb phvesd m=1 w=15.50 l=0.55 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pudrvr_strong nghs_h<4> nghs_h<3> nghs_h<2> pad 
+ pghs_h<4> pghs_h<3> pghs_h<2> pu_csd_h pu_h_n<3> pu_h_n<2> pug_h<4> pug_h<3> 
+ pug_h<2> tie_hi_esd vddio vddio_amx vpb_drvr vssd vssio
*.PININFO nghs_h<4>:I nghs_h<3>:I nghs_h<2>:I pghs_h<4>:I pghs_h<3>:I 
*.PININFO pghs_h<2>:I pu_csd_h:I pu_h_n<3>:I pu_h_n<2>:I vddio:I vssd:I 
*.PININFO vssio:I tie_hi_esd:O pad:B pug_h<4>:B pug_h<3>:B pug_h<2>:B 
*.PININFO vddio_amx:B vpb_drvr:B
XI155<0> vpb_drvr / icecap
XI155<1> vpb_drvr / icecap
XICEtie_hi_vpbdrvr tie_hi_vpbdrvr / icecap
XICEpug_h<2> pug_h<2> / icecap
XICEnet83 net83 / icecap
XICEvddio_amx vddio_amx / icecap
XICEpu_h_n<3> pu_h_n<3> / icecap
XICEpug_h<3> pug_h<3> / icecap
XICEpghs_h<3> pghs_h<3> / icecap
XICEnet81 net81 / icecap
XICEpug_h<4> pug_h<4> / icecap
XICEpghs_h<4> pghs_h<4> / icecap
XICEnghs_h<4> nghs_h<4> / icecap
XICEpu_csd_h pu_csd_h / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XICEpghs_h<2> pghs_h<2> / icecap
XICEnghs_h<2> nghs_h<2> / icecap
XICEnet079 net079 / icecap
XICEpu_h_n<2> pu_h_n<2> / icecap
XICEnghs_h<3> nghs_h<3> / icecap
XICEnet79 net79 / icecap
XICEpad pad / icecap
XI49 vddio tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
XI133 vpb_drvr tie_hi_vpbdrvr / sky130_fd_io__tk_tie_r_out_esd
XI112 pug_h<2> net83 / sky130_fd_io__tk_em2o
XI111 pug_h<4> net81 / sky130_fd_io__tk_em2o
XI141 pug_h<3> net79 / sky130_fd_io__tk_em2o
XI152 pug_h<4> net079 / sky130_fd_io__tk_em2o
XI142 tie_hi_vpbdrvr net79 / sky130_fd_io__tk_em2s
XI82 tie_hi_vpbdrvr net83 / sky130_fd_io__tk_em2s
XI109 tie_hi_vpbdrvr net81 / sky130_fd_io__tk_em2s
XI153 tie_hi_vpbdrvr net079 / sky130_fd_io__tk_em2s
Xn7 vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn6 vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<2> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<1> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn5<0> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn4 vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<3> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<2> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<1> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn2<0> vpb_drvr pad net83 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<1> vpb_drvr pad net79 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn9<0> vpb_drvr pad net79 vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<1> vpb_drvr pad pug_h<4> vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn11<0> vpb_drvr pad pug_h<4> vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<1> vpb_drvr pad net81 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn12<0> vpb_drvr pad net81 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<1> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn1<0> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<1> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn3<0> vpb_drvr pad pug_h<2> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<1> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn8<0> vpb_drvr pad pug_h<3> vddio / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<1> vpb_drvr pad net079 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
Xn10<0> vpb_drvr pad net079 vddio_amx / sky130_fd_io__gpio_ovtv2_pudrvr_unit_2_5
mI136 pug_h<4> nghs_h<4> pu_csd_h vssio nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI127 pug_h<2> nghs_h<2> pu_h_n<2> vssio nhv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 pug_h<3> nghs_h<3> pu_h_n<3> vssio nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI137 pu_csd_h pghs_h<4> pug_h<4> vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI128 pu_h_n<2> pghs_h<2> pug_h<2> vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 pu_h_n<3> pghs_h<3> pug_h<3> vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_sub nghs_h pad pad_esd pd_csd_h pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pghs_h pu_csd_h pu_h_n<3> pu_h_n<2> pu_h_n<1> 
+ pu_h_n<0> pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> tie_hi_esd tie_lo_esd 
+ vddio vddio_amx vpb_drvr vssd vssio vssio_amx
*.PININFO nghs_h:I pd_csd_h:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pghs_h:I 
*.PININFO pu_csd_h:I pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vddio:I 
*.PININFO vssd:I vssio:I vssio_amx:I pad:B pad_esd:B pug_h<4>:B pug_h<3>:B 
*.PININFO pug_h<2>:B pug_h<1>:B pug_h<0>:B tie_hi_esd:B tie_lo_esd:B 
*.PININFO vddio_amx:B vpb_drvr:B
Xpddrvr_strong_slow strong_slow_pad pd_h<1> vddio vssio / 
+ sky130_fd_io__gpio_pddrvr_strong_slow
XI73 weak_pad pd_h<0> vddio vssio / sky130_fd_io__gpio_pddrvr_weak
Xres strong_slow_pad pad_esd vssio / sky130_fd_io__com_res_strong_slow
Xres_weak weak_pad pad_esd vssio / sky130_fd_io__com_res_weak
Xpd_drvr pad pd_csd_h pd_h<3> pd_h<2> tie_lo_esd vddio vssio vssio_amx / 
+ sky130_fd_io__gpio_ovtv2_pddrvr
Xpudrvr_weak nghs_h weak_pad pghs_h pu_h_n<0> pug_h<0> vddio vpb_drvr vssd 
+ vssio / sky130_fd_io__gpio_ovtv2_pudrvr_weak
Xstrong_slow_pudrvr nghs_h strong_slow_pad pghs_h pu_h_n<1> pug_h<1> vddio 
+ vpb_drvr vssd vssio / sky130_fd_io__gpio_ovtv2_pudrvr_strong_slow
Xpudrvr_strong nghs_h nghs_h nghs_h pad pghs_h pghs_h pghs_h pu_csd_h 
+ pu_h_n<3> pu_h_n<2> pug_h<4> pug_h<3> pug_h<2> tie_hi_esd vddio vddio_amx 
+ vpb_drvr vssd vssio / sky130_fd_io__gpio_ovtv2_pudrvr_strong
Xres_esd pad_esd pad / s8_esd_res75only_small
xI72 vssio vddio condiode
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix force_h<1> nga_pad_vpmp_h 
+ ngb_pad_vpmp_h nghs_h od_i_h_n oe_hs_h pad pd_csd_h pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pghs_h pu_csd_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<7> 
+ pug_h<6> pug_h<5> tie_hi_esd tie_lo_esd vddio vddio_amx vpb_drvr vssa vssd 
+ vssio vssio_amx
*.PININFO force_h<1>:I nga_pad_vpmp_h:I ngb_pad_vpmp_h:I od_i_h_n:I oe_hs_h:I 
*.PININFO pd_csd_h:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pu_csd_h:I 
*.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vddio:I vssa:I 
*.PININFO vssd:I vssio:I vssio_amx:I nghs_h:O pad:O pghs_h:O tie_hi_esd:O 
*.PININFO tie_lo_esd:O pug_h<7>:B pug_h<6>:B pug_h<5>:B vddio_amx:B vpb_drvr:B
XICEnghs_h nghs_h / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XICEpad_esd pad_esd / icecap
XICEpd_csd_h pd_csd_h / icecap
XICEpghs_h pghs_h / icecap
XICEoe_hs_h oe_hs_h / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEpu_csd_h pu_csd_h / icecap
XICEnet74 net74 / icecap
XI196<0> pu_h_n<3> / icecap
XI196<1> pu_h_n<2> / icecap
XI196<2> pu_h_n<1> / icecap
XI196<3> pu_h_n<0> / icecap
XICEp2g p2g / icecap
XI195<0> pd_h<3> / icecap
XI195<1> pd_h<2> / icecap
XI195<2> pd_h<1> / icecap
XI199<0> pug_h<4> / icecap
XI199<1> pug_h<3> / icecap
XI199<2> pug_h<2> / icecap
XI199<3> pug_h<1> / icecap
XI199<4> pug_h<0> / icecap
XICEforce_h<1> force_h<1> / icecap
XICEpad pad / icecap
XI194<0> pd_h<3> / icecap
XI194<1> pd_h<2> / icecap
XI194<2> pd_h<1> / icecap
XI194<3> pd_h<0> / icecap
XI197<0> pd_csd_h / icecap
XI197<1> nga_pad_vpmp_h / icecap
XI197<2> ngb_pad_vpmp_h / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XI198<0> pug_h<7> / icecap
XI198<1> pug_h<6> / icecap
XI198<2> pug_h<5> / icecap
XI198<3> pug_h<4> / icecap
XI198<4> pug_h<3> / icecap
XI198<5> pug_h<2> / icecap
XI198<6> pug_h<1> / icecap
XI198<7> pug_h<0> / icecap
Xhotswap force_h<1> nghs_h od_i_h_n oe_hs_h p2g pad pad_esd pghs_h pug_h<7> 
+ pug_h<6> pug_h<5> pug_h<4> pug_h<3> pug_h<2> pug_h<1> pug_h<0> net74 vddio 
+ vpb_drvr vddio vssd / sky130_fd_io__gpio_ovtv2_hotswap_i2c_fix_leak_fix
Xbondpad pad vssio / sky130_fd_io__com_pad
Xodrvr tie_hi_esd pad pad_esd pd_csd_h pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h 
+ pu_csd_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<4> pug_h<3> pug_h<2> 
+ pug_h<1> pug_h<0> tie_hi_esd tie_lo_esd vddio vddio_amx vpb_drvr vssd vssio 
+ vssio_amx / sky130_fd_io__gpio_ovtv2_odrvr_sub
mI122<2> pd_h<3> pghs_h net106<0> vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI122<1> pd_h<2> pghs_h net106<1> vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI122<0> pd_h<1> pghs_h net106<2> vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI85<2> net106<0> pghs_h vssio vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI85<1> net106<1> pghs_h vssio vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI85<0> net106<2> pghs_h vssio vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI104<2> net102<0> pghs_h vssa vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI104<1> net102<1> pghs_h vssa vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI104<0> net102<2> pghs_h vssa vssio nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI103<2> pd_csd_h pghs_h net102<0> vssio nhv m=1 w=0.42 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI103<1> nga_pad_vpmp_h pghs_h net102<1> vssio nhv m=1 w=0.42 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI103<0> ngb_pad_vpmp_h pghs_h net102<2> vssio nhv m=1 w=0.42 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nor3_dnw in0 in1 in2 out vgnd vpwr
*.PININFO in0:I in1:I in2:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
XICEin2 in2 / icecap
mI3 net43 in0 vpwr vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 net39 in1 net43 vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 out in2 net39 vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in0 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out in1 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 out in2 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_inv_x1_dnw in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEin in / icecap
XICEout out / icecap
mI1 out in vpwr vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 out in vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_nand2_dnw in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out in1 vpwr vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net25 vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net25 in0 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_nor2_dnw in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEin1 in1 / icecap
XICEin0 in0 / icecap
XICEout out / icecap
mI3 net17 in0 vpwr vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out in1 net17 vpwr phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in0 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out in1 vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_predrvr_switch nmos_en pmos_en sig1 sig2 vcc_io 
+ vgnd_io
*.PININFO nmos_en:I pmos_en:I vcc_io:I vgnd_io:I sig1:B sig2:B
XICEpmos_en pmos_en / icecap
XICEsig1 sig1 / icecap
XICEnmos_en nmos_en / icecap
XICEsig2 sig2 / icecap
mI374 sig1 nmos_en sig2 vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI375 sig2 pmos_en sig1 vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix drvlo_h_n en_cmos_b 
+ i2c_mode_h_n nghs_h nsw_en_int oe_i_h_n pad_cap pd_dis_h pd_h<3> pd_h<2> 
+ pden_h_n<1> pghs_h pug_h slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> 
+ slew_ctl_h_n<0> slow_h_n vcc_io vgnd_io vpb_drvr vssd
*.PININFO drvlo_h_n:I i2c_mode_h_n:I nghs_h:I oe_i_h_n:I pd_dis_h:I 
*.PININFO pden_h_n<1>:I pghs_h:I pug_h:I slew_ctl_h<1>:I slew_ctl_h<0>:I 
*.PININFO slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I slow_h_n:I vcc_io:I vgnd_io:I 
*.PININFO vpb_drvr:I vssd:I en_cmos_b:O nsw_en_int:O pd_h<3>:O pd_h<2>:O 
*.PININFO pad_cap:B
XICEnsw_en_int nsw_en_int / icecap
XICEpug_h pug_h / icecap
XI319<0> cas3 / icecap
XI319<1> cas10 / icecap
XICEen_cmos_b en_cmos_b / icecap
XICEcas4 cas4 / icecap
XICEnet200 net200 / icecap
XICEna na / icecap
XICEnet519 net519 / icecap
XICEvdiode vdiode / icecap
XICEslew_ctl_h_n<1> slew_ctl_h_n<1> / icecap
XICEnet400 net400 / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEcas2 cas2 / icecap
XICEslew_ctl_h<0> slew_ctl_h<0> / icecap
XICEne ne / icecap
XICEnet336 net336 / icecap
XICEpd_h<3> pd_h<3> / icecap
XICEdrvlo_h_n_i2c_4 drvlo_h_n_i2c_4 / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEcas5 cas5 / icecap
XICEslew_ctl_h<1> slew_ctl_h<1> / icecap
XICEnet278 net278 / icecap
XICEnet352 net352 / icecap
XICEnet404 net404 / icecap
XICEbiasp biasp / icecap
XI318<0> na / icecap
XI318<1> nb / icecap
XI318<2> nc / icecap
XI318<3> nd / icecap
XI318<4> ne / icecap
XI318<5> nf / icecap
XICEenb enb / icecap
XICEnet263 net263 / icecap
XICEcas10 cas10 / icecap
XICEnet303 net303 / icecap
XICEnet369 net369 / icecap
XICEnet288 net288 / icecap
XICEmode2b mode2b / icecap
XICEpad_cap pad_cap / icecap
XICEdrvlo_h_n_i2c_1 drvlo_h_n_i2c_1 / icecap
XICEnet313 net313 / icecap
XICEdrvlo_h_n_buf drvlo_h_n_buf / icecap
XICEen en / icecap
XICEnet531 net531 / icecap
XICEnet298 net298 / icecap
XICEnet193 net193 / icecap
XICEnet420 net420 / icecap
XICEvr vr / icecap
XICEnet388 net388 / icecap
XICEnc nc / icecap
XICEnet552 pd_h<3> / icecap
XICEnet318 net318 / icecap
XICEnet535 net535 / icecap
XICEslew_ctl_h_n<0> slew_ctl_h_n<0> / icecap
XICEpd_h<2> pd_h<2> / icecap
XICEnsw_en nsw_en / icecap
XICEdrvlo_h_n_i2c_2 drvlo_h_n_i2c_2 / icecap
XICEnet499 vcc_io / icecap
XICEnet283 net283 / icecap
XICEnghs_h nghs_h / icecap
XICEpd_dis_h pd_dis_h / icecap
XICE2vtn N0 / icecap
XICEvdelay vdelay / icecap
XICEnsw_enb nsw_enb / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEdrvlo_h drvlo_h / icecap
XICEmode3b mode3b / icecap
XICEnet613 net352 / icecap
XICEnf nf / icecap
XICEpghs_h pghs_h / icecap
XICEnet190 net190 / icecap
XICEbiasp1 biasp1 / icecap
XICEpden_h<1> pden_h<1> / icecap
XICEmode1b mode1b / icecap
XICEnb nb / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEdrvlo_h_n_i2c drvlo_h_n_i2c / icecap
XICEslow_h_n slow_h_n / icecap
XICEcas3 cas3 / icecap
XICEdrvlo_h_n_i2c_3 drvlo_h_n_i2c_3 / icecap
XICEnet293 net293 / icecap
XICEnd nd / icecap
rI288 N0 net193 mrdn_hv m=1 w=0.5 l=113.375 isHV=TRUE
rI287 vdiode net190 mrdn_hv m=1 w=0.5 l=113.375 isHV=TRUE
XI123 pd_dis_h nsw_enb oe_i_h_n net200 vgnd_io vcc_io / sky130_fd_io__nor3_dnw
xI208 vgnd_io vcc_io condiode
XI161 net293 drvlo_h_n_i2c_2 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI159 net298 drvlo_h_n_i2c_1 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI224 net288 net247 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI605 en enb vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI176 net318 drvlo_h_n_i2c_4 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI191 nsw_en nsw_enb vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI198 net303 drvlo_h_n_i2c vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI179 net283 nsw_en_int vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI168 net263 mode1b vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI122 drvlo_h drvlo_h_n_buf vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI170 net278 mode3b vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI715 pden_h_n<1> pden_h<1> vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI162 net313 drvlo_h_n_i2c_3 vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI254 drvlo_h_n drvlo_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
XI602 vdelay net200 en vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
XI112 pden_h<1> nsw_enb en_cmos_b vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
XI430 slew_ctl_h<1> slew_ctl_h_n<0> net263 vgnd_io vcc_io / 
+ sky130_fd_io__com_nand2_dnw
XI175 drvlo_h_n_i2c mode4b net318 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI163 drvlo_h_n_i2c mode3b net313 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI109 slow_h_n i2c_mode_h_n nsw_en vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI197 nsw_enb drvlo_h_n_buf net303 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI158 drvlo_h_n_i2c mode1b net298 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI160 drvlo_h_n_i2c mode2b net293 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI225 slew_ctl_h<1> slew_ctl_h<0> net288 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI181 pden_h_n<1> nsw_en net283 vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
XI169 slew_ctl_h<1> slew_ctl_h_n<0> net278 vgnd_io vcc_io / 
+ sky130_fd_io__com_nor2_dnw
xI99 net0101 net0100 net099 net098 xcmvpp8p6x7p9_m3shield m=18
mI206 N0 en vgnd_io vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI190 net531 en vgnd_io vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI220 net420 enb vgnd_io vgnd_io nhv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI153 pd_h<2> pden_h_n<1> vgnd_io vgnd_io nhv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI182 vgnd_io vdelay vgnd_io vgnd_io nhv m=4 w=5.00 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI201 net352 N0 net190 vgnd_io nhvnative m=10 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI625 net404 pd_h<3> net348 vgnd_io nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI339 net400 pden_h<1> vgnd_io vgnd_io nhv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI125 pd_h<3> drvlo_h_n_buf net400 vgnd_io nhv m=4 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI344 pd_h<3> pden_h_n<1> vgnd_io vgnd_io nhv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI63 net388 vdiode pd_h<3> vgnd_io nhvnative m=2 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI189 net388 vgnd_io vgnd_io vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI10 biasp vdiode net336 vgnd_io nhvnative m=5 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI374 net519 nsw_en pd_h<3> vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI137 biasp1 vdiode vgnd_io vgnd_io nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 net369 net369 vgnd_io vgnd_io nhv m=5 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 vdiode vdiode vgnd_io vgnd_io nhv m=5 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI165 vdiode en vgnd_io vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 N0 N0 net369 vgnd_io nhv m=5 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 net352 N0 net190 vgnd_io nhvnative m=4 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI755 net348 pd_h<3> vgnd_io vgnd_io nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI579 vdelay drvlo_h net404 vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI192 net519 vgnd_io vgnd_io vgnd_io nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI219 net336 vdiode vr vgnd_io nlowvt m=5 w=7.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI232<1> cas3 pghs_h pd_h<3> vgnd_io nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI232<0> cas10 pghs_h pd_h<3> vgnd_io nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI278 vgnd_io vgnd_io vgnd_io vgnd_io nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 pug_h nghs_h nsw_enb vgnd_io nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI245 cas10 vcc_io cas4 vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI196 nc biasp vcc_io vcc_io pshort m=5 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI200 cas3 biasp1 nc vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI199 pd_h<3> drvlo_h_n_i2c_2 cas3 vcc_io phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI205 net352 en vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI156 cas5 biasp1 ne vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI580 vdelay drvlo_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI136 biasp biasp1 na vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI144 cas4 biasp1 nd vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI84 pd_h<3> drvlo_h_n_i2c cas2 vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI230 nc vcc_io vcc_io vcc_io pshort m=1 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI79 nb biasp vcc_io vcc_io pshort m=17 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI260 net535 enb vcc_io vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI228 pd_h<3> drvlo_h_n_i2c net535 vcc_io phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI73 net388 drvlo_h_n_i2c net531 vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI561 pd_h<3> drvlo_h_n_i2c_1 cas4 vcc_io phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI560 nd biasp vcc_io vcc_io pshort m=14 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI375 pd_h<3> pug_h net519 vpb_drvr phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI164 biasp enb vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI167 biasp1 enb vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI138 biasp1 biasp1 vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI145 cas2 biasp1 nb vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI141 na biasp vcc_io vcc_io pshort m=10 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI154 ne biasp vcc_io vcc_io pshort m=14 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI178 net193 en vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI155 pd_h<3> drvlo_h_n_i2c_3 cas5 vcc_io phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI241 cas10 biasp1 nf vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI240 nf biasp vcc_io vcc_io pshort m=8 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI229 ne vcc_io vcc_io vcc_io pshort m=2 w=0.55 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI217 nb vcc_io vcc_io vcc_io pshort m=3 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI216 nd vcc_io vcc_io vcc_io pshort m=2 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI215 cas3 vcc_io cas2 vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI214 cas5 vcc_io cas2 vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI239 pd_h<3> drvlo_h_n_i2c_3 cas10 vcc_io phv m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI213 cas3 vcc_io cas4 vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI212 na vcc_io vcc_io vcc_io pshort m=2 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI211 vcc_io vcc_io vcc_io vcc_io pshort m=4 w=0.55 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI210 vcc_io vcc_io vcc_io vcc_io pshort m=6 w=0.55 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI248<5> na enb vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI248<4> nb enb vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI248<3> nc enb vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI248<2> nd enb vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI248<1> ne enb vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI248<0> nf enb vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 nsw_enb pghs_h pug_h vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI70 net531 en vcc_io vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
XI94 nsw_en nsw_enb pd_h<2> pd_h<3> vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_predrvr_switch
rI221 net420 vr mrp1 m=1 w=0.75 l=513.445
rI186 slew_ctl_h_n<0> mode4b short
rI157 net247 mode2b short
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix drvlo_h_n en_cmos_b 
+ i2c_mode_h_n nghs_h nsw_en oe_i_h_n pad pd_dis_h pd_h<3> pd_h<2> pden_h_n<1> 
+ pghs_h pug_h slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> 
+ slow_h_n vcc_io vgnd_io vpb_drvr vssd
*.PININFO drvlo_h_n:I i2c_mode_h_n:I nghs_h:I oe_i_h_n:I pd_dis_h:I 
*.PININFO pden_h_n<1>:I pghs_h:I pug_h:I slew_ctl_h<1>:I slew_ctl_h<0>:I 
*.PININFO slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I slow_h_n:I vcc_io:I vgnd_io:I 
*.PININFO vpb_drvr:I vssd:I en_cmos_b:O nsw_en:O pd_h<3>:O pd_h<2>:O pad:B
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEpad pad / icecap
XICEvssd vssd / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEpug_h pug_h / icecap
XICEpghs_h pghs_h / icecap
XICEen_cmos_b en_cmos_b / icecap
XI89<0> slew_ctl_h<1> / icecap
XI89<1> slew_ctl_h<0> / icecap
XICEnghs_h nghs_h / icecap
XI88<0> pd_h<3> / icecap
XI88<1> pd_h<2> / icecap
XICEslow_h_n slow_h_n / icecap
XICEnsw_en nsw_en / icecap
XICEpd_dis_h pd_dis_h / icecap
XI90<0> slew_ctl_h_n<1> / icecap
XI90<1> slew_ctl_h_n<0> / icecap
XICEvpb_drvr vpb_drvr / icecap
Xpd_strong drvlo_h_n en_cmos_b i2c_mode_h_n nghs_h nsw_en oe_i_h_n pad 
+ pd_dis_h pd_h<3> pd_h<2> pden_h_n<1> pghs_h pug_h slew_ctl_h<1> 
+ slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> slow_h_n vcc_io vgnd_io 
+ vpb_drvr vssd / sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_leak_fix
.ENDS
.SUBCKT sky130_fd_io__com_pupredrvr_strong_slow drvhi_h pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XICEnet17 net17 / icecap
XICEdrvhi_h drvhi_h / icecap
XICEpu_h_n pu_h_n / icecap
XICEpuen_h puen_h / icecap
mI3 pu_h_n drvhi_h net17 vgnd_io nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI39 net17 puen_h vgnd_io vgnd_io nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI38 pu_h_n puen_h vcc_io vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI37 pu_h_n drvhi_h vcc_io vcc_io phv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_pupredrvr_weak drvhi_h pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XICEpu_h_n pu_h_n / icecap
XICEpuen_h puen_h / icecap
XICEdrvhi_h drvhi_h / icecap
mI3 pu_h_n drvhi_h net21 vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI39 net21 puen_h vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI38 pu_h_n puen_h vcc_io vcc_io phv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI37 pu_h_n drvhi_h vcc_io vcc_io phv m=2 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_pdpredrvr_weak drvlo_h_n pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
XICEdrvlo_h_n drvlo_h_n / icecap
XICEpd_h pd_h / icecap
XICEnet25 net25 / icecap
XICEpden_h_n pden_h_n / icecap
mI26 pd_h pden_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 pd_h drvlo_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 net25 pden_h_n vcc_io vcc_io phv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI23 pd_h drvlo_h_n net25 vcc_io phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_pdpredrvr_strong_slow drvlo_h_n pd_h pden_h_n vcc_io 
+ vgnd_io
*.PININFO drvlo_h_n:I pden_h_n:I vcc_io:I vgnd_io:I pd_h:O
XICEdrvlo_h_n drvlo_h_n / icecap
XICEpd_h pd_h / icecap
XICEnet25 net25 / icecap
XICEpden_h_n pden_h_n / icecap
mI26 pd_h pden_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 pd_h drvlo_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 net25 pden_h_n vcc_io vcc_io phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI23 pd_h drvlo_h_n net25 vcc_io phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__tk_opto out spd spu
*.PININFO out:B spd:B spu:B
Xe1 spu out / sky130_fd_io__tk_em1o
Xe2 out spd / sky130_fd_io__tk_em1s
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias drvlo_h_n en_h en_h_n pbias pd_h 
+ pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_h:I en_h_n:I pd_h:I pden_h_n:I vcc_io:I vgnd_io:I 
*.PININFO pbias:O
XICEbias_g bias_g / icecap
XICEpbias pbias / icecap
XICEnet183 net183 / icecap
XICEpden_h_n pden_h_n / icecap
XICEen_h en_h / icecap
XICEn<101> n<101> / icecap
XICEnet157 net157 / icecap
XICEnet108 net108 / icecap
XICEnet171 net171 / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEdrvlo_i_h drvlo_i_h / icecap
XICEen_h_n en_h_n / icecap
XICEnet84 net84 / icecap
XICEpbias1 pbias1 / icecap
XICE2vtp N0 / icecap
XICEn<0> n<0> / icecap
XICEpd_h pd_h / icecap
XICEnet88 net88 / icecap
XICEn<1> n<1> / icecap
XICEnet161 net161 / icecap
XE1 n<1> n<0> / sky130_fd_io__tk_em1o
XE2 pbias pbias1 / sky130_fd_io__tk_em1o
XE3 pbias1 net88 / sky130_fd_io__tk_em1s
XE4 net108 pbias / sky130_fd_io__tk_em1s
XE6 pbias net84 / sky130_fd_io__tk_em1s
XE5 n<101> bias_g / sky130_fd_io__tk_em1s
XI27 n<0> pd_h en_h_n / sky130_fd_io__tk_opto
mI47 pbias bias_g vgnd_io vgnd_io nhv m=2 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 n<1> drvlo_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 bias_g drvlo_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI23 n<0> n<0> n<1> vgnd_io nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 drvlo_i_h drvlo_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 bias_g n<1> vgnd_io vgnd_io nhv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 bias_g en_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI34 net157 bias_g vgnd_io vgnd_io nhv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 net108 bias_g vgnd_io vgnd_io nhv m=2 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI38 n<1> pden_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI48 n<100> pd_h vgnd_io vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI41 n<101> pd_h n<100> vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI44 pbias pbias pbias1 vcc_io phv m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI45 pbias1 pbias1 vcc_io vcc_io phv m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 net183 en_h_n vcc_io vcc_io phv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 net171 n<0> net183 vcc_io phv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 pbias en_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 drvlo_i_h drvlo_h_n vcc_io vcc_io phv m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI17 bias_g drvlo_h_n net171 vcc_io phv m=3 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 pbias drvlo_i_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI33 N0 vgnd_io vcc_io vcc_io phv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI32 net161 net161 N0 vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 net157 net157 net161 vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 net88 N0 vcc_io vcc_io phv m=8 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI43 net84 bias_g vcc_io vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI40 N0 drvlo_i_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
XICEpd_h pd_h / icecap
XICEen_fast_n<0> en_fast_n<0> / icecap
XICEpden_h_n pden_h_n / icecap
XICEint_nor<1> int_nor<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEen_fast_n<1> en_fast_n<1> / icecap
XICEint_slow int_slow / icecap
XICEint_nor<0> int_nor<0> / icecap
XI373<0> int_nor<1> / icecap
XI373<1> int_nor<0> / icecap
mmnin pd_h drvlo_h_n vgnd_io vgnd_io nhv m=5 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI56 int_slow pden_h_n vcc_io vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_slow pd_h drvlo_h_n int_slow vcc_io phv m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_slow int_slow pden_h_n vcc_io vcc_io phv m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<1> pd_h drvlo_h_n int_nor<1> net19<0> phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<0> pd_h drvlo_h_n int_nor<0> net19<1> phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io phv m=4 w=1.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io phv m=2 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I pden_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h:O
XICEpd_h pd_h / icecap
XICEen_fast_n<0> en_fast_n<0> / icecap
XICEpden_h_n pden_h_n / icecap
XICEint_nor<1> int_nor<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEen_fast_n<1> en_fast_n<1> / icecap
XICEint_slow int_slow / icecap
XICEint_nor<0> int_nor<0> / icecap
XI361<0> int_nor<1> / icecap
XI361<1> int_nor<0> / icecap
mmnin pd_h drvlo_h_n vgnd_io vgnd_io nhv m=5 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI56 int_slow pden_h_n vcc_io vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_slow pd_h drvlo_h_n int_slow vcc_io phv m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_slow int_slow pden_h_n vcc_io vcc_io phv m=1 w=1.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<1> pd_h drvlo_h_n int_nor<1> net19<0> phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<0> pd_h drvlo_h_n int_nor<0> net19<1> phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io phv m=4 w=1.00 l=1.00 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io phv m=2 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__tk_opti out spd spu
*.PININFO out:B spd:B spu:B
Xe2 spd out / sky130_fd_io__tk_em1o
Xe1 out spu / sky130_fd_io__tk_em1s
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos drvhi_h drvlo_h_n en_cmos_b 
+ nsw_en_int pd_h<3> pd_h<2> pden_h_n slow_h vcc_io vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I en_cmos_b:I nsw_en_int:I pden_h_n:I slow_h:I 
*.PININFO vcc_io:I vgnd_io:I pd_h<3>:O pd_h<2>:O
Xbias drvhi_h en_fast_h en_fast_h_n pbias_out pd_h<2> pden_h_n vcc_io vgnd_io 
+ / sky130_fd_io__gpio_ovtv2_pdpredrvr_pbias
Xnr3 drvlo_h_n net76 net76 pd_h<2> nsw_en_int vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr2
Xnr2 drvlo_h_n en_fast2_n<1> en_fast2_n<0> pd_h<3> nsw_en_int vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI76 net76 pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> vcc_io / sky130_fd_io__tk_opti
Xinv en_fast_h en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xnor slow_h en_cmos_b en_fast_h vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XICEnet30 net30 / icecap
XICEint<0> int<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XICEen_fast<0> en_fast<0> / icecap
XICEpu_h_n pu_h_n / icecap
XICEpuen_h puen_h / icecap
XI152<0> int<3> / icecap
XI152<1> int<2> / icecap
XI152<2> int<1> / icecap
XICEint_res int_res / icecap
XICEn<2> n<2> / icecap
XI150<0> en_fast<3> / icecap
XI150<1> en_fast<2> / icecap
XI150<2> en_fast<1> / icecap
XI151<0> int<3> / icecap
XI151<1> int<2> / icecap
XI151<2> int<1> / icecap
XI151<3> int<0> / icecap
XE1 net30 pu_h_n / sky130_fd_io__tk_em1s
rrespu1 int_res net30 mrp1 m=1 w=0.33 l=11
rrespu2 pu_h_n int_res mrp1 m=1 w=0.33 l=4
mmnin_fast<3> net30 drvhi_h int<3> net017<0> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<2> net30 drvhi_h int<2> net017<1> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<1> net30 drvhi_h int<1> net017<2> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<0> net30 drvhi_h int<0> net017<3> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_slow1 n<2> puen_h vgnd_io vgnd_io nhv m=1 w=0.75 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_slow pu_h_n drvhi_h n<2> vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<3> int<3> en_fast<3> vgnd_io net018<0> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<2> int<2> en_fast<2> vgnd_io net018<1> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<1> int<1> en_fast<1> vgnd_io net018<2> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen pu_h_n puen_h vcc_io vcc_io phv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin pu_h_n drvhi_h vcc_io vcc_io phv m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XI148<0> int<3> / icecap
XI148<1> int<2> / icecap
XI148<2> int<1> / icecap
XI148<3> int<0> / icecap
XI147<0> en_fast<3> / icecap
XI147<1> en_fast<2> / icecap
XI147<2> en_fast<1> / icecap
XICEn<2> n<2> / icecap
XICEpu_h_n pu_h_n / icecap
XICEnet30 net30 / icecap
XICEpuen_h puen_h / icecap
XICEint<0> int<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XI149<0> int<3> / icecap
XI149<1> int<2> / icecap
XI149<2> int<1> / icecap
XICEen_fast<0> en_fast<0> / icecap
XICEint_res int_res / icecap
XE1 net30 pu_h_n / sky130_fd_io__tk_em1s
rrespu1 int_res net30 mrp1 m=1 w=0.33 l=11
rrespu2 pu_h_n int_res mrp1 m=1 w=0.33 l=4
mmnin_fast<3> net30 drvhi_h int<3> net017<0> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<2> net30 drvhi_h int<2> net017<1> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<1> net30 drvhi_h int<1> net017<2> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<0> net30 drvhi_h int<0> net017<3> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_slow1 n<2> puen_h vgnd_io vgnd_io nhv m=1 w=0.75 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_slow pu_h_n drvhi_h n<2> vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<3> int<3> en_fast<3> vgnd_io net018<0> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<2> int<2> en_fast<2> vgnd_io net018<1> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<1> int<1> en_fast<1> vgnd_io net018<2> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<0> int<0> en_fast<0> vgnd_io vgnd_io nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen pu_h_n puen_h vcc_io vcc_io phv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin pu_h_n drvhi_h vcc_io vcc_io phv m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_pupredrvr_nbias drvhi_h en_h en_h_n nbias pu_h_n puen_h 
+ vcc_io vgnd_io
*.PININFO drvhi_h:I en_h:I en_h_n:I pu_h_n:I puen_h:I vcc_io:I vgnd_io:I 
*.PININFO nbias:O
XICEn<6> n<6> / icecap
XICEdrvhi_i_h_n drvhi_i_h_n / icecap
XICEen_h_n en_h_n / icecap
XICEbias_g bias_g / icecap
XICEn<2> n<2> / icecap
XICEn<8> n<8> / icecap
XICEdrvhi_h drvhi_h / icecap
XICEen_h en_h / icecap
XICEnet141 net141 / icecap
XICEvccio_2vtn vccio_2vtn / icecap
XICEnbias nbias / icecap
XICEnet153 net153 / icecap
XICEpu_h_n pu_h_n / icecap
XICEnet88 net88 / icecap
XICEn<7> n<7> / icecap
XICEn<1> n<1> / icecap
XICEnet90 net90 / icecap
XICEpuen_h puen_h / icecap
XI36 n<2> pu_h_n en_h / sky130_fd_io__tk_opto
XE5 nbias net88 / sky130_fd_io__tk_em1s
XE4 n<6> net153 / sky130_fd_io__tk_em1s
XE7 bias_g net90 / sky130_fd_io__tk_em1s
XE6 net141 nbias / sky130_fd_io__tk_em1s
XE1 n<2> n<1> / sky130_fd_io__tk_em1o
XE2 n<6> nbias / sky130_fd_io__tk_em1o
mI34 n<1> drvhi_h vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI32 n<1> n<2> n<2> vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 bias_g n<1> vcc_io vcc_io phv m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 bias_g drvhi_h vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 bias_g en_h vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 nbias bias_g vcc_io vcc_io phv m=4 w=1.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 drvhi_i_h_n drvhi_h vcc_io vcc_io phv m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI47 n<7> bias_g vcc_io vcc_io phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI49 net88 bias_g vcc_io vcc_io phv m=4 w=1.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI50 n<1> puen_h vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI56 vcc_io pu_h_n net90 vcc_io phv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 n<6> n<6> vgnd_io vgnd_io nhv m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 nbias nbias n<6> vgnd_io nhv m=4 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI28 bias_g drvhi_h n<3> vgnd_io nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI27 n<3> n<2> n<4> vgnd_io nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI26 n<4> en_h vgnd_io vgnd_io nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 drvhi_i_h_n drvhi_h vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 nbias en_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI53 vccio_2vtn drvhi_i_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 nbias drvhi_i_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI40 vccio_2vtn vcc_io vgnd_io vgnd_io nhv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI39 net153 vccio_2vtn vgnd_io vgnd_io nhv m=4 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI44 n<8> n<8> vccio_2vtn vgnd_io nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI41 n<7> n<7> n<8> vgnd_io nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI54 net141 bias_g vgnd_io vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> 
+ puen_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O
Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> 
+ pu_h_n<3> puen_h vcc_io vgnd_io / sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd3
Xnd2a drvhi_h net54 net54 net54 net54 pu_h_n<2> puen_h vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h / sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h / sky130_fd_io__tk_opto
Xinv en_fast_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io 
+ / sky130_fd_io__com_pupredrvr_nbias
Xnand puen_h slow_h_n en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_old drvhi_h drvlo_h_n en_cmos_b nsw_en 
+ pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> slow_h slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I en_cmos_b:I nsw_en:I pden_h_n<1>:I 
*.PININFO pden_h_n<0>:I puen_h<1>:I puen_h<0>:I slow_h:I slow_h_n:I vcc_io:I 
*.PININFO vgnd_io:I pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O
XICEpden_h_n<0> pden_h_n<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XICEpd_h<0> pd_h<0> / icecap
XICEpuen_h<1> puen_h<1> / icecap
XICEslow_h slow_h / icecap
XICEpd_h<1> pd_h<1> / icecap
XICEpu_h_n<0> pu_h_n<0> / icecap
XICEslow_h_n slow_h_n / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEen_cmos_b en_cmos_b / icecap
XICEnsw_en nsw_en / icecap
XI23<0> pd_h<3> / icecap
XI23<1> pd_h<2> / icecap
XI22<0> pu_h_n<3> / icecap
XI22<1> pu_h_n<2> / icecap
XICEpuen_h<0> puen_h<0> / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEpu_h_n<1> pu_h_n<1> / icecap
xI19 vgnd_io vcc_io condiode
Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io / 
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io / 
+ sky130_fd_io__com_pupredrvr_weak
XI151 drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io / 
+ sky130_fd_io__com_pdpredrvr_weak
Xpd_strong_slow drvlo_h_n pd_h<1> en_cmos_b vcc_io vgnd_io / 
+ sky130_fd_io__com_pdpredrvr_strong_slow
XI150 drvlo_h_n drvlo_h_n en_cmos_b nsw_en pd_h<3> pd_h<2> pden_h_n<1> slow_h 
+ vcc_io vgnd_io / sky130_fd_io__gpio_ovtv2_pdpredrvr_strong_cmos
Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io / 
+ sky130_fd_io__gpio_ovtv2_pupredrvr_strong
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix drvhi_h drvlo_h_n i2c_mode_h_n 
+ nghs_h oe_i_h_n pad pd_dis_h pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> 
+ pden_h_n<0> pghs_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
+ puen_h<0> pug_h slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> 
+ slow_h slow_h_n vcc_io vgnd_io vpb_drvr vssd
*.PININFO drvhi_h:I drvlo_h_n:I i2c_mode_h_n:I nghs_h:I oe_i_h_n:I pd_dis_h:I 
*.PININFO pden_h_n<1>:I pden_h_n<0>:I pghs_h:I puen_h<1>:I puen_h<0>:I pug_h:I 
*.PININFO slew_ctl_h<1>:I slew_ctl_h<0>:I slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I 
*.PININFO slow_h:I slow_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I vssd:I pd_h<3>:O 
*.PININFO pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O 
*.PININFO pu_h_n<0>:O pad:B
XICEpad pad / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEdrvhi_h drvhi_h / icecap
XI375<0> pu_h_n<3> / icecap
XI375<1> pu_h_n<2> / icecap
XI375<2> pu_h_n<1> / icecap
XI375<3> pu_h_n<0> / icecap
XICEvssd vssd / icecap
XI374<0> pd_h<3> / icecap
XI374<1> pd_h<2> / icecap
XI374<2> pd_h<1> / icecap
XI374<3> pd_h<0> / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEpug_h pug_h / icecap
XI376<0> puen_h<1> / icecap
XI376<1> puen_h<0> / icecap
XI377<0> pden_h_n<1> / icecap
XI377<1> pden_h_n<0> / icecap
XICEpd_dis_h pd_dis_h / icecap
XICEnsw_en nsw_en / icecap
XICEslow_h slow_h / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XI380<0> slew_ctl_h_n<1> / icecap
XI380<1> slew_ctl_h_n<0> / icecap
XICEslow_h_n slow_h_n / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEpghs_h pghs_h / icecap
XI379<0> pd_h<3> / icecap
XI379<1> pd_h<2> / icecap
XI378<0> slew_ctl_h<1> / icecap
XI378<1> slew_ctl_h<0> / icecap
XICEen_cmos_b en_cmos_b / icecap
XICEnghs_h nghs_h / icecap
XI192 drvlo_h_n en_cmos_b i2c_mode_h_n nghs_h nsw_en oe_i_h_n pad pd_dis_h 
+ pd_h<3> pd_h<2> pden_h_n<1> pghs_h pug_h slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow_h_n vcc_io vgnd_io vpb_drvr vssd / 
+ sky130_fd_io__gpio_ovtv2_obpredrvr_new_leak_fix
XI191 drvhi_h drvlo_h_n en_cmos_b nsw_en pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
+ puen_h<0> slow_h slow_h_n vcc_io vgnd_io / sky130_fd_io__gpio_ovtv2_obpredrvr_old
.ENDS
.SUBCKT sky130_fd_io__gpio_dat_ls hld_h_n in out_h out_h_n rst_h set_h vcc_io vgnd 
+ vpwr_ka
*.PININFO hld_h_n:I in:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr_ka:I out_h:O 
*.PININFO out_h_n:O
XICEnet107 net107 / icecap
XICEhld_h_n hld_h_n / icecap
XICEset_h set_h / icecap
XICEnet79 net79 / icecap
XICEnet83 net83 / icecap
XICEout_h out_h / icecap
XICErst_h rst_h / icecap
XICEnet103 net103 / icecap
XICEin in / icecap
XICEout_h_n out_h_n / icecap
XICEin_i in_i / icecap
XICEfbk fbk / icecap
XICEin_i_n in_i_n / icecap
XICEfbk_n fbk_n / icecap
mI3 fbk fbk_n vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI4 fbk_n fbk vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 fbk hld_h_n net79 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 fbk_n hld_h_n net83 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 net107 in_i_n vgnd vgnd nlowvt m=8 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 net103 in_i vgnd vgnd nlowvt m=8 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out_h fbk_n vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h_n fbk vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmnset fbk_n set_h vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmnrst fbk rst_h vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI34 in_i_n in vgnd vgnd nshort m=2 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI35 in_i in_i_n vgnd vgnd nshort m=2 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 net83 vpwr_ka net103 vgnd nhvnative m=8 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 net79 vpwr_ka net107 vgnd nhvnative m=8 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk_n fbk vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk fbk_n vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI33 in_i in_i_n vpwr_ka vpwr_ka phighvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI11 out_h fbk_n vcc_io vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 out_h_n fbk vcc_io vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI32 in_i_n in vpwr_ka vpwr_ka phighvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_cclat_hvnor3 in0 in1 in2 out vcc_io vgnd vnb
*.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
XICEin0 in0 / icecap
XICEin2 in2 / icecap
XICEout out / icecap
XICEn<1> n<1> / icecap
XICEin1 in1 / icecap
XICEn<0> n<0> / icecap
mmp0 n<0> in0 vcc_io vcc_io phv m=8 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmp2 out in2 n<1> vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmp1 n<1> in1 n<0> vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmn0 out in0 vgnd vnb nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmn2 out in2 vgnd vnb nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmn1 out in1 vgnd vnb nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_cclat_hvnand3 in0 in1 in2 out vcc_io vgnd vnb
*.PININFO in0:I in1:I in2:I vcc_io:I vgnd:I vnb:I out:O
XICEin0 in0 / icecap
XICEn0 n0 / icecap
XICEin2 in2 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
XICEn1 n1 / icecap
mmp0 out in0 vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmp2 out in2 vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmp1 out in1 vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmn2 out in2 n1 vnb nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mmn0 n0 in0 vgnd vnb nhv m=4 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmn1 n1 in1 n0 vnb nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_cclat_inv_in in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XICEin in / icecap
XICEout out / icecap
mmp1 out in vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmn1 out in vgnd vnb nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_cclat_inv_out in out vcc_io vgnd vnb
*.PININFO in:I vcc_io:I vgnd:I vnb:I out:O
XICEin in / icecap
XICEout out / icecap
mI1 out in vcc_io vcc_io phv m=6 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 out in vgnd vnb nhv m=6 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_cclat_i2c_fix drvhi_h drvlo_h_n oe_h pd_dis_h pu_dis_h 
+ vcc_io vgnd
*.PININFO oe_h:I pd_dis_h:I pu_dis_h:I vcc_io:I vgnd:I drvhi_h:O drvlo_h_n:O
XICEpd_dis_h pd_dis_h / icecap
XICEoe_h oe_h / icecap
XICEdrvhi_h drvhi_h / icecap
XICEn0 n0 / icecap
XICEn1 n1 / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEpu_dis_h pu_dis_h / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEpu_dis_h_n pu_dis_h_n / icecap
Xnor3 oe_i_h_n drvhi_h pd_dis_h n1 vcc_io vgnd vgnd / sky130_fd_io__com_cclat_hvnor3
Xnand3 oe_h drvlo_h_n pu_dis_h_n n0 vcc_io vgnd vgnd / 
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe2 oe_h oe_i_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_pudis pu_dis_h pu_dis_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_out n1 drvlo_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
Xinv_out_1 n0 drvhi_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
.ENDS
.SUBCKT sky130_fd_io__hvsbt_inv_x1 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEin in / icecap
XICEout out / icecap
mI1 out in vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 out in vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_dat_ls_i2c_fix hld_h_n in out_h_n set_h set_h_n vcc_io 
+ vgnd vpwr_ka
*.PININFO hld_h_n:I in:I set_h:I set_h_n:I vcc_io:I vgnd:I vpwr_ka:I out_h_n:O
XICEnet76 net76 / icecap
XICEin_i_n in_i_n / icecap
XICEset_h set_h / icecap
XICEin in / icecap
XICEnet96 net96 / icecap
XICEout_h_n out_h_n / icecap
XICEhld_h_n hld_h_n / icecap
XICEnet100 net100 / icecap
XICEfbk_n fbk_n / icecap
XICEfbk fbk / icecap
XICEin_i in_i / icecap
XICEnet80 net80 / icecap
XICEset_h_n set_h_n / icecap
mI3 fbk fbk_n vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI4 fbk_n fbk vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 fbk hld_h_n net76 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 fbk_n hld_h_n net80 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 net100 in_i_n vgnd vgnd nlowvt m=8 w=1.00 l=0.15 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 net96 in_i vgnd vgnd nlowvt m=8 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h_n fbk vgnd vgnd nhv m=2 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmnset fbk_n set_h vgnd vgnd nhv m=4 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI34 in_i_n in vgnd vgnd nshort m=2 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI35 in_i in_i_n vgnd vgnd nshort m=2 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 net80 vpwr_ka net96 vgnd nhvnative m=8 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 net76 vpwr_ka net100 vgnd nhvnative m=8 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk_n fbk vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk fbk_n vcc_io vcc_io phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI33 in_i in_i_n vpwr_ka vpwr_ka phighvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 out_h_n fbk vcc_io vcc_io phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 fbk set_h_n vcc_io vcc_io phv m=3 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI32 in_i_n in vpwr_ka vpwr_ka phighvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix drvhi_h drvlo_h_n hld_h_n 
+ hld_i_ovr_h od_i_h_n oe_h oe_n out pd_dis_h vcc_io vgnd vpwr_ka
*.PININFO hld_h_n:I hld_i_ovr_h:I od_i_h_n:I oe_n:I out:I vcc_io:I vgnd:I 
*.PININFO vpwr_ka:I drvhi_h:O drvlo_h_n:O oe_h:O pd_dis_h:O
XICEhld_h_n hld_h_n / icecap
XICEnet56 net56 / icecap
XICEoe_h oe_h / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEout out / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XICEpu_dis_h pu_dis_h / icecap
XICEpd_dis_h pd_dis_h / icecap
XICEdrvhi_h drvhi_h / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEnet60 net60 / icecap
XICEoe_n oe_n / icecap
Xdat_ls hld_i_ovr_h out pd_dis_h pu_dis_h vgnd net60 vcc_io vgnd vpwr_ka / 
+ sky130_fd_io__gpio_dat_ls
Xcclat drvhi_h drvlo_h_n oe_h pd_dis_h pu_dis_h vcc_io vgnd / 
+ sky130_fd_io__com_cclat_i2c_fix
XI36 od_i_h_n net60 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI37 od_i_h_n net56 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xoe_ls hld_i_ovr_h oe_n oe_h net56 od_i_h_n vcc_io vgnd vpwr_ka / 
+ sky130_fd_io__gpio_dat_ls_i2c_fix
.ENDS
.SUBCKT sky130_fd_io__hvsbt_nor in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
mI3 net16 in0 vpwr vpwr phv m=1 w=1.00 l=0.60 mult=2 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out in1 net16 vpwr phv m=1 w=1.00 l=0.60 mult=2 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out in1 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__hvsbt_xor in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEin0 in0 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
XICEnet54 net54 / icecap
XICEnet29 net29 / icecap
XICEnet70 net70 / icecap
XICEnet45 net45 / icecap
mI3 net29 in0 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out net54 net45 vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI17 net70 in1 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 net54 in0 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 net45 in1 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out net70 net29 vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net58 vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 net70 in1 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out net70 net62 vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 net62 net54 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 net58 in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 net54 in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__hvsbt_inv_x2 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vgnd nhv m=2 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in vpwr vpwr phv m=4 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_ctl_ls hld_h_n in out_h out_h_n rst_h set_h vcc_io vgnd 
+ vpwr
*.PININFO hld_h_n:I in:I rst_h:I set_h:I vcc_io:I vgnd:I vpwr:I out_h:O 
*.PININFO out_h_n:O
XICEout_h_n out_h_n / icecap
XICEset_h set_h / icecap
XICEfbk_n fbk_n / icecap
XICErst_h rst_h / icecap
XICEnet122 net122 / icecap
XICEnet130 net130 / icecap
XICEnet94 net94 / icecap
XICEhld_h_n hld_h_n / icecap
XICEfbk fbk / icecap
XICEout_h out_h / icecap
XICEnet98 net98 / icecap
XICEin in / icecap
XICEin_i in_i / icecap
XICEin_i_n in_i_n / icecap
mI14 out_h_n fbk vcc_io vcc_io phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI34 in_i in_i_n vpwr vpwr phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 in_i_n in vpwr vpwr phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI11 out_h fbk_n vcc_io vcc_io phv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk fbk_n vcc_io vcc_io phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk_n fbk vcc_io vcc_io phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h_n fbk vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmnset fbk_n set_h vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI32 in_i in_i_n vgnd vgnd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out_h fbk_n vgnd vgnd nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI58 net130 vpwr net94 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnrst fbk rst_h vgnd vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI59 net122 vpwr net98 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 fbk_n hld_h_n net122 vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI27 in_i_n in vgnd vgnd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 fbk hld_h_n net130 vgnd nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI4 fbk_n fbk vgnd vgnd nhv m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI3 fbk fbk_n vgnd vgnd nhv m=1 w=0.75 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 net98 in_i vgnd vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 net94 in_i_n vgnd vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_octl_i2c_fix dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> 
+ dm_h_n<1> dm_h_n<0> hld_i_h_n od_i_h_n pden_h_n<2> pden_h_n<1> pden_h_n<0> 
+ puen_0_h puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd 
+ vpwr vreg_en_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I od_i_h_n:I slow:I vcc_io:I vgnd:I vpwr:I vreg_en_h_n:I 
*.PININFO pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O puen_2or1_h:O 
*.PININFO puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O
XI211 n<8> dm_h_n<1> puen_0_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI366 dm_h<1> dm_h<0> net87 vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI210 dm_h<2> dm_h<0> n<8> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI200 dm_h<2> dm_h<1> n<10> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI185 dm_h_n<0> n<4> net207 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI187 dm_h<1> dm_h<0> n<3> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI203 n<10> dm_h<0> n<1> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI204 n<9> dm_h_n<0> n<0> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> puen_2or1_h vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI365 net87 dm_h<2> pden_h_n<2> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n puen_h<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n puen_h<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 pden_h_n<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 pden_h_n<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI377 puen_0_h puen_h0_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI374 net207 pden_h1 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI381 od_i_h_n n9 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xls_slow hld_i_h_n slow slow_h slow_h_n n9 vgnd vcc_io vgnd vpwr / 
+ sky130_fd_io__com_ctl_ls
XICEn<0> n<0> / icecap
XICEn<4> n<4> / icecap
XICEpuen_2or1_h puen_2or1_h / icecap
XICEdm_h<2> dm_h<2> / icecap
XICEpden_h1 pden_h1 / icecap
XICEn<10> n<10> / icecap
XICEslow_h_n slow_h_n / icecap
XICEdm_h_n<1> dm_h_n<1> / icecap
XICEpden_h0 pden_h0 / icecap
XICEdm_h<1> dm_h<1> / icecap
XICEn<8> n<8> / icecap
XICEslow slow / icecap
XICEdm_h<0> dm_h<0> / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEn<9> n<9> / icecap
XICEpuen_0_h puen_0_h / icecap
XICEpuen_h1_n puen_h1_n / icecap
XICEpuen_h<0> puen_h<0> / icecap
XICEpuen_h0_n puen_h0_n / icecap
XICEdm_h_n<2> dm_h_n<2> / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEnet177 net207 / icecap
XICEn<3> n<3> / icecap
XICEvreg_en_h_n vreg_en_h_n / icecap
XICEdm_h_n<0> dm_h_n<0> / icecap
XICEpden_h_n<0> pden_h_n<0> / icecap
XICEn<1> n<1> / icecap
XICEn<2> n<2> / icecap
XICEpuen_h<1> puen_h<1> / icecap
XICEslow_h slow_h / icecap
XICEn<5> n<5> / icecap
XICEnet198 net87 / icecap
.ENDS
.SUBCKT sky130_fd_io__sio_hvsbt_inv_x2 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEin in / icecap
XICEout out / icecap
mI1 out in vpwr vpb phv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI2 out in vgnd vnb nhv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h nghs_h od_i_h_n 
+ oe_hs_h oe_n out pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow slow_h_n vccd vddio vpb_drvr vpwr_ka 
+ vssd vssio
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I nghs_h:I od_i_h_n:I oe_n:I out:I pghs_h:I 
*.PININFO pug_h:I slew_ctl_h<1>:I slew_ctl_h<0>:I slew_ctl_h_n<1>:I 
*.PININFO slew_ctl_h_n<0>:I slow:I vccd:I vddio:I vpb_drvr:I vpwr_ka:I vssd:I 
*.PININFO vssio:I drvhi_h:O oe_hs_h:O pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O 
*.PININFO pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O slow_h_n:O pad:B
XI425<0> pd_h<3> / icecap
XI425<1> pd_h<2> / icecap
XI425<2> pd_h<1> / icecap
XI425<3> pd_h<0> / icecap
XICEpden_h_n<2> pden_h_n<2> / icecap
XICEoe_h oe_h / icecap
XICEvpb_drvr vpb_drvr / icecap
XICEod_i_h_n od_i_h_n / icecap
XI431<0> pden_h_n<1> / icecap
XI431<1> pden_h_n<0> / icecap
XICEoe_hs_i_h_n oe_hs_i_h_n / icecap
XICEoe_hs_i_h oe_hs_i_h / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XICEn<1> n<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEslow_h_n slow_h_n / icecap
XICEnghs_h nghs_h / icecap
XI422<0> pu_h_n<3> / icecap
XI422<1> pu_h_n<2> / icecap
XI422<2> pu_h_n<1> / icecap
XI422<3> pu_h_n<0> / icecap
XI424<0> dm_h<2> / icecap
XI424<1> dm_h<1> / icecap
XI424<2> dm_h<0> / icecap
XI430<0> puen_h<1> / icecap
XI430<1> puen_h<0> / icecap
XI423<0> pd_h<3> / icecap
XI423<1> pd_h<2> / icecap
XI423<2> pd_h<1> / icecap
XI423<3> pd_h<0> / icecap
XICEnet85 net85 / icecap
XICEpad pad / icecap
XI429<0> pu_h_n<3> / icecap
XI429<1> pu_h_n<2> / icecap
XI429<2> pu_h_n<1> / icecap
XI429<3> pu_h_n<0> / icecap
XI432<0> slew_ctl_h_n<1> / icecap
XI432<1> slew_ctl_h_n<0> / icecap
XICEdrvhi_h drvhi_h / icecap
XI426<0> dm_h_n<2> / icecap
XI426<1> dm_h_n<1> / icecap
XI426<2> dm_h_n<0> / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEslow_h slow_h / icecap
XICEoe_n oe_n / icecap
XICEpug_h pug_h / icecap
XICEnet86 net86 / icecap
XICEslow slow / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEoe_hs_h oe_hs_h / icecap
XICEpghs_h pghs_h / icecap
XICEnet72 net72 / icecap
XI427<0> slew_ctl_h<1> / icecap
XI427<1> slew_ctl_h<0> / icecap
XICEout out / icecap
XI428<0> pden_h_n<2> / icecap
XI428<1> pden_h_n<1> / icecap
XI428<2> pden_h_n<0> / icecap
Xpredrvr drvhi_h drvlo_h_n pden_h_n<2> nghs_h oe_i_h_n pad net72 pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pghs_h pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> pug_h slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow_h slow_h_n vddio vssio vpb_drvr vssd / 
+ sky130_fd_io__gpio_ovtv2_obpredrvr_leak_fix
Xdatoe drvhi_h drvlo_h_n hld_i_h_n hld_i_ovr_h od_i_h_n oe_h oe_n out net72 
+ vddio vssd vpwr_ka / sky130_fd_io__gpio_ovtv2_opath_datoe_i2c_fix
Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_i_h_n 
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> net86 net85 puen_h<1> puen_h<0> slow 
+ slow_h slow_h_n vddio vssd vccd vddio / sky130_fd_io__gpio_ovtv2_octl_i2c_fix
XI354 oe_hs_i_h oe_hs_i_h_n vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x1
XI353 oe_h oe_i_h_n vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x2
XI355 oe_hs_i_h_n oe_hs_h vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_inv_x2
XI351 net86 net85 n<1> vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_nor
XI352 n<1> oe_i_h_n oe_hs_i_h vssd vssd vddio vddio / sky130_fd_io__sio_hvsbt_nor
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n hld_i_ovr_h nga_pad_vpmp_h 
+ ngb_pad_vpmp_h od_i_h_n oe_n out pad pd_csd_h pghs_h pu_csd_h pug_h<6> 
+ pug_h<5> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> slow 
+ tie_hi_esd tie_lo_esd vccd vddio vddio_amx vpb_drvr vpwr_ka vssa vssd vssio 
+ vssio_amx
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I nga_pad_vpmp_h:I ngb_pad_vpmp_h:I 
*.PININFO od_i_h_n:I oe_n:I out:I pd_csd_h:I pu_csd_h:I slew_ctl_h<1>:I 
*.PININFO slew_ctl_h<0>:I slew_ctl_h_n<1>:I slew_ctl_h_n<0>:I slow:I vccd:I 
*.PININFO vddio:I vpwr_ka:I vssa:I vssd:I vssio:I vssio_amx:I pad:O pghs_h:O 
*.PININFO tie_hi_esd:O tie_lo_esd:O pug_h<6>:B pug_h<5>:B vddio_amx:B 
*.PININFO vpb_drvr:B
Xodrvr tie_lo_esd nga_pad_vpmp_h ngb_pad_vpmp_h nghs_h od_i_h_n oe_hs_h pad 
+ pd_csd_h pd_h<3> pd_h<2> pd_h<1> pd_h<0> pghs_h pu_csd_h pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> pug_h<7> pug_h<6> pug_h<5> tie_hi_esd tie_lo_esd vddio 
+ vddio_amx vpb_drvr vssa vssd vssio vssio_amx / 
+ sky130_fd_io__gpio_ovtv2_odrvr_i2c_fix_leak_fix
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n 
+ hld_i_ovr_h nghs_h od_i_h_n oe_hs_h oe_n out pad pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pghs_h pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> pug_h<7> 
+ slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> slow slow_h_n 
+ vccd vddio vpb_drvr vpwr_ka vssd vssio / 
+ sky130_fd_io__gpio_ovtv2_octl_dat_i2c_fix_leak_fix
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix in in_b out_h rst_h rst_h_n vgnd 
+ vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O
XICEnet70 net70 / icecap
XICEnet75 net75 / icecap
XICErst_h_n rst_h_n / icecap
XICEfbk_n fbk_n / icecap
XICEin in / icecap
XICEnet71 net71 / icecap
XICEin_b in_b / icecap
XICEout_h out_h / icecap
XICErst_h rst_h / icecap
XICEfbk fbk / icecap
mI14 fbk_n rst_h_n vpwr_hv vpwr_hv phv m=2 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI11 out_h fbk_n vpwr_hv vpwr_hv phv m=2 w=0.75 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk_n fbk vpwr_hv vpwr_hv phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk fbk_n vpwr_hv vpwr_hv phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 net70 rst_h_n vgnd vgnd nhv m=4 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out_h fbk_n vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI58 fbk vpwr_lv net71 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnrst fbk rst_h vgnd vgnd nhv m=3 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI59 fbk_n vpwr_lv net75 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 net75 in net70 vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 net71 in_b net70 vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ls_inv_x1 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in vpwr vpwr phv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_lshv2hv in in_b out_h out_h_n rst_h rst_h_n 
+ vgnd vpwr_hv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I out_h:O out_h_n:O
XICEnet64 net64 / icecap
XICEin in / icecap
XICErst_h_n rst_h_n / icecap
XICEout_h out_h / icecap
XICEfbk fbk / icecap
XICEin_b in_b / icecap
XICEfbk_n fbk_n / icecap
XICErst_h rst_h / icecap
XICEout_h_n out_h_n / icecap
mI14 out_h_n fbk vpwr_hv vpwr_hv phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI11 out_h fbk_n vpwr_hv vpwr_hv phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk fbk_n vpwr_hv vpwr_hv phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk_n fbk vpwr_hv vpwr_hv phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI64 net64 rst_h_n vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h_n fbk vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out_h fbk_n vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmnrst fbk rst_h vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 fbk_n in net64 vgnd nhv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 fbk in_b net64 vgnd nhv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_inv_1 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI27 out in vgnd vgnd nshort m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 out in vpwr vpwr phighvt m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ls_i2c_fix amux_en_vdda_h amux_en_vdda_h_n 
+ amux_en_vddio_h amux_en_vswitch_h amux_en_vswitch_h_n analog_en 
+ enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h_n vccd vdda vddio_q 
+ vssa vssd vswitch
*.PININFO analog_en:I enable_vdda_h:I enable_vswitch_h:I hld_i_h_n:I vccd:I 
*.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I amux_en_vdda_h:O 
*.PININFO amux_en_vdda_h_n:O amux_en_vddio_h:O amux_en_vswitch_h:O 
*.PININFO amux_en_vswitch_h_n:O enable_vdda_h_n:O
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEanalog_en analog_en / icecap
XICEnet028 net028 / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEnet83 net83 / icecap
XICEana_en_i_n ana_en_i_n / icecap
XICEnet082 net082 / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEana_en_i ana_en_i / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
Xpd_vddio_ls ana_en_i ana_en_i_n amux_en_vddio_h net082 hld_i_h_n vssd vddio_q 
+ vccd / sky130_fd_io__gpiov2_amux_ctl_ls_i2c_fix
XI32 enable_vdda_h enable_vdda_h_n vssa vdda / sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls amux_en_vddio_h net028 amux_en_vswitch_h amux_en_vswitch_h_n 
+ net83 enable_vswitch_h vssa vswitch / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls amux_en_vddio_h net028 amux_en_vdda_h amux_en_vdda_h_n 
+ enable_vdda_h_n enable_vdda_h vssa vdda / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 analog_en ana_en_i_n vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 enable_vswitch_h net83 vssa vswitch / sky130_fd_io__hvsbt_inv_x1
XI36 amux_en_vddio_h net028 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI35 hld_i_h_n net082 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2 in in_b out_h out_h_n 
+ rst2_h rst2_h_n rst_h rst_h_n vgnd vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst2_h:I rst2_h_n:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I 
*.PININFO vpwr_lv:I out_h:O out_h_n:O
XICEin_b in_b / icecap
XICEnet76 net76 / icecap
XICEout_h out_h / icecap
XICEnet56 net56 / icecap
XICErst_h rst_h / icecap
XICErst2_h_n rst2_h_n / icecap
XICErst_h_n rst_h_n / icecap
XICEnet52 net52 / icecap
XICEin in / icecap
XICEout_h_n out_h_n / icecap
XICErst2_h rst2_h / icecap
XICEnet72 net72 / icecap
mI11 out_h_n out_h vpwr_hv vpwr_hv phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI9 out_h out_h_n vpwr_hv vpwr_hv phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 out_h_n rst2_h_n vpwr_hv vpwr_hv phv m=3 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI28 out_h_n rst_h_n vpwr_hv vpwr_hv phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 net56 vpwr_lv net76 vgnd nhvnative m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 net52 vpwr_lv net72 vgnd nhvnative m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI17 out_h rst_h vgnd vgnd nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net76 in vgnd vgnd nlowvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 net72 in_b vgnd vgnd nlowvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 out_h rst2_h vgnd vgnd nhv m=3 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 out_h rst_h_n net52 vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 out_h_n rst_h_n net56 vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_buf A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XICEA A / icecap
XICEY Y / icecap
XICEint int / icecap
mI75 int A vssa vssa nhv m=4 w=0.42 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 Y int vssa vssa nhv m=3 w=0.42 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI74 int A vda vda phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI5 Y int vda vda phv m=5 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3 in in_b out_h out_h_n rst2_h_n 
+ rst_h_n vgnd vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst2_h_n:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O 
*.PININFO out_h_n:O
XICEout_h_n out_h_n / icecap
XICErst2_h_n rst2_h_n / icecap
XICErst_h_n rst_h_n / icecap
XICEnet074 net074 / icecap
XICEout_h out_h / icecap
XICEnet75 net75 / icecap
XICEnet51 net51 / icecap
XICEnet086 net086 / icecap
XICEin in / icecap
XICEnet55 net55 / icecap
XICEin_b in_b / icecap
XICEnet79 net79 / icecap
XI34 rst_h_n net086 vgnd vpwr_hv / sky130_fd_io__hvsbt_inv_x1
XI33 rst2_h_n net074 vgnd vpwr_hv / sky130_fd_io__hvsbt_inv_x1
mI11 out_h_n out_h vpwr_hv vpwr_hv phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI9 out_h out_h_n vpwr_hv vpwr_hv phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 out_h_n rst2_h_n vpwr_hv vpwr_hv phv m=3 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI28 out_h_n rst_h_n vpwr_hv vpwr_hv phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 net55 vpwr_lv net79 vgnd nhvnative m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 net51 vpwr_lv net75 vgnd nhvnative m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI17 out_h net086 vgnd vgnd nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net79 in vgnd vgnd nlowvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 net75 in_b vgnd vgnd nlowvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 out_h net074 vgnd vgnd nhv m=3 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 out_h rst_h_n net51 vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 out_h_n rst_h_n net55 vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_lshv2hv in in_b out_h_n rst_h rst_h_n vgnd 
+ vpwr_hv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I out_h_n:O
XICErst_h rst_h / icecap
XICEout_h_n out_h_n / icecap
XICEin in / icecap
XICEfbk fbk / icecap
XICEin_b in_b / icecap
XICEnet52 net52 / icecap
XICEfbk_n fbk_n / icecap
XICErst_h_n rst_h_n / icecap
mI14 out_h_n fbk vpwr_hv vpwr_hv phv m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk fbk_n vpwr_hv vpwr_hv phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk_n fbk vpwr_hv vpwr_hv phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI64 net52 rst_h_n vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h_n fbk vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mmnrst fbk rst_h vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 fbk_n in net52 vgnd nhv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 fbk in_b net52 vgnd nhv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amx_inv4 A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XICEA A / icecap
XICEY Y / icecap
mI75 Y A vssa vssa nhv m=2 w=0.42 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI74 Y A vda vda phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amx_pdcsd_inv A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XICEA A / icecap
XICEY Y / icecap
mI414 Y A vssa vssa nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI519 Y vssa vssa vssa nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI517 Y A vda vda phv m=1 w=0.75 l=2.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI429 Y A vda vda phv m=1 w=0.75 l=2.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__amx_inv1 A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XICEA A / icecap
XICEY Y / icecap
mI92 Y A vssa vssa nhv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI54 Y A vda vda phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_ls in in_b out_h out_h_n rst_h rst_h_n vgnd 
+ vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O 
*.PININFO out_h_n:O
XICEin_b in_b / icecap
XICErst_h_n rst_h_n / icecap
XICEnet42 net42 / icecap
XICErst_h rst_h / icecap
XICEnet38 net38 / icecap
XICEin in / icecap
XICEnet54 net54 / icecap
XICEout_h_n out_h_n / icecap
XICEout_h out_h / icecap
XICEnet58 net58 / icecap
mI11 out_h_n out_h vpwr_hv vpwr_hv phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI9 out_h out_h_n vpwr_hv vpwr_hv phv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 net42 vpwr_lv net58 vgnd nhvnative m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 net38 vpwr_lv net54 vgnd nhvnative m=2 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI17 out_h rst_h vgnd vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net58 in vgnd vgnd nlowvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 net54 in_b vgnd vgnd nlowvt m=2 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 out_h rst_h_n net38 vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 out_h_n rst_h_n net42 vgnd nhv m=2 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr_i2c_fix amux_en_vdda_h amux_en_vdda_h_n 
+ amux_en_vddio_h amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on 
+ amuxbusa_on_n amuxbusb_on amuxbusb_on_n hld_i_h_n nga_amx_vswitch_h 
+ nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h 
+ ngb_pad_vswitch_h_n nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd 
+ nmidb_vccd_n pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n 
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
+ pu_csd_vddioq_h_n pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO amux_en_vdda_h:I amux_en_vdda_h_n:I amux_en_vddio_h:I 
*.PININFO amux_en_vswitch_h:I amux_en_vswitch_h_n:I amuxbusa_on:I 
*.PININFO amuxbusa_on_n:I amuxbusb_on:I amuxbusb_on_n:I hld_i_h_n:I 
*.PININFO nmida_on_n:I nmidb_on_n:I pd_on:I pd_on_n:I pu_on:I pu_on_n:I vccd:I 
*.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I nga_amx_vswitch_h:O 
*.PININFO nga_pad_vswitch_h:O nga_pad_vswitch_h_n:O ngb_amx_vswitch_h:O 
*.PININFO ngb_pad_vswitch_h:O ngb_pad_vswitch_h_n:O nmida_vccd:O 
*.PININFO nmida_vccd_n:O nmidb_vccd:O nmidb_vccd_n:O pd_csd_vswitch_h:O 
*.PININFO pd_csd_vswitch_h_n:O pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O 
*.PININFO pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
XICEhld_i_h_n hld_i_h_n / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEpu_on_n pu_on_n / icecap
XICEnet295 net295 / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEnet278 net278 / icecap
XICEnet160 net160 / icecap
XICEnet154 net154 / icecap
XICEhld_i_h hld_i_h / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEnet149 net149 / icecap
XICEpd_on pd_on / icecap
XICEnet284 net284 / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEnet296 net296 / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEpd_on_n pd_on_n / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
XICEnet167 net167 / icecap
XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
XICEnet293 net293 / icecap
XICEnet168 net168 / icecap
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
XICEnet287 net287 / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEpu_on pu_on / icecap
XICEnet144 net144 / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
Xpga_pad_ls amuxbusa_on amuxbusa_on_n net154 net160 hld_i_h hld_i_h_n 
+ amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q vccd / 
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
Xpgb_pad_ls amuxbusb_on amuxbusb_on_n net144 net149 hld_i_h hld_i_h_n 
+ amux_en_vddio_h_n amux_en_vddio_h vssd vddio_q vccd / 
+ sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3_ver2
XI38 net168 pu_csd_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_pucsd_buf
Xpu_csd_ls pu_on pu_on_n net167 net168 hld_i_h_n amux_en_vddio_h vssd vddio_q 
+ vccd / sky130_fd_io__gpiov2_amux_drvr_ls_i2c_fix3
XI111 hld_i_h_n hld_i_h vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI110 amux_en_vddio_h amux_en_vddio_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI93 nmida_vccd nmida_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
XI105 nmidb_vccd nmidb_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
Xpga_amx_ls net154 net160 pga_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h 
+ vssa vdda / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net144 net149 pgb_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h vssa vdda 
+ / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net295 nga_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI42 net154 pga_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI47 net295 nga_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI62 net144 pgb_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI63 net284 ngb_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI64 net284 ngb_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI53 nmidb_on_n nmidb_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
XI89 nmida_on_n nmida_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv net293 pd_csd_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_pdcsd_inv
XI87 nga_pad_vswitch_h nga_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI85 ngb_pad_vswitch_h ngb_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI90 pd_csd_vswitch_h pd_csd_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
mI76 ngb_amx_vswitch_h amux_en_vdda_h_n vssa vssa nhv m=1 w=1.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI77 ngb_pad_vswitch_h amux_en_vddio_h_n vssa vssa nhv m=1 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI75 nga_amx_vswitch_h amux_en_vdda_h_n vssa vssa nhv m=1 w=1.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI78 nga_pad_vswitch_h amux_en_vddio_h_n vssa vssa nhv m=1 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI104 pd_csd_vswitch_h amux_en_vddio_h_n vssa vssa nhv m=1 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xnga_ls amuxbusa_on amuxbusa_on_n net296 net295 amux_en_vswitch_h_n 
+ amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls pd_on pd_on_n net287 net293 amux_en_vswitch_h_n amux_en_vswitch_h 
+ vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls amuxbusb_on amuxbusb_on_n net278 net284 amux_en_vswitch_h_n 
+ amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
.ENDS
.SUBCKT sky130_fd_io__nor2_1 A B Y vgnd vnb vpb vpwr
*.PININFO A:I B:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XICEY Y / icecap
XICEA A / icecap
XICEB B / icecap
mMP0 vpwr A sndPA vpb phighvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMP1 sndPA B Y vpb phighvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMN0 Y A vgnd vnb nshort m=1 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMN1 Y B vgnd vnb nshort m=1 w=740e-3 l=150e-3 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nand2_1 A B Y vgnd vnb vpb vpwr
*.PININFO A:I B:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XICEA A / icecap
XICEB B / icecap
XICEY Y / icecap
mMP0 Y A vpwr vpb phighvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMP1 Y B vpwr vpb phighvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMN0 Y A sndA vnb nshort m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMN1 sndA B vgnd vnb nshort m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_nand5 in0 in1 in2 in3 in4 out vgnd vpwr
*.PININFO in0:I in1:I in2:I in3:I in4:I vgnd:I vpwr:I out:O
XICEin4 in4 / icecap
XICEin3 in3 / icecap
XICEin1 in1 / icecap
XICEout out / icecap
XICEin2 in2 / icecap
XICEin0 in0 / icecap
XICEout_n out_n / icecap
mI3 out in0 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 out out_n vpwr vpwr phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 out_n out vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net51 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 net63 in4 net59 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net59 in0 vgnd vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 net55 in3 net63 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 net51 in2 net55 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI22 out_n out vgnd vgnd nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI23 vgnd out_n vgnd vgnd nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_nand4 in0 in1 in2 in3 out vgnd vpwr
*.PININFO in0:I in1:I in2:I in3:I vgnd:I vpwr:I out:O
XICEout_n out_n / icecap
XICEin1 in1 / icecap
XICEout out / icecap
XICEin3 in3 / icecap
XICEin0 in0 / icecap
XICEin2 in2 / icecap
mI3 out in0 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 out_n out vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 out out_n vpwr vpwr phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net50 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net58 in0 vgnd vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 net54 in3 net58 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 net50 in2 net54 vgnd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 out_n out vgnd vgnd nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI21 vgnd out_n vgnd vgnd nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__xor2_1 A B X vgnd vpwr
*.PININFO A:I B:I vgnd:I vpwr:I X:O
XICEpmid pmid / icecap
XICEinor inor / icecap
XICEX X / icecap
XICEA A / icecap
XICEB B / icecap
mMNnor0 inor A vgnd vgnd nshort m=1 w=840e-3 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMNnor1 inor B vgnd vgnd nshort m=1 w=840e-3 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMNaoi10 vgnd A sndNA vgnd nshort m=1 w=840e-3 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMNaoi11 sndNA B X vgnd nshort m=1 w=840e-3 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMNaoi20 X inor vgnd vgnd nshort m=1 w=840e-3 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMPnor0 vpwr A sndPA vpwr phighvt m=1 w=1.26 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMPnor1 sndPA B inor vpwr phighvt m=1 w=1.26 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMPaoi10 pmid A vpwr vpwr phighvt m=1 w=1.26 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMPaoi11 pmid B vpwr vpwr phighvt m=1 w=1.26 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMPaoi20 X inor pmid vpwr phighvt m=1 w=1.26 l=150e-3 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__inv_1 A Y vgnd vnb vpb vpwr
*.PININFO A:I vgnd:I vnb:I vpb:I vpwr:I Y:O
XICEA A / icecap
XICEY Y / icecap
mMIN1 Y A vgnd vnb nshort m=1 w=0.74 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mMIP1 Y A vpwr vpb phighvt m=1 w=1.12 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on 
+ amuxbusb_on_n analog_en analog_pol analog_sel nga_pad_vswitch_h 
+ nga_pad_vswitch_h_n ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n 
+ nmida_vccd_n nmidb_on_n nmidb_vccd_n out pd_on pd_on_n pd_vswitch_h_n 
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
+ pu_on pu_on_n pu_vddioq_h_n vccd vssd
*.PININFO analog_en:I analog_pol:I analog_sel:I nga_pad_vswitch_h:I 
*.PININFO nga_pad_vswitch_h_n:I ngb_pad_vswitch_h:I ngb_pad_vswitch_h_n:I 
*.PININFO nmida_vccd_n:I nmidb_vccd_n:I out:I pd_vswitch_h_n:I 
*.PININFO pga_amx_vdda_h_n:I pga_pad_vddioq_h_n:I pgb_amx_vdda_h_n:I 
*.PININFO pgb_pad_vddioq_h_n:I pu_vddioq_h_n:I vccd:I vssd:I amuxbusa_on:O 
*.PININFO amuxbusa_on_n:O amuxbusb_on:O amuxbusb_on_n:O nmida_on_n:O 
*.PININFO nmidb_on_n:O pd_on:O pd_on_n:O pu_on:O pu_on_n:O
XICEint_pu_on int_pu_on / icecap
XICEout_i_n out_i_n / icecap
XICEpd_vswitch_h_n pd_vswitch_h_n / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEnet167 net167 / icecap
XICEanalog_pol analog_pol / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
XICEint_pd_on int_pd_on / icecap
XICEout out / icecap
XICEana_en_i_n ana_en_i_n / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEint_amuxb_on int_amuxb_on / icecap
XICEint_pd_on_n int_pd_on_n / icecap
XICEpu_on pu_on / icecap
XICEpu_vddioq_h_n pu_vddioq_h_n / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEnet212 net212 / icecap
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEpd_on_n pd_on_n / icecap
XICEint_amuxa_on int_amuxa_on / icecap
XICEint_amux_a_on_n int_amux_a_on_n / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEint_amux_b_on_n int_amux_b_on_n / icecap
XICEint_fbk_puon_n int_fbk_puon_n / icecap
XICEnet222 net222 / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEana_pol_i ana_pol_i / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEint_fbk_pdon_n int_fbk_pdon_n / icecap
XICEnet137 net137 / icecap
XICEanalog_en analog_en / icecap
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEana_sel_i ana_sel_i / icecap
XICEnet144 net144 / icecap
XICEpd_on pd_on / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEanalog_sel analog_sel / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEpol_xor_out pol_xor_out / icecap
XICEana_sel_i_n ana_sel_i_n / icecap
XICEout_i out_i / icecap
XICEpu_on_n pu_on_n / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEint_pu_on_n int_pu_on_n / icecap
XICEnet172 net172 / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEana_pol_i_n ana_pol_i_n / icecap
XI116 ana_en_i_n int_pd_on_n int_pd_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI113 ana_en_i_n net144 int_amuxa_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI115 ana_en_i_n int_pu_on_n int_pu_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI114 ana_en_i_n net137 int_amuxb_on vssd vssd vccd vccd / sky130_fd_io__nor2_1
XI111 ana_pol_i out_i int_pu_on_n vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI112 ana_pol_i_n out_i_n int_pd_on_n vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI109 ana_sel_i_n pol_xor_out net144 vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI110 pol_xor_out ana_sel_i net137 vssd vssd vccd vccd / sky130_fd_io__nand2_1
XI106 ngb_pad_vswitch_h net212 net172 vssd vccd / sky130_fd_io__hvsbt_nor
XI102 nga_pad_vswitch_h net222 net167 vssd vccd / sky130_fd_io__hvsbt_nor
XI79 int_pu_on pga_pad_vddioq_h_n pgb_pad_vddioq_h_n nga_pad_vswitch_h_n 
+ ngb_pad_vswitch_h_n int_fbk_puon_n vssd vccd / sky130_fd_io__gpiov2_amux_nand5
XI80 int_pd_on pga_pad_vddioq_h_n pgb_pad_vddioq_h_n nga_pad_vswitch_h_n 
+ ngb_pad_vswitch_h_n int_fbk_pdon_n vssd vccd / sky130_fd_io__gpiov2_amux_nand5
XI78 int_amuxb_on pu_vddioq_h_n pd_vswitch_h_n nmidb_vccd_n amuxbusb_on_n vssd 
+ vccd / sky130_fd_io__gpiov2_amux_nand4
XI77 int_amuxa_on pu_vddioq_h_n pd_vswitch_h_n nmida_vccd_n amuxbusa_on_n vssd 
+ vccd / sky130_fd_io__gpiov2_amux_nand4
XI101 pga_pad_vddioq_h_n pga_amx_vdda_h_n net222 vssd vccd / 
+ sky130_fd_io__hvsbt_nand2
XI121 int_amux_b_on_n net172 nmidb_on_n vssd vccd / sky130_fd_io__hvsbt_nand2
XI105 pgb_pad_vddioq_h_n pgb_amx_vdda_h_n net212 vssd vccd / 
+ sky130_fd_io__hvsbt_nand2
XI120 int_amux_a_on_n net167 nmida_on_n vssd vccd / sky130_fd_io__hvsbt_nand2
XI45 ana_pol_i out_i pol_xor_out vssd vccd / sky130_fd_io__xor2_1
XI41 ana_pol_i_n ana_pol_i vssd vssd vccd vccd / sky130_fd_io__inv_1
XI89 int_amuxa_on int_amux_a_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI39 analog_sel ana_sel_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI40 ana_sel_i_n ana_sel_i vssd vssd vccd vccd / sky130_fd_io__inv_1
XI35 analog_pol ana_pol_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI74 amuxbusb_on_n amuxbusb_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI73 amuxbusa_on_n amuxbusa_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI76 int_fbk_pdon_n pd_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI58 analog_en ana_en_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI75 int_fbk_puon_n pu_on vssd vssd vccd vccd / sky130_fd_io__inv_1
XI43 out out_i_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI44 out_i_n out_i vssd vssd vccd vccd / sky130_fd_io__inv_1
XI91 int_amuxb_on int_amux_b_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI93 pu_on pu_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
XI95 pd_on pd_on_n vssd vssd vccd vccd / sky130_fd_io__inv_1
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix analog_en analog_pol analog_sel 
+ enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h_n nga_amx_vswitch_h 
+ nga_pad_vswitch_h ngb_amx_vswitch_h ngb_pad_vswitch_h nmida_vccd nmidb_vccd 
+ out pd_csd_vswitch_h pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n 
+ pgb_pad_vddioq_h_n pu_csd_vddioq_h_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
*.PININFO enable_vswitch_h:I hld_i_h_n:I out:I vccd:I vdda:I vddio_q:I vssa:I 
*.PININFO vssd:I vswitch:I enable_vdda_h_n:O nga_amx_vswitch_h:O 
*.PININFO nga_pad_vswitch_h:O ngb_amx_vswitch_h:O ngb_pad_vswitch_h:O 
*.PININFO nmida_vccd:O nmidb_vccd:O pd_csd_vswitch_h:O pga_amx_vdda_h_n:O 
*.PININFO pga_pad_vddioq_h_n:O pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O 
*.PININFO pu_csd_vddioq_h_n:O
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEpu_on pu_on / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
XICEpd_on pd_on / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEout out / icecap
XICEpu_on_n pu_on_n / icecap
XICEanalog_en analog_en / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEpd_on_n pd_on_n / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEanalog_pol analog_pol / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEanalog_sel analog_sel / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
Xamux_ls amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vswitch_h 
+ amux_en_vswitch_h_n analog_en enable_vdda_h enable_vdda_h_n enable_vswitch_h 
+ hld_i_h_n vccd vdda vddio_q vssa vssd vswitch / 
+ sky130_fd_io__gpiov2_amux_ls_i2c_fix
Xamux_sw_drvr amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h 
+ amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on amuxbusa_on_n amuxbusb_on 
+ amuxbusb_on_n hld_i_h_n nga_amx_vswitch_h nga_pad_vswitch_h 
+ nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h ngb_pad_vswitch_h_n 
+ nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd nmidb_vccd_n 
+ pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n 
+ pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch / 
+ sky130_fd_io__gpiov2_amux_drvr_i2c_fix
Xamux_lv_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n analog_en 
+ analog_pol analog_sel nga_pad_vswitch_h nga_pad_vswitch_h_n 
+ ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n 
+ nmidb_vccd_n out pd_on pd_on_n pd_csd_vswitch_h_n pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_on pu_on_n 
+ pu_csd_vddioq_h_n vccd vssd / sky130_fd_io__gpiov2_amux_decoder
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_amux_switch ag_hv ng_ag_vpmp ng_pad_vpmp nghs_h 
+ nmid_vdda pad_hv_n0 pad_hv_n1 pad_hv_n2 pad_hv_n3 pad_hv_p0 pad_hv_p1 
+ pd_h_vdda pd_h_vddio pg_ag_vdda pg_pad_vddioq pghs_h pug_h vdda vddio 
+ vpb_drvr vssa vssd vssio
*.PININFO ng_ag_vpmp:I ng_pad_vpmp:I nghs_h:I nmid_vdda:I pd_h_vdda:I 
*.PININFO pd_h_vddio:I pg_ag_vdda:I pg_pad_vddioq:I pghs_h:I vdda:I vddio:I 
*.PININFO vssa:I vssd:I vssio:I ag_hv:B pad_hv_n0:B pad_hv_n1:B pad_hv_n2:B 
*.PININFO pad_hv_n3:B pad_hv_p0:B pad_hv_p1:B pug_h:B vpb_drvr:B
XICEnmid_vdda nmid_vdda / icecap
XICEpad_hv_n1 pad_hv_n1 / icecap
XICEpug_h pug_h / icecap
XICEnet85 net85 / icecap
XICEpad_hv_n3 pad_hv_n3 / icecap
XI78<0> mid / icecap
XI78<1> mid1 / icecap
XICEpg_pad_vddioq pg_pad_vddioq / icecap
XICEpd_h_vddio pd_h_vddio / icecap
XICEnghs_h nghs_h / icecap
XICEpg_ag_vdda pg_ag_vdda / icecap
XICEag_hv ag_hv / icecap
XICEvddio vddio / icecap
XICEpad_hv_p1 pad_hv_p1 / icecap
XICEpad_hv_n2 pad_hv_n2 / icecap
XICEmid1 mid1 / icecap
XICEmid mid / icecap
XICEnet83 net83 / icecap
XICEpad_hv_n0 pad_hv_n0 / icecap
XICEpghs_h pghs_h / icecap
XICEpd_h_vdda pd_h_vdda / icecap
XICEng_ag_vpmp ng_ag_vpmp / icecap
XICEng_pad_vpmp ng_pad_vpmp / icecap
XICEpad_hv_p0 pad_hv_p0 / icecap
xI72 vssa vddio condiode
xI71 mid1 vddio condiode
xI70 mid vddio condiode
XI56 vssa net85 / s8_esd_res75only_small
XI12 vssa net83 / s8_esd_res75only_small
mI46 pad_hv_n3 ng_pad_vpmp mid1 mid1 nhv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI35 mid ng_pad_vpmp pad_hv_n1 mid nhv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 pad_hv_n0 ng_pad_vpmp mid mid nhv m=3 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI45 mid1 ng_pad_vpmp pad_hv_n2 mid1 nhv m=3 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI28 mid ng_ag_vpmp ag_hv mid nhv m=5 w=10.0 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI57 mid1 nmid_vdda net85 vssa nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI63 pug_h nghs_h pg_pad_vddioq vssio nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI47 mid1 ng_ag_vpmp ag_hv mid1 nhv m=5 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI75<1> mid pd_h_vdda vssa net050<0> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI75<0> mid1 pd_h_vdda vssa net050<1> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI74<1> mid pd_h_vddio vssa net051<0> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI74<0> mid1 pd_h_vddio vssa net051<1> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 mid nmid_vdda net83 vssa nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI22 mid pug_h pad_hv_p1 vpb_drvr phv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 mid pug_h pad_hv_p0 vpb_drvr phv m=2 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI62 pg_pad_vddioq pghs_h pug_h vpb_drvr phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI26 mid pg_ag_vdda ag_hv vdda phv m=4 w=10.0 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_amux_i2c_fix amuxbus_a amuxbus_b analog_en 
+ analog_pol analog_sel enable_vdda_h enable_vswitch_h hld_i_h_n 
+ nga_pad_vpmp_h ngb_pad_vpmp_h nghs_h out pad pd_csd_h pghs_h pu_csd_h 
+ pug_h<1> pug_h<0> vccd vdda vddio vddio_q vpb_drvr vssa vssd vssio vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
*.PININFO enable_vswitch_h:I hld_i_h_n:I nghs_h:I out:I pghs_h:I vccd:I vdda:I 
*.PININFO vddio:I vddio_q:I vssa:I vssd:I vssio:I vswitch:I nga_pad_vpmp_h:O 
*.PININFO ngb_pad_vpmp_h:O pd_csd_h:O pu_csd_h:O amuxbus_a:B amuxbus_b:B pad:B 
*.PININFO pug_h<1>:B pug_h<0>:B vpb_drvr:B
XICEpghs_h pghs_h / icecap
XICEnga_pad_vpmp_h nga_pad_vpmp_h / icecap
XICEngb_amx_vpmp_h ngb_amx_vpmp_h / icecap
XICEanalog_pol analog_pol / icecap
XICEvssio vssio / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEpad pad / icecap
XICEnet128 net128 / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEnet126 net126 / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEpug_h<1> pug_h<1> / icecap
XICEamuxbus_a amuxbus_a / icecap
XICEpu_csd_h pu_csd_h / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEhld_i_h_amux_sw hld_i_h_amux_sw / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEnet120 net120 / icecap
XICEout out / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEnga_amx_vpmp_h nga_amx_vpmp_h / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEnet142 net142 / icecap
XICEnghs_h nghs_h / icecap
XICEnet139 net139 / icecap
XICEnet124 net124 / icecap
XICEpug_h<0> pug_h<0> / icecap
XICEngb_pad_vpmp_h ngb_pad_vpmp_h / icecap
XICEamuxbus_b amuxbus_b / icecap
XICEnet143 net143 / icecap
XICEanalog_sel analog_sel / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEpd_csd_h pd_csd_h / icecap
XICEnet144 net144 / icecap
XICEanalog_en analog_en / icecap
XI78 hld_i_h_n hld_i_h_amux_sw vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XBBM_logic analog_en analog_pol analog_sel enable_vdda_h enable_vdda_h_n 
+ enable_vswitch_h hld_i_h_n nga_amx_vpmp_h nga_pad_vpmp_h ngb_amx_vpmp_h 
+ ngb_pad_vpmp_h nmida_vccd nmidb_vccd out pd_csd_h pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_h vccd vdda 
+ vddio_q vssa vssd vswitch / sky130_fd_io__gpiov2_amux_ctl_logic_i2c_fix
xI77 vssa vdda condiode
XI26 net128 net142 / s8_esd_res75only_small
XI58 net126 net139 / s8_esd_res75only_small
XI28 net124 net144 / s8_esd_res75only_small
XI57 pad net126 / s8_esd_res75only_small
XI27 net120 net143 / s8_esd_res75only_small
XI55 pad net128 / s8_esd_res75only_small
XI54 pad net124 / s8_esd_res75only_small
XI53 pad net120 / s8_esd_res75only_small
Xmux_a amuxbus_a nga_amx_vpmp_h nga_pad_vpmp_h nghs_h nmida_vccd net144 net144 
+ net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pghs_h pug_h<0> vdda vddio vpb_drvr vssa vssd vssio / 
+ sky130_fd_io__gpio_ovtv2_amux_switch
Xmux_b amuxbus_b ngb_amx_vpmp_h ngb_pad_vpmp_h nghs_h nmidb_vccd net144 net144 
+ net139 net139 net143 net142 enable_vdda_h_n hld_i_h_amux_sw pgb_amx_vdda_h_n 
+ pgb_pad_vddioq_h_n pghs_h pug_h<1> vdda vddio vpb_drvr vssa vssd vssio / 
+ sky130_fd_io__gpio_ovtv2_amux_switch
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix dm<2> dm<1> dm<0> dm_h<2> 
+ dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n hyst_trim 
+ hyst_trim_h hyst_trim_h_n ib_mode_sel<1> ib_mode_sel<0> ib_mode_sel_h<1> 
+ ib_mode_sel_h<0> ib_mode_sel_h_n<1> ib_mode_sel_h_n<0> inp_dis inp_dis_h 
+ inp_dis_h_n od_i_h_n slew_ctl<1> slew_ctl<0> slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> startup_rst_h startup_st_h vcc_io vgnd vpwr 
+ vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I hld_i_h_n:I hyst_trim:I ib_mode_sel<1>:I 
*.PININFO ib_mode_sel<0>:I inp_dis:I od_i_h_n:I slew_ctl<1>:I slew_ctl<0>:I 
*.PININFO startup_rst_h:I startup_st_h:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I 
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
*.PININFO hyst_trim_h:O hyst_trim_h_n:O ib_mode_sel_h<1>:O ib_mode_sel_h<0>:O 
*.PININFO ib_mode_sel_h_n<1>:O ib_mode_sel_h_n<0>:O inp_dis_h:O inp_dis_h_n:O 
*.PININFO slew_ctl_h<1>:O slew_ctl_h<0>:O slew_ctl_h_n<1>:O slew_ctl_h_n<0>:O 
*.PININFO vtrip_sel_h:O vtrip_sel_h_n:O
XICEdm_h_n<0> dm_h_n<0> / icecap
XI851<0> ib_mode_sel<1> / icecap
XI851<1> ib_mode_sel<0> / icecap
XI837<0> ib_mode_sel_rst_h<1> / icecap
XI837<1> ib_mode_sel_rst_h<0> / icecap
XI843<0> dm_h<2> / icecap
XI843<1> dm_h<1> / icecap
XICEod_i_h od_i_h / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEdm_h<0> dm_h<0> / icecap
XICEie_n_st_h ie_n_st_h / icecap
XICEhyst_trim_st_h hyst_trim_st_h / icecap
XICEvtrip_sel vtrip_sel / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XICEinp_dis inp_dis / icecap
XICEdm<0> dm<0> / icecap
XICEdm_rst_h<2> dm_rst_h<2> / icecap
XI844<0> slew_ctl<1> / icecap
XI844<1> slew_ctl<0> / icecap
XI846<0> slew_ctl_h<1> / icecap
XI846<1> slew_ctl_h<0> / icecap
XICEhyst_trim_h_n hyst_trim_h_n / icecap
XICEdm_st_h<2> dm_st_h<2> / icecap
XICEhyst_trim_rst_h hyst_trim_rst_h / icecap
XICEdm_rst_h<0> dm_rst_h<0> / icecap
XI845<0> slew_ctl_rst_h<1> / icecap
XI845<1> slew_ctl_rst_h<0> / icecap
XI839<0> dm<2> / icecap
XI839<1> dm<1> / icecap
XICEie_n_rst_h ie_n_rst_h / icecap
XI840<0> dm_h_n<2> / icecap
XI840<1> dm_h_n<1> / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEdm_st_h<0> dm_st_h<0> / icecap
XICEhyst_trim_h hyst_trim_h / icecap
XI838<0> dm_st_h<2> / icecap
XI838<1> dm_st_h<1> / icecap
XICEinp_dis_h inp_dis_h / icecap
XICEdm_rst_h<1> dm_rst_h<1> / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEstartup_rst_h startup_rst_h / icecap
XICEstartup_st_h startup_st_h / icecap
XICEhyst_trim hyst_trim / icecap
XI841<0> ib_mode_sel_h<1> / icecap
XI841<1> ib_mode_sel_h<0> / icecap
XI848<0> ib_mode_sel_st_h<1> / icecap
XI848<1> ib_mode_sel_st_h<0> / icecap
XICEdm_st_h<1> dm_st_h<1> / icecap
XI847<0> slew_ctl_st_h<1> / icecap
XI847<1> slew_ctl_st_h<0> / icecap
XICEtrip_sel_st_h trip_sel_st_h / icecap
XICEtrip_sel_rst_h trip_sel_rst_h / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XI850<0> slew_ctl_h_n<1> / icecap
XI850<1> slew_ctl_h_n<0> / icecap
XI849<0> ib_mode_sel_h_n<1> / icecap
XI849<1> ib_mode_sel_h_n<0> / icecap
XI842<0> dm_rst_h<2> / icecap
XI842<1> dm_rst_h<1> / icecap
XI836 od_i_h_n od_i_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
Xtrip_sel_st trip_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> od_i_h vgnd / sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> vgnd od_i_h / sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> startup_st_h startup_rst_h / sky130_fd_io__tk_opti
XI615 hyst_trim_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI614 hyst_trim_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
XI598<1> ib_mode_sel_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
XI598<0> ib_mode_sel_st_h<0> od_i_h vgnd / sky130_fd_io__tk_opti
XI597<1> ib_mode_sel_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI597<0> ib_mode_sel_rst_h<0> vgnd od_i_h / sky130_fd_io__tk_opti
XI337<1> dm_st_h<0> startup_rst_h startup_st_h / sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI666<1> slew_ctl_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
XI666<0> slew_ctl_st_h<0> od_i_h vgnd / sky130_fd_io__tk_opti
XI665<1> slew_ctl_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI665<0> slew_ctl_rst_h<0> vgnd od_i_h / sky130_fd_io__tk_opti
XI687 ie_n_st_h startup_st_h startup_rst_h / sky130_fd_io__tk_opti
XI686 ie_n_rst_h startup_rst_h startup_st_h / sky130_fd_io__tk_opti
Xdm_ls_0 hld_i_h_n dm<0> dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
Xinp_dis_ls hld_i_h_n inp_dis inp_dis_h inp_dis_h_n ie_n_rst_h ie_n_st_h 
+ vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
Xtrip_sel_ls hld_i_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n trip_sel_rst_h 
+ trip_sel_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
XI616 hld_i_h_n hyst_trim hyst_trim_h hyst_trim_h_n hyst_trim_rst_h 
+ hyst_trim_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
XI595<1> hld_i_h_n ib_mode_sel<1> ib_mode_sel_h<1> ib_mode_sel_h_n<1> 
+ ib_mode_sel_rst_h<1> ib_mode_sel_st_h<1> net58<0> net56<0> net57<0> / 
+ sky130_fd_io__com_ctl_ls
XI595<0> hld_i_h_n ib_mode_sel<0> ib_mode_sel_h<0> ib_mode_sel_h_n<0> 
+ ib_mode_sel_rst_h<0> ib_mode_sel_st_h<0> net58<1> net56<1> net57<1> / 
+ sky130_fd_io__com_ctl_ls
XI667<1> hld_i_h_n slew_ctl<1> slew_ctl_h<1> slew_ctl_h_n<1> slew_ctl_rst_h<1> 
+ slew_ctl_st_h<1> net61<0> net59<0> net60<0> / sky130_fd_io__com_ctl_ls
XI667<0> hld_i_h_n slew_ctl<0> slew_ctl_h<0> slew_ctl_h_n<0> slew_ctl_rst_h<0> 
+ slew_ctl_st_h<0> net61<1> net59<1> net60<1> / sky130_fd_io__com_ctl_ls
Xdm_ls<2> hld_i_h_n dm<2> dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
Xdm_ls<1> hld_i_h_n dm<1> dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
.ENDS
.SUBCKT sky130_fd_io__enh_nand2_1_sp in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpwr phv m=4 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out in1 vpwr vpwr phv m=2 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net25 vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net25 in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__enh_nor2_x1 in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEnet16 net16 / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 net16 in0 vpwr vpwr phv m=1 w=1.00 l=0.60 mult=2 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out in1 net16 vpwr phv m=1 w=1.00 l=0.60 mult=2 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out in1 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__enh_nand2_1 in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 out in0 vpwr vpwr phv m=3 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out in1 vpwr vpwr phv m=3 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net25 vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net25 in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nor2_4_enhpath in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEnet16 net16 / icecap
XICEin0 in0 / icecap
XICEin1 in1 / icecap
mI3 net16 in0 vpwr vpwr phv m=16 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out in1 net16 vpwr phv m=16 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in0 vgnd vgnd nhv m=8 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out in1 vgnd vgnd nhv m=8 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__nand2_2_enhpath in0 in1 out vgnd vpwr
*.PININFO in0:I in1:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin1 in1 / icecap
XICEin0 in0 / icecap
mI3 out in0 vpwr vpwr phv m=4 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 out in1 vpwr vpwr phv m=4 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in1 net25 vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 net25 in0 vgnd vgnd nhv m=1 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix enable_h hld_h_n hld_i_h_n 
+ hld_i_ovr_h hld_ovr od_i_h_n vcc_io vgnd vpwr
*.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h_n:O 
*.PININFO hld_i_ovr_h:O od_i_h_n:O
Xhld_nand enable_h hld_h_n n1 vgnd vcc_io / sky130_fd_io__enh_nand2_1_sp
XI50 od_i_h_n net45 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI46 n1 n1 n2 vgnd vcc_io / sky130_fd_io__enh_nor2_x1
XI49 od_h od_h od_i_h_n vgnd vcc_io / sky130_fd_io__enh_nor2_x1
XI48 enable_h enable_h od_h vgnd vcc_io / sky130_fd_io__enh_nand2_1
XI155 n3 n3 hld_i_h_n vgnd vcc_io / sky130_fd_io__nor2_4_enhpath
XI154 n2 n2 n3 vgnd vcc_io / sky130_fd_io__nand2_2_enhpath
Xhld_ovr_ls n2 hld_ovr hld_ovr_h net79 od_h vgnd vcc_io vgnd vpwr / 
+ sky130_fd_io__com_ctl_ls
XI30 net45 hld_i_ovr_h_n hld_i_ovr_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI26 n2 hld_ovr_h hld_i_ovr_h_n vgnd vcc_io / sky130_fd_io__hvsbt_nor
.ENDS
.SUBCKT sky130_fd_io__gpio_ctlv2_i2c_fix dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_h enable_inp_h hld_h_n hld_i_h_n 
+ hld_i_ovr_h hld_ovr hyst_trim hyst_trim_h hyst_trim_h_n ib_mode_sel<1> 
+ ib_mode_sel<0> ib_mode_sel_h<1> ib_mode_sel_h<0> ib_mode_sel_h_n<1> 
+ ib_mode_sel_h_n<0> inp_dis inp_dis_h_n od_i_h_n slew_ctl<1> slew_ctl<0> 
+ slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> vccd vddio_q 
+ vssd vtrip_sel vtrip_sel_h
*.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I enable_inp_h:I hld_h_n:I 
*.PININFO hld_ovr:I hyst_trim:I ib_mode_sel<1>:I ib_mode_sel<0>:I inp_dis:I 
*.PININFO slew_ctl<1>:I slew_ctl<0>:I vccd:I vddio_q:I vssd:I vtrip_sel:I 
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
*.PININFO hld_i_h_n:O hld_i_ovr_h:O hyst_trim_h:O hyst_trim_h_n:O 
*.PININFO ib_mode_sel_h<1>:O ib_mode_sel_h<0>:O ib_mode_sel_h_n<1>:O 
*.PININFO ib_mode_sel_h_n<0>:O inp_dis_h_n:O od_i_h_n:O slew_ctl_h<1>:O 
*.PININFO slew_ctl_h<0>:O slew_ctl_h_n<1>:O slew_ctl_h_n<0>:O vtrip_sel_h:O
Xls_bank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hyst_trim hyst_trim_h hyst_trim_h_n ib_mode_sel<1> 
+ ib_mode_sel<0> ib_mode_sel_h<1> ib_mode_sel_h<0> ib_mode_sel_h_n<1> 
+ ib_mode_sel_h_n<0> inp_dis net83 inp_dis_h_n od_i_h_n slew_ctl<1> 
+ slew_ctl<0> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> slew_ctl_h_n<0> 
+ startup_rst_h inp_startup_en_h vddio_q vssd vccd vtrip_sel vtrip_sel_h net77 
+ / sky130_fd_io__gpio_ovtv2_ctl_lsbank_i2c_fix
Xhld_dis_blk enable_h hld_h_n hld_i_h_n hld_i_ovr_h hld_ovr od_i_h_n vddio_q 
+ vssd vccd / sky130_fd_io__gpio_ovtv2_ctl_hld_i2c_fix
XI75 enable_inp_h enable_h startup_rst_h vssd vddio_q / sky130_fd_io__hvsbt_nor
XI56 net109 enable_inp_h net108 vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI77 od_i_h_n net109 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI57 net108 inp_startup_en_h vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_lvls enable_vddio_lv in out out_b vcchib vssd
*.PININFO enable_vddio_lv:I in:I vcchib:I vssd:I out:O out_b:O
XICEin in / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEout out / icecap
XICEfbk fbk / icecap
XICEout_b out_b / icecap
XICEfbk_n fbk_n / icecap
mI248 fbk_n in vcchib vcchib phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI271 out out_b vcchib vcchib phighvt m=2 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI281 fbk_n enable_vddio_lv vcchib vcchib phv m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI272 out_b fbk vcchib vcchib phighvt m=1 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI277 fbk fbk_n vcchib vcchib phighvt m=1 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI273 out out_b vssd vssd nshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI278 fbk fbk_n vssd vssd nshort m=1 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI305 out_b fbk vssd vssd nshort m=1 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI535 fbk_n in vssd_1 vssd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI279 vssd_1 enable_vddio_lv vssd vssd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ipath_hvls en_h_n in inb out out_b vddio_q vssd
*.PININFO en_h_n:I in:I inb:I vddio_q:I vssd:I out:O out_b:O
XICEfbk_b fbk_b / icecap
XICEout out / icecap
XICEinb inb / icecap
XICEout_b out_b / icecap
XICEen_h_n en_h_n / icecap
XICEfbk fbk / icecap
XICEin in / icecap
mI250 fbk fbk_b vddio_q vddio_q phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI253 out out_b vddio_q vddio_q phv m=5 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI249 fbk_b fbk vddio_q vddio_q phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI248 out_b fbk vddio_q vddio_q phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI247 out_b fbk vssd vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI252 out out_b vssd vssd nhv m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI304 fbk inb vssd vssd nhv m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI262 fbk en_h_n vssd vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI246 fbk_b in vssd vssd nhv m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_in_buf en_h en_h_n enable_vddio_lv in_h in_vt 
+ mode_normal_n mode_ref_3v_n mode_ref_n mode_vccd_n out out_n vcchib vddio_q 
+ vrefin vssd vtrip_sel_h vtrip_sel_h_n
*.PININFO en_h:I en_h_n:I enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I 
*.PININFO mode_ref_3v_n:I mode_ref_n:I mode_vccd_n:I vcchib:I vddio_q:I 
*.PININFO vrefin:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I out:O out_n:O
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEvirt_pwr virt_pwr / icecap
XICEvddio_ref vddio_ref / icecap
XICEvcchib_int1 vcchib_int1 / icecap
XICEvddio_ref1 vddio_ref1 / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEfbk fbk / icecap
XICEin_h in_h / icecap
XICEen_h en_h / icecap
XICEen_h_n en_h_n / icecap
XICEout out / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEvrefin vrefin / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEvcchib_int vcchib_int / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEvirt_pwr2 virt_pwr2 / icecap
XICEin_b in_b / icecap
XICEmode_normal_cmos_h mode_normal_cmos_h / icecap
XICEout_n out_n / icecap
XICEenable_vddio_lv_n enable_vddio_lv_n / icecap
XICEmode_normal_cmos_h_n mode_normal_cmos_h_n / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEvirt_pwr1 virt_pwr1 / icecap
XICEin_vt in_vt / icecap
XICEfbk1 fbk1 / icecap
XICEfbk2 fbk2 / icecap
XI35 enable_vddio_lv en_h enable_vddio_lv_n vssd vcchib / sky130_fd_io__hvsbt_nand2
xI405 virt_pwr1 vddio_q condiode
xI404 virt_pwr vddio_q condiode
XI488 vtrip_sel_h mode_normal_n mode_normal_cmos_h vssd vddio_q / 
+ sky130_fd_io__hvsbt_nor
XI43 mode_normal_cmos_h mode_normal_cmos_h_n vssd vddio_q / 
+ sky130_fd_io__hvsbt_inv_x1
mI630 vssd vssd vssd vssd nhv m=3 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI105 fbk1 in_b fbk vssd nhv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI620 vssd vssd vssd vssd nhv m=3 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI441 in_vt vtrip_sel_h_n vssd vssd nhv m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI417 out en_h_n vssd vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI419 out_n en_h_n vssd vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI394 vssd vssd vssd vssd nhv m=3 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI494 fbk in_h vssd vssd nhv m=6 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 fbk2 in_b fbk vssd nhv m=3 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI26 out in_b vssd vssd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI49 vddio_ref vrefin virt_pwr virt_pwr nhvnative m=3 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI451 fbk in_vt vssd vssd nhv m=12 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI453 in_b in_h fbk vssd nhv m=6 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI111 vddio_ref1 vrefin virt_pwr1 virt_pwr1 nhvnative m=3 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI446 out_n out vssd vssd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI389 virt_pwr vssd vssd vssd nhv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI450 in_b in_vt fbk vssd nhv m=6 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI274 fbk1 mode_ref_n virt_pwr1 virt_pwr1 phv m=4 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI116 virt_pwr mode_normal_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI109 in_b in_h virt_pwr virt_pwr phv m=3 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI25 out in_b virt_pwr1 virt_pwr1 phv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 fbk2 mode_normal_cmos_h_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI611 fbk1 mode_normal_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI396 vddio_ref1 mode_ref_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI115 virt_pwr mode_vccd_n vcchib_int virt_pwr phv m=4 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI478 vcchib_int1 enable_vddio_lv_n vcchib vcchib pshort m=8 w=5.00 l=0.25 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI373 vddio_ref mode_ref_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI403 out in_b virt_pwr2 virt_pwr2 phv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI376 fbk2 mode_ref_3v_n virt_pwr1 virt_pwr1 phv m=4 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI477 vcchib_int enable_vddio_lv_n vcchib vcchib pshort m=8 w=5.00 l=0.25 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI401 in_b in_h virt_pwr2 virt_pwr2 phv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI457 out_n out virt_pwr1 virt_pwr1 phv m=5 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI486 fbk1 mode_vccd_n vcchib_int virt_pwr1 phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI400 virt_pwr2 mode_vccd_n vcchib_int virt_pwr2 phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI381 virt_pwr1 mode_vccd_n vcchib_int1 virt_pwr1 phv m=6 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI380 virt_pwr1 mode_normal_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ibuf_se en_h en_h_n enable_vddio_lv ibufmux_out 
+ ibufmux_out_h in_h in_vt mode_normal_n mode_ref_3v_n mode_ref_n mode_vccd_n 
+ vcchib vddio_q vrefin vssd vtrip_sel_h vtrip_sel_h_n
*.PININFO en_h:I en_h_n:I enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I 
*.PININFO mode_ref_3v_n:I mode_ref_n:I mode_vccd_n:I vcchib:I vddio_q:I 
*.PININFO vrefin:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I ibufmux_out:O 
*.PININFO ibufmux_out_h:O
XICEnet43 net43 / icecap
XICEin_h in_h / icecap
XICEout_n out_n / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEin_vt in_vt / icecap
XICEvrefin vrefin / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEen_h_n en_h_n / icecap
XICEibufmux_out_h ibufmux_out_h / icecap
XICEibufmux_out ibufmux_out / icecap
XICEen_h en_h / icecap
XICEout out / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEnet49 net49 / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
Xlvls enable_vddio_lv out ibufmux_out net43 vcchib vssd / 
+ sky130_fd_io__gpio_ovtv2_ipath_lvls
Xhvls en_h_n out out_n ibufmux_out_h net49 vddio_q vssd / 
+ sky130_fd_io__gpio_ovtv2_ipath_hvls
Xbuf en_h en_h_n enable_vddio_lv in_h in_vt mode_normal_n mode_ref_3v_n 
+ mode_ref_n mode_vccd_n out out_n vcchib vddio_q vrefin vssd vtrip_sel_h 
+ vtrip_sel_h_n / sky130_fd_io__gpio_ovtv2_in_buf
.ENDS
.SUBCKT s8_esd_res250only_small pad rout
*.PININFO pad:B rout:B
rI175 net12 net16 mrp1 m=1 w=2 l=10.07
rI229 net16 rout mrp1 m=1 w=2 l=0.17
rI228 pad net12 mrp1 m=1 w=2 l=0.17
rI237<1> net16 rout short
rI237<2> net16 rout short
rI234<1> pad net12 short
rI234<2> pad net12 short
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_buf_localesd in_h out_h out_vt vddio_q vssd 
+ vtrip_sel_h
*.PININFO in_h:I vtrip_sel_h:I out_h:O out_vt:O vddio_q:B vssd:B
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEin_h in_h / icecap
XICEout_vt out_vt / icecap
XICEout_h out_h / icecap
mhv_passgate out_h vtrip_sel_h out_vt vssd nhv m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xesd_res in_h out_h / s8_esd_res250only_small
Xggnfet6 vssd vddio_q vssd vddio_q out_h / s8_esd_signal_5_sym_hv_local_5term
Xggnfet1 vssd out_h vssd vddio_q vssd / s8_esd_signal_5_sym_hv_local_5term
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ictl_logic dm_h_n<2> dm_h_n<1> dm_h_n<0> hys_trim 
+ ibuf_mode_sel<0> ibuf_mode_sel<1> inp_dis_h_n inp_dis_i_h inp_dis_i_h_n 
+ mode_normal_n mode_ref_3v_n mode_ref_n mode_vccd_n tripsel_i_h tripsel_i_h_n 
+ vddio_q vssd vtrip_sel_h
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I hys_trim:I ibuf_mode_sel<0>:I 
*.PININFO ibuf_mode_sel<1>:I inp_dis_h_n:I vddio_q:I vssd:I vtrip_sel_h:I 
*.PININFO inp_dis_i_h:O inp_dis_i_h_n:O mode_normal_n:O mode_ref_3v_n:O 
*.PININFO mode_ref_n:O mode_vccd_n:O tripsel_i_h:O tripsel_i_h_n:O
XICEtripsel_i_h_n tripsel_i_h_n / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEibuf_mode_sel<1> ibuf_mode_sel<1> / icecap
XICEinp_dis_i_h_n inp_dis_i_h_n / icecap
XICEnet55 net55 / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XICEinp_dis_i_h inp_dis_i_h / icecap
XICEibuf_mode_sel<0> ibuf_mode_sel<0> / icecap
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEtripsel_i_h tripsel_i_h / icecap
XICEnand_dm01 nand_dm01 / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEdm_h_n<0> dm_h_n<0> / icecap
XICEand_dm01 and_dm01 / icecap
XICEnet60 net60 / icecap
XICEnet66 net66 / icecap
XICEdm_buf_dis dm_buf_dis / icecap
XICEdm_h_n<1> dm_h_n<1> / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEmode_ref mode_ref / icecap
XICEnet70 net70 / icecap
XICEhys_trim hys_trim / icecap
XICEdm_h_n<2> dm_h_n<2> / icecap
XI41 net66 mode_normal_n tripsel_i_h vssd vddio_q / sky130_fd_io__hvsbt_nor
XI34 ibuf_mode_sel<1> net70 net60 vssd vddio_q / sky130_fd_io__hvsbt_nor
XI33 ibuf_mode_sel<1> ibuf_mode_sel<0> net55 vssd vddio_q / sky130_fd_io__hvsbt_nor
Xdm10nand_inv nand_dm01 and_dm01 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI68 inp_dis_i_h inp_dis_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI43 tripsel_i_h tripsel_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI50 mode_ref_n mode_ref vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI39 ibuf_mode_sel<0> net70 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI61 vtrip_sel_h net66 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
Xinpdis dm_buf_dis inp_dis_h_n inp_dis_i_h vssd vddio_q / sky130_fd_io__hvsbt_nand2
Xdm210 dm_h_n<2> and_dm01 dm_buf_dis vssd vddio_q / sky130_fd_io__hvsbt_nand2
Xdm10 dm_h_n<1> dm_h_n<0> nand_dm01 vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI40 inp_dis_i_h_n ibuf_mode_sel<1> mode_ref_n vssd vddio_q / 
+ sky130_fd_io__hvsbt_nand2
XI36 inp_dis_i_h_n net60 mode_vccd_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI35 inp_dis_i_h_n net55 mode_normal_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI52 mode_ref hys_trim mode_ref_3v_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
.ENDS
.SUBCKT sky130_fd_io__gpio_ovtv2_ipath dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ enable_vddio_lv hys_trim_h ib_mode_sel_h<1> ib_mode_sel_h<0> inp_dis_h_n out 
+ out_h pad vcchib vddio_q vinref vssd vtrip_sel_h
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I enable_vddio_lv:I hys_trim_h:I 
*.PININFO ib_mode_sel_h<1>:I ib_mode_sel_h<0>:I inp_dis_h_n:I vcchib:I 
*.PININFO vddio_q:I vssd:I vtrip_sel_h:I out:O out_h:O pad:B vinref:B
XICEib_mode_sel_h<0> ib_mode_sel_h<0> / icecap
XICEmode_ref_n mode_ref_n / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEhys_trim_h hys_trim_h / icecap
XICEib_mode_sel_h<1> ib_mode_sel_h<1> / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XI111<0> dm_h_n<2> / icecap
XI111<1> dm_h_n<1> / icecap
XI111<2> dm_h_n<0> / icecap
XICEin_vt in_vt / icecap
XICEen_h_n en_h_n / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEpad pad / icecap
XICEtripsel_i_h_n tripsel_i_h_n / icecap
XICEout out / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEen_h en_h / icecap
XICEvinref vinref / icecap
XICEmode_ref_3v_n mode_ref_3v_n / icecap
XICEmode_vccd_n mode_vccd_n / icecap
XICEtripsel_i_h tripsel_i_h / icecap
XICEin_h in_h / icecap
XICEout_h out_h / icecap
Xibuf_se en_h en_h_n enable_vddio_lv out out_h in_h in_vt mode_normal_n 
+ mode_ref_3v_n mode_ref_n mode_vccd_n vcchib vddio_q vinref vssd tripsel_i_h 
+ tripsel_i_h_n / sky130_fd_io__gpio_ovtv2_ibuf_se
Xesd pad in_h in_vt vddio_q vssd tripsel_i_h / sky130_fd_io__gpio_ovtv2_buf_localesd
Xlogic dm_h_n<2> dm_h_n<1> dm_h_n<0> hys_trim_h ib_mode_sel_h<0> 
+ ib_mode_sel_h<1> inp_dis_h_n en_h_n en_h mode_normal_n mode_ref_3v_n 
+ mode_ref_n mode_vccd_n tripsel_i_h tripsel_i_h_n vddio_q vssd vtrip_sel_h / 
+ sky130_fd_io__gpio_ovtv2_ictl_logic
.ENDS
.SUBCKT sky130_fd_io__top_gpio_ovtv2 amuxbus_a amuxbus_b analog_en analog_pol 
+ analog_sel dm<2> dm<1> dm<0> enable_h enable_inp_h enable_vdda_h 
+ enable_vddio enable_vswitch_h hld_h_n hld_ovr hys_trim ib_mode_sel<1> 
+ ib_mode_sel<0> in in_h inp_dis oe_n out pad pad_a_esd_0_h pad_a_esd_1_h 
+ pad_a_noesd_h slew_ctl<1> slew_ctl<0> slow tie_hi_esd tie_lo_esd vccd vcchib 
+ vdda vddio vddio_q vinref vssa vssd vssio vssio_q vswitch vtrip_sel
*.PININFO analog_en:I analog_pol:I analog_sel:I dm<2>:I dm<1>:I dm<0>:I 
*.PININFO enable_h:I enable_inp_h:I enable_vdda_h:I enable_vddio:I 
*.PININFO enable_vswitch_h:I hld_h_n:I hld_ovr:I hys_trim:I ib_mode_sel<1>:I 
*.PININFO ib_mode_sel<0>:I inp_dis:I oe_n:I out:I slew_ctl<1>:I slew_ctl<0>:I 
*.PININFO slow:I vinref:I vtrip_sel:I in:O in_h:O tie_hi_esd:O tie_lo_esd:O 
*.PININFO amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_0_h:B pad_a_esd_1_h:B 
*.PININFO pad_a_noesd_h:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B 
*.PININFO vssd:B vssio:B vssio_q:B vswitch:B
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_ovr_h nga_pad_vpmp_h ngb_pad_vpmp_h od_i_h_n oe_n out pad pd_csd_h 
+ pghs_h pu_csd_h pug_h<6> pug_h<5> slew_ctl_h<1> slew_ctl_h<0> 
+ slew_ctl_h_n<1> slew_ctl_h_n<0> slow tie_hi_esd tie_lo_esd vccd vddio 
+ vddio_q vpb_drvr vcchib vssa vssd vssio vssio_q / 
+ sky130_fd_io__gpio_ovtv2_opath_i2c_fix_leak_fix
Xovt_amux amuxbus_a amuxbus_b analog_en analog_pol analog_sel enable_vdda_h 
+ enable_vswitch_h hld_i_h_n nga_pad_vpmp_h ngb_pad_vpmp_h tie_hi_esd out pad 
+ pd_csd_h pghs_h pu_csd_h pug_h<6> pug_h<5> vccd vdda vddio vddio_q vpb_drvr 
+ vssa vssd vssio vswitch / sky130_fd_io__gpio_ovtv2_amux_i2c_fix
Xctrl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ enable_h enable_inp_h hld_h_n hld_i_h_n hld_i_ovr_h hld_ovr hys_trim 
+ hyst_trim_h net164 ib_mode_sel<1> ib_mode_sel<0> ib_mode_sel_h<1> 
+ ib_mode_sel_h<0> net166<0> net166<1> inp_dis inp_dis_h_n od_i_h_n 
+ slew_ctl<1> slew_ctl<0> slew_ctl_h<1> slew_ctl_h<0> slew_ctl_h_n<1> 
+ slew_ctl_h_n<0> vccd vddio_q vssd vtrip_sel vtrip_sel_h / 
+ sky130_fd_io__gpio_ctlv2_i2c_fix
XI336 net193 pad_a_esd_1_h / s8_esd_res75only_small
XI335 pad net193 / s8_esd_res75only_small
XI334 net189 pad_a_esd_0_h / s8_esd_res75only_small
Xresd4 pad net189 / s8_esd_res75only_small
rS0 pad pad_a_noesd_h short
Xipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio hyst_trim_h ib_mode_sel_h<1> 
+ ib_mode_sel_h<0> inp_dis_h_n in in_h pad vcchib vddio_q vinref vssd 
+ vtrip_sel_h / sky130_fd_io__gpio_ovtv2_ipath
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_switch amuxbus_hv ng_amx_vpmp_h ng_pad_vpmp_h 
+ nmid_vccd pad_hv_n0 pad_hv_n1 pad_hv_n2 pad_hv_n3 pad_hv_p0 pad_hv_p1 
+ pd_h_vdda pd_h_vddio pg_amx_vdda_h_n pg_pad_vddioq_h_n vdda vddio vssa vssd
*.PININFO ng_amx_vpmp_h:I ng_pad_vpmp_h:I nmid_vccd:I pd_h_vdda:I pd_h_vddio:I 
*.PININFO pg_amx_vdda_h_n:I pg_pad_vddioq_h_n:I vdda:I vddio:I vssa:I vssd:I 
*.PININFO amuxbus_hv:B pad_hv_n0:B pad_hv_n1:B pad_hv_n2:B pad_hv_n3:B 
*.PININFO pad_hv_p0:B pad_hv_p1:B
XICEnet79 net79 / icecap
XICEpad_hv_n1 pad_hv_n1 / icecap
XICEpad_hv_n3 pad_hv_n3 / icecap
XICEpd_h_vdda pd_h_vdda / icecap
XICEng_pad_vpmp_h ng_pad_vpmp_h / icecap
XICEpg_pad_vddioq_h_n pg_pad_vddioq_h_n / icecap
XICEpg_amx_vdda_h_n pg_amx_vdda_h_n / icecap
XICEpad_hv_n0 pad_hv_n0 / icecap
XICEpad_hv_n2 pad_hv_n2 / icecap
XICEng_amx_vpmp_h ng_amx_vpmp_h / icecap
XICEnet77 net77 / icecap
XICEpad_hv_p0 pad_hv_p0 / icecap
XI85<0> mid / icecap
XI85<1> mid1 / icecap
XICEpad_hv_p1 pad_hv_p1 / icecap
XICEamuxbus_hv amuxbus_hv / icecap
XICEmid1 mid1 / icecap
XICEpd_h_vddio pd_h_vddio / icecap
XICEmid mid / icecap
XICEnmid_vccd nmid_vccd / icecap
xI72 vssa vdda condiode
xI71 mid1 vdda condiode
xI70 mid vdda condiode
XI56 vssa net79 / s8_esd_res75only_small
XI12 vssa net77 / s8_esd_res75only_small
mI46 pad_hv_n3 ng_pad_vpmp_h mid1 mid1 nhv m=4 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI35 mid ng_pad_vpmp_h pad_hv_n1 mid nhv m=4 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 pad_hv_n0 ng_pad_vpmp_h mid mid nhv m=3 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI45 mid1 ng_pad_vpmp_h pad_hv_n2 mid1 nhv m=4 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI28 mid ng_amx_vpmp_h amuxbus_hv mid nhv m=7 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI57 mid1 nmid_vccd net79 vssa nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI47 mid1 ng_amx_vpmp_h amuxbus_hv mid1 nhv m=7 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI78<1> mid pd_h_vdda vssa net043<0> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI78<0> mid1 pd_h_vdda vssa net043<1> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI77<1> mid pd_h_vddio vssa net044<0> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI77<0> mid1 pd_h_vddio vssa net044<1> nhv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 mid nmid_vccd net77 vssa nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI26 mid pg_amx_vdda_h_n amuxbus_hv vdda phv m=5 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI22 mid pg_pad_vddioq_h_n pad_hv_p1 vddio phv m=3 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 mid pg_pad_vddioq_h_n pad_hv_p0 vddio phv m=3 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amx_pucsd_inv A Y vda vssa
*.PININFO A:I vda:I vssa:I Y:O
XICEA A / icecap
XICEY Y / icecap
mI75 Y A vssa vssa nhv m=7 w=0.42 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
mI74 Y A vda vda phv m=7 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_drvr amux_en_vdda_h amux_en_vdda_h_n 
+ amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n 
+ amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n nga_amx_vswitch_h 
+ nga_pad_vswitch_h nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h 
+ ngb_pad_vswitch_h_n nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd 
+ nmidb_vccd_n pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n 
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
+ pu_csd_vddioq_h_n pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch
*.PININFO amux_en_vdda_h:I amux_en_vdda_h_n:I amux_en_vddio_h:I 
*.PININFO amux_en_vddio_h_n:I amux_en_vswitch_h:I amux_en_vswitch_h_n:I 
*.PININFO amuxbusa_on:I amuxbusa_on_n:I amuxbusb_on:I amuxbusb_on_n:I 
*.PININFO nmida_on_n:I nmidb_on_n:I pd_on:I pd_on_n:I pu_on:I pu_on_n:I vccd:I 
*.PININFO vdda:I vddio_q:I vssa:I vssd:I vswitch:I nga_amx_vswitch_h:O 
*.PININFO nga_pad_vswitch_h:O nga_pad_vswitch_h_n:O ngb_amx_vswitch_h:O 
*.PININFO ngb_pad_vswitch_h:O ngb_pad_vswitch_h_n:O nmida_vccd:O 
*.PININFO nmida_vccd_n:O nmidb_vccd:O nmidb_vccd_n:O pd_csd_vswitch_h:O 
*.PININFO pd_csd_vswitch_h_n:O pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O 
*.PININFO pgb_amx_vdda_h_n:O pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
XICEnmidb_vccd nmidb_vccd / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
XICEpu_on_n pu_on_n / icecap
XICEnet272 net272 / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEpd_on_n pd_on_n / icecap
XICEnet236 net236 / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
XICEnet239 net239 / icecap
XICEnet256 net256 / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEpu_on pu_on / icecap
XICEnet265 net265 / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEnet274 net274 / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEnet254 net254 / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
XICEnet275 net275 / icecap
XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEnet248 net248 / icecap
XICEnet257 net257 / icecap
XICEpd_on pd_on / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEnet230 net230 / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEnet245 net245 / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XI93 nmida_vccd nmida_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
XI105 nmidb_vccd nmidb_vccd_n vssd vccd / sky130_fd_io__hvsbt_inv_x1
XI38 net274 pu_csd_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_pucsd_inv
Xpga_amx_ls net265 net272 pga_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h 
+ vssa vdda / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI103 net239 net245 pgb_amx_vdda_h_n amux_en_vdda_h_n amux_en_vdda_h vssa vdda 
+ / sky130_fd_io__gpiov2_amux_drvr_lshv2hv
XI45 net256 nga_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI42 net265 pga_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI47 net256 nga_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI62 net239 pgb_pad_vddioq_h_n vddio_q vssd / sky130_fd_io__gpiov2_amx_inv4
XI63 net236 ngb_amx_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI64 net236 ngb_pad_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_inv4
XI53 nmidb_on_n nmidb_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
XI89 nmida_on_n nmida_vccd vssd vccd / sky130_fd_io__hvsbt_inv_x2
Xpdcsd_inv net254 pd_csd_vswitch_h vswitch vssa / sky130_fd_io__gpiov2_amx_pdcsd_inv
XI90 pd_csd_vswitch_h pd_csd_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI85 ngb_pad_vswitch_h ngb_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
XI87 nga_pad_vswitch_h nga_pad_vswitch_h_n vswitch vssa / sky130_fd_io__amx_inv1
mI76 ngb_amx_vswitch_h amux_en_vdda_h_n vssa vssa nhv m=1 w=1.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI77 ngb_pad_vswitch_h amux_en_vddio_h_n vssa vssa nhv m=1 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI75 nga_amx_vswitch_h amux_en_vdda_h_n vssa vssa nhv m=1 w=1.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI78 nga_pad_vswitch_h amux_en_vddio_h_n vssa vssa nhv m=1 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI104 pd_csd_vswitch_h amux_en_vddio_h_n vssa vssa nhv m=1 w=1.00 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xpu_csd_ls pu_on pu_on_n net274 net275 amux_en_vddio_h_n amux_en_vddio_h vssd 
+ vddio_q vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpga_pad_ls amuxbusa_on amuxbusa_on_n net265 net272 amux_en_vddio_h_n 
+ amux_en_vddio_h vssd vddio_q vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xnga_ls amuxbusa_on amuxbusa_on_n net257 net256 amux_en_vswitch_h_n 
+ amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpd_csd_ls pd_on pd_on_n net248 net254 amux_en_vswitch_h_n amux_en_vswitch_h 
+ vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xpgb_pad_ls amuxbusb_on amuxbusb_on_n net239 net245 amux_en_vddio_h_n 
+ amux_en_vddio_h vssd vddio_q vccd / sky130_fd_io__gpiov2_amux_drvr_ls
Xngb_ls amuxbusb_on amuxbusb_on_n net230 net236 amux_en_vswitch_h_n 
+ amux_en_vswitch_h vssa vswitch vccd / sky130_fd_io__gpiov2_amux_drvr_ls
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_ls in in_b out_h out_h_n rst_h rst_h_n vgnd 
+ vpwr_hv vpwr_lv
*.PININFO in:I in_b:I rst_h:I rst_h_n:I vgnd:I vpwr_hv:I vpwr_lv:I out_h:O 
*.PININFO out_h_n:O
XICEout_h out_h / icecap
XICEout_h_n out_h_n / icecap
XICEnet61 net61 / icecap
XICEfbk_n fbk_n / icecap
XICEfbk fbk / icecap
XICEin_b in_b / icecap
XICErst_h rst_h / icecap
XICEnet66 net66 / icecap
XICEnet62 net62 / icecap
XICEin in / icecap
XICErst_h_n rst_h_n / icecap
mI14 out_h fbk_n vpwr_hv vpwr_hv phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI11 out_h_n fbk vpwr_hv vpwr_hv phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 fbk_n fbk vpwr_hv vpwr_hv phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 fbk fbk_n vpwr_hv vpwr_hv phv m=1 w=0.75 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 net61 rst_h_n vgnd vgnd nhv m=4 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 out_h fbk_n vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 out_h_n fbk vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI58 fbk vpwr_lv net62 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnrst fbk rst_h vgnd vgnd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI59 fbk_n vpwr_lv net66 vgnd nhvnative m=4 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 net66 in net61 vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 net62 in_b net61 vgnd nlowvt m=4 w=1.00 l=0.15 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ls amux_en_vdda_h amux_en_vdda_h_n 
+ amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n 
+ analog_en enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n 
+ vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I enable_vdda_h:I enable_vswitch_h:I hld_i_h:I hld_i_h_n:I 
*.PININFO vccd:I vdda:I vddio_q:I vssa:I vssd:I vswitch:I amux_en_vdda_h:O 
*.PININFO amux_en_vdda_h_n:O amux_en_vddio_h:O amux_en_vddio_h_n:O 
*.PININFO amux_en_vswitch_h:O amux_en_vswitch_h_n:O enable_vdda_h_n:O
XICEanalog_en analog_en / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEana_en_i_n ana_en_i_n / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEhld_i_h hld_i_h / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEana_en_i ana_en_i / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
XICEnet74 net74 / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XI32 enable_vdda_h enable_vdda_h_n vssa vdda / sky130_fd_io__gpiov2_amux_ls_inv_x1
Xpd_vswitch_ls amux_en_vddio_h amux_en_vddio_h_n amux_en_vswitch_h 
+ amux_en_vswitch_h_n net74 enable_vswitch_h vssa vswitch / 
+ sky130_fd_io__gpiov2_amux_ctl_lshv2hv
Xpd_vdda_ls amux_en_vddio_h amux_en_vddio_h_n amux_en_vdda_h amux_en_vdda_h_n 
+ enable_vdda_h_n enable_vdda_h vssa vdda / sky130_fd_io__gpiov2_amux_ctl_lshv2hv
XI15 analog_en ana_en_i_n vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI16 ana_en_i_n ana_en_i vssd vccd / sky130_fd_io__gpiov2_amux_ctl_inv_1
XI18 enable_vswitch_h net74 vssa vswitch / sky130_fd_io__hvsbt_inv_x1
Xpd_vddio_ls ana_en_i ana_en_i_n amux_en_vddio_h amux_en_vddio_h_n hld_i_h 
+ hld_i_h_n vssd vddio_q vccd / sky130_fd_io__gpiov2_amux_ctl_ls
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux_ctl_logic analog_en analog_pol analog_sel 
+ enable_vdda_h enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n 
+ nga_amx_vswitch_h nga_pad_vswitch_h ngb_amx_vswitch_h ngb_pad_vswitch_h 
+ nmida_vccd nmidb_vccd out pd_csd_vswitch_h pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n 
+ vccd vdda vddio_q vssa vssd vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
*.PININFO enable_vswitch_h:I hld_i_h:I hld_i_h_n:I out:I vccd:I vdda:I 
*.PININFO vddio_q:I vssa:I vssd:I vswitch:I enable_vdda_h_n:O 
*.PININFO nga_amx_vswitch_h:O nga_pad_vswitch_h:O ngb_amx_vswitch_h:O 
*.PININFO ngb_pad_vswitch_h:O nmida_vccd:O nmidb_vccd:O pd_csd_vswitch_h:O 
*.PININFO pga_amx_vdda_h_n:O pga_pad_vddioq_h_n:O pgb_amx_vdda_h_n:O 
*.PININFO pgb_pad_vddioq_h_n:O pu_csd_vddioq_h_n:O
XICEngb_pad_vswitch_h_n ngb_pad_vswitch_h_n / icecap
XICEnga_pad_vswitch_h nga_pad_vswitch_h / icecap
XICEnmida_vccd_n nmida_vccd_n / icecap
XICEanalog_pol analog_pol / icecap
XICEamux_en_vswitch_h_n amux_en_vswitch_h_n / icecap
XICEnga_pad_vswitch_h_n nga_pad_vswitch_h_n / icecap
XICEamux_en_vddio_h amux_en_vddio_h / icecap
XICEngb_pad_vswitch_h ngb_pad_vswitch_h / icecap
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEamuxbusa_on_n amuxbusa_on_n / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEpd_on_n pd_on_n / icecap
XICEanalog_en analog_en / icecap
XICEngb_amx_vswitch_h ngb_amx_vswitch_h / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEamuxbusb_on_n amuxbusb_on_n / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEamux_en_vswitch_h amux_en_vswitch_h / icecap
XICEhld_i_h hld_i_h / icecap
XICEnmida_on_n nmida_on_n / icecap
XICEamuxbusa_on amuxbusa_on / icecap
XICEout out / icecap
XICEnga_amx_vswitch_h nga_amx_vswitch_h / icecap
XICEpd_csd_vswitch_h_n pd_csd_vswitch_h_n / icecap
XICEpu_on_n pu_on_n / icecap
XICEnmidb_on_n nmidb_on_n / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEpd_on pd_on / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEnmidb_vccd_n nmidb_vccd_n / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEamux_en_vddio_h_n amux_en_vddio_h_n / icecap
XICEamuxbusb_on amuxbusb_on / icecap
XICEpu_on pu_on / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEamux_en_vdda_h_n amux_en_vdda_h_n / icecap
XICEamux_en_vdda_h amux_en_vdda_h / icecap
XICEanalog_sel analog_sel / icecap
Xamux_sw_drvr amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h 
+ amux_en_vddio_h_n amux_en_vswitch_h amux_en_vswitch_h_n amuxbusa_on 
+ amuxbusa_on_n amuxbusb_on amuxbusb_on_n nga_amx_vswitch_h nga_pad_vswitch_h 
+ nga_pad_vswitch_h_n ngb_amx_vswitch_h ngb_pad_vswitch_h ngb_pad_vswitch_h_n 
+ nmida_on_n nmida_vccd nmida_vccd_n nmidb_on_n nmidb_vccd nmidb_vccd_n 
+ pd_csd_vswitch_h pd_csd_vswitch_h_n pd_on pd_on_n pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_csd_vddioq_h_n 
+ pu_on pu_on_n vccd vdda vddio_q vssa vssd vswitch / sky130_fd_io__gpiov2_amux_drvr
Xamux_lv_decoder amuxbusa_on amuxbusa_on_n amuxbusb_on amuxbusb_on_n analog_en 
+ analog_pol analog_sel nga_pad_vswitch_h nga_pad_vswitch_h_n 
+ ngb_pad_vswitch_h ngb_pad_vswitch_h_n nmida_on_n nmida_vccd_n nmidb_on_n 
+ nmidb_vccd_n out pd_on pd_on_n pd_csd_vswitch_h_n pga_amx_vdda_h_n 
+ pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n pu_on pu_on_n 
+ pu_csd_vddioq_h_n vccd vssd / sky130_fd_io__gpiov2_amux_decoder
Xamux_ls amux_en_vdda_h amux_en_vdda_h_n amux_en_vddio_h amux_en_vddio_h_n 
+ amux_en_vswitch_h amux_en_vswitch_h_n analog_en enable_vdda_h 
+ enable_vdda_h_n enable_vswitch_h hld_i_h hld_i_h_n vccd vdda vddio_q vssa 
+ vssd vswitch / sky130_fd_io__gpiov2_amux_ls
.ENDS
.SUBCKT sky130_fd_io__gpiov2_amux amuxbus_a amuxbus_b analog_en analog_pol 
+ analog_sel enable_vdda_h enable_vswitch_h hld_i_h hld_i_h_n out pad vccd 
+ vdda vddio_q vssa vssd vssio_q vswitch
*.PININFO analog_en:I analog_pol:I analog_sel:I enable_vdda_h:I 
*.PININFO enable_vswitch_h:I hld_i_h:I hld_i_h_n:I out:I vccd:I vdda:I 
*.PININFO vddio_q:I vssa:I vssd:I vssio_q:I vswitch:I amuxbus_a:B amuxbus_b:B 
*.PININFO pad:B
XICEnet168 net168 / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEamuxbus_a amuxbus_a / icecap
XICEnet101 net101 / icecap
XICEpga_pad_vddioq_h_n pga_pad_vddioq_h_n / icecap
XICEanalog_pol analog_pol / icecap
XICEpgb_pad_vddioq_h_n pgb_pad_vddioq_h_n / icecap
XICEnet0127 net0127 / icecap
XICEnet166 net166 / icecap
XICEnmidb_vccd nmidb_vccd / icecap
XICEanalog_en analog_en / icecap
XICEnet99 net99 / icecap
XICEenable_vdda_h enable_vdda_h / icecap
XICEnet85 net85 / icecap
XICEpgb_amx_vdda_h_n pgb_amx_vdda_h_n / icecap
XICEpga_amx_vdda_h_n pga_amx_vdda_h_n / icecap
XICEenable_vswitch_h enable_vswitch_h / icecap
XICEpad pad / icecap
XICEanalog_sel analog_sel / icecap
XICEnet97 net97 / icecap
XICEamuxbus_b amuxbus_b / icecap
XICEnga_amx_vpmp_h nga_amx_vpmp_h / icecap
XICEnet81 net81 / icecap
XICEpd_csd_vswitch_h pd_csd_vswitch_h / icecap
XICEout out / icecap
XICEnet100 net100 / icecap
XICEpu_csd_vddioq_h_n pu_csd_vddioq_h_n / icecap
XICEnga_pad_vpmp_h nga_pad_vpmp_h / icecap
XICEnmida_vccd nmida_vccd / icecap
XICEngb_pad_vpmp_h ngb_pad_vpmp_h / icecap
XICEhld_i_h hld_i_h / icecap
XICEngb_amx_vpmp_h ngb_amx_vpmp_h / icecap
xI43 vssio_q vdda condiode
xI78 vssa vswitch condiode
mI52 net81 pu_csd_vddioq_h_n vddio_q vddio_q phv m=3 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMP_PU net85 pu_csd_vddioq_h_n vddio_q vddio_q phv m=4 w=15.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI49 net81 pd_csd_vswitch_h vssio_q vssio_q nhv m=6 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mMN_PD net85 pd_csd_vswitch_h vssio_q vssio_q nhv m=8 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xmux_a amuxbus_a nga_amx_vpmp_h nga_pad_vpmp_h nmida_vccd net101 net101 net97 
+ net97 net100 net99 net0127 hld_i_h pga_amx_vdda_h_n pga_pad_vddioq_h_n vdda 
+ vddio_q vssa vssd / sky130_fd_io__gpiov2_amux_switch
Xmux_b amuxbus_b ngb_amx_vpmp_h ngb_pad_vpmp_h nmidb_vccd net101 net101 net97 
+ net97 net100 net99 net0127 hld_i_h pgb_amx_vdda_h_n pgb_pad_vddioq_h_n vdda 
+ vddio_q vssa vssd / sky130_fd_io__gpiov2_amux_switch
XBBM_logic analog_en analog_pol analog_sel enable_vdda_h net0127 
+ enable_vswitch_h hld_i_h hld_i_h_n nga_amx_vpmp_h nga_pad_vpmp_h 
+ ngb_amx_vpmp_h ngb_pad_vpmp_h nmida_vccd nmidb_vccd out pd_csd_vswitch_h 
+ pga_amx_vdda_h_n pga_pad_vddioq_h_n pgb_amx_vdda_h_n pgb_pad_vddioq_h_n 
+ pu_csd_vddioq_h_n vccd vdda vddio_q vssa vssd vswitch / 
+ sky130_fd_io__gpiov2_amux_ctl_logic
XI26 pad net99 / s8_esd_res75only_small
XI58 net168 net97 / s8_esd_res75only_small
XI28 net166 net101 / s8_esd_res75only_small
XI57 pad net168 / s8_esd_res75only_small
XI27 pad net100 / s8_esd_res75only_small
XI55 pad pad / s8_esd_res75only_small
XI54 pad net166 / s8_esd_res75only_small
XI53 pad pad / s8_esd_res75only_small
XI39 pad net81 / s8_esd_res75only_small
XI40 pad net85 / s8_esd_res75only_small
.ENDS
.SUBCKT sky130_fd_io__com_pddrvr_unit_2_5 nd ngin ns
*.PININFO ngin:I nd:B ns:B
XICEngin ngin / icecap
XICEnet10 ngin / icecap
XICEnd nd / icecap
mndrv nd ngin ns ns nhv m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_pddrvr_strong pad pd_h<3> pd_h<2> pd_h_i2c tie_lo_esd 
+ vcc_io vgnd_io
*.PININFO pd_h<3>:I pd_h<2>:I pd_h_i2c:I vcc_io:I vgnd_io:I pad:O tie_lo_esd:O
XICEpd_h<2> pd_h<2> / icecap
XICEpad pad / icecap
XICEpd_h<3> pd_h<3> / icecap
XICEnet78 net78 / icecap
XICEnet80 net80 / icecap
XICEpd_h_i2c pd_h_i2c / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XICEnet66 net66 / icecap
XICEnet76 net76 / icecap
XICEnet68 net68 / icecap
XICEnet72 net72 / icecap
XICEnet46 net46 / icecap
XI97 pd_h<3> net80 / sky130_fd_io__tk_em2s
XI108 pd_h<3> net78 / sky130_fd_io__tk_em2s
XI109 tie_lo_esd net76 / sky130_fd_io__tk_em2s
XI102 pd_h<3> net72 / sky130_fd_io__tk_em2s
XI104 pd_h<3> net68 / sky130_fd_io__tk_em2s
XI96 pd_h<3> net66 / sky130_fd_io__tk_em2s
XI113 pd_h<2> net46 / sky130_fd_io__tk_em2s
XI99 tie_lo_esd net80 / sky130_fd_io__tk_em2o
XI98 pd_h<2> net80 / sky130_fd_io__tk_em2o
XI106 pd_h<2> net78 / sky130_fd_io__tk_em2o
XI107 tie_lo_esd net78 / sky130_fd_io__tk_em2o
XI110 pd_h<3> net76 / sky130_fd_io__tk_em2o
XI111 pd_h<2> net76 / sky130_fd_io__tk_em2o
XI100 tie_lo_esd net72 / sky130_fd_io__tk_em2o
XI101 pd_h<2> net72 / sky130_fd_io__tk_em2o
XI103 tie_lo_esd net68 / sky130_fd_io__tk_em2o
XI105 pd_h<2> net68 / sky130_fd_io__tk_em2o
XI95 pd_h<2> net66 / sky130_fd_io__tk_em2o
XI94 tie_lo_esd net66 / sky130_fd_io__tk_em2o
XI88 pd_h<3> net46 / sky130_fd_io__tk_em2o
XI87 tie_lo_esd net46 / sky130_fd_io__tk_em2o
XI49 vgnd_io tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
Xn24<2> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0> pad net80 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0> pad net66 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn12 pad pd_h_i2c vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0> pad net68 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0> pad net78 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0> pad net76 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn13 pad net46 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn31 pad net72 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
xI72 vgnd_io vcc_io condiode
.ENDS
.SUBCKT sky130_fd_io__gpio_pudrvr_unit_2_5 pd pgin ps
*.PININFO pgin:I pd:B ps:B
XICEnet10 pgin / icecap
XICEpgin pgin / icecap
XICEpd pd / icecap
mpdrv pd pgin ps ps phv m=2 w=5.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 
+ topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_pudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io 
+ vnb
*.PININFO pu_h_n<3>:I pu_h_n<2>:I vcc_io:I vnb:I pad:O tie_hi_esd:O
XI112 pu_h_n<2> net43 / sky130_fd_io__tk_em2s
XI108 tie_hi_esd net59 / sky130_fd_io__tk_em2s
XI109 tie_hi_esd net53 / sky130_fd_io__tk_em2s
XI104 pu_h_n<3> net49 / sky130_fd_io__tk_em2s
XI125 pu_h_n<3> net45 / sky130_fd_io__tk_em2s
XI83 pu_h_n<3> net43 / sky130_fd_io__tk_em2o
XI82 tie_hi_esd net43 / sky130_fd_io__tk_em2o
XI106 pu_h_n<2> net59 / sky130_fd_io__tk_em2o
XI107 pu_h_n<3> net59 / sky130_fd_io__tk_em2o
XI110 pu_h_n<3> net53 / sky130_fd_io__tk_em2o
XI111 pu_h_n<2> net53 / sky130_fd_io__tk_em2o
XI103 tie_hi_esd net49 / sky130_fd_io__tk_em2o
XI105 pu_h_n<2> net49 / sky130_fd_io__tk_em2o
XI124 tie_hi_esd net45 / sky130_fd_io__tk_em2o
XI123 pu_h_n<2> net45 / sky130_fd_io__tk_em2o
XI49 vcc_io tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
Xn24<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn24<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn23<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn22 pad net45 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn21 pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<2> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<1> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn12<0> pad net43 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<2> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<1> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn32<0> pad net49 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<1> pad net59 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn33<0> pad net59 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<2> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<1> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn34<0> pad net53 vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<2> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<1> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn11<0> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<2> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<1> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn13<0> pad pu_h_n<2> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<2> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<1> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
Xn31<0> pad pu_h_n<3> vcc_io / sky130_fd_io__gpio_pudrvr_unit_2_5
.ENDS
.SUBCKT sky130_fd_io__com_pudrvr_weak pad pu_h_n vcc_io vgnd_io vpb_drvr
*.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
XICEpad pad / icecap
XICEpu_h_n pu_h_n / icecap
mpdrv pad pu_h_n vcc_io vpb_drvr phv m=4 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI29 pad pu_h_n vcc_io vpb_drvr phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_pudrvr_strong_slow pad pu_h_n vcc_io vgnd_io vpb_drvr
*.PININFO pu_h_n:I vcc_io:I vgnd_io:I vpb_drvr:I pad:O
XICEpu_h_n pu_h_n / icecap
XICEpad pad / icecap
mpdrv pad pu_h_n vcc_io vpb_drvr phv m=8 w=7.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_odrvr_sub force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> 
+ pd_h<0> pd_h_i2c pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd 
+ tie_lo_esd vcc_io vgnd vgnd_io
*.PININFO force_hi_h_n:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pd_h_i2c:I 
*.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I pad:O tie_hi_esd:B tie_lo_esd:B
XICEpad pad / icecap
XICEpu_h_n<0> pu_h_n<0> / icecap
XICEpad_r250 pad_r250 / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XICEweak_pad weak_pad / icecap
XI75<0> pu_h_n<3> / icecap
XI75<1> pu_h_n<2> / icecap
XICEvgnd vgnd / icecap
XI74<0> pd_h<3> / icecap
XI74<1> pd_h<2> / icecap
XICEpu_h_n<1> pu_h_n<1> / icecap
XICEpd_h<1> pd_h<1> / icecap
XICEpd_h_i2c pd_h_i2c / icecap
XICEforce_hi_h_n force_hi_h_n / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XICEstrong_slow_pad strong_slow_pad / icecap
XICEpd_h<0> pd_h<0> / icecap
Xpddrvr_strong pad pd_h<3> pd_h<2> pd_h_i2c tie_lo_esd vcc_io vgnd_io / 
+ sky130_fd_io__gpiov2_pddrvr_strong
Xpudrvr_strong pad pu_h_n<3> pu_h_n<2> tie_hi_esd vcc_io vgnd / 
+ sky130_fd_io__gpio_pudrvr_strong
Xpudrvr_weak weak_pad pu_h_n<0> vcc_io vgnd vcc_io / sky130_fd_io__com_pudrvr_weak
Xpddrvr_weak weak_pad pd_h<0> vcc_io vgnd_io / sky130_fd_io__gpio_pddrvr_weak
Xstrong_slow_pddrvr strong_slow_pad pd_h<1> vcc_io vgnd_io / 
+ sky130_fd_io__gpio_pddrvr_strong_slow
Xstrong_slow_pudrvr strong_slow_pad pu_h_n<1> vcc_io vgnd vcc_io / 
+ sky130_fd_io__com_pudrvr_strong_slow
Xres strong_slow_pad pad_r250 vgnd_io / sky130_fd_io__com_res_strong_slow
Xres_weak weak_pad pad_r250 vgnd_io / sky130_fd_io__com_res_weak
Xresd pad pad_r250 / s8_esd_res250only_small
xI60 vgnd_io vcc_io condiode
xI59 vgnd_io vcc_io condiode
xI58 vgnd_io vcc_io condiode
xI72 vgnd_io vcc_io condiode
.ENDS
.SUBCKT sky130_fd_io__gpiov2_odrvr force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pd_h_i2c pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd 
+ vcc_io vgnd vgnd_io
*.PININFO force_hi_h_n:I pd_h<3>:I pd_h<2>:I pd_h<1>:I pd_h<0>:I pd_h_i2c:I 
*.PININFO pu_h_n<3>:I pu_h_n<2>:I pu_h_n<1>:I pu_h_n<0>:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I pad:O tie_hi_esd:O tie_lo_esd:O
Xodrvr force_hi_h_n pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h_i2c pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io / 
+ sky130_fd_io__gpiov2_odrvr_sub
Xbondpad pad vgnd_io / sky130_fd_io__com_pad
.ENDS
.SUBCKT sky130_fd_io__com_cclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io 
+ vgnd
*.PININFO oe_h_n:I pd_dis_h:I pu_dis_h:I vcc_io:I vgnd:I drvhi_h:O drvlo_h_n:O
XICEpu_dis_h_n pu_dis_h_n / icecap
XICEn0 n0 / icecap
XICEn1 n1 / icecap
XICEoe_i_h_n oe_i_h_n / icecap
XICEpu_dis_h pu_dis_h / icecap
XICEoe_h_n oe_h_n / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEoe_i_h oe_i_h / icecap
XICEpd_dis_h pd_dis_h / icecap
XICEdrvhi_h drvhi_h / icecap
Xnor3 oe_i_h_n drvhi_h pd_dis_h n1 vcc_io vgnd vgnd / sky130_fd_io__com_cclat_hvnor3
Xnand3 oe_i_h drvlo_h_n pu_dis_h_n n0 vcc_io vgnd vgnd / 
+ sky130_fd_io__com_cclat_hvnand3
Xinv_oe1 oe_h_n oe_i_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_oe2 oe_i_h oe_i_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_pudis pu_dis_h pu_dis_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_in
Xinv_out n1 drvlo_h_n vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
Xinv_out_1 n0 drvhi_h vcc_io vgnd vgnd / sky130_fd_io__com_cclat_inv_out
.ENDS
.SUBCKT sky130_fd_io__gpiov2_opath_datoe drvhi_h drvlo_h_n hld_h_n hld_i_ovr_h od_h 
+ oe_h oe_n out vcc_io vgnd vpwr_ka
*.PININFO hld_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I vcc_io:I vgnd:I 
*.PININFO vpwr_ka:I drvhi_h:O drvlo_h_n:O oe_h:O
XICEhld_h_n hld_h_n / icecap
XICEdrvhi_h drvhi_h / icecap
XICEout out / icecap
XICEod_h od_h / icecap
XICEoe_n oe_n / icecap
XICEoe_h oe_h / icecap
XICEoe_h_n oe_h_n / icecap
XICEpd_dis_h pd_dis_h / icecap
XICEpu_dis_h pu_dis_h / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
Xdat_ls hld_i_ovr_h out pd_dis_h pu_dis_h vgnd od_h vcc_io vgnd vpwr_ka / 
+ sky130_fd_io__gpio_dat_ls
Xoe_ls hld_i_ovr_h oe_n oe_h_n oe_h vgnd od_h vcc_io vgnd vpwr_ka / 
+ sky130_fd_io__gpio_dat_ls
Xcclat drvhi_h drvlo_h_n oe_h_n pd_dis_h pu_dis_h vcc_io vgnd / 
+ sky130_fd_io__com_cclat
.ENDS
.SUBCKT sky130_fd_io__gpiov2_octl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n od_h pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h 
+ puen_2or1_h puen_h<1> puen_h<0> slow slow_h slow_h_n vcc_io vgnd vpwr 
+ vreg_en_h_n
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I od_h:I slow:I vcc_io:I vgnd:I vpwr:I vreg_en_h_n:I 
*.PININFO pden_h_n<2>:O pden_h_n<1>:O pden_h_n<0>:O puen_0_h:O puen_2or1_h:O 
*.PININFO puen_h<1>:O puen_h<0>:O slow_h:O slow_h_n:O
XICEn<5> n<5> / icecap
XICEpuen_h<1> puen_h<1> / icecap
XICEod_h od_h / icecap
XICEvreg_en_h_n vreg_en_h_n / icecap
XICEn<4> n<4> / icecap
XICEpden_h0 pden_h0 / icecap
XICEn<1> n<1> / icecap
XICEn<2> n<2> / icecap
XICEdm_h_n<0> dm_h_n<0> / icecap
XICEpuen_h1_n puen_h1_n / icecap
XICEn<3> n<3> / icecap
XICEdm_h_n<2> dm_h_n<2> / icecap
XICEnet70 net70 / icecap
XICEpden_h_n<0> pden_h_n<0> / icecap
XICEslow_h slow_h / icecap
XICEslow slow / icecap
XICEpuen_h0_n puen_h0_n / icecap
XICEslow_h_n slow_h_n / icecap
XICEn<9> n<9> / icecap
XICEpuen_0_h puen_0_h / icecap
XICEpuen_2or1_h puen_2or1_h / icecap
XICEn<0> n<0> / icecap
XICEn<8> n<8> / icecap
XICEdm_h_n<1> dm_h_n<1> / icecap
XICEdm_h<1> dm_h<1> / icecap
XICEdm_h<2> dm_h<2> / icecap
XICEpden_h_n<2> pden_h_n<2> / icecap
XICEdm_h<0> dm_h<0> / icecap
XICEpuen_h<0> puen_h<0> / icecap
XICEnet130 net130 / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEn<10> n<10> / icecap
XICEpden_h1 pden_h1 / icecap
XI211 n<8> dm_h_n<1> puen_0_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI201 dm_h_n<2> dm_h_n<1> n<9> vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI381 dm_h<1> dm_h<0> net70 vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI210 dm_h<2> dm_h<0> n<8> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI200 dm_h<2> dm_h<1> n<10> vgnd vcc_io / sky130_fd_io__hvsbt_xor
XI185 dm_h_n<0> n<4> net130 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI186 dm_h_n<2> dm_h_n<1> n<4> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI187 dm_h<1> dm_h<0> n<3> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI208 puen_2or1_h vreg_en_h_n n<5> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI203 n<10> dm_h<0> n<1> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI204 n<9> dm_h_n<0> n<0> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI205 n<1> n<0> puen_2or1_h vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI382 dm_h<2> net70 pden_h_n<2> vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI254 puen_h1_n puen_h<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI256 puen_h0_n puen_h<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI249 pden_h0 pden_h_n<0> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI247 pden_h1 pden_h_n<1> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x2
XI377 puen_0_h puen_h0_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI209 n<5> n<2> vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI376 n<2> puen_h1_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI374 net130 pden_h1 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI375 n<3> pden_h0 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xls_slow hld_i_h_n slow slow_h slow_h_n od_h vgnd vcc_io vgnd vpwr / 
+ sky130_fd_io__com_ctl_ls
.ENDS
.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong_nd2 drvhi_h en_fast<3> en_fast<2> 
+ en_fast<1> en_fast<0> pu_h_n puen_h vcc_io vgnd_io
*.PININFO drvhi_h:I en_fast<3>:I en_fast<2>:I en_fast<1>:I en_fast<0>:I 
*.PININFO puen_h:I vcc_io:I vgnd_io:I pu_h_n:O
XICEpuen_h puen_h / icecap
XICEpu_h_n pu_h_n / icecap
XI134<0> en_fast<3> / icecap
XI134<1> en_fast<2> / icecap
XI134<2> en_fast<1> / icecap
XI134<3> en_fast<0> / icecap
XICEint_res int_res / icecap
XICEnet24 net24 / icecap
XICEdrvhi_h drvhi_h / icecap
XE1 net24 pu_h_n / sky130_fd_io__tk_em1s
rrespu1 int_res net24 mrp1 m=1 w=0.33 l=11
rrespu2 pu_h_n int_res mrp1 m=1 w=0.33 l=4
mmnin_fast<3> net24 drvhi_h int<3> net013<0> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<2> net24 drvhi_h int<2> net013<1> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<1> net24 drvhi_h int<1> net013<2> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_fast<0> net24 drvhi_h int<0> net013<3> nhv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_slow1 n<2> puen_h vgnd_io vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin_slow pu_h_n drvhi_h n<2> vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<3> int<3> en_fast<3> vgnd_io net014<0> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<2> int<2> en_fast<2> vgnd_io net014<1> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<1> int<1> en_fast<1> vgnd_io net014<2> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen_fast<0> int<0> en_fast<0> vgnd_io net014<3> nhv m=1 w=1.50 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen pu_h_n puen_h vcc_io vcc_io phv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin pu_h_n drvhi_h vcc_io vcc_io phv m=3 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_pupredrvr_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h 
+ slow_h_n vcc_io vgnd_io
*.PININFO drvhi_h:I puen_h:I slow_h_n:I vcc_io:I vgnd_io:I pu_h_n<3>:O 
*.PININFO pu_h_n<2>:O
Xnd2b drvhi_h en_fast_h_3<3> en_fast_h_3<2> en_fast_h_3<1> en_fast_h_3<0> 
+ pu_h_n<3> puen_h vcc_io vgnd_io / sky130_fd_io__gpiov2_pupredrvr_strong_nd2
Xnd2a drvhi_h net54 net54 net54 net54 pu_h_n<2> puen_h vcc_io vgnd_io / 
+ sky130_fd_io__gpiov2_pupredrvr_strong_nd2
XI98 en_fast_h_3<0> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI97 en_fast_h_3<1> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opti
XI92 en_fast_h_3<3> nbias_out en_fast_h / sky130_fd_io__tk_opto
XI96 en_fast_h_3<2> en_fast_h_3<3> vgnd_io / sky130_fd_io__tk_opto
XI93 net54 nbias_out en_fast_h / sky130_fd_io__tk_opto
Xinv en_fast_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xnbias drvhi_h en_fast_h en_fast_h_n nbias_out pu_h_n<2> puen_h vcc_io vgnd_io 
+ / sky130_fd_io__com_pupredrvr_nbias
Xnand puen_h slow_h_n en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_nand2_dnw
.ENDS
.SUBCKT sky130_fd_io__gpiov2_octl_mux a_h b_h sel_h sel_h_n vccio vssio y_h
*.PININFO a_h:I b_h:I sel_h:I sel_h_n:I vccio:I vssio:I y_h:O
XICEsel_h sel_h / icecap
XICEy_h y_h / icecap
XICEa_h a_h / icecap
XICEsel_h_n sel_h_n / icecap
XICEb_h b_h / icecap
mI2 y_h sel_h b_h vccio phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI3 y_h sel_h_n a_h vccio phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 b_h sel_h_n y_h vssio nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI4 a_h sel_h y_h vssio nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr2 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> i2c_mode_h pd_h pd_i2c_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I i2c_mode_h:I pden_h_n:I 
*.PININFO vcc_io:I vgnd_io:I pd_h:O pd_i2c_h:O
XICEpden_h_n pden_h_n / icecap
XI105<0> net53<0> / icecap
XI105<1> net53<1> / icecap
XICEnet62 net62 / icecap
XICEpd_i2c_h pd_i2c_h / icecap
XICEi2c_mode_h i2c_mode_h / icecap
XICEpd_h pd_h / icecap
XI104<0> en_fast_n<1> / icecap
XI104<1> en_fast_n<0> / icecap
XICEen_fast_n<1> en_fast_n<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEnet42 net42 / icecap
mmpin_slow pd_i2c_h drvlo_h_n int_slow vcc_io phv m=1 w=0.42 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_slow int_slow pden_h_n vcc_io vcc_io phv m=1 w=0.42 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<1> pd_i2c_h drvlo_h_n net62 net030<0> phv m=1 w=0.42 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<0> pd_i2c_h drvlo_h_n net62 net030<1> phv m=1 w=0.42 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast1 net62 en_fast_n<1> vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI72<1> net53<0> en_fast_n<1> net42 net031<0> phv m=1 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI72<0> net53<1> en_fast_n<0> net42 net031<1> phv m=1 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI74<1> pd_h drvlo_h_n net53<0> net032<0> phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI74<0> pd_h drvlo_h_n net53<1> net032<1> phv m=2 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI75 net039 pden_h_n net42 vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI76 pd_h drvlo_h_n net45 vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI73 net42 i2c_mode_h vcc_io vcc_io phv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI101 net45 pden_h_n net039 vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI94 pd_h i2c_mode_h vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin pd_i2c_h drvlo_h_n vgnd_io vgnd_io nhv m=2 w=3.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen pd_i2c_h pden_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI78 pd_h pden_h_n vgnd_io vgnd_io nhv m=1 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI77 pd_h drvlo_h_n vgnd_io vgnd_io nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong_nr3 drvlo_h_n en_fast_n<1> 
+ en_fast_n<0> i2c_mode_h pd_h pden_h_n vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_fast_n<1>:I en_fast_n<0>:I i2c_mode_h:I pden_h_n:I 
*.PININFO vcc_io:I vgnd_io:I pd_h:O
XI110<0> en_fast_n<1> / icecap
XI110<1> en_fast_n<0> / icecap
XICEint1 int1 / icecap
XICEpden_h_n pden_h_n / icecap
XICEpd_h pd_h / icecap
XICEi2c_mode_h i2c_mode_h / icecap
XICEint2 int2 / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
mI85 int1 i2c_mode_h vcc_io vcc_io phv m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_slow pd_h drvlo_h_n int_slow vcc_io phv m=1 w=0.42 l=2.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_slow int_slow pden_h_n vcc_io vcc_io phv m=1 w=0.42 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<1> pd_h drvlo_h_n int_nor<1> vcc_io phv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpin_fast<0> pd_h drvlo_h_n int_nor<0> vcc_io phv m=1 w=1.50 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast<1> int_nor<1> en_fast_n<1> vcc_io vcc_io phv m=1 w=1.50 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmpen_fast<0> int_nor<0> en_fast_n<0> vcc_io vcc_io phv m=1 w=1.50 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI90 pd_h drvlo_h_n net43 vcc_io phv m=1 w=0.42 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI56 net43 pden_h_n int1 vcc_io phv m=1 w=0.42 l=2.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI87<1> pd_h drvlo_h_n int2 vcc_io phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI87<0> pd_h drvlo_h_n int2 vcc_io phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI86<1> int2 en_fast_n<1> int1 vcc_io phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI86<0> int2 en_fast_n<0> int1 vcc_io phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnin pd_h drvlo_h_n vgnd_io vgnd_io nhv m=5 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mmnen pd_h pden_h_n vgnd_io vgnd_io nhv m=2 w=3.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__com_pdpredrvr_pbias drvlo_h_n en_h en_h_n pbias pd_h pden_h_n 
+ vcc_io vgnd_io
*.PININFO drvlo_h_n:I en_h:I en_h_n:I pd_h:I pden_h_n:I vcc_io:I vgnd_io:I 
*.PININFO pbias:O
XICEpbias pbias / icecap
XICEpden_h_n pden_h_n / icecap
XICEbias_g bias_g / icecap
XICEnet157 net157 / icecap
XICEnet108 net108 / icecap
XICEn<101> n<101> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEdrvlo_i_h drvlo_i_h / icecap
XICEen_h en_h / icecap
XICEpbias1 pbias1 / icecap
XICEnet84 net84 / icecap
XICEn<0> n<0> / icecap
XICEn<1> n<1> / icecap
XICE2vtp N0 / icecap
XICEen_h_n en_h_n / icecap
XICEpd_h pd_h / icecap
XICEnet88 net88 / icecap
XICEnet161 net161 / icecap
XI27 n<0> pd_h en_h_n / sky130_fd_io__tk_opto
XE1 n<1> n<0> / sky130_fd_io__tk_em1o
XE2 pbias pbias1 / sky130_fd_io__tk_em1o
XE3 pbias1 net88 / sky130_fd_io__tk_em1s
XE4 net108 pbias / sky130_fd_io__tk_em1s
XE6 pbias net84 / sky130_fd_io__tk_em1s
XE5 n<101> bias_g / sky130_fd_io__tk_em1s
mI47 pbias bias_g vgnd_io vgnd_io nhv m=2 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI24 n<1> drvlo_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI18 bias_g drvlo_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI23 n<0> n<0> n<1> vgnd_io nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI13 drvlo_i_h drvlo_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI20 bias_g n<1> vgnd_io vgnd_io nhv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI19 bias_g en_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI34 net157 bias_g vgnd_io vgnd_io nhv m=1 w=5.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI36 net108 bias_g vgnd_io vgnd_io nhv m=2 w=1.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI38 n<1> pden_h_n vgnd_io vgnd_io nhv m=1 w=1.00 l=0.60 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI48 n<100> pd_h vgnd_io vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI41 n<101> pd_h n<100> vgnd_io nhv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI44 pbias pbias pbias1 vcc_io phv m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI45 pbias1 pbias1 vcc_io vcc_io phv m=8 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI15 net183 en_h_n vcc_io vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI16 net171 n<0> net183 vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 pbias en_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI12 drvlo_i_h drvlo_h_n vcc_io vcc_io phv m=2 w=1.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI17 bias_g drvlo_h_n net171 vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 pbias drvlo_i_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI33 N0 vgnd_io vcc_io vcc_io phv m=1 w=0.42 l=8.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI32 net161 net161 N0 vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI31 net157 net157 net161 vcc_io phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI30 net88 N0 vcc_io vcc_io phv m=8 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI43 net84 bias_g vcc_io vcc_io phv m=1 w=0.42 l=4.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI40 N0 drvlo_i_h vcc_io vcc_io phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_pdpredrvr_strong drvlo_h_n i2c_mode_h_n pd_h<4> 
+ pd_h<3> pd_h<2> pden_h_n slow_h tie_hi_esd vcc_io vgnd vgnd_io
*.PININFO drvlo_h_n:I i2c_mode_h_n:I pden_h_n:I slow_h:I tie_hi_esd:I vcc_io:I 
*.PININFO vgnd:I vgnd_io:I pd_h<4>:O pd_h<3>:O pd_h<2>:O
XICEpd_h<2> pd_h<2> / icecap
XI162<0> en_fast2_n<1> / icecap
XI162<1> en_fast2_n<0> / icecap
XICEpden_h_n pden_h_n / icecap
XICEmod_drvlo_h_n mod_drvlo_h_n / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XICEnet142 net142 / icecap
XICEen_fast2_n<0> en_fast2_n<0> / icecap
XICEpd_h<3> pd_h<3> / icecap
XICEmod_slow_h mod_slow_h / icecap
XICEi2c_mode_h i2c_mode_h / icecap
XICEnet75 net75 / icecap
XICEen_fast_h_n en_fast_h_n / icecap
XICEen_fast2_n<1> en_fast2_n<1> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEslow_h slow_h / icecap
XICEen_fast_h en_fast_h / icecap
XI163<0> pbias_out / icecap
XI163<1> pbias_out / icecap
XICEint_slow1 int_slow1 / icecap
XICEpbias_out pbias_out / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEpd_h<4> pd_h<4> / icecap
XICEmod_drvlo_h_n_i2c mod_drvlo_h_n_i2c / icecap
XICEnet118 net118 / icecap
mI87 mod_drvlo_h_n_i2c pd_h<4> vcc_io vcc_io phv m=1 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI88 mod_drvlo_h_n_i2c pd_h<4> vgnd vgnd nhv m=1 w=0.42 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI160 i2c_mode_h_n slow_h net75 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI98 i2c_mode_h slow_h int_slow1 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI161 net75 net142 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI97 int_slow1 mod_slow_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI93 i2c_mode_h_n i2c_mode_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xmux mod_drvlo_h_n_i2c drvlo_h_n i2c_mode_h i2c_mode_h_n vcc_io vgnd_io 
+ mod_drvlo_h_n / sky130_fd_io__gpiov2_octl_mux
Xnr3 drvlo_h_n pbias_out pbias_out mod_slow_h pd_h<2> pd_h<4> pden_h_n vcc_io 
+ vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong_nr2
Xnr2 mod_drvlo_h_n en_fast2_n<1> en_fast2_n<0> mod_slow_h pd_h<3> pden_h_n 
+ vcc_io vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong_nr3
XI77 en_fast2_n<1> pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI76 net118 pbias_out en_fast_h_n / sky130_fd_io__tk_opto
XI79 en_fast2_n<0> en_fast2_n<1> vcc_io / sky130_fd_io__tk_opti
Xinv en_fast_h en_fast_h_n vgnd_io vcc_io / sky130_fd_io__com_inv_x1_dnw
Xbias drvlo_h_n en_fast_h en_fast_h_n pbias_out pd_h<4> pden_h_n vcc_io 
+ vgnd_io / sky130_fd_io__com_pdpredrvr_pbias
Xnor net142 pden_h_n en_fast_h vgnd_io vcc_io / sky130_fd_io__com_nor2_dnw
.ENDS
.SUBCKT sky130_fd_io__gpiov2_obpredrvr drvhi_h drvlo_h_n i2c_mode_h_n pd_h<4> 
+ pd_h<3> pd_h<2> pd_h<1> pd_h<0> pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> puen_h<1> puen_h<0> slow_h slow_h_n tie_hi_esd vcc_io 
+ vgnd vgnd_io
*.PININFO drvhi_h:I drvlo_h_n:I i2c_mode_h_n:I pden_h_n<1>:I pden_h_n<0>:I 
*.PININFO puen_h<1>:I puen_h<0>:I slow_h:I slow_h_n:I tie_hi_esd:I vcc_io:I 
*.PININFO vgnd:I vgnd_io:I pd_h<4>:O pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O 
*.PININFO pu_h_n<3>:O pu_h_n<2>:O pu_h_n<1>:O pu_h_n<0>:O
XICEtie_hi_esd tie_hi_esd / icecap
XICEpden_h_n<1> pden_h_n<1> / icecap
XICEpu_h_n<0> pu_h_n<0> / icecap
XICEpuen_h<1> puen_h<1> / icecap
XICEslow_h slow_h / icecap
XICEslow_h_n slow_h_n / icecap
XICEpden_h_n<0> pden_h_n<0> / icecap
XI125<0> pu_h_n<3> / icecap
XI125<1> pu_h_n<2> / icecap
XI126<0> pd_h<4> / icecap
XI126<1> pd_h<3> / icecap
XI126<2> pd_h<2> / icecap
XICEi2c_mode_h_n i2c_mode_h_n / icecap
XICEdrvhi_h drvhi_h / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XICEpu_h_n<1> pu_h_n<1> / icecap
XICEpd_h<1> pd_h<1> / icecap
XICEpuen_h<0> puen_h<0> / icecap
XICEpd_h<0> pd_h<0> / icecap
Xpu_strong drvhi_h pu_h_n<3> pu_h_n<2> puen_h<1> slow_h_n vcc_io vgnd_io / 
+ sky130_fd_io__gpiov2_pupredrvr_strong
Xpd_strong drvlo_h_n i2c_mode_h_n pd_h<4> pd_h<3> pd_h<2> pden_h_n<1> slow_h 
+ tie_hi_esd vcc_io vgnd vgnd_io / sky130_fd_io__gpiov2_pdpredrvr_strong
Xpu_weak drvhi_h pu_h_n<0> puen_h<0> vcc_io vgnd_io / 
+ sky130_fd_io__com_pupredrvr_weak
Xpd_weak drvlo_h_n pd_h<0> pden_h_n<0> vcc_io vgnd_io / 
+ sky130_fd_io__com_pdpredrvr_weak
Xpu_strong_slow drvhi_h pu_h_n<1> puen_h<1> vcc_io vgnd_io / 
+ sky130_fd_io__com_pupredrvr_strong_slow
Xpd_strong_slow drvlo_h_n pd_h<1> pden_h_n<1> vcc_io vgnd_io / 
+ sky130_fd_io__com_pdpredrvr_strong_slow
xI15 vgnd_io vcc_io condiode
.ENDS
.SUBCKT sky130_fd_io__gpiov2_octl_dat dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> drvhi_h hld_i_h_n hld_i_ovr_h od_h oe_n out pd_h<4> pd_h<3> 
+ pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> slow 
+ slow_h_n tie_hi_esd vcc_io vgnd vgnd_io vpwr vpwr_ka
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I tie_hi_esd:I 
*.PININFO vcc_io:I vgnd:I vgnd_io:I vpwr:I vpwr_ka:I drvhi_h:O pd_h<4>:O 
*.PININFO pd_h<3>:O pd_h<2>:O pd_h<1>:O pd_h<0>:O pu_h_n<3>:O pu_h_n<2>:O 
*.PININFO pu_h_n<1>:O pu_h_n<0>:O slow_h_n:O
XICEhld_i_h_n hld_i_h_n / icecap
XI204<0> pden_h_n<2> / icecap
XI204<1> pden_h_n<1> / icecap
XI204<2> pden_h_n<0> / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XI202<0> pd_h<4> / icecap
XI202<1> pd_h<3> / icecap
XI202<2> pd_h<2> / icecap
XI202<3> pd_h<1> / icecap
XI202<4> pd_h<0> / icecap
XICEdrvlo_h_n drvlo_h_n / icecap
XI200<0> pu_h_n<3> / icecap
XI200<1> pu_h_n<2> / icecap
XI200<2> pu_h_n<1> / icecap
XI200<3> pu_h_n<0> / icecap
XI203<0> pd_h<4> / icecap
XI203<1> pd_h<3> / icecap
XI203<2> pd_h<2> / icecap
XI203<3> pd_h<1> / icecap
XI203<4> pd_h<0> / icecap
XI205<0> pu_h_n<3> / icecap
XI205<1> pu_h_n<2> / icecap
XI205<2> pu_h_n<1> / icecap
XI205<3> pu_h_n<0> / icecap
XICEpuen_0_h puen_0_h / icecap
XI207<0> pden_h_n<1> / icecap
XI207<1> pden_h_n<0> / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XI201<0> dm_h_n<2> / icecap
XI201<1> dm_h_n<1> / icecap
XI201<2> dm_h_n<0> / icecap
XICEod_h od_h / icecap
XI206<0> puen_h<1> / icecap
XI206<1> puen_h<0> / icecap
XICEoe_n oe_n / icecap
XICEout out / icecap
XI199<0> dm_h<2> / icecap
XI199<1> dm_h<1> / icecap
XI199<2> dm_h<0> / icecap
XICEpden_h_n<2> pden_h_n<2> / icecap
XICEslow_h_n slow_h_n / icecap
XICEpuen_2or1_h puen_2or1_h / icecap
XICEslow_h slow_h / icecap
XICEdrvhi_h drvhi_h / icecap
XICEslow slow / icecap
XICEoe_h oe_h / icecap
Xdatoe drvhi_h drvlo_h_n hld_i_h_n hld_i_ovr_h od_h oe_h oe_n out vcc_io vgnd 
+ vpwr_ka / sky130_fd_io__gpiov2_opath_datoe
Xctl dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n od_h 
+ pden_h_n<2> pden_h_n<1> pden_h_n<0> puen_0_h puen_2or1_h puen_h<1> puen_h<0> 
+ slow slow_h slow_h_n vcc_io vgnd vpwr vcc_io / sky130_fd_io__gpiov2_octl
Xpredrvr drvhi_h drvlo_h_n pden_h_n<2> pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> 
+ pden_h_n<1> pden_h_n<0> pu_h_n<3> pu_h_n<2> pu_h_n<1> pu_h_n<0> puen_h<1> 
+ puen_h<0> slow_h slow_h_n tie_hi_esd vcc_io vgnd vgnd_io / 
+ sky130_fd_io__gpiov2_obpredrvr
.ENDS
.SUBCKT sky130_fd_io__gpiov2_opath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n hld_i_ovr_h od_h oe_n out pad slow tie_hi_esd tie_lo_esd 
+ vcc_io vgnd vgnd_io vpwr vpwr_ka
*.PININFO dm_h<2>:I dm_h<1>:I dm_h<0>:I dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I 
*.PININFO hld_i_h_n:I hld_i_ovr_h:I od_h:I oe_n:I out:I slow:I vcc_io:I vgnd:I 
*.PININFO vgnd_io:I vpwr:I vpwr_ka:I pad:O tie_hi_esd:O tie_lo_esd:O
Xodrvr net70 pad pd_h<3> pd_h<2> pd_h<1> pd_h<0> pd_h<4> pu_h_n<3> pu_h_n<2> 
+ pu_h_n<1> pu_h_n<0> tie_hi_esd tie_lo_esd vcc_io vgnd vgnd_io / 
+ sky130_fd_io__gpiov2_odrvr
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> drvhi_h hld_i_h_n 
+ hld_i_ovr_h od_h oe_n out pd_h<4> pd_h<3> pd_h<2> pd_h<1> pd_h<0> pu_h_n<3> 
+ pu_h_n<2> pu_h_n<1> pu_h_n<0> slow slow_h_n tie_hi_esd vcc_io vgnd vgnd_io 
+ vpwr vpwr_ka / sky130_fd_io__gpiov2_octl_dat
.ENDS
.SUBCKT sky130_fd_io__hvsbt_inv_x4 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEin in / icecap
XICEout out / icecap
mI1 out in vpwr vpwr phv m=8 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 out in vgnd vgnd nhv m=4 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__hvsbt_inv_x8 in out vgnd vpwr
*.PININFO in:I vgnd:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vgnd nhv m=8 w=0.70 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in vpwr vpwr phv m=16 w=1.00 l=0.60 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ctl_hld enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h 
+ hld_ovr od_i_h vcc_io vgnd vpwr
*.PININFO enable_h:I hld_h_n:I hld_ovr:I vcc_io:I vgnd:I vpwr:I hld_i_h:O 
*.PININFO hld_i_h_n:O hld_i_ovr_h:O od_i_h:O
XICEenable_vdda_h_n enable_vdda_h_n / icecap
XICEhld_ovr hld_ovr / icecap
XICEod_i_h od_i_h / icecap
XICEhld_h_n hld_h_n / icecap
XICEod_h od_h / icecap
XICEhld_ovr_h hld_ovr_h / icecap
XICEod_i_h_n od_i_h_n / icecap
XICEnet37 net37 / icecap
XICEhld_i_ovr_h_n hld_i_ovr_h_n / icecap
XICEnet65 net65 / icecap
XICEenable_h enable_h / icecap
XICEnet64 net64 / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
Xhld_ovr_ls net65 hld_ovr hld_ovr_h net37 od_h vgnd vcc_io vgnd vpwr / 
+ sky130_fd_io__com_ctl_ls
XI30 od_i_h hld_i_ovr_h_n hld_i_ovr_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
XI26 net65 hld_ovr_h hld_i_ovr_h_n vgnd vcc_io / sky130_fd_io__hvsbt_nor
Xhld_i_h_inv4 net65 enable_vdda_h_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x4
XI31 od_i_h_n od_i_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x4
Xhld_nand enable_h hld_h_n net64 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
Xod_h_inv enable_h od_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv1 net64 net65 vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
XI32 od_h od_i_h_n vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
Xhld_i_h_inv8<1> enable_vdda_h_n hld_i_h_n_net<1> net019<0> net018<0> / 
+ sky130_fd_io__hvsbt_inv_x8
Xhld_i_h_inv8<0> enable_vdda_h_n hld_i_h_n_net<0> net019<1> net018<1> / 
+ sky130_fd_io__hvsbt_inv_x8
rshort<1> hld_i_h_n_net<1> hld_i_h_n short
rshort<0> hld_i_h_n_net<0> hld_i_h_n short
rshort_hld_i_h enable_vdda_h_n hld_i_h short
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ctl_lsbank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n ib_mode_sel ib_mode_sel_h 
+ ib_mode_sel_h_n inp_dis inp_dis_h inp_dis_h_n od_i_h startup_rst_h 
+ startup_st_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I hld_i_h_n:I ib_mode_sel:I inp_dis:I od_i_h:I 
*.PININFO startup_rst_h:I startup_st_h:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I 
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
*.PININFO ib_mode_sel_h:O ib_mode_sel_h_n:O inp_dis_h:O inp_dis_h_n:O 
*.PININFO vtrip_sel_h:O vtrip_sel_h_n:O
XICEdm_h_n<0> dm_h_n<0> / icecap
XICEie_n_rst_h ie_n_rst_h / icecap
XICEdm_st_h<2> dm_st_h<2> / icecap
XI660<0> dm_h_n<2> / icecap
XI660<1> dm_h_n<1> / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEinp_dis inp_dis / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
XICEdm_rst_h<2> dm_rst_h<2> / icecap
XICEinp_dis_h inp_dis_h / icecap
XICEtrip_sel_rst_h trip_sel_rst_h / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEstartup_rst_h startup_rst_h / icecap
XI659<0> dm_st_h<2> / icecap
XI659<1> dm_st_h<1> / icecap
XICEib_mode_sel_rst_h ib_mode_sel_rst_h / icecap
XI663<0> dm_h<2> / icecap
XI663<1> dm_h<1> / icecap
XI662<0> dm_rst_h<2> / icecap
XI662<1> dm_rst_h<1> / icecap
XICEdm_st_h<1> dm_st_h<1> / icecap
XICEvtrip_sel vtrip_sel / icecap
XICEdm<0> dm<0> / icecap
XICEib_mode_sel ib_mode_sel / icecap
XICEdm_rst_h<1> dm_rst_h<1> / icecap
XICEstartup_st_h startup_st_h / icecap
XICEdm_h<0> dm_h<0> / icecap
XICEdm_rst_h<0> dm_rst_h<0> / icecap
XICEod_i_h od_i_h / icecap
XICEib_mode_sel_h ib_mode_sel_h / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XICEib_mode_sel_st_h ib_mode_sel_st_h / icecap
XICEie_n_st_h ie_n_st_h / icecap
XI661<0> dm<2> / icecap
XI661<1> dm<1> / icecap
XICEdm_st_h<0> dm_st_h<0> / icecap
XICEtrip_sel_st_h trip_sel_st_h / icecap
Xtrip_sel_st trip_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
Xtrip_sel_rst trip_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
Xie_n_rst ie_n_rst_h startup_rst_h startup_st_h / sky130_fd_io__tk_opti
Xie_n_st ie_n_st_h startup_st_h startup_rst_h / sky130_fd_io__tk_opti
XI338<1> dm_rst_h<0> startup_st_h startup_rst_h / sky130_fd_io__tk_opti
XI803<1> dm_st_h<1> od_i_h vgnd / sky130_fd_io__tk_opti
XI802<1> dm_st_h<2> od_i_h vgnd / sky130_fd_io__tk_opti
XI804<1> dm_rst_h<2> vgnd od_i_h / sky130_fd_io__tk_opti
XI805<1> dm_rst_h<1> vgnd od_i_h / sky130_fd_io__tk_opti
XI598 ib_mode_sel_st_h od_i_h vgnd / sky130_fd_io__tk_opti
XI597 ib_mode_sel_rst_h vgnd od_i_h / sky130_fd_io__tk_opti
XI337<1> dm_st_h<0> startup_rst_h startup_st_h / sky130_fd_io__tk_opti
Xdm_ls<0> hld_i_h_n dm<0> dm_h<0> dm_h_n<0> dm_rst_h<0> dm_st_h<0> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
Xinp_dis_ls hld_i_h_n inp_dis inp_dis_h inp_dis_h_n ie_n_rst_h ie_n_st_h 
+ vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
Xtrip_sel_ls hld_i_h_n vtrip_sel vtrip_sel_h vtrip_sel_h_n trip_sel_rst_h 
+ trip_sel_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
Xdm_ls<2> hld_i_h_n dm<2> dm_h<2> dm_h_n<2> dm_rst_h<2> dm_st_h<2> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
Xdm_ls<1> hld_i_h_n dm<1> dm_h<1> dm_h_n<1> dm_rst_h<1> dm_st_h<1> vcc_io vgnd 
+ vpwr / sky130_fd_io__com_ctl_ls
XI595 hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n ib_mode_sel_rst_h 
+ ib_mode_sel_st_h vcc_io vgnd vpwr / sky130_fd_io__com_ctl_ls
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ctl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> 
+ dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_h enable_inp_h hld_h_n hld_i_h 
+ hld_i_h_n hld_i_ovr_h hld_ovr ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n 
+ inp_dis inp_dis_h_n od_i_h vcc_io vgnd vpwr vtrip_sel vtrip_sel_h 
+ vtrip_sel_h_n
*.PININFO dm<2>:I dm<1>:I dm<0>:I enable_h:I enable_inp_h:I hld_h_n:I 
*.PININFO hld_ovr:I ib_mode_sel:I inp_dis:I vcc_io:I vgnd:I vpwr:I vtrip_sel:I 
*.PININFO dm_h<2>:O dm_h<1>:O dm_h<0>:O dm_h_n<2>:O dm_h_n<1>:O dm_h_n<0>:O 
*.PININFO hld_i_h:O hld_i_h_n:O hld_i_ovr_h:O ib_mode_sel_h:O 
*.PININFO ib_mode_sel_h_n:O inp_dis_h_n:O od_i_h:O vtrip_sel_h:O 
*.PININFO vtrip_sel_h_n:O
XICEnet92 net92 / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEvtrip_sel vtrip_sel / icecap
XICEstartup_rst_h startup_rst_h / icecap
XICEinp_startup_en_h inp_startup_en_h / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEib_mode_sel_h ib_mode_sel_h / icecap
XI78<0> dm_h_n<2> / icecap
XI78<1> dm_h_n<1> / icecap
XI78<2> dm_h_n<0> / icecap
XICEenable_h enable_h / icecap
XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
XICEib_mode_sel ib_mode_sel / icecap
XICEhld_ovr hld_ovr / icecap
XI76<0> dm_h<2> / icecap
XI76<1> dm_h<1> / icecap
XI76<2> dm_h<0> / icecap
XICEinp_dis inp_dis / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEnet80 net80 / icecap
XICEhld_i_h hld_i_h / icecap
XICEenable_inp_h enable_inp_h / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XI77<0> dm<2> / icecap
XI77<1> dm<1> / icecap
XI77<2> dm<0> / icecap
XICEod_i_h od_i_h / icecap
XICEhld_h_n hld_h_n / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XI75 enable_inp_h enable_h startup_rst_h vgnd vcc_io / sky130_fd_io__hvsbt_nor
Xhld_dis_blk enable_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr od_i_h 
+ vcc_io vgnd vpwr / sky130_fd_io__gpiov2_ctl_hld
Xls_bank dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> 
+ dm_h_n<0> hld_i_h_n ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n inp_dis net80 
+ inp_dis_h_n od_i_h startup_rst_h inp_startup_en_h vcc_io vgnd vpwr vtrip_sel 
+ vtrip_sel_h vtrip_sel_h_n / sky130_fd_io__gpiov2_ctl_lsbank
XI56 od_i_h enable_inp_h net92 vgnd vcc_io / sky130_fd_io__hvsbt_nand2
XI57 net92 inp_startup_en_h vgnd vcc_io / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpiov2_inbuf_lvinv_x1 in out vgnd vnb vpb vpwr
*.PININFO in:I vgnd:I vnb:I vpb:I vpwr:I out:O
XICEout out / icecap
XICEin in / icecap
mI2 out in vgnd vnb nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI1 out in vpwr vpb phighvt m=1 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ipath_lvls in_vcchib in_vddio mode_normal_lv 
+ mode_normal_lv_n mode_vcchib_lv mode_vcchib_lv_n out out_b vcchib vssd
*.PININFO in_vcchib:I in_vddio:I mode_normal_lv:I mode_normal_lv_n:I 
*.PININFO mode_vcchib_lv:I mode_vcchib_lv_n:I vcchib:I vssd:I out:O out_b:O
XICEin_vcchib in_vcchib / icecap
XICEout out / icecap
XICEmode_normal_lv mode_normal_lv / icecap
XICEfbk_n fbk_n / icecap
XICEmode_vcchib_lv mode_vcchib_lv / icecap
XICEnet50 net50 / icecap
XICEnet78 net78 / icecap
XICEfbk fbk / icecap
XICEmode_normal_lv_n mode_normal_lv_n / icecap
XICEin_vddio in_vddio / icecap
XICEnet95 net95 / icecap
XICEmode_vcchib_lv_n mode_vcchib_lv_n / icecap
XICEnet115 net115 / icecap
XICEnet111 net111 / icecap
XICEout_b out_b / icecap
mI345 fbk_n in_vddio vcchib vcchib phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI344 net70 mode_vcchib_lv vcchib vcchib pshort m=1 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI343 out_b fbk net78 vcchib pshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI342 net78 mode_normal_lv_n vcchib vcchib pshort m=2 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI341 out_b mode_normal_lv net70 vcchib pshort m=1 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI340 net50 mode_vcchib_lv_n vcchib vcchib pshort m=2 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI339 fbk_n mode_normal_lv vcchib vcchib pshort m=1 w=5.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI338 fbk fbk_n vcchib vcchib pshort m=1 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI337 out out_b vcchib vcchib pshort m=4 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI336 out_b in_vcchib net50 vcchib pshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI351 net111 mode_normal_lv vssd vssd nshort m=2 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI350 out_b fbk net111 vssd nshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI349 out out_b vssd vssd nshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI348 fbk fbk_n vssd vssd nshort m=1 w=3.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI347 net95 mode_vcchib_lv vssd vssd nshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI346 out_b in_vcchib net95 vssd nshort m=2 w=3.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI353 fbk_n in_vddio net115 vssd nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI352 net115 mode_normal_lv vssd vssd nshort m=1 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ipath_hvls in_vcchib in_vddio inb_vcchib mode_normal 
+ mode_normal_n mode_vcchib mode_vcchib_n out out_b vddio_q vssd
*.PININFO in_vcchib:I in_vddio:I inb_vcchib:I mode_normal:I mode_normal_n:I 
*.PININFO mode_vcchib:I mode_vcchib_n:I vddio_q:I vssd:I out:O out_b:O
XICEinb_vcchib inb_vcchib / icecap
XICEin_vcchib in_vcchib / icecap
XICEnet75 net75 / icecap
XICEin_vddio in_vddio / icecap
XICEnet84 net84 / icecap
XICEout out / icecap
XICEout_b out_b / icecap
XICEmode_vcchib_n mode_vcchib_n / icecap
XICEnet92 net92 / icecap
XICEfbk fbk / icecap
XICEmode_normal mode_normal / icecap
XICEfbk_b fbk_b / icecap
XICEnet116 net116 / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEnet55 net55 / icecap
XICEmode_vcchib mode_vcchib / icecap
mI325 fbk fbk_b vddio_q vddio_q phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI324 fbk_b fbk vddio_q vddio_q phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI323 net63 mode_normal vddio_q vddio_q phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI322 out_b in_vddio net75 vddio_q phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI321 net75 mode_normal_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI320 out out_b vddio_q vddio_q phv m=5 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI319 out_b mode_vcchib net63 vddio_q phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI318 net55 mode_vcchib_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI317 out_b net84 net55 vddio_q phv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI336 net84 fbk_b vddio_q vddio_q phv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI335 out_b net84 net88 vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI334 fbk inb_vcchib net116 vssd nhv m=3 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI333 net116 mode_vcchib vssd vssd nhv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI332 net112 mode_normal vssd vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI331 out out_b vssd vssd nhv m=3 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI330 out_b in_vddio net112 vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI329 fbk_b in_vcchib net92 vssd nhv m=3 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI328 fbk mode_vcchib_n vssd vssd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI327 net92 mode_vcchib vssd vssd nhv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI326 net88 mode_vcchib vssd vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI337 net84 fbk_b vssd vssd nhv m=1 w=1.50 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_vcchib_in_buf in_h mode_vcchib_lv_n out out_n vcchib 
+ vssd
*.PININFO in_h:I mode_vcchib_lv_n:I vcchib:I vssd:I out:O out_n:O
XICEnet57 net57 / icecap
XICEnet81 net81 / icecap
XICEnet112 net112 / icecap
XICEmode_vcchib_lv_n mode_vcchib_lv_n / icecap
XICEout out / icecap
XICEout_n out_n / icecap
XICEnet108 net108 / icecap
XICEin_b in_b / icecap
XICEfbk fbk / icecap
XICEin_h in_h / icecap
mI420 net57 in_b fbk vssd nhv m=3 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI552 vssd vssd vssd vssd nhv m=1 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI544 fbk in_h vssd vssd nhv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI551 vssd vssd vssd vssd nhv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI424 net81 in_b vssd vssd nshort m=2 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI423 out_n net81 vssd vssd nshort m=1 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI545 in_b in_h fbk vssd nhv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI487 out out_n vssd vssd nshort m=3 w=1.00 l=0.25 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI541 net81 mode_vcchib_lv_n vssd vssd nshort m=2 w=1.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI549 net57 mode_vcchib_lv_n vcchib vcchib pshort m=1 w=5.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI436 net81 in_b net112 vcchib pshort m=2 w=1.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI543 in_b in_h net108 vcchib phv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI429 out_n net81 vcchib vcchib pshort m=1 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI538 net112 mode_vcchib_lv_n vcchib vcchib pshort m=1 w=3.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI489 out out_n vcchib vcchib pshort m=1 w=5.00 l=0.25 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI547 net108 mode_vcchib_lv_n vcchib vcchib pshort m=3 w=5.00 l=0.25 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_in_buf in_h in_vt mode_normal_n out out_n vddio_q vssd 
+ vtrip_sel_h vtrip_sel_h_n
*.PININFO in_h:I in_vt:I mode_normal_n:I vddio_q:I vssd:I vtrip_sel_h:I 
*.PININFO vtrip_sel_h_n:I out:O out_n:O
XICEmode_normal_n mode_normal_n / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEnet122 net122 / icecap
XICEin_h in_h / icecap
XICEin_vt in_vt / icecap
XICEnet158 net158 / icecap
XICEnet103 net103 / icecap
XICEmode_normal_cmos_h_n mode_normal_cmos_h_n / icecap
XICEnet138 net138 / icecap
XICEmode_normal_cmos_h mode_normal_cmos_h / icecap
XICEnet91 net91 / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEout out / icecap
XICEfbk fbk / icecap
XICEfbk2 fbk2 / icecap
XICEout_n out_n / icecap
XICEin_b in_b / icecap
XI43 mode_normal_cmos_h mode_normal_cmos_h_n vssd vddio_q / 
+ sky130_fd_io__hvsbt_inv_x1
XI488 vtrip_sel_h mode_normal_n mode_normal_cmos_h vssd vddio_q / 
+ sky130_fd_io__hvsbt_nor
mI583 in_vt vtrip_sel_h_n vssd vssd nhv m=1 w=3.00 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI644 vssd vssd vssd vssd nhv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI646 vssd vssd vssd vssd nhv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI593 net91 mode_normal_n vssd vssd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI592 net103 in_b fbk vssd nhv m=4 w=1.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI591 fbk in_h vssd vssd nhv m=6 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI590 fbk2 in_b fbk vssd nhv m=4 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI589 net91 in_b vssd vssd nhv m=2 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI588 fbk in_vt vssd vssd nhv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI587 in_b in_h fbk vssd nhv m=5 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI586 out_n net91 vssd vssd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI642 out out_n vssd vssd nhv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI629 in_b in_h net158 vddio_q phv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI636 net158 mode_normal_cmos_h_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI632 net122 mode_normal_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI647 vddio_q vddio_q vddio_q vddio_q phv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI600 net103 mode_normal_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI598 net91 in_b net138 vddio_q phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI597 fbk2 mode_normal_cmos_h_n vddio_q vddio_q phv m=2 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI596 out_n net91 vddio_q vddio_q phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI595 net138 mode_normal_n vddio_q vddio_q phv m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI631 in_b in_h net122 vddio_q phv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI643 out out_n vddio_q vddio_q phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ibuf_se enable_vddio_lv ibufmux_out ibufmux_out_h in_h 
+ in_vt mode_normal_n mode_vcchib_n vcchib vddio_q vssd vtrip_sel_h 
+ vtrip_sel_h_n
*.PININFO enable_vddio_lv:I in_h:I in_vt:I mode_normal_n:I mode_vcchib_n:I 
*.PININFO vcchib:I vddio_q:I vssd:I vtrip_sel_h:I vtrip_sel_h_n:I 
*.PININFO ibufmux_out:O ibufmux_out_h:O
XICEvtrip_sel_h vtrip_sel_h / icecap
XICEout_n_vddio out_n_vddio / icecap
XICEmode_vcchib mode_vcchib / icecap
XICEmode_vcchib_lv_n mode_vcchib_lv_n / icecap
XICEout_n_vcchib out_n_vcchib / icecap
XICEmode_normal_lv_n mode_normal_lv_n / icecap
XICEmode_normal mode_normal / icecap
XICEin_h in_h / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEout_vcchib out_vcchib / icecap
XICEnet57 net57 / icecap
XICEibufmux_out ibufmux_out / icecap
XICEmode_vcchib_n mode_vcchib_n / icecap
XICEibufmux_out_h ibufmux_out_h / icecap
XICEmode_normal_lv mode_normal_lv / icecap
XICEnet68 net68 / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEout_vddio out_vddio / icecap
XICEmode_vcchib_lv mode_vcchib_lv / icecap
XICEin_vt in_vt / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XI148 enable_vddio_lv mode_vcchib mode_vcchib_lv_n vssd vcchib / 
+ sky130_fd_io__hvsbt_nand2
XI149 enable_vddio_lv mode_normal mode_normal_lv_n vssd vcchib / 
+ sky130_fd_io__hvsbt_nand2
XI112 mode_normal_lv_n mode_normal_lv vssd vssd vcchib vcchib / 
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1
XI111 mode_vcchib_lv_n mode_vcchib_lv vssd vssd vcchib vcchib / 
+ sky130_fd_io__gpiov2_inbuf_lvinv_x1
Xlvls out_vcchib out_vddio mode_normal_lv mode_normal_lv_n mode_vcchib_lv 
+ mode_vcchib_lv_n ibufmux_out net57 vcchib vssd / sky130_fd_io__gpiov2_ipath_lvls
Xhvls out_vcchib out_vddio out_n_vcchib mode_normal mode_normal_n mode_vcchib 
+ mode_vcchib_n ibufmux_out_h net68 vddio_q vssd / sky130_fd_io__gpiov2_ipath_hvls
XI88 in_h mode_vcchib_lv_n out_vcchib out_n_vcchib vcchib vssd / 
+ sky130_fd_io__gpiov2_vcchib_in_buf
Xbuf in_h in_vt mode_normal_n out_vddio out_n_vddio vddio_q vssd vtrip_sel_h 
+ vtrip_sel_h_n / sky130_fd_io__gpiov2_in_buf
XI491 mode_normal_n mode_normal vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI105 mode_vcchib_n mode_vcchib vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ictl_logic dm_h_n<2> dm_h_n<1> dm_h_n<0> ib_mode_sel_h 
+ ib_mode_sel_h_n inp_dis_h_n inp_dis_i_h inp_dis_i_h_n mode_normal_n 
+ mode_vcchib_n tripsel_i_h tripsel_i_h_n vddio_q vssd vtrip_sel_h_n
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I ib_mode_sel_h:I 
*.PININFO ib_mode_sel_h_n:I inp_dis_h_n:I vddio_q:I vssd:I vtrip_sel_h_n:I 
*.PININFO inp_dis_i_h:O inp_dis_i_h_n:O mode_normal_n:O mode_vcchib_n:O 
*.PININFO tripsel_i_h:O tripsel_i_h_n:O
XICEdm_buf_dis_n dm_buf_dis_n / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEand_dm01 and_dm01 / icecap
XICEdm_h_n<1> dm_h_n<1> / icecap
XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
XICEinp_dis_i_h inp_dis_i_h / icecap
XICEnand_dm01 nand_dm01 / icecap
XICEtripsel_i_h_n tripsel_i_h_n / icecap
XICEinp_dis_h_n inp_dis_h_n / icecap
XICEinp_dis_i_h_n inp_dis_i_h_n / icecap
XICEtripsel_i_h tripsel_i_h / icecap
XICEdm_h_n<2> dm_h_n<2> / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEmode_vcchib_n mode_vcchib_n / icecap
XICEdm_h_n<0> dm_h_n<0> / icecap
XICEib_mode_sel_h ib_mode_sel_h / icecap
XI71 vtrip_sel_h_n mode_normal_n tripsel_i_h vssd vddio_q / sky130_fd_io__hvsbt_nor
XI80 dm_buf_dis_n inp_dis_h_n inp_dis_i_h vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI79 dm_h_n<2> and_dm01 dm_buf_dis_n vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI78 dm_h_n<1> dm_h_n<0> nand_dm01 vssd vddio_q / sky130_fd_io__hvsbt_nand2
XI36 inp_dis_i_h_n ib_mode_sel_h mode_vcchib_n vssd vddio_q / 
+ sky130_fd_io__hvsbt_nand2
XI35 inp_dis_i_h_n ib_mode_sel_h_n mode_normal_n vssd vddio_q / 
+ sky130_fd_io__hvsbt_nand2
XI111 inp_dis_i_h inp_dis_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI75 nand_dm01 and_dm01 vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI74 tripsel_i_h tripsel_i_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
.ENDS
.SUBCKT sky130_fd_io__gpiov2_ipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio_lv 
+ ib_mode_sel_h ib_mode_sel_h_n inp_dis_h_n out out_h pad vcchib vddio_q vssd 
+ vtrip_sel_h_n
*.PININFO dm_h_n<2>:I dm_h_n<1>:I dm_h_n<0>:I enable_vddio_lv:I 
*.PININFO ib_mode_sel_h:I ib_mode_sel_h_n:I inp_dis_h_n:I vcchib:I vddio_q:I 
*.PININFO vssd:I vtrip_sel_h_n:I out:O out_h:O pad:B
XICEinp_dis_h_n inp_dis_h_n / icecap
XICEin_h in_h / icecap
XICEmode_normal_n mode_normal_n / icecap
XICEen_h_n en_h_n / icecap
XICEpad pad / icecap
XICEen_h en_h / icecap
XICEout_h out_h / icecap
XICEin_vt in_vt / icecap
XICEvtrip_sel_h_n vtrip_sel_h_n / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEtripsel_i_h tripsel_i_h / icecap
XICEib_mode_sel_h_n ib_mode_sel_h_n / icecap
XI152<0> dm_h_n<2> / icecap
XI152<1> dm_h_n<1> / icecap
XI152<2> dm_h_n<0> / icecap
XICEtripsel_i_h_n tripsel_i_h_n / icecap
XICEib_mode_sel_h ib_mode_sel_h / icecap
XICEmode_vcchib_n mode_vcchib_n / icecap
XICEout out / icecap
XI106 enable_vddio_lv out out_h in_h in_vt mode_normal_n mode_vcchib_n vcchib 
+ vddio_q vssd tripsel_i_h tripsel_i_h_n / sky130_fd_io__gpiov2_ibuf_se
XI107 dm_h_n<2> dm_h_n<1> dm_h_n<0> ib_mode_sel_h ib_mode_sel_h_n inp_dis_h_n 
+ en_h_n en_h mode_normal_n mode_vcchib_n tripsel_i_h tripsel_i_h_n vddio_q 
+ vssd vtrip_sel_h_n / sky130_fd_io__gpiov2_ictl_logic
XI120 pad in_h in_vt vddio_q vssd tripsel_i_h / 
+ sky130_fd_io__gpio_ovtv2_buf_localesd
.ENDS
.SUBCKT sky130_fd_io__top_gpiov2 amuxbus_a amuxbus_b analog_en analog_pol 
+ analog_sel dm<2> dm<1> dm<0> enable_h enable_inp_h enable_vdda_h 
+ enable_vddio enable_vswitch_h hld_h_n hld_ovr ib_mode_sel in in_h inp_dis 
+ oe_n out pad pad_a_esd_0_h pad_a_esd_1_h pad_a_noesd_h slow tie_hi_esd 
+ tie_lo_esd vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q vswitch 
+ vtrip_sel
*.PININFO analog_en:I analog_pol:I analog_sel:I dm<2>:I dm<1>:I dm<0>:I 
*.PININFO enable_h:I enable_inp_h:I enable_vdda_h:I enable_vddio:I 
*.PININFO enable_vswitch_h:I hld_h_n:I hld_ovr:I ib_mode_sel:I inp_dis:I 
*.PININFO oe_n:I out:I slow:I vtrip_sel:I in:O in_h:O tie_hi_esd:O 
*.PININFO tie_lo_esd:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_0_h:B 
*.PININFO pad_a_esd_1_h:B pad_a_noesd_h:B vccd:B vcchib:B vdda:B vddio:B 
*.PININFO vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xamux amuxbus_a amuxbus_b analog_en analog_pol analog_sel enable_vdda_h 
+ enable_vswitch_h hld_i_h hld_i_h_n out pad vccd vdda vddio_q vssa vssd 
+ vssio_q vswitch / sky130_fd_io__gpiov2_amux
Xopath dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> hld_i_h_n 
+ hld_i_ovr_h od_i_h oe_n out pad slow tie_hi_esd tie_lo_esd vddio vssd vssio 
+ vccd vcchib / sky130_fd_io__gpiov2_opath
Xctrl dm<2> dm<1> dm<0> dm_h<2> dm_h<1> dm_h<0> dm_h_n<2> dm_h_n<1> dm_h_n<0> 
+ enable_h enable_inp_h hld_h_n hld_i_h hld_i_h_n hld_i_ovr_h hld_ovr 
+ ib_mode_sel ib_mode_sel_h ib_mode_sel_h_n inp_dis inp_dis_h_n od_i_h vddio_q 
+ vssd vccd vtrip_sel vtrip_sel_h vtrip_sel_h_n / sky130_fd_io__gpiov2_ctl
Xipath dm_h_n<2> dm_h_n<1> dm_h_n<0> enable_vddio ib_mode_sel_h 
+ ib_mode_sel_h_n inp_dis_h_n in in_h pad vcchib vddio_q vssd vtrip_sel_h_n / 
+ sky130_fd_io__gpiov2_ipath
Xresd3 pad_a_esd_1_h net210 / s8_esd_res75only_small
Xresd1 net204 pad / s8_esd_res75only_small
Xresd4 net210 pad / s8_esd_res75only_small
Xresd2 pad_a_esd_0_h net204 / s8_esd_res75only_small
XICEoe_n oe_n / icecap
XICEhld_h_n hld_h_n / icecap
XICEslow slow / icecap
XICEpad pad / icecap
XICEtie_hi_esd tie_hi_esd / icecap
XI259<0> dm_h_n<2> / icecap
XI259<1> dm_h_n<1> / icecap
XI259<2> dm_h_n<0> / icecap
XI257<0> dm_h<2> / icecap
XI257<1> dm_h<1> / icecap
XI257<2> dm_h<0> / icecap
XICEhld_i_h_n hld_i_h_n / icecap
XICEtie_lo_esd tie_lo_esd / icecap
XI258<0> dm<2> / icecap
XI258<1> dm<1> / icecap
XI258<2> dm<0> / icecap
XICEinp_dis inp_dis / icecap
XICEhld_i_ovr_h hld_i_ovr_h / icecap
XICEhld_ovr hld_ovr / icecap
XICEout out / icecap
XICEvtrip_sel vtrip_sel / icecap
XICEod_h od_i_h / icecap
rS0<2> pad pad_a_noesd_h short
rS0<1> pad pad_a_noesd_h short
rS0<0> pad pad_a_noesd_h short
.ENDS

.SUBCKT s8_esd_gnd2gnd_120x2_lv_isosub vssi vssn vsub
*.PININFO vssi:B vssn:B vsub:B
dI9 vssn vssi pdiode m=4 area=22.5 pj=33
dI10 vssi vssn pdiode m=4 area=22.5 pj=33
.ENDS

.SUBCKT sky130_fd_io__top_power_lvc_wpad amuxbus_a amuxbus_b bdy2_b2b drn_lvc1 
+ drn_lvc2 ogc_lvc p_core p_pad src_bdy_lvc1 src_bdy_lvc2 vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B bdy2_b2b:B drn_lvc1:B drn_lvc2:B ogc_lvc:B 
*.PININFO p_core:B p_pad:B src_bdy_lvc1:B src_bdy_lvc2:B vccd:B vcchib:B 
*.PININFO vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xesd bdy2_b2b src_bdy_lvc1 vssd / s8_esd_gnd2gnd_120x2_lv_isosub
xI54 src_bdy_lvc2 vddio condiode
xI50 src_bdy_lvc1 vddio condiode
rI21 p_pad p_core short
mpre_p1 g_nclamp_lvc1 g_pdpre_lvc1 drn_lvc1 drn_lvc1 pshort m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI40 g_nclamp_lvc2 g_pdpre_lvc2 drn_lvc2 drn_lvc2 pshort m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mclamp_xtor drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=166 
+ w=7.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ area=0.063 perim=1.14
mI42 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=152 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI61 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=38 w=5.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI62 drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=20 w=5.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mncap src_bdy_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=15 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mpre_n1 g_nclamp_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=3 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI43 g_nclamp_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=2 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI58 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=6 w=5.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI60 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=1 w=5.00 
+ l=4.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI59 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=10 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
rrc_res g_pdpre_lvc1 drn_lvc1 mrp1 m=1 w=0.33 l=1950
rI44 drn_lvc2 net161 mrp1 m=1 w=0.33 l=900
rI47 net161 net155 mrp1 m=1 w=0.33 l=300
rI46 g_pdpre_lvc2 net157 mrp1 m=1 w=0.33 l=200
rI45 net157 net155 mrp1 m=1 w=0.33 l=720
.ENDS

.SUBCKT sky130_fd_io__top_ground_lvc_wpad amuxbus_a amuxbus_b bdy2_b2b drn_lvc1 
+ drn_lvc2 g_core g_pad ogc_lvc src_bdy_lvc1 src_bdy_lvc2 vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B bdy2_b2b:B drn_lvc1:B drn_lvc2:B g_core:B 
*.PININFO g_pad:B ogc_lvc:B src_bdy_lvc1:B src_bdy_lvc2:B vccd:B vcchib:B 
*.PININFO vdda:B vddio:B vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
Xesd bdy2_b2b src_bdy_lvc1 vssd / s8_esd_gnd2gnd_120x2_lv_isosub
xI54 src_bdy_lvc2 vddio condiode
xI50 src_bdy_lvc1 vddio condiode
rI21 g_pad g_core short
mpre_p1 g_nclamp_lvc1 g_pdpre_lvc1 drn_lvc1 drn_lvc1 pshort m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI40 g_nclamp_lvc2 g_pdpre_lvc2 drn_lvc2 drn_lvc2 pshort m=20 w=7.00 l=0.18 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mclamp_xtor drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=166 
+ w=7.00 l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal 
+ area=0.063 perim=1.14
mI42 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=152 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI61 drn_lvc2 g_nclamp_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=38 w=5.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI62 drn_lvc1 g_nclamp_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=20 w=5.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mncap src_bdy_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=15 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mpre_n1 g_nclamp_lvc1 g_pdpre_lvc1 src_bdy_lvc1 src_bdy_lvc1 nshort m=3 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI43 g_nclamp_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=2 w=7.00 
+ l=0.18 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI58 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=6 w=5.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI60 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=1 w=5.00 
+ l=4.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
mI59 src_bdy_lvc2 g_pdpre_lvc2 src_bdy_lvc2 src_bdy_lvc2 nshort m=10 w=7.00 
+ l=8.00 mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 
+ perim=1.14
rrc_res g_pdpre_lvc1 drn_lvc1 mrp1 m=1 w=0.33 l=1950
rI44 drn_lvc2 net161 mrp1 m=1 w=0.33 l=900
rI47 net161 net155 mrp1 m=1 w=0.33 l=300
rI46 g_pdpre_lvc2 net157 mrp1 m=1 w=0.33 l=200
rI45 net157 net155 mrp1 m=1 w=0.33 l=720
.ENDS

.SUBCKT sky130_fd_io__top_ground_hvc_wpad amuxbus_a amuxbus_b drn_hvc g_core g_pad 
+ ogc_hvc src_bdy_hvc vccd vcchib vdda vddio vddio_q vssa vssd vssio vssio_q 
+ vswitch
*.PININFO amuxbus_a:B amuxbus_b:B drn_hvc:B g_core:B g_pad:B ogc_hvc:B 
*.PININFO src_bdy_hvc:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B 
*.PININFO vssio:B vssio_q:B vswitch:B
mcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc nhv m=22 w=10.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc nhv m=5 w=5.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc nhv m=15 w=5.00 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc nhv m=15 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc nhv m=120 w=20.0 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
rrc_res g_pdpre net94 mrp1 m=1 w=0.33 l=470
rI38 net90 drn_hvc mrp1 m=1 w=0.33 l=700
rI37 net94 net90 mrp1 m=1 w=0.33 l=1550
mpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc phv m=50 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
xI39 src_bdy_hvc vddio condiode
rI13 g_pad g_core short
.ENDS
.SUBCKT sky130_fd_io__top_hvclamp_wopadv2 drn_hvc ogc_hvc src_bdy_hvc vssd
*.PININFO drn_hvc:B ogc_hvc:B src_bdy_hvc:B vssd:B
xI39 src_bdy_hvc ogc_hvc condiode
mpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc phv m=50 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
rrc_res g_pdpre net41 mrp1 m=1 w=0.33 l=470
rI38 net37 drn_hvc mrp1 m=1 w=0.33 l=700
rI37 net41 net37 mrp1 m=1 w=0.33 l=1550
mclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc nhv m=120 w=20.0 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc nhv m=15 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc nhv m=15 w=5.00 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc nhv m=5 w=5.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc nhv m=22 w=10.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 amuxbus_a amuxbus_b drn_hvc ogc_hvc 
+ p_core p_pad src_bdy_hvc vccd vcchib vdda vddio vddio_q vssa vssd vssio 
+ vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B drn_hvc:B ogc_hvc:B p_core:B p_pad:B 
*.PININFO src_bdy_hvc:B vccd:B vcchib:B vdda:B vddio:B vddio_q:B vssa:B vssd:B 
*.PININFO vssio:B vssio_q:B vswitch:B
xI39 src_bdy_hvc vddio condiode
mpre_p1 g_nclamp g_pdpre drn_hvc drn_hvc phv m=50 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
rrc_res g_pdpre net67 mrp1 m=1 w=0.33 l=470
rI38 net63 drn_hvc mrp1 m=1 w=0.33 l=700
rI37 net67 net63 mrp1 m=1 w=0.33 l=1550
mclamp_xtor drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc nhv m=120 w=20.0 l=0.50 
+ mult=1 sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mpre_n1 g_nclamp g_pdpre src_bdy_hvc src_bdy_hvc nhv m=15 w=7.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnc1 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc nhv m=15 w=5.00 l=8.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mnc2 src_bdy_hvc g_pdpre src_bdy_hvc src_bdy_hvc nhv m=5 w=5.00 l=4.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mcxtor2 drn_hvc g_nclamp src_bdy_hvc src_bdy_hvc nhv m=22 w=10.0 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
rI13 p_pad p_core short
.ENDS
.SUBCKT sky130_fd_io__top_vrefcapv2 amuxbus_a amuxbus_b cneg cpos vccd vcchib vdda 
+ vddio vddio_q vssa vssd vssio vssio_q vswitch
*.PININFO amuxbus_a:B amuxbus_b:B cneg:B cpos:B vccd:B vcchib:B vdda:B vddio:B 
*.PININFO vddio_q:B vssa:B vssd:B vssio:B vssio_q:B vswitch:B
xI271 cneg vddio_q condiode
mI334 cneg cpos cneg cneg nhvnative m=180 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__xres4v2_in_buf enable_hv enable_vddio_lv in_h in_h_n pad 
+ vcchib vddio vgnd vnormal vnormal_b
*.PININFO enable_hv:I enable_vddio_lv:I pad:I vcchib:I vddio:I vgnd:I 
*.PININFO vnormal:I vnormal_b:I in_h:O in_h_n:O
XICEnet152 net152 / icecap
XICEnet193 net193 / icecap
XICEenable_vddio_lv_n enable_vddio_lv_n / icecap
XICEnet110 net110 / icecap
XICEpad_inv pad_inv / icecap
XICEvnormal_b vnormal_b / icecap
XICEpad1 pad1 / icecap
XICEvcchib_int vcchib_int / icecap
XICEnet116 net116 / icecap
XICEnet124 net124 / icecap
XICEenable_vddio_lv enable_vddio_lv / icecap
XICEnet106 net106 / icecap
XICEmode_vcchib mode_vcchib / icecap
XICEnet235 net235 / icecap
XICEin_h in_h / icecap
XICEin_h_n in_h_n / icecap
XICEenable_hv_b enable_hv_b / icecap
XICEpad pad / icecap
XICEnet140 net140 / icecap
XICEnet112 net112 / icecap
XICEvcchib vcchib / icecap
XICEnet207 net207 / icecap
XICEnet206 net206 / icecap
XICEvnormal vnormal / icecap
XICEenable_hv enable_hv / icecap
XICEfbk fbk / icecap
XICEnet120 net120 / icecap
XICEnet108 net108 / icecap
XI165 enable_vddio_lv enable_vddio_lv_n vgnd vgnd vcchib vcchib / 
+ sky130_fd_io__inv_1
XI61 net106 mode_vcchib vgnd vddio / sky130_fd_io__hvsbt_inv_x1
XI35 vnormal_b enable_hv net106 vgnd vddio / sky130_fd_io__hvsbt_nand2
rI132 net207 net110 mrdn_hv m=1 w=0.29 l=1077.19
rI159 net235 net108 mrp1 m=1 w=0.4 l=713.695
mI8 net193 pad1 vgnd vgnd nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI86 pad1 pad_inv vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI85 pad_inv pad net140 vgnd nhv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI114 net152 pad_inv net140 vgnd nhv m=4 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI145 enable_hv_b enable_hv vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI251 in_h in_h_n vgnd vgnd nhv m=3 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI83 net140 pad vgnd vgnd nhv m=2 w=5.00 l=0.80 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI7 fbk pad_inv vgnd vgnd nhv m=2 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI213 in_h_n fbk vgnd vgnd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI152 vgnd vgnd vgnd vgnd nhvnative m=1 w=10.0 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI113 net124 pad net152 vgnd nhvnative m=1 w=1.00 l=0.90 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI154 net120 mode_vcchib net206 vgnd nhvnative m=1 w=1.00 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI151 net116 mode_vcchib vcchib_int vgnd nhvnative m=1 w=10.0 l=0.90 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI150 net112 pad_inv net140 vgnd nhv m=1 w=5.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI116 pad1 pad_inv net235 vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI143 net124 vnormal vddio vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI156 net116 enable_vddio_lv_n vcchib vcchib phv m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI252 in_h in_h_n vddio vddio phv m=3 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI107 net108 mode_vcchib vddio vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI146 enable_hv_b enable_hv vddio vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI88 pad_inv pad vcchib_int vcchib_int phv m=1 w=1.00 l=0.80 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI89 pad_inv pad net207 vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI90 pad1 pad_inv net206 net206 phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI133 net110 mode_vcchib vddio vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI2 net193 fbk vddio vddio phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI219 fbk net193 vddio vddio phv m=1 w=0.42 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI14 in_h_n fbk vddio vddio phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI158 net120 enable_vddio_lv_n vcchib vcchib phv m=1 w=5.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI139 net207 vnormal_b net110 vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI136 net112 vnormal_b vddio vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI153 vcchib_int vcchib_int vcchib_int vcchib_int phv m=1 w=1.00 l=0.80 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI160 net235 vnormal_b net108 vddio phv m=1 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__gpio_buf_localesd in_h out_h out_vt vcc_io vgnd vtrip_sel_h
*.PININFO in_h:I vtrip_sel_h:I out_h:O out_vt:O vcc_io:B vgnd:B
XICEout_vt out_vt / icecap
XICEin_h in_h / icecap
XICEout_h out_h / icecap
XICEvtrip_sel_h vtrip_sel_h / icecap
mhv_passgate out_h vtrip_sel_h out_vt vgnd nhv m=1 w=3.00 l=1.00 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
Xesd_res in_h out_h / s8_esd_res250only_small
Xggnfet2 vgnd out_vt vgnd vcc_io vgnd / s8_esd_signal_5_sym_hv_local_5term
Xggnfet6 vgnd vcc_io vgnd vcc_io out_h / s8_esd_signal_5_sym_hv_local_5term
Xggnfet5 vgnd vcc_io vgnd vcc_io out_vt / s8_esd_signal_5_sym_hv_local_5term
Xggnfet1 vgnd out_h vgnd vcc_io vgnd / s8_esd_signal_5_sym_hv_local_5term
.ENDS
.SUBCKT sky130_fd_io__gpio_pddrvr_strong force_lo_h force_lovol_h pad pd_h<3> 
+ pd_h<2> tie_lo_esd vcc_io vgnd_io vssio_amx
*.PININFO force_lo_h:I force_lovol_h:I pd_h<3>:I pd_h<2>:I vcc_io:I vgnd_io:I 
*.PININFO vssio_amx:I pad:O tie_lo_esd:O
XI112 pd_h<2> net61 / sky130_fd_io__tk_em2s
XI113 pd_h<2> net59 / sky130_fd_io__tk_em2s
XI97 pd_h<3> net85 / sky130_fd_io__tk_em2s
XI108 tie_lo_esd net83 / sky130_fd_io__tk_em2s
XI109 tie_lo_esd net77 / sky130_fd_io__tk_em2s
XI102 pd_h<3> net73 / sky130_fd_io__tk_em2s
XI104 pd_h<3> net69 / sky130_fd_io__tk_em2s
XI96 pd_h<3> net67 / sky130_fd_io__tk_em2s
XI87 tie_lo_esd net59 / sky130_fd_io__tk_em2o
XI83 pd_h<3> net61 / sky130_fd_io__tk_em2o
XI99 tie_lo_esd net85 / sky130_fd_io__tk_em2o
XI82 tie_lo_esd net61 / sky130_fd_io__tk_em2o
XI98 pd_h<2> net85 / sky130_fd_io__tk_em2o
XI106 pd_h<2> net83 / sky130_fd_io__tk_em2o
XI107 pd_h<3> net83 / sky130_fd_io__tk_em2o
XI110 pd_h<3> net77 / sky130_fd_io__tk_em2o
XI111 pd_h<2> net77 / sky130_fd_io__tk_em2o
XI100 tie_lo_esd net73 / sky130_fd_io__tk_em2o
XI101 pd_h<2> net73 / sky130_fd_io__tk_em2o
XI103 tie_lo_esd net69 / sky130_fd_io__tk_em2o
XI105 pd_h<2> net69 / sky130_fd_io__tk_em2o
XI95 pd_h<2> net67 / sky130_fd_io__tk_em2o
XI94 tie_lo_esd net67 / sky130_fd_io__tk_em2o
XI88 pd_h<3> net59 / sky130_fd_io__tk_em2o
XI49 vgnd_io tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
Xn24<2> pad net85 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<1> pad net85 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn24<0> pad net85 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<2> pad net67 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<1> pad net67 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn23<0> pad net67 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn22<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<2> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<1> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn21<0> pad pd_h<3> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn12 pad net61 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<2> pad net69 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<1> pad net69 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn32<0> pad net69 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<2> pad net83 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<1> pad net83 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn33<0> pad net83 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<3> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<2> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<1> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn34<0> pad net77 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<2> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<1> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn11<0> pad pd_h<2> vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn13 pad net59 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
Xn31 pad net73 vgnd_io / sky130_fd_io__com_pddrvr_unit_2_5
xI72 vgnd_io vcc_io condiode
.ENDS
.SUBCKT sky130_fd_io__xres_esd out_h out_vt pad vddio vssd vssio
*.PININFO out_h:B out_vt:B pad:B vddio:B vssd:B vssio:B
Xesd pad out_h out_vt vddio vssd vssd / sky130_fd_io__gpio_buf_localesd
Xpddrvr_strong tie_lo_esd tie_lo_esd pad tie_lo_esd tie_lo_esd tie_lo_esd 
+ vddio vssio vssio / sky130_fd_io__gpio_pddrvr_strong
Xpudrvr_strong pad tie_hi_esd tie_hi_esd tie_hi_esd vddio vssd / 
+ sky130_fd_io__gpio_pudrvr_strong
xI271 vssio vddio condiode
.ENDS
.SUBCKT sky130_fd_io__xres_wpu pad vddio vssd
*.PININFO pad:B vddio:B vssd:B
Xesdr pad net15 / s8_esd_res250only_small
X5kres vddio net15 vssd / sky130_fd_io__com_res_weak
.ENDS
.SUBCKT sky130_fd_io__com_xres_weak_pu ra rb vgnd_io
*.PININFO vgnd_io:I ra:B rb:B
XICEn<3> n<3> / icecap
XICEn<2> n<2> / icecap
XICErb rb / icecap
XICEn<0> n<0> / icecap
XICEn<4> n<4> / icecap
XICEra ra / icecap
XICEnet64 net64 / icecap
XICEn<1> n<1> / icecap
XICEn<5> n<5> / icecap
Xe9 n<0> n<1> / sky130_fd_io__tk_em1s
Xe11 n<2> n<3> / sky130_fd_io__tk_em1s
Xe10 n<1> n<2> / sky130_fd_io__tk_em1s
Xe12 n<3> rb / sky130_fd_io__tk_em1s
Xe13 n<4> n<0> / sky130_fd_io__tk_em1s
Xe14 n<5> n<4> / sky130_fd_io__tk_em1o
rI84 n<0> n<1> mrp1 m=1 w=0.8 l=1.5
rI62 n<3> rb mrp1 m=1 w=0.8 l=1.5
rI82 n<2> n<3> mrp1 m=1 w=0.8 l=1.5
rI85 ra net64 mrp1 m=1 w=0.8 l=50
rI83 n<1> n<2> mrp1 m=1 w=0.8 l=1.5
rI116 net64 n<5> mrp1 m=1 w=0.8 l=12
rI104 n<4> n<0> mrp1 m=1 w=0.8 l=6
rI134 n<5> n<4> mrp1 m=1 w=0.8 l=6
.ENDS
.SUBCKT sky130_fd_io__xres_tk_emlo a b
*.PININFO a:B b:B
rI2 b net8 short
rI1 a net3 short
.ENDS
.SUBCKT sky130_fd_io__xres_tk_emlc a
*.PININFO a:B
rI2 a net7 short
rI1 a net2 short
.ENDS
.SUBCKT sky130_fd_io__xres_rcfilter_lpf_res_sub in out vgnd
*.PININFO in:I out:O vgnd:B
Xe1 in / sky130_fd_io__xres_tk_emlc
Xe2 out net30 / sky130_fd_io__xres_tk_emlo
rropti out net30 mrdn m=1 w=0.5 l=14 isHV=FALSE
rr1 net30 in mrdn m=1 w=0.5 l=47 isHV=FALSE
rropto in in mrdn m=1 w=0.5 l=14 isHV=FALSE
.ENDS
.SUBCKT sky130_fd_io__xres_rcfilter_lpf_rcunit in out vgnd vnb vpwr
*.PININFO in:I out:O vgnd:B vnb:B vpwr:B
Xr1b net14 out vnb / sky130_fd_io__xres_rcfilter_lpf_res_sub
Xr1a in net14 vnb / sky130_fd_io__xres_rcfilter_lpf_res_sub
mI242 vgnd out vgnd vnb nhv m=1 w=7.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI244 vpwr out vpwr vpwr phv m=1 w=7.00 l=4.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__xres_rcfilter_lpf in out vcc_io vssd
*.PININFO in:I out:O vcc_io:B vssd:B
Xe5 net65 net40 / sky130_fd_io__xres_tk_emlo
Xe1 net135 net67 / sky130_fd_io__xres_tk_emlo
Xe4 net43 net65 / sky130_fd_io__xres_tk_emlo
XI200 net59 out / sky130_fd_io__xres_tk_emlo
XI199 net62 out / sky130_fd_io__xres_tk_emlo
XI198 vssd net59 / sky130_fd_io__xres_tk_emlo
XI197 vssd net57 / sky130_fd_io__xres_tk_emlo
XI194 net57 out / sky130_fd_io__xres_tk_emlo
XI193 net45 out / sky130_fd_io__xres_tk_emlo
XI191 net42 out / sky130_fd_io__xres_tk_emlo
XI190 net40 out / sky130_fd_io__xres_tk_emlo
XI187 vssd out / sky130_fd_io__xres_tk_emlo
XI186 vssd net45 / sky130_fd_io__xres_tk_emlo
Xe2 net67 net43 / sky130_fd_io__xres_tk_emlo
XI183 net42 vssd / sky130_fd_io__xres_tk_emlo
XI181 net40 vssd / sky130_fd_io__xres_tk_emlo
XI202 vssd / sky130_fd_io__xres_tk_emlc
XI201 vssd / sky130_fd_io__xres_tk_emlc
XI192 out / sky130_fd_io__xres_tk_emlc
XI189 vssd / sky130_fd_io__xres_tk_emlc
XI188 vssd / sky130_fd_io__xres_tk_emlc
XI180 net40 / sky130_fd_io__xres_tk_emlc
XI182 net42 / sky130_fd_io__xres_tk_emlc
Xe3 net43 / sky130_fd_io__xres_tk_emlc
XI172 in net135 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI184 vssd net57 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI185 vssd net45 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI196 vssd net62 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI195 vssd net59 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI179 net43 net65 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI178 net65 net40 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI177 net40 net42 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI176 net42 out vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI175 net67 net43 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI174 net43 net43 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
XI173 net135 net67 vssd vssd vcc_io / sky130_fd_io__xres_rcfilter_lpf_rcunit
.ENDS
.SUBCKT sky130_fd_io__xres_inv_hys in_h out_h vcc_io vssd
*.PININFO in_h:I vcc_io:I vssd:I out_h:O
XICEpmid1 pmid1 / icecap
XICEout_h_n out_h_n / icecap
XICEout_h out_h / icecap
XICEin_h in_h / icecap
XICEnmid1 nmid1 / icecap
mI7 pmid1 in_h vcc_io vcc_io phv m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI8 out_h_n in_h pmid1 vcc_io phv m=1 w=3.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI9 out_h out_h_n vcc_io vcc_io phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI10 pmid1 out_h vcc_io vcc_io phv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI4 out_h_n in_h nmid1 vssd nhv m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI5 nmid1 in_h vssd vssd nhv m=1 w=1.00 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI6 out_h out_h_n vssd vssd nhv m=1 w=1.00 l=0.50 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
mI11 nmid1 out_h vssd vssd nhv m=1 w=0.42 l=1.00 mult=1 sa=265e-3 sb=265e-3 
+ sd=280e-3 topography=normal area=0.063 perim=1.14
.ENDS
.SUBCKT sky130_fd_io__top_xres4v2 amuxbus_a amuxbus_b disable_pullup_h 
+ en_vddio_sig_h enable_h enable_vddio filt_in_h inp_sel_h pad pad_a_esd_h 
+ pullup_h tie_hi_esd tie_lo_esd tie_weak_hi_h vccd vcchib vdda vddio vddio_q 
+ vssa vssd vssio vssio_q vswitch xres_h_n
*.PININFO disable_pullup_h:I en_vddio_sig_h:I enable_h:I enable_vddio:I 
*.PININFO filt_in_h:I inp_sel_h:I vccd:I vcchib:I vdda:I vddio:I vddio_q:I 
*.PININFO vssa:I vssd:I vssio:I vssio_q:I vswitch:I tie_hi_esd:O tie_lo_esd:O 
*.PININFO xres_h_n:O amuxbus_a:B amuxbus_b:B pad:B pad_a_esd_h:B pullup_h:B 
*.PININFO tie_weak_hi_h:B
XI326 vssio tie_lo_esd / sky130_fd_io__tk_tie_r_out_esd
XI49 vddio tie_hi_esd / sky130_fd_io__tk_tie_r_out_esd
Xgpio_inbuf enable_h enable_vddio net79 net83 in_h vcchib vddio_q vssd 
+ en_vddio_sig_h en_vddio_sig_h_n / sky130_fd_io__xres4v2_in_buf
Xxresesd in_h net86 pad vddio vssd vssio / sky130_fd_io__xres_esd
Xweakpullup tie_weak_hi_h vddio vssd / sky130_fd_io__xres_wpu
Xesd_res pad pad_a_esd_h / s8_esd_res250only_small
XI335 net97 pullup_h vssd / sky130_fd_io__com_xres_weak_pu
XI363 inp_sel_h inp_sel_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x2
XI334 net103 net107 vssd vddio / sky130_fd_io__hvsbt_inv_x2
XI333 disable_pullup_h net103 vssd vddio / sky130_fd_io__hvsbt_inv_x2
XI374 en_vddio_sig_h en_vddio_sig_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x2
mI361 net124 inp_sel_h_n filt_in_h vddio_q phv m=1 w=3.00 l=0.50 mult=1 
+ sa=265e-3 sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI358 net124 inp_sel_h net79 vddio_q phv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI332 net97 net107 vddio vddio phv m=4 w=5.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI360 net124 inp_sel_h filt_in_h vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
mI357 net124 inp_sel_h_n net79 vssd nhv m=1 w=3.00 l=0.50 mult=1 sa=265e-3 
+ sb=265e-3 sd=280e-3 topography=normal area=0.063 perim=1.14
XI368 net124 out_rcfilt_h vddio_q vssd / sky130_fd_io__xres_rcfilter_lpf
XI367 out_rcfilt_h out_hysbuf_h vddio_q vssd / sky130_fd_io__xres_inv_hys
XI365 out_hysbuf_h out_h_n vssd vddio_q / sky130_fd_io__hvsbt_inv_x1
XI364<1> out_h_n xres_h_n net039<0> net038<0> / sky130_fd_io__hvsbt_inv_x4
XI364<0> out_h_n xres_h_n net039<1> net038<1> / sky130_fd_io__hvsbt_inv_x4
.ENDS

.SUBCKT condiode pin0 pin1
.ENDS condiode
