DFFRAM.extracted.ngspice