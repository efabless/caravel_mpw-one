*** UC SPICE *** , MIN_RESIST 4.0, MIN_CAPAC 0.1FF

* Most models come from here:

 .lib ~/foss/pdks/sky130A/libs.tech/ngspice/sky130.lib.spice tt

* This device is also missing from the libraries:

* .include ./sky130_fd_io__condiode.spice
 .include ./sky130_fd_pr__model__parasitic__diode_ps2nw.spice 
 .include ./sky130_fd_pr__model__parasitic__diode_pw2dn.spice
 .include ./sky130_fd_pr__model__parasitic__diode_ps2dn.spice

vvss		VSS		0 		dc 	0
vvdd3v3		VDD3V3		0 		pwl	0 0 2u 3.3  1m 3.3

RL		VDD3V3		0		1

X1 		VSS 		VDD3V3 		sky130_fd_pr__model__parasitic__diode_ps2dn  
X2 		VSS 		VDD3V3 		sky130_fd_pr__model__parasitic__diode_ps2nw  
X3 		VSS 		VDD3V3 		sky130_fd_pr__model__parasitic__diode_pw2dn  

.SAVE i(vvdd3v3) v(vdd3v3) 
.TRAN 10n 15u

.END

