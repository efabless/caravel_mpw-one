*SPICE netlist created from verilog structural netlist module ring_osc2x13 by vlog2Spice (qflow)
* Warning: This file contains <> array delimiters in net names_
* Note: Library sky130_fd_sc_hd_spice has been removed;  reference library as an
* include file from the testbench instead_

.subckt ring_osc2x13 VPB VGND clockp<0> clockp<1> reset trim<0> trim<1>
+ trim<2> trim<3> trim<4> trim<5> trim<6> trim<7> trim<8> trim<9>
+ trim<10> trim<11> trim<12> trim<13> trim<14> trim<15> trim<16> trim<17>
+ trim<18> trim<19> trim<20> trim<21> trim<22> trim<23> trim<24> trim<25>
+ 

X_1_ _0_<0> VGND VGND VPB VPB clockp<0> sky130_fd_sc_hd__buf_2
X_2_ _0_<1> VGND VGND VPB VPB clockp<1> sky130_fd_sc_hd__buf_2
Xdstage<0>_id_delaybuf0  dstage<0>_id_in VGND VGND VPB VPB dstage<0>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<0>_id_delaybuf1  dstage<0>_id_ts VGND VGND VPB VPB dstage<0>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<0>_id_delayen0  dstage<0>_id_d2 trim<0> VGND VGND VPB VPB 
+ dstage<0>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<0>_id_delayen1  dstage<0>_id_d0 trim<13> VGND VGND VPB VPB 
+ dstage<0>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<0>_id_delayenb0  dstage<0>_id_ts trim<0> VGND VGND VPB VPB 
+ dstage<0>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<0>_id_delayenb1  dstage<0>_id_ts trim<13> VGND VGND VPB VPB 
+ dstage<0>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<0>_id_delayint0  dstage<0>_id_d1 VGND VGND VPB VPB dstage<0>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<10>_id_delaybuf0  dstage<10>_id_in VGND VGND VPB VPB dstage<10>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<10>_id_delaybuf1  dstage<10>_id_ts VGND VGND VPB VPB dstage<10>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<10>_id_delayen0  dstage<10>_id_d2 trim<10> VGND VGND VPB VPB 
+ dstage<10>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<10>_id_delayen1  dstage<10>_id_d0 trim<23> VGND VGND VPB VPB 
+ dstage<10>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<10>_id_delayenb0  dstage<10>_id_ts trim<10> VGND VGND VPB VPB 
+ dstage<10>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<10>_id_delayenb1  dstage<10>_id_ts trim<23> VGND VGND VPB VPB 
+ dstage<10>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<10>_id_delayint0  dstage<10>_id_d1 VGND VGND VPB VPB dstage<10>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<11>_id_delaybuf0  dstage<10>_id_out VGND VGND VPB VPB dstage<11>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<11>_id_delaybuf1  dstage<11>_id_ts VGND VGND VPB VPB dstage<11>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<11>_id_delayen0  dstage<11>_id_d2 trim<11> VGND VGND VPB VPB 
+ dstage<11>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<11>_id_delayen1  dstage<11>_id_d0 trim<24> VGND VGND VPB VPB 
+ dstage<11>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<11>_id_delayenb0  dstage<11>_id_ts trim<11> VGND VGND VPB VPB 
+ dstage<11>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<11>_id_delayenb1  dstage<11>_id_ts trim<24> VGND VGND VPB VPB 
+ dstage<11>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<11>_id_delayint0  dstage<11>_id_d1 VGND VGND VPB VPB dstage<11>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<1>_id_delaybuf0  dstage<0>_id_out VGND VGND VPB VPB dstage<1>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<1>_id_delaybuf1  dstage<1>_id_ts VGND VGND VPB VPB dstage<1>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<1>_id_delayen0  dstage<1>_id_d2 trim<1> VGND VGND VPB VPB 
+ dstage<1>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<1>_id_delayen1  dstage<1>_id_d0 trim<14> VGND VGND VPB VPB 
+ dstage<1>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<1>_id_delayenb0  dstage<1>_id_ts trim<1> VGND VGND VPB VPB 
+ dstage<1>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<1>_id_delayenb1  dstage<1>_id_ts trim<14> VGND VGND VPB VPB 
+ dstage<1>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<1>_id_delayint0  dstage<1>_id_d1 VGND VGND VPB VPB dstage<1>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<2>_id_delaybuf0  dstage<1>_id_out VGND VGND VPB VPB dstage<2>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<2>_id_delaybuf1  dstage<2>_id_ts VGND VGND VPB VPB dstage<2>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<2>_id_delayen0  dstage<2>_id_d2 trim<2> VGND VGND VPB VPB 
+ dstage<2>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<2>_id_delayen1  dstage<2>_id_d0 trim<15> VGND VGND VPB VPB 
+ dstage<2>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<2>_id_delayenb0  dstage<2>_id_ts trim<2> VGND VGND VPB VPB 
+ dstage<2>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<2>_id_delayenb1  dstage<2>_id_ts trim<15> VGND VGND VPB VPB 
+ dstage<2>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<2>_id_delayint0  dstage<2>_id_d1 VGND VGND VPB VPB dstage<2>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<3>_id_delaybuf0  dstage<2>_id_out VGND VGND VPB VPB dstage<3>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<3>_id_delaybuf1  dstage<3>_id_ts VGND VGND VPB VPB dstage<3>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<3>_id_delayen0  dstage<3>_id_d2 trim<3> VGND VGND VPB VPB 
+ dstage<3>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<3>_id_delayen1  dstage<3>_id_d0 trim<16> VGND VGND VPB VPB 
+ dstage<3>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<3>_id_delayenb0  dstage<3>_id_ts trim<3> VGND VGND VPB VPB 
+ dstage<3>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<3>_id_delayenb1  dstage<3>_id_ts trim<16> VGND VGND VPB VPB 
+ dstage<3>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<3>_id_delayint0  dstage<3>_id_d1 VGND VGND VPB VPB dstage<3>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<4>_id_delaybuf0  dstage<3>_id_out VGND VGND VPB VPB dstage<4>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<4>_id_delaybuf1  dstage<4>_id_ts VGND VGND VPB VPB dstage<4>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<4>_id_delayen0  dstage<4>_id_d2 trim<4> VGND VGND VPB VPB 
+ dstage<4>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<4>_id_delayen1  dstage<4>_id_d0 trim<17> VGND VGND VPB VPB 
+ dstage<4>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<4>_id_delayenb0  dstage<4>_id_ts trim<4> VGND VGND VPB VPB 
+ dstage<4>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<4>_id_delayenb1  dstage<4>_id_ts trim<17> VGND VGND VPB VPB 
+ dstage<4>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<4>_id_delayint0  dstage<4>_id_d1 VGND VGND VPB VPB dstage<4>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<5>_id_delaybuf0  dstage<4>_id_out VGND VGND VPB VPB dstage<5>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<5>_id_delaybuf1  dstage<5>_id_ts VGND VGND VPB VPB dstage<5>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<5>_id_delayen0  dstage<5>_id_d2 trim<5> VGND VGND VPB VPB 
+ dstage<5>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<5>_id_delayen1  dstage<5>_id_d0 trim<18> VGND VGND VPB VPB 
+ dstage<5>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<5>_id_delayenb0  dstage<5>_id_ts trim<5> VGND VGND VPB VPB 
+ dstage<5>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<5>_id_delayenb1  dstage<5>_id_ts trim<18> VGND VGND VPB VPB 
+ dstage<5>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<5>_id_delayint0  dstage<5>_id_d1 VGND VGND VPB VPB dstage<5>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<6>_id_delaybuf0  dstage<5>_id_out VGND VGND VPB VPB dstage<6>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<6>_id_delaybuf1  dstage<6>_id_ts VGND VGND VPB VPB dstage<6>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<6>_id_delayen0  dstage<6>_id_d2 trim<6> VGND VGND VPB VPB 
+ dstage<6>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<6>_id_delayen1  dstage<6>_id_d0 trim<19> VGND VGND VPB VPB 
+ dstage<6>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<6>_id_delayenb0  dstage<6>_id_ts trim<6> VGND VGND VPB VPB 
+ dstage<6>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<6>_id_delayenb1  dstage<6>_id_ts trim<19> VGND VGND VPB VPB 
+ dstage<6>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<6>_id_delayint0  dstage<6>_id_d1 VGND VGND VPB VPB dstage<6>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<7>_id_delaybuf0  dstage<6>_id_out VGND VGND VPB VPB dstage<7>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<7>_id_delaybuf1  dstage<7>_id_ts VGND VGND VPB VPB dstage<7>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<7>_id_delayen0  dstage<7>_id_d2 trim<7> VGND VGND VPB VPB 
+ dstage<7>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<7>_id_delayen1  dstage<7>_id_d0 trim<20> VGND VGND VPB VPB 
+ dstage<7>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<7>_id_delayenb0  dstage<7>_id_ts trim<7> VGND VGND VPB VPB 
+ dstage<7>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<7>_id_delayenb1  dstage<7>_id_ts trim<20> VGND VGND VPB VPB 
+ dstage<7>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<7>_id_delayint0  dstage<7>_id_d1 VGND VGND VPB VPB dstage<7>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<8>_id_delaybuf0  dstage<7>_id_out VGND VGND VPB VPB dstage<8>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<8>_id_delaybuf1  dstage<8>_id_ts VGND VGND VPB VPB dstage<8>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<8>_id_delayen0  dstage<8>_id_d2 trim<8> VGND VGND VPB VPB 
+ dstage<8>_id_out
+ sky130_fd_sc_hd__einvp_2
Xdstage<8>_id_delayen1  dstage<8>_id_d0 trim<21> VGND VGND VPB VPB 
+ dstage<8>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<8>_id_delayenb0  dstage<8>_id_ts trim<8> VGND VGND VPB VPB 
+ dstage<8>_id_out
+ sky130_fd_sc_hd__einvn_8
Xdstage<8>_id_delayenb1  dstage<8>_id_ts trim<21> VGND VGND VPB VPB 
+ dstage<8>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<8>_id_delayint0  dstage<8>_id_d1 VGND VGND VPB VPB dstage<8>_id_d2 sky130_fd_sc_hd__clkinv_1
Xdstage<9>_id_delaybuf0  dstage<8>_id_out VGND VGND VPB VPB dstage<9>_id_ts sky130_fd_sc_hd__clkbuf_2
Xdstage<9>_id_delaybuf1  dstage<9>_id_ts VGND VGND VPB VPB dstage<9>_id_d0 sky130_fd_sc_hd__clkbuf_1
Xdstage<9>_id_delayen0  dstage<9>_id_d2 trim<9> VGND VGND VPB VPB 
+ dstage<10>_id_in
+ sky130_fd_sc_hd__einvp_2
Xdstage<9>_id_delayen1  dstage<9>_id_d0 trim<22> VGND VGND VPB VPB 
+ dstage<9>_id_d1
+ sky130_fd_sc_hd__einvp_2
Xdstage<9>_id_delayenb0  dstage<9>_id_ts trim<9> VGND VGND VPB VPB 
+ dstage<10>_id_in
+ sky130_fd_sc_hd__einvn_8
Xdstage<9>_id_delayenb1  dstage<9>_id_ts trim<22> VGND VGND VPB VPB 
+ dstage<9>_id_d1
+ sky130_fd_sc_hd__einvn_4
Xdstage<9>_id_delayint0  dstage<9>_id_d1 VGND VGND VPB VPB dstage<9>_id_d2 sky130_fd_sc_hd__clkinv_1
Xibufp00 dstage<0>_id_in VGND VGND VPB VPB c<0> sky130_fd_sc_hd__clkinv_2
Xibufp01 c<0> VGND VGND VPB VPB _0_<0> sky130_fd_sc_hd__clkinv_8
Xibufp10 dstage<5>_id_out VGND VGND VPB VPB c<1> sky130_fd_sc_hd__clkinv_2
Xibufp11 c<1> VGND VGND VPB VPB _0_<1> sky130_fd_sc_hd__clkinv_8
Xiss_const1  VGND VGND VPB VPB iss_one _noconnect_1_ sky130_fd_sc_hd__conb_1
Xiss_ctrlen0  reset trim<12> VGND VGND VPB VPB 
+ iss_ctrl0
+ sky130_fd_sc_hd__or2_2
Xiss_delaybuf0  dstage<11>_id_out VGND VGND VPB VPB iss_d0 sky130_fd_sc_hd__clkbuf_1
Xiss_delayen0  iss_d2 trim<12> VGND VGND VPB VPB 
+ dstage<0>_id_in
+ sky130_fd_sc_hd__einvp_2
Xiss_delayen1  iss_d0 trim<25> VGND VGND VPB VPB 
+ iss_d1
+ sky130_fd_sc_hd__einvp_2
Xiss_delayenb0  dstage<11>_id_out iss_ctrl0 VGND VGND VPB VPB 
+ dstage<0>_id_in
+ sky130_fd_sc_hd__einvn_8
Xiss_delayenb1  dstage<11>_id_out trim<25> VGND VGND VPB VPB 
+ iss_d1
+ sky130_fd_sc_hd__einvn_4
Xiss_delayint0  iss_d1 VGND VGND VPB VPB iss_d2 sky130_fd_sc_hd__clkinv_1
Xiss_reseten0  iss_one reset VGND VGND VPB VPB 
+ dstage<0>_id_in
+ sky130_fd_sc_hd__einvp_1
Xantenna_0 reset VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<25> trim<25> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<24> trim<24> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<23> trim<23> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<22> trim<22> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<21> trim<21> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<20> trim<20> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<19> trim<19> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<18> trim<18> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<17> trim<17> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<16> trim<16> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<15> trim<15> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<14> trim<14> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<13> trim<13> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<12> trim<12> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<11> trim<11> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<10> trim<10> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<9> trim<9> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<8> trim<8> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<7> trim<7> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<6> trim<6> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<5> trim<5> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<4> trim<4> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<3> trim<3> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<2> trim<2> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<1> trim<1> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2
Xantenna_1<0> trim<0> VGND VGND VPB VPB sky130_fd_sc_hd__diode_2

.ends
.end
