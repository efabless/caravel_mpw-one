* SKY130 Spice File.
* RF MOS Parameters
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_b__wafer.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt_b__wafer.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_g5v0d10v5_b__wafer.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_b__wafer.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_01v8_lvt__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_nfet_g5v0d10v5__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8__mismatch.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_mvt__wafer_discrete.corner.spice"
.include "../../../../libs.ref/sky130_fd_pr/spice/sky130_fd_pr__rf_pfet_01v8_mvt__mismatch.corner.spice"
