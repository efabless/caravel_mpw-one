magic
tech sky130A
magscale 1 2
timestamp 1606789161
<< checkpaint >>
rect -1260 -1260 42396 42300
<< locali >>
rect 19585 28595 19619 28697
rect 18481 11187 18515 11425
<< viali >>
rect 20597 29853 20631 29887
rect 14985 29785 15019 29819
rect 15445 29785 15479 29819
rect 18941 29785 18975 29819
rect 19861 29785 19895 29819
rect 20413 29785 20447 29819
rect 22621 29785 22655 29819
rect 26393 29785 26427 29819
rect 28969 29785 29003 29819
rect 21149 29717 21183 29751
rect 21701 29717 21735 29751
rect 22713 29717 22747 29751
rect 21609 29649 21643 29683
rect 14801 29581 14835 29615
rect 15537 29581 15571 29615
rect 19033 29581 19067 29615
rect 19677 29581 19711 29615
rect 26209 29581 26243 29615
rect 29061 29581 29095 29615
rect 18849 29309 18883 29343
rect 20045 29309 20079 29343
rect 14525 29241 14559 29275
rect 16089 29241 16123 29275
rect 20137 29241 20171 29275
rect 20781 29241 20815 29275
rect 21609 29241 21643 29275
rect 13605 29173 13639 29207
rect 14433 29173 14467 29207
rect 15169 29173 15203 29207
rect 15997 29173 16031 29207
rect 17561 29173 17595 29207
rect 19033 29173 19067 29207
rect 19585 29173 19619 29207
rect 20689 29173 20723 29207
rect 21517 29173 21551 29207
rect 22713 29173 22747 29207
rect 23357 29173 23391 29207
rect 24277 29173 24311 29207
rect 25473 29173 25507 29207
rect 26209 29173 26243 29207
rect 29245 29173 29279 29207
rect 13697 29105 13731 29139
rect 15261 29105 15295 29139
rect 23633 29105 23667 29139
rect 24829 29105 24863 29139
rect 26393 29105 26427 29139
rect 24093 29037 24127 29071
rect 24921 29037 24955 29071
rect 27129 29037 27163 29071
rect 27221 29037 27255 29071
rect 29061 29037 29095 29071
rect 24461 28833 24495 28867
rect 28141 28833 28175 28867
rect 14801 28765 14835 28799
rect 18481 28765 18515 28799
rect 19677 28765 19711 28799
rect 22897 28765 22931 28799
rect 25565 28765 25599 28799
rect 27497 28765 27531 28799
rect 11673 28697 11707 28731
rect 14065 28697 14099 28731
rect 14985 28697 15019 28731
rect 15445 28697 15479 28731
rect 16733 28697 16767 28731
rect 19585 28697 19619 28731
rect 19861 28697 19895 28731
rect 20689 28697 20723 28731
rect 22161 28697 22195 28731
rect 23633 28697 23667 28731
rect 24369 28697 24403 28731
rect 26301 28697 26335 28731
rect 26945 28697 26979 28731
rect 27405 28697 27439 28731
rect 27957 28697 27991 28731
rect 29153 28697 29187 28731
rect 17929 28629 17963 28663
rect 22805 28629 22839 28663
rect 23725 28629 23759 28663
rect 25473 28629 25507 28663
rect 26393 28629 26427 28663
rect 16733 28561 16767 28595
rect 18389 28561 18423 28595
rect 19585 28561 19619 28595
rect 21977 28561 22011 28595
rect 11765 28493 11799 28527
rect 19953 28493 19987 28527
rect 29245 28493 29279 28527
rect 20873 28289 20907 28323
rect 23265 28221 23299 28255
rect 25749 28221 25783 28255
rect 26945 28221 26979 28255
rect 14157 28153 14191 28187
rect 14617 28153 14651 28187
rect 15445 28153 15479 28187
rect 15905 28153 15939 28187
rect 18665 28153 18699 28187
rect 22805 28153 22839 28187
rect 14709 28085 14743 28119
rect 15997 28085 16031 28119
rect 17193 28085 17227 28119
rect 17745 28085 17779 28119
rect 18573 28085 18607 28119
rect 19217 28085 19251 28119
rect 19861 28085 19895 28119
rect 20137 28085 20171 28119
rect 20781 28085 20815 28119
rect 23357 28085 23391 28119
rect 24461 28085 24495 28119
rect 25381 28085 25415 28119
rect 26485 28085 26519 28119
rect 27037 28085 27071 28119
rect 17009 28017 17043 28051
rect 17837 28017 17871 28051
rect 20597 28017 20631 28051
rect 28049 28017 28083 28051
rect 28785 28017 28819 28051
rect 28141 27949 28175 27983
rect 28877 27949 28911 27983
rect 16733 27745 16767 27779
rect 19585 27677 19619 27711
rect 19861 27677 19895 27711
rect 19953 27677 19987 27711
rect 20321 27677 20355 27711
rect 27405 27677 27439 27711
rect 12225 27609 12259 27643
rect 14709 27609 14743 27643
rect 16641 27609 16675 27643
rect 17285 27609 17319 27643
rect 17929 27609 17963 27643
rect 18297 27609 18331 27643
rect 18481 27609 18515 27643
rect 19769 27609 19803 27643
rect 21793 27609 21827 27643
rect 22621 27609 22655 27643
rect 23449 27609 23483 27643
rect 24185 27609 24219 27643
rect 25381 27609 25415 27643
rect 25841 27609 25875 27643
rect 26761 27609 26795 27643
rect 27865 27609 27899 27643
rect 29153 27609 29187 27643
rect 18021 27541 18055 27575
rect 21885 27541 21919 27575
rect 22713 27541 22747 27575
rect 23357 27541 23391 27575
rect 24277 27541 24311 27575
rect 29153 27473 29187 27507
rect 12409 27405 12443 27439
rect 14893 27405 14927 27439
rect 25197 27405 25231 27439
rect 18205 27201 18239 27235
rect 27129 27133 27163 27167
rect 13789 27065 13823 27099
rect 19677 27065 19711 27099
rect 23817 27065 23851 27099
rect 24645 27065 24679 27099
rect 26669 27065 26703 27099
rect 27221 27065 27255 27099
rect 28417 27065 28451 27099
rect 28969 27065 29003 27099
rect 11305 26997 11339 27031
rect 17009 26997 17043 27031
rect 18113 26997 18147 27031
rect 22713 26997 22747 27031
rect 23081 26997 23115 27031
rect 23725 26997 23759 27031
rect 24553 26997 24587 27031
rect 25565 26997 25599 27031
rect 11581 26929 11615 26963
rect 13329 26929 13363 26963
rect 14065 26929 14099 26963
rect 15813 26929 15847 26963
rect 16733 26929 16767 26963
rect 17101 26929 17135 26963
rect 17469 26929 17503 26963
rect 17929 26929 17963 26963
rect 18941 26929 18975 26963
rect 19125 26929 19159 26963
rect 19309 26929 19343 26963
rect 20137 26929 20171 26963
rect 20505 26929 20539 26963
rect 20873 26929 20907 26963
rect 22529 26929 22563 26963
rect 28877 26929 28911 26963
rect 16917 26861 16951 26895
rect 19217 26861 19251 26895
rect 20321 26861 20355 26895
rect 20413 26861 20447 26895
rect 25657 26861 25691 26895
rect 20321 26657 20355 26691
rect 22805 26657 22839 26691
rect 26393 26657 26427 26691
rect 28601 26657 28635 26691
rect 11949 26589 11983 26623
rect 17837 26589 17871 26623
rect 20413 26589 20447 26623
rect 20505 26589 20539 26623
rect 21517 26589 21551 26623
rect 22069 26589 22103 26623
rect 23725 26589 23759 26623
rect 27681 26589 27715 26623
rect 27957 26589 27991 26623
rect 28509 26589 28543 26623
rect 12501 26521 12535 26555
rect 12685 26521 12719 26555
rect 12869 26521 12903 26555
rect 13237 26521 13271 26555
rect 15261 26521 15295 26555
rect 15905 26521 15939 26555
rect 17653 26521 17687 26555
rect 17745 26521 17779 26555
rect 20137 26521 20171 26555
rect 21701 26521 21735 26555
rect 22529 26521 22563 26555
rect 22713 26521 22747 26555
rect 23909 26521 23943 26555
rect 25381 26521 25415 26555
rect 25933 26521 25967 26555
rect 26117 26521 26151 26555
rect 27037 26521 27071 26555
rect 29153 26521 29187 26555
rect 13329 26453 13363 26487
rect 17469 26453 17503 26487
rect 18205 26453 18239 26487
rect 20873 26453 20907 26487
rect 24277 26453 24311 26487
rect 25197 26453 25231 26487
rect 29245 26385 29279 26419
rect 15353 26317 15387 26351
rect 15997 26317 16031 26351
rect 12593 26113 12627 26147
rect 24921 26113 24955 26147
rect 15997 26045 16031 26079
rect 26945 26045 26979 26079
rect 28877 26045 28911 26079
rect 13973 25977 14007 26011
rect 15261 25977 15295 26011
rect 15353 25977 15387 26011
rect 25381 25977 25415 26011
rect 26485 25977 26519 26011
rect 27037 25977 27071 26011
rect 28969 25977 29003 26011
rect 11673 25909 11707 25943
rect 12777 25909 12811 25943
rect 13237 25909 13271 25943
rect 14433 25909 14467 25943
rect 14617 25909 14651 25943
rect 14801 25909 14835 25943
rect 15905 25909 15939 25943
rect 16917 25909 16951 25943
rect 17929 25909 17963 25943
rect 18113 25909 18147 25943
rect 18665 25909 18699 25943
rect 19309 25909 19343 25943
rect 20321 25909 20355 25943
rect 21425 25909 21459 25943
rect 23173 25909 23207 25943
rect 23357 25909 23391 25943
rect 25289 25909 25323 25943
rect 25657 25909 25691 25943
rect 25749 25909 25783 25943
rect 28417 25909 28451 25943
rect 16733 25841 16767 25875
rect 17101 25841 17135 25875
rect 17469 25841 17503 25875
rect 18297 25841 18331 25875
rect 19125 25841 19159 25875
rect 20137 25841 20171 25875
rect 20689 25841 20723 25875
rect 21241 25841 21275 25875
rect 21793 25841 21827 25875
rect 23725 25841 23759 25875
rect 11765 25773 11799 25807
rect 17009 25773 17043 25807
rect 18205 25773 18239 25807
rect 19401 25773 19435 25807
rect 13053 25569 13087 25603
rect 15721 25569 15755 25603
rect 18849 25569 18883 25603
rect 19861 25569 19895 25603
rect 24461 25569 24495 25603
rect 25841 25569 25875 25603
rect 26853 25569 26887 25603
rect 12777 25501 12811 25535
rect 13973 25501 14007 25535
rect 17377 25501 17411 25535
rect 18205 25501 18239 25535
rect 20045 25501 20079 25535
rect 28969 25501 29003 25535
rect 29245 25501 29279 25535
rect 11949 25433 11983 25467
rect 12961 25433 12995 25467
rect 14801 25433 14835 25467
rect 15445 25433 15479 25467
rect 15629 25433 15663 25467
rect 17193 25433 17227 25467
rect 17285 25433 17319 25467
rect 18352 25433 18386 25467
rect 19953 25433 19987 25467
rect 21333 25433 21367 25467
rect 21517 25433 21551 25467
rect 22345 25433 22379 25467
rect 22529 25433 22563 25467
rect 23817 25433 23851 25467
rect 25197 25433 25231 25467
rect 25344 25433 25378 25467
rect 27221 25433 27255 25467
rect 27589 25433 27623 25467
rect 27681 25433 27715 25467
rect 28325 25433 28359 25467
rect 14525 25365 14559 25399
rect 14985 25365 15019 25399
rect 17009 25365 17043 25399
rect 17745 25365 17779 25399
rect 18573 25365 18607 25399
rect 19677 25365 19711 25399
rect 20413 25365 20447 25399
rect 21885 25365 21919 25399
rect 22897 25365 22931 25399
rect 24185 25365 24219 25399
rect 25565 25365 25599 25399
rect 27037 25365 27071 25399
rect 18481 25297 18515 25331
rect 12133 25229 12167 25263
rect 23955 25229 23989 25263
rect 24093 25229 24127 25263
rect 25473 25229 25507 25263
rect 21241 25025 21275 25059
rect 22621 25025 22655 25059
rect 24001 25025 24035 25059
rect 24369 25025 24403 25059
rect 28049 25025 28083 25059
rect 17009 24957 17043 24991
rect 20873 24957 20907 24991
rect 22510 24957 22544 24991
rect 14341 24889 14375 24923
rect 16880 24889 16914 24923
rect 17101 24889 17135 24923
rect 18205 24889 18239 24923
rect 18941 24889 18975 24923
rect 19401 24889 19435 24923
rect 20965 24889 20999 24923
rect 22713 24889 22747 24923
rect 23081 24889 23115 24923
rect 24093 24889 24127 24923
rect 25933 24889 25967 24923
rect 29061 24889 29095 24923
rect 11305 24821 11339 24855
rect 14249 24821 14283 24855
rect 14525 24821 14559 24855
rect 15813 24821 15847 24855
rect 20137 24821 20171 24855
rect 20744 24821 20778 24855
rect 22345 24821 22379 24855
rect 23872 24821 23906 24855
rect 25105 24821 25139 24855
rect 26025 24821 26059 24855
rect 27957 24821 27991 24855
rect 28601 24821 28635 24855
rect 11581 24753 11615 24787
rect 13329 24753 13363 24787
rect 15629 24753 15663 24787
rect 16181 24753 16215 24787
rect 16733 24753 16767 24787
rect 18481 24753 18515 24787
rect 18573 24753 18607 24787
rect 19769 24753 19803 24787
rect 20597 24753 20631 24787
rect 23725 24753 23759 24787
rect 24921 24753 24955 24787
rect 25473 24753 25507 24787
rect 26485 24753 26519 24787
rect 29153 24753 29187 24787
rect 17377 24685 17411 24719
rect 18389 24685 18423 24719
rect 19585 24685 19619 24719
rect 19677 24685 19711 24719
rect 26945 24685 26979 24719
rect 27037 24685 27071 24719
rect 21517 24481 21551 24515
rect 25197 24481 25231 24515
rect 27773 24481 27807 24515
rect 15261 24413 15295 24447
rect 17101 24413 17135 24447
rect 18297 24413 18331 24447
rect 19033 24413 19067 24447
rect 20781 24413 20815 24447
rect 24461 24413 24495 24447
rect 29429 24413 29463 24447
rect 12041 24345 12075 24379
rect 12225 24345 12259 24379
rect 13973 24345 14007 24379
rect 15169 24345 15203 24379
rect 15813 24345 15847 24379
rect 17285 24345 17319 24379
rect 18636 24345 18670 24379
rect 19585 24345 19619 24379
rect 20229 24345 20263 24379
rect 20413 24345 20447 24379
rect 21241 24345 21275 24379
rect 21425 24345 21459 24379
rect 23173 24345 23207 24379
rect 25381 24345 25415 24379
rect 26301 24345 26335 24379
rect 26485 24345 26519 24379
rect 26853 24345 26887 24379
rect 26945 24345 26979 24379
rect 27957 24345 27991 24379
rect 28141 24345 28175 24379
rect 28509 24345 28543 24379
rect 29245 24345 29279 24379
rect 15960 24277 15994 24311
rect 16181 24277 16215 24311
rect 17653 24277 17687 24311
rect 23320 24277 23354 24311
rect 23541 24277 23575 24311
rect 28417 24277 28451 24311
rect 16273 24209 16307 24243
rect 18573 24209 18607 24243
rect 24553 24209 24587 24243
rect 12317 24141 12351 24175
rect 14065 24141 14099 24175
rect 16089 24141 16123 24175
rect 18435 24141 18469 24175
rect 19677 24141 19711 24175
rect 23449 24141 23483 24175
rect 23817 24141 23851 24175
rect 26117 24141 26151 24175
rect 14433 23937 14467 23971
rect 16089 23937 16123 23971
rect 21222 23937 21256 23971
rect 29245 23937 29279 23971
rect 17239 23869 17273 23903
rect 17377 23869 17411 23903
rect 21333 23869 21367 23903
rect 11581 23801 11615 23835
rect 12869 23801 12903 23835
rect 14709 23801 14743 23835
rect 17469 23801 17503 23835
rect 18389 23801 18423 23835
rect 18941 23801 18975 23835
rect 20045 23801 20079 23835
rect 21425 23801 21459 23835
rect 23909 23801 23943 23835
rect 24645 23801 24679 23835
rect 25197 23801 25231 23835
rect 25657 23801 25691 23835
rect 28509 23801 28543 23835
rect 12041 23733 12075 23767
rect 12225 23733 12259 23767
rect 12409 23733 12443 23767
rect 13053 23733 13087 23767
rect 13513 23733 13547 23767
rect 14801 23733 14835 23767
rect 15169 23733 15203 23767
rect 15353 23733 15387 23767
rect 15997 23733 16031 23767
rect 18481 23733 18515 23767
rect 20137 23733 20171 23767
rect 20597 23733 20631 23767
rect 21793 23733 21827 23767
rect 22529 23733 22563 23767
rect 22897 23733 22931 23767
rect 23541 23733 23575 23767
rect 25473 23733 25507 23767
rect 26117 23733 26151 23767
rect 26945 23733 26979 23767
rect 27037 23733 27071 23767
rect 27957 23733 27991 23767
rect 29153 23733 29187 23767
rect 17101 23665 17135 23699
rect 21057 23665 21091 23699
rect 22345 23665 22379 23699
rect 23357 23665 23391 23699
rect 28417 23665 28451 23699
rect 13605 23597 13639 23631
rect 17745 23597 17779 23631
rect 26209 23597 26243 23631
rect 16273 23393 16307 23427
rect 17285 23393 17319 23427
rect 18205 23393 18239 23427
rect 19677 23393 19711 23427
rect 20873 23393 20907 23427
rect 25473 23393 25507 23427
rect 12225 23325 12259 23359
rect 16365 23325 16399 23359
rect 20229 23325 20263 23359
rect 22345 23325 22379 23359
rect 24001 23325 24035 23359
rect 25197 23325 25231 23359
rect 26761 23325 26795 23359
rect 28969 23325 29003 23359
rect 12869 23257 12903 23291
rect 13237 23257 13271 23291
rect 13421 23257 13455 23291
rect 14525 23257 14559 23291
rect 14617 23257 14651 23291
rect 14893 23257 14927 23291
rect 15445 23257 15479 23291
rect 16181 23257 16215 23291
rect 17193 23257 17227 23291
rect 18021 23257 18055 23291
rect 18389 23257 18423 23291
rect 19585 23257 19619 23291
rect 22989 23257 23023 23291
rect 23357 23257 23391 23291
rect 23541 23257 23575 23291
rect 24185 23257 24219 23291
rect 25381 23257 25415 23291
rect 27405 23257 27439 23291
rect 28325 23257 28359 23291
rect 12961 23189 12995 23223
rect 13973 23189 14007 23223
rect 15077 23189 15111 23223
rect 15997 23189 16031 23223
rect 16733 23189 16767 23223
rect 20376 23189 20410 23223
rect 20597 23189 20631 23223
rect 22897 23189 22931 23223
rect 20505 23053 20539 23087
rect 24277 23053 24311 23087
rect 26853 23053 26887 23087
rect 13973 22849 14007 22883
rect 20459 22849 20493 22883
rect 22897 22849 22931 22883
rect 25657 22849 25691 22883
rect 20597 22781 20631 22815
rect 12225 22713 12259 22747
rect 15629 22713 15663 22747
rect 18297 22713 18331 22747
rect 19125 22713 19159 22747
rect 19861 22713 19895 22747
rect 20689 22713 20723 22747
rect 22989 22713 23023 22747
rect 23909 22713 23943 22747
rect 24001 22713 24035 22747
rect 24829 22713 24863 22747
rect 26393 22713 26427 22747
rect 26945 22713 26979 22747
rect 12133 22645 12167 22679
rect 12409 22645 12443 22679
rect 13881 22645 13915 22679
rect 15261 22645 15295 22679
rect 16733 22645 16767 22679
rect 16917 22645 16951 22679
rect 17101 22645 17135 22679
rect 17469 22645 17503 22679
rect 17722 22645 17756 22679
rect 19309 22645 19343 22679
rect 20321 22645 20355 22679
rect 21057 22645 21091 22679
rect 22621 22645 22655 22679
rect 22768 22645 22802 22679
rect 23357 22645 23391 22679
rect 24737 22645 24771 22679
rect 25381 22645 25415 22679
rect 25565 22645 25599 22679
rect 28417 22645 28451 22679
rect 29061 22645 29095 22679
rect 15077 22577 15111 22611
rect 19477 22577 19511 22611
rect 26853 22577 26887 22611
rect 29337 22577 29371 22611
rect 19401 22509 19435 22543
rect 19677 22305 19711 22339
rect 24277 22305 24311 22339
rect 13973 22237 14007 22271
rect 15445 22237 15479 22271
rect 18573 22237 18607 22271
rect 20873 22237 20907 22271
rect 21609 22237 21643 22271
rect 28509 22237 28543 22271
rect 11857 22169 11891 22203
rect 14801 22169 14835 22203
rect 14985 22169 15019 22203
rect 15629 22169 15663 22203
rect 16825 22169 16859 22203
rect 18113 22169 18147 22203
rect 18389 22169 18423 22203
rect 19585 22169 19619 22203
rect 20321 22169 20355 22203
rect 20505 22169 20539 22203
rect 22805 22169 22839 22203
rect 22952 22169 22986 22203
rect 24001 22169 24035 22203
rect 24185 22169 24219 22203
rect 25197 22169 25231 22203
rect 25933 22169 25967 22203
rect 26853 22169 26887 22203
rect 29245 22169 29279 22203
rect 14525 22101 14559 22135
rect 16733 22101 16767 22135
rect 21977 22101 22011 22135
rect 23173 22101 23207 22135
rect 23541 22101 23575 22135
rect 28417 22101 28451 22135
rect 29337 22101 29371 22135
rect 21774 22033 21808 22067
rect 23081 22033 23115 22067
rect 27405 22033 27439 22067
rect 12041 21965 12075 21999
rect 15721 21965 15755 21999
rect 17009 21965 17043 21999
rect 21885 21965 21919 21999
rect 22069 21965 22103 21999
rect 25289 21965 25323 21999
rect 17009 21761 17043 21795
rect 18021 21761 18055 21795
rect 21701 21761 21735 21795
rect 23955 21761 23989 21795
rect 20505 21693 20539 21727
rect 21333 21693 21367 21727
rect 22897 21693 22931 21727
rect 24093 21693 24127 21727
rect 13237 21625 13271 21659
rect 14065 21625 14099 21659
rect 15169 21625 15203 21659
rect 19217 21625 19251 21659
rect 21425 21625 21459 21659
rect 22768 21625 22802 21659
rect 22989 21625 23023 21659
rect 24185 21625 24219 21659
rect 28509 21625 28543 21659
rect 12317 21557 12351 21591
rect 12593 21557 12627 21591
rect 12685 21557 12719 21591
rect 13145 21557 13179 21591
rect 14525 21557 14559 21591
rect 14801 21557 14835 21591
rect 14985 21557 15019 21591
rect 15537 21557 15571 21591
rect 16917 21557 16951 21591
rect 17929 21557 17963 21591
rect 19493 21557 19527 21591
rect 20413 21557 20447 21591
rect 21204 21557 21238 21591
rect 22621 21557 22655 21591
rect 25565 21557 25599 21591
rect 26485 21557 26519 21591
rect 27221 21557 27255 21591
rect 27957 21557 27991 21591
rect 28417 21557 28451 21591
rect 11857 21489 11891 21523
rect 16733 21489 16767 21523
rect 17745 21489 17779 21523
rect 19585 21489 19619 21523
rect 19953 21489 19987 21523
rect 21057 21489 21091 21523
rect 23357 21489 23391 21523
rect 23817 21489 23851 21523
rect 26301 21489 26335 21523
rect 27037 21489 27071 21523
rect 29061 21489 29095 21523
rect 29245 21489 29279 21523
rect 19401 21421 19435 21455
rect 24461 21421 24495 21455
rect 18573 21217 18607 21251
rect 11581 21149 11615 21183
rect 15169 21149 15203 21183
rect 15721 21149 15755 21183
rect 18665 21149 18699 21183
rect 19033 21149 19067 21183
rect 23725 21149 23759 21183
rect 27129 21149 27163 21183
rect 29429 21149 29463 21183
rect 11305 21081 11339 21115
rect 13329 21081 13363 21115
rect 14433 21081 14467 21115
rect 15353 21081 15387 21115
rect 16273 21081 16307 21115
rect 16457 21081 16491 21115
rect 16641 21081 16675 21115
rect 16917 21081 16951 21115
rect 17170 21081 17204 21115
rect 18481 21081 18515 21115
rect 20229 21081 20263 21115
rect 20597 21081 20631 21115
rect 20781 21081 20815 21115
rect 21885 21081 21919 21115
rect 22253 21081 22287 21115
rect 23633 21081 23667 21115
rect 24461 21081 24495 21115
rect 24553 21081 24587 21115
rect 25657 21081 25691 21115
rect 26669 21081 26703 21115
rect 27865 21081 27899 21115
rect 29153 21081 29187 21115
rect 17745 21013 17779 21047
rect 18297 21013 18331 21047
rect 20137 21013 20171 21047
rect 21701 21013 21735 21047
rect 22161 21013 22195 21047
rect 26209 21013 26243 21047
rect 27221 21013 27255 21047
rect 26117 20945 26151 20979
rect 14525 20877 14559 20911
rect 19677 20877 19711 20911
rect 21517 20877 21551 20911
rect 15445 20673 15479 20707
rect 19217 20673 19251 20707
rect 20597 20673 20631 20707
rect 22621 20673 22655 20707
rect 24001 20673 24035 20707
rect 20229 20605 20263 20639
rect 24737 20605 24771 20639
rect 12225 20537 12259 20571
rect 13145 20537 13179 20571
rect 18389 20537 18423 20571
rect 20100 20537 20134 20571
rect 20321 20537 20355 20571
rect 21701 20537 21735 20571
rect 26853 20537 26887 20571
rect 11857 20469 11891 20503
rect 13329 20469 13363 20503
rect 13697 20469 13731 20503
rect 13881 20469 13915 20503
rect 14525 20469 14559 20503
rect 15353 20469 15387 20503
rect 17929 20469 17963 20503
rect 18113 20469 18147 20503
rect 19125 20469 19159 20503
rect 19953 20469 19987 20503
rect 21149 20469 21183 20503
rect 21241 20469 21275 20503
rect 22345 20469 22379 20503
rect 22529 20469 22563 20503
rect 24185 20469 24219 20503
rect 24645 20469 24679 20503
rect 25289 20469 25323 20503
rect 26485 20469 26519 20503
rect 27957 20469 27991 20503
rect 11673 20401 11707 20435
rect 14341 20401 14375 20435
rect 14893 20401 14927 20435
rect 18941 20401 18975 20435
rect 28693 20401 28727 20435
rect 28877 20401 28911 20435
rect 12777 20333 12811 20367
rect 18389 20129 18423 20163
rect 18481 20129 18515 20163
rect 21425 20129 21459 20163
rect 27221 20129 27255 20163
rect 15813 20061 15847 20095
rect 17009 20061 17043 20095
rect 17561 20061 17595 20095
rect 18573 20061 18607 20095
rect 18941 20061 18975 20095
rect 19585 20061 19619 20095
rect 19769 20061 19803 20095
rect 19953 20061 19987 20095
rect 24093 20061 24127 20095
rect 26393 20061 26427 20095
rect 29061 20061 29095 20095
rect 11673 19993 11707 20027
rect 12685 19993 12719 20027
rect 12961 19993 12995 20027
rect 14249 19993 14283 20027
rect 14617 19993 14651 20027
rect 17193 19993 17227 20027
rect 19861 19993 19895 20027
rect 21793 19993 21827 20027
rect 22161 19993 22195 20027
rect 22253 19993 22287 20027
rect 23357 19993 23391 20027
rect 23541 19993 23575 20027
rect 24001 19993 24035 20027
rect 25473 19993 25507 20027
rect 26117 19993 26151 20027
rect 27129 19993 27163 20027
rect 27957 19993 27991 20027
rect 28601 19993 28635 20027
rect 12777 19925 12811 19959
rect 14341 19925 14375 19959
rect 16181 19925 16215 19959
rect 18205 19925 18239 19959
rect 20321 19925 20355 19959
rect 21701 19925 21735 19959
rect 29153 19925 29187 19959
rect 11765 19857 11799 19891
rect 15951 19857 15985 19891
rect 16089 19789 16123 19823
rect 16457 19789 16491 19823
rect 27773 19789 27807 19823
rect 27129 19585 27163 19619
rect 20229 19517 20263 19551
rect 24277 19517 24311 19551
rect 28693 19517 28727 19551
rect 13329 19449 13363 19483
rect 13789 19449 13823 19483
rect 14709 19449 14743 19483
rect 15445 19449 15479 19483
rect 17837 19449 17871 19483
rect 18941 19449 18975 19483
rect 19677 19449 19711 19483
rect 20873 19449 20907 19483
rect 13605 19381 13639 19415
rect 15353 19381 15387 19415
rect 15721 19381 15755 19415
rect 15905 19381 15939 19415
rect 16733 19381 16767 19415
rect 17745 19381 17779 19415
rect 19217 19381 19251 19415
rect 20137 19381 20171 19415
rect 20413 19381 20447 19415
rect 22989 19381 23023 19415
rect 24461 19381 24495 19415
rect 25473 19381 25507 19415
rect 25657 19381 25691 19415
rect 25841 19381 25875 19415
rect 26209 19381 26243 19415
rect 26485 19381 26519 19415
rect 28877 19381 28911 19415
rect 29245 19381 29279 19415
rect 29337 19381 29371 19415
rect 12777 19313 12811 19347
rect 19309 19313 19343 19347
rect 25013 19313 25047 19347
rect 27037 19313 27071 19347
rect 16825 19245 16859 19279
rect 19125 19245 19159 19279
rect 20321 19041 20355 19075
rect 21425 19041 21459 19075
rect 24369 19041 24403 19075
rect 26945 19041 26979 19075
rect 29245 19041 29279 19075
rect 13237 18973 13271 19007
rect 14249 18973 14283 19007
rect 16825 18973 16859 19007
rect 18573 18973 18607 19007
rect 19677 18973 19711 19007
rect 22713 18973 22747 19007
rect 22897 18973 22931 19007
rect 23817 18973 23851 19007
rect 26025 18973 26059 19007
rect 26117 18973 26151 19007
rect 12685 18905 12719 18939
rect 12961 18905 12995 18939
rect 14709 18905 14743 18939
rect 14893 18905 14927 18939
rect 15077 18905 15111 18939
rect 15353 18905 15387 18939
rect 21333 18905 21367 18939
rect 21977 18905 22011 18939
rect 23357 18905 23391 18939
rect 25565 18905 25599 18939
rect 27957 18905 27991 18939
rect 29429 18905 29463 18939
rect 12317 18837 12351 18871
rect 15629 18837 15663 18871
rect 16549 18837 16583 18871
rect 19824 18837 19858 18871
rect 20045 18837 20079 18871
rect 23909 18837 23943 18871
rect 24461 18837 24495 18871
rect 26577 18837 26611 18871
rect 26945 18769 26979 18803
rect 27773 18769 27807 18803
rect 19953 18701 19987 18735
rect 27957 18497 27991 18531
rect 15721 18429 15755 18463
rect 15905 18429 15939 18463
rect 17469 18429 17503 18463
rect 18297 18429 18331 18463
rect 22805 18429 22839 18463
rect 27313 18429 27347 18463
rect 28877 18429 28911 18463
rect 13329 18361 13363 18395
rect 15592 18361 15626 18395
rect 15813 18361 15847 18395
rect 18757 18361 18791 18395
rect 22345 18361 22379 18395
rect 25657 18361 25691 18395
rect 12869 18293 12903 18327
rect 13053 18293 13087 18327
rect 13421 18293 13455 18327
rect 14157 18293 14191 18327
rect 17285 18293 17319 18327
rect 18665 18293 18699 18327
rect 19033 18293 19067 18327
rect 19217 18293 19251 18327
rect 20045 18293 20079 18327
rect 20229 18293 20263 18327
rect 23541 18293 23575 18327
rect 24185 18293 24219 18327
rect 24369 18293 24403 18327
rect 25013 18293 25047 18327
rect 26485 18293 26519 18327
rect 27221 18293 27255 18327
rect 27957 18293 27991 18327
rect 28785 18293 28819 18327
rect 15445 18225 15479 18259
rect 20137 18225 20171 18259
rect 20689 18225 20723 18259
rect 22897 18225 22931 18259
rect 26301 18225 26335 18259
rect 26669 18225 26703 18259
rect 12685 18157 12719 18191
rect 14249 18157 14283 18191
rect 23357 18157 23391 18191
rect 24829 18157 24863 18191
rect 14249 17953 14283 17987
rect 15721 17953 15755 17987
rect 16917 17953 16951 17987
rect 13973 17885 14007 17919
rect 15629 17885 15663 17919
rect 15813 17885 15847 17919
rect 16641 17885 16675 17919
rect 24369 17885 24403 17919
rect 29245 17885 29279 17919
rect 12225 17817 12259 17851
rect 12409 17817 12443 17851
rect 12593 17817 12627 17851
rect 12869 17817 12903 17851
rect 13053 17817 13087 17851
rect 14157 17817 14191 17851
rect 16825 17817 16859 17851
rect 19953 17817 19987 17851
rect 20689 17817 20723 17851
rect 21149 17817 21183 17851
rect 23449 17817 23483 17851
rect 24093 17817 24127 17851
rect 26485 17817 26519 17851
rect 27773 17817 27807 17851
rect 28509 17817 28543 17851
rect 29429 17817 29463 17851
rect 11673 17749 11707 17783
rect 15445 17749 15479 17783
rect 16181 17749 16215 17783
rect 20321 17749 20355 17783
rect 25197 17749 25231 17783
rect 25749 17749 25783 17783
rect 25657 17681 25691 17715
rect 27773 17681 27807 17715
rect 21333 17613 21367 17647
rect 13513 17409 13547 17443
rect 16825 17341 16859 17375
rect 25565 17341 25599 17375
rect 12593 17273 12627 17307
rect 14617 17273 14651 17307
rect 14985 17273 15019 17307
rect 15445 17273 15479 17307
rect 22529 17273 22563 17307
rect 23449 17273 23483 17307
rect 26209 17273 26243 17307
rect 28509 17273 28543 17307
rect 29337 17273 29371 17307
rect 12501 17205 12535 17239
rect 12777 17205 12811 17239
rect 13421 17205 13455 17239
rect 15169 17205 15203 17239
rect 15537 17205 15571 17239
rect 16733 17205 16767 17239
rect 17009 17205 17043 17239
rect 17929 17205 17963 17239
rect 19309 17205 19343 17239
rect 23357 17205 23391 17239
rect 24093 17205 24127 17239
rect 25013 17205 25047 17239
rect 27037 17205 27071 17239
rect 27129 17205 27163 17239
rect 28417 17205 28451 17239
rect 29245 17205 29279 17239
rect 17469 17137 17503 17171
rect 19585 17137 19619 17171
rect 21333 17137 21367 17171
rect 22621 17137 22655 17171
rect 26301 17137 26335 17171
rect 18113 17069 18147 17103
rect 19953 16865 19987 16899
rect 26025 16865 26059 16899
rect 11581 16797 11615 16831
rect 13329 16797 13363 16831
rect 14249 16797 14283 16831
rect 24093 16797 24127 16831
rect 27589 16797 27623 16831
rect 11305 16729 11339 16763
rect 13973 16729 14007 16763
rect 16733 16729 16767 16763
rect 19677 16729 19711 16763
rect 19861 16729 19895 16763
rect 23541 16729 23575 16763
rect 25197 16729 25231 16763
rect 25933 16729 25967 16763
rect 27129 16729 27163 16763
rect 28601 16729 28635 16763
rect 15997 16661 16031 16695
rect 17009 16661 17043 16695
rect 18757 16661 18791 16695
rect 20873 16661 20907 16695
rect 21149 16661 21183 16695
rect 22897 16661 22931 16695
rect 24001 16661 24035 16695
rect 27681 16661 27715 16695
rect 29153 16661 29187 16695
rect 29061 16593 29095 16627
rect 25381 16525 25415 16559
rect 12133 16321 12167 16355
rect 14617 16321 14651 16355
rect 15353 16321 15387 16355
rect 15997 16321 16031 16355
rect 19585 16321 19619 16355
rect 22529 16321 22563 16355
rect 27129 16321 27163 16355
rect 18021 16253 18055 16287
rect 20965 16185 20999 16219
rect 25657 16185 25691 16219
rect 11949 16117 11983 16151
rect 14433 16117 14467 16151
rect 15261 16117 15295 16151
rect 15905 16117 15939 16151
rect 17101 16117 17135 16151
rect 17193 16117 17227 16151
rect 17653 16117 17687 16151
rect 17837 16117 17871 16151
rect 19125 16117 19159 16151
rect 19401 16117 19435 16151
rect 20597 16117 20631 16151
rect 21425 16117 21459 16151
rect 22345 16117 22379 16151
rect 23633 16117 23667 16151
rect 26117 16117 26151 16151
rect 27037 16117 27071 16151
rect 27957 16117 27991 16151
rect 28601 16117 28635 16151
rect 19309 16049 19343 16083
rect 20413 16049 20447 16083
rect 21517 16049 21551 16083
rect 23909 16049 23943 16083
rect 26301 15981 26335 16015
rect 28049 15981 28083 16015
rect 28785 15981 28819 16015
rect 24093 15777 24127 15811
rect 11765 15641 11799 15675
rect 13053 15641 13087 15675
rect 14709 15641 14743 15675
rect 14801 15641 14835 15675
rect 15261 15641 15295 15675
rect 15445 15641 15479 15675
rect 17193 15641 17227 15675
rect 17745 15641 17779 15675
rect 18389 15641 18423 15675
rect 18573 15641 18607 15675
rect 20045 15641 20079 15675
rect 20137 15641 20171 15675
rect 21885 15641 21919 15675
rect 22253 15641 22287 15675
rect 23081 15641 23115 15675
rect 23633 15641 23667 15675
rect 23817 15641 23851 15675
rect 25473 15641 25507 15675
rect 25565 15641 25599 15675
rect 26025 15641 26059 15675
rect 26209 15641 26243 15675
rect 11673 15573 11707 15607
rect 18941 15573 18975 15607
rect 22345 15573 22379 15607
rect 22989 15573 23023 15607
rect 27405 15573 27439 15607
rect 27681 15573 27715 15607
rect 29429 15573 29463 15607
rect 13145 15505 13179 15539
rect 19861 15505 19895 15539
rect 21701 15505 21735 15539
rect 11949 15437 11983 15471
rect 15721 15437 15755 15471
rect 17101 15437 17135 15471
rect 20321 15437 20355 15471
rect 26485 15437 26519 15471
rect 19125 15233 19159 15267
rect 19953 15233 19987 15267
rect 24185 15233 24219 15267
rect 29153 15233 29187 15267
rect 21609 15165 21643 15199
rect 11949 15097 11983 15131
rect 12961 15097 12995 15131
rect 13237 15097 13271 15131
rect 14985 15097 15019 15131
rect 23357 15097 23391 15131
rect 23909 15097 23943 15131
rect 25565 15097 25599 15131
rect 27313 15097 27347 15131
rect 11673 15029 11707 15063
rect 11857 15029 11891 15063
rect 15445 15029 15479 15063
rect 17285 15029 17319 15063
rect 17561 15029 17595 15063
rect 17745 15029 17779 15063
rect 18205 15029 18239 15063
rect 19033 15029 19067 15063
rect 20505 15029 20539 15063
rect 20597 15029 20631 15063
rect 20873 15029 20907 15063
rect 20965 15029 20999 15063
rect 21517 15029 21551 15063
rect 22437 15029 22471 15063
rect 23265 15029 23299 15063
rect 24001 15029 24035 15063
rect 25289 15029 25323 15063
rect 27957 15029 27991 15063
rect 28141 15029 28175 15063
rect 28601 15029 28635 15063
rect 28693 15029 28727 15063
rect 16733 14961 16767 14995
rect 18849 14961 18883 14995
rect 22529 14961 22563 14995
rect 15537 14893 15571 14927
rect 18297 14893 18331 14927
rect 14157 14689 14191 14723
rect 18205 14689 18239 14723
rect 18941 14689 18975 14723
rect 23541 14689 23575 14723
rect 26485 14689 26519 14723
rect 26577 14621 26611 14655
rect 26945 14621 26979 14655
rect 11949 14553 11983 14587
rect 12317 14553 12351 14587
rect 12969 14553 13003 14587
rect 13973 14553 14007 14587
rect 15169 14553 15203 14587
rect 15353 14553 15387 14587
rect 15905 14553 15939 14587
rect 16089 14553 16123 14587
rect 17193 14553 17227 14587
rect 17653 14553 17687 14587
rect 17745 14553 17779 14587
rect 18849 14553 18883 14587
rect 19769 14553 19803 14587
rect 22437 14553 22471 14587
rect 22805 14553 22839 14587
rect 22989 14553 23023 14587
rect 23449 14553 23483 14587
rect 25289 14553 25323 14587
rect 26393 14553 26427 14587
rect 29429 14553 29463 14587
rect 12041 14485 12075 14519
rect 12409 14485 12443 14519
rect 17009 14485 17043 14519
rect 19677 14485 19711 14519
rect 22529 14485 22563 14519
rect 25197 14485 25231 14519
rect 26209 14485 26243 14519
rect 27405 14485 27439 14519
rect 27681 14485 27715 14519
rect 16273 14417 16307 14451
rect 11397 14349 11431 14383
rect 13053 14349 13087 14383
rect 19953 14349 19987 14383
rect 22069 14349 22103 14383
rect 25473 14349 25507 14383
rect 13053 14145 13087 14179
rect 14893 14145 14927 14179
rect 22621 14145 22655 14179
rect 28233 14145 28267 14179
rect 28969 14145 29003 14179
rect 24645 14009 24679 14043
rect 11581 13941 11615 13975
rect 11949 13941 11983 13975
rect 12317 13941 12351 13975
rect 13605 13941 13639 13975
rect 13697 13941 13731 13975
rect 13973 13941 14007 13975
rect 14157 13941 14191 13975
rect 14801 13941 14835 13975
rect 15629 13941 15663 13975
rect 16825 13941 16859 13975
rect 17561 13941 17595 13975
rect 19585 13941 19619 13975
rect 20045 13941 20079 13975
rect 20229 13941 20263 13975
rect 20781 13941 20815 13975
rect 22345 13941 22379 13975
rect 22529 13941 22563 13975
rect 24185 13941 24219 13975
rect 24829 13941 24863 13975
rect 25105 13941 25139 13975
rect 25381 13941 25415 13975
rect 28141 13941 28175 13975
rect 29153 13941 29187 13975
rect 12501 13873 12535 13907
rect 14617 13873 14651 13907
rect 17837 13873 17871 13907
rect 20413 13873 20447 13907
rect 27957 13873 27991 13907
rect 15721 13805 15755 13839
rect 17009 13805 17043 13839
rect 20321 13805 20355 13839
rect 15813 13601 15847 13635
rect 19677 13601 19711 13635
rect 23541 13601 23575 13635
rect 29245 13601 29279 13635
rect 12317 13533 12351 13567
rect 12869 13533 12903 13567
rect 14709 13533 14743 13567
rect 17745 13533 17779 13567
rect 12501 13465 12535 13499
rect 13973 13465 14007 13499
rect 16181 13465 16215 13499
rect 16549 13465 16583 13499
rect 18389 13465 18423 13499
rect 18757 13465 18791 13499
rect 18941 13465 18975 13499
rect 19861 13465 19895 13499
rect 20137 13465 20171 13499
rect 21425 13465 21459 13499
rect 21885 13465 21919 13499
rect 21977 13465 22011 13499
rect 23449 13465 23483 13499
rect 24093 13465 24127 13499
rect 24277 13465 24311 13499
rect 24645 13465 24679 13499
rect 25381 13465 25415 13499
rect 25473 13465 25507 13499
rect 26577 13465 26611 13499
rect 29061 13465 29095 13499
rect 14341 13397 14375 13431
rect 16273 13397 16307 13431
rect 16457 13397 16491 13431
rect 18297 13397 18331 13431
rect 21241 13397 21275 13431
rect 25197 13397 25231 13431
rect 26853 13397 26887 13431
rect 28601 13397 28635 13431
rect 14249 13329 14283 13363
rect 14111 13261 14145 13295
rect 22437 13261 22471 13295
rect 25657 13261 25691 13295
rect 25197 13057 25231 13091
rect 28141 13057 28175 13091
rect 14525 12989 14559 13023
rect 21057 12989 21091 13023
rect 12961 12921 12995 12955
rect 13421 12921 13455 12955
rect 18941 12921 18975 12955
rect 19493 12921 19527 12955
rect 28785 12921 28819 12955
rect 12409 12853 12443 12887
rect 12501 12853 12535 12887
rect 13605 12853 13639 12887
rect 14065 12853 14099 12887
rect 14157 12853 14191 12887
rect 15261 12853 15295 12887
rect 19033 12853 19067 12887
rect 19401 12853 19435 12887
rect 21241 12853 21275 12887
rect 21609 12853 21643 12887
rect 21701 12853 21735 12887
rect 22345 12853 22379 12887
rect 23909 12853 23943 12887
rect 24921 12853 24955 12887
rect 25105 12853 25139 12887
rect 25933 12853 25967 12887
rect 26025 12853 26059 12887
rect 27957 12853 27991 12887
rect 28693 12853 28727 12887
rect 18389 12785 18423 12819
rect 15353 12717 15387 12751
rect 22437 12717 22471 12751
rect 23909 12717 23943 12751
rect 29153 12513 29187 12547
rect 13145 12445 13179 12479
rect 18665 12445 18699 12479
rect 20505 12445 20539 12479
rect 27497 12445 27531 12479
rect 12041 12377 12075 12411
rect 12593 12377 12627 12411
rect 12869 12377 12903 12411
rect 13973 12377 14007 12411
rect 14157 12377 14191 12411
rect 14709 12377 14743 12411
rect 14893 12377 14927 12411
rect 15905 12377 15939 12411
rect 16641 12377 16675 12411
rect 19585 12377 19619 12411
rect 21149 12377 21183 12411
rect 21517 12377 21551 12411
rect 21701 12377 21735 12411
rect 25473 12377 25507 12411
rect 27957 12377 27991 12411
rect 28141 12377 28175 12411
rect 28693 12377 28727 12411
rect 28877 12377 28911 12411
rect 16917 12309 16951 12343
rect 21241 12309 21275 12343
rect 22253 12309 22287 12343
rect 22529 12309 22563 12343
rect 24277 12309 24311 12343
rect 25749 12309 25783 12343
rect 15077 12241 15111 12275
rect 16089 12173 16123 12207
rect 19677 12173 19711 12207
rect 11765 11969 11799 12003
rect 12777 11969 12811 12003
rect 21517 11969 21551 12003
rect 26577 11969 26611 12003
rect 28049 11969 28083 12003
rect 13237 11833 13271 11867
rect 16181 11833 16215 11867
rect 17193 11833 17227 11867
rect 18665 11833 18699 11867
rect 18941 11833 18975 11867
rect 20689 11833 20723 11867
rect 21241 11833 21275 11867
rect 22437 11833 22471 11867
rect 23909 11833 23943 11867
rect 25933 11833 25967 11867
rect 11673 11765 11707 11799
rect 13145 11765 13179 11799
rect 13513 11765 13547 11799
rect 13697 11765 13731 11799
rect 14157 11765 14191 11799
rect 17745 11765 17779 11799
rect 18021 11765 18055 11799
rect 18205 11765 18239 11799
rect 21333 11765 21367 11799
rect 22345 11765 22379 11799
rect 26393 11765 26427 11799
rect 27957 11765 27991 11799
rect 14433 11697 14467 11731
rect 24185 11697 24219 11731
rect 16089 11425 16123 11459
rect 17561 11425 17595 11459
rect 18481 11425 18515 11459
rect 18757 11425 18791 11459
rect 19861 11425 19895 11459
rect 25565 11425 25599 11459
rect 15077 11289 15111 11323
rect 15629 11289 15663 11323
rect 15813 11289 15847 11323
rect 17377 11289 17411 11323
rect 14985 11221 15019 11255
rect 21885 11357 21919 11391
rect 18665 11289 18699 11323
rect 19677 11289 19711 11323
rect 20781 11289 20815 11323
rect 20873 11289 20907 11323
rect 21333 11289 21367 11323
rect 21517 11289 21551 11323
rect 23909 11289 23943 11323
rect 25381 11289 25415 11323
rect 18481 11153 18515 11187
rect 23081 11153 23115 11187
<< metal1 >>
rect 11000 30066 30136 30088
rect 11000 30014 19142 30066
rect 19194 30014 19206 30066
rect 19258 30014 19270 30066
rect 19322 30014 19334 30066
rect 19386 30014 29142 30066
rect 29194 30014 29206 30066
rect 29258 30014 29270 30066
rect 29322 30014 29334 30066
rect 29386 30014 30136 30066
rect 11000 29992 30136 30014
rect 20585 29887 20643 29893
rect 20585 29884 20597 29887
rect 19864 29856 20597 29884
rect 19864 29828 19892 29856
rect 20585 29853 20597 29856
rect 20631 29853 20643 29887
rect 20585 29847 20643 29853
rect 14970 29816 14976 29828
rect 14931 29788 14976 29816
rect 14970 29776 14976 29788
rect 15028 29776 15034 29828
rect 15062 29776 15068 29828
rect 15120 29816 15126 29828
rect 15433 29819 15491 29825
rect 15433 29816 15445 29819
rect 15120 29788 15445 29816
rect 15120 29776 15126 29788
rect 15433 29785 15445 29788
rect 15479 29785 15491 29819
rect 15433 29779 15491 29785
rect 18929 29819 18987 29825
rect 18929 29785 18941 29819
rect 18975 29816 18987 29819
rect 19754 29816 19760 29828
rect 18975 29788 19760 29816
rect 18975 29785 18987 29788
rect 18929 29779 18987 29785
rect 19754 29776 19760 29788
rect 19812 29776 19818 29828
rect 19846 29776 19852 29828
rect 19904 29816 19910 29828
rect 20401 29819 20459 29825
rect 19904 29788 19997 29816
rect 19904 29776 19910 29788
rect 20401 29785 20413 29819
rect 20447 29785 20459 29819
rect 20401 29779 20459 29785
rect 22609 29819 22667 29825
rect 22609 29785 22621 29819
rect 22655 29816 22667 29819
rect 23342 29816 23348 29828
rect 22655 29788 23348 29816
rect 22655 29785 22667 29788
rect 22609 29779 22667 29785
rect 20416 29680 20444 29779
rect 23342 29776 23348 29788
rect 23400 29776 23406 29828
rect 26378 29816 26384 29828
rect 26339 29788 26384 29816
rect 26378 29776 26384 29788
rect 26436 29776 26442 29828
rect 28678 29776 28684 29828
rect 28736 29816 28742 29828
rect 28957 29819 29015 29825
rect 28957 29816 28969 29819
rect 28736 29788 28969 29816
rect 28736 29776 28742 29788
rect 28957 29785 28969 29788
rect 29003 29785 29015 29819
rect 28957 29779 29015 29785
rect 21134 29748 21140 29760
rect 21095 29720 21140 29748
rect 21134 29708 21140 29720
rect 21192 29708 21198 29760
rect 21689 29751 21747 29757
rect 21689 29717 21701 29751
rect 21735 29748 21747 29751
rect 22701 29751 22759 29757
rect 22701 29748 22713 29751
rect 21735 29720 22713 29748
rect 21735 29717 21747 29720
rect 21689 29711 21747 29717
rect 22701 29717 22713 29720
rect 22747 29717 22759 29751
rect 22701 29711 22759 29717
rect 21597 29683 21655 29689
rect 21597 29680 21609 29683
rect 20416 29652 21609 29680
rect 21597 29649 21609 29652
rect 21643 29680 21655 29683
rect 21962 29680 21968 29692
rect 21643 29652 21968 29680
rect 21643 29649 21655 29652
rect 21597 29643 21655 29649
rect 21962 29640 21968 29652
rect 22020 29640 22026 29692
rect 14694 29572 14700 29624
rect 14752 29612 14758 29624
rect 14789 29615 14847 29621
rect 14789 29612 14801 29615
rect 14752 29584 14801 29612
rect 14752 29572 14758 29584
rect 14789 29581 14801 29584
rect 14835 29581 14847 29615
rect 14789 29575 14847 29581
rect 15525 29615 15583 29621
rect 15525 29581 15537 29615
rect 15571 29612 15583 29615
rect 15982 29612 15988 29624
rect 15571 29584 15988 29612
rect 15571 29581 15583 29584
rect 15525 29575 15583 29581
rect 15982 29572 15988 29584
rect 16040 29572 16046 29624
rect 19018 29612 19024 29624
rect 18979 29584 19024 29612
rect 19018 29572 19024 29584
rect 19076 29572 19082 29624
rect 19662 29612 19668 29624
rect 19623 29584 19668 29612
rect 19662 29572 19668 29584
rect 19720 29572 19726 29624
rect 26197 29615 26255 29621
rect 26197 29581 26209 29615
rect 26243 29612 26255 29615
rect 27482 29612 27488 29624
rect 26243 29584 27488 29612
rect 26243 29581 26255 29584
rect 26197 29575 26255 29581
rect 27482 29572 27488 29584
rect 27540 29572 27546 29624
rect 28862 29572 28868 29624
rect 28920 29612 28926 29624
rect 29049 29615 29107 29621
rect 29049 29612 29061 29615
rect 28920 29584 29061 29612
rect 28920 29572 28926 29584
rect 29049 29581 29061 29584
rect 29095 29581 29107 29615
rect 29049 29575 29107 29581
rect 11000 29522 30136 29544
rect 11000 29470 14142 29522
rect 14194 29470 14206 29522
rect 14258 29470 14270 29522
rect 14322 29470 14334 29522
rect 14386 29470 24142 29522
rect 24194 29470 24206 29522
rect 24258 29470 24270 29522
rect 24322 29470 24334 29522
rect 24386 29470 30136 29522
rect 11000 29448 30136 29470
rect 21318 29408 21324 29420
rect 13424 29380 21324 29408
rect 13424 29204 13452 29380
rect 21318 29368 21324 29380
rect 21376 29368 21382 29420
rect 18374 29300 18380 29352
rect 18432 29340 18438 29352
rect 18837 29343 18895 29349
rect 18837 29340 18849 29343
rect 18432 29312 18849 29340
rect 18432 29300 18438 29312
rect 18837 29309 18849 29312
rect 18883 29309 18895 29343
rect 18837 29303 18895 29309
rect 19754 29300 19760 29352
rect 19812 29340 19818 29352
rect 20033 29343 20091 29349
rect 20033 29340 20045 29343
rect 19812 29312 20045 29340
rect 19812 29300 19818 29312
rect 20033 29309 20045 29312
rect 20079 29309 20091 29343
rect 20033 29303 20091 29309
rect 13498 29232 13504 29284
rect 13556 29272 13562 29284
rect 14513 29275 14571 29281
rect 14513 29272 14525 29275
rect 13556 29244 14525 29272
rect 13556 29232 13562 29244
rect 14513 29241 14525 29244
rect 14559 29241 14571 29275
rect 16077 29275 16135 29281
rect 14513 29235 14571 29241
rect 14988 29244 16028 29272
rect 13593 29207 13651 29213
rect 13593 29204 13605 29207
rect 13424 29176 13605 29204
rect 13593 29173 13605 29176
rect 13639 29173 13651 29207
rect 13593 29167 13651 29173
rect 14421 29207 14479 29213
rect 14421 29173 14433 29207
rect 14467 29204 14479 29207
rect 14988 29204 15016 29244
rect 15154 29204 15160 29216
rect 14467 29176 15016 29204
rect 15115 29176 15160 29204
rect 14467 29173 14479 29176
rect 14421 29167 14479 29173
rect 15154 29164 15160 29176
rect 15212 29164 15218 29216
rect 16000 29213 16028 29244
rect 16077 29241 16089 29275
rect 16123 29272 16135 29275
rect 16350 29272 16356 29284
rect 16123 29244 16356 29272
rect 16123 29241 16135 29244
rect 16077 29235 16135 29241
rect 16350 29232 16356 29244
rect 16408 29232 16414 29284
rect 19662 29232 19668 29284
rect 19720 29272 19726 29284
rect 20125 29275 20183 29281
rect 20125 29272 20137 29275
rect 19720 29244 20137 29272
rect 19720 29232 19726 29244
rect 20125 29241 20137 29244
rect 20171 29241 20183 29275
rect 20125 29235 20183 29241
rect 20769 29275 20827 29281
rect 20769 29241 20781 29275
rect 20815 29272 20827 29275
rect 21134 29272 21140 29284
rect 20815 29244 21140 29272
rect 20815 29241 20827 29244
rect 20769 29235 20827 29241
rect 21134 29232 21140 29244
rect 21192 29232 21198 29284
rect 21597 29275 21655 29281
rect 21597 29241 21609 29275
rect 21643 29272 21655 29275
rect 22054 29272 22060 29284
rect 21643 29244 22060 29272
rect 21643 29241 21655 29244
rect 21597 29235 21655 29241
rect 22054 29232 22060 29244
rect 22112 29232 22118 29284
rect 23526 29272 23532 29284
rect 22256 29244 23532 29272
rect 15985 29207 16043 29213
rect 15985 29173 15997 29207
rect 16031 29173 16043 29207
rect 15985 29167 16043 29173
rect 17549 29207 17607 29213
rect 17549 29173 17561 29207
rect 17595 29204 17607 29207
rect 17638 29204 17644 29216
rect 17595 29176 17644 29204
rect 17595 29173 17607 29176
rect 17549 29167 17607 29173
rect 13685 29139 13743 29145
rect 13685 29105 13697 29139
rect 13731 29136 13743 29139
rect 14050 29136 14056 29148
rect 13731 29108 14056 29136
rect 13731 29105 13743 29108
rect 13685 29099 13743 29105
rect 14050 29096 14056 29108
rect 14108 29096 14114 29148
rect 15249 29139 15307 29145
rect 15249 29105 15261 29139
rect 15295 29136 15307 29139
rect 15430 29136 15436 29148
rect 15295 29108 15436 29136
rect 15295 29105 15307 29108
rect 15249 29099 15307 29105
rect 15430 29096 15436 29108
rect 15488 29096 15494 29148
rect 16000 29136 16028 29167
rect 17638 29164 17644 29176
rect 17696 29164 17702 29216
rect 19021 29207 19079 29213
rect 19021 29173 19033 29207
rect 19067 29173 19079 29207
rect 19021 29167 19079 29173
rect 19573 29207 19631 29213
rect 19573 29173 19585 29207
rect 19619 29204 19631 29207
rect 20030 29204 20036 29216
rect 19619 29176 20036 29204
rect 19619 29173 19631 29176
rect 19573 29167 19631 29173
rect 18558 29136 18564 29148
rect 16000 29108 18564 29136
rect 18558 29096 18564 29108
rect 18616 29096 18622 29148
rect 19036 29136 19064 29167
rect 20030 29164 20036 29176
rect 20088 29164 20094 29216
rect 20674 29204 20680 29216
rect 20635 29176 20680 29204
rect 20674 29164 20680 29176
rect 20732 29164 20738 29216
rect 21505 29207 21563 29213
rect 21505 29204 21517 29207
rect 20784 29176 21517 29204
rect 19846 29136 19852 29148
rect 19036 29108 19852 29136
rect 19846 29096 19852 29108
rect 19904 29096 19910 29148
rect 18576 29068 18604 29096
rect 20784 29068 20812 29176
rect 21505 29173 21517 29176
rect 21551 29204 21563 29207
rect 22256 29204 22284 29244
rect 23526 29232 23532 29244
rect 23584 29232 23590 29284
rect 22698 29204 22704 29216
rect 21551 29176 22284 29204
rect 22659 29176 22704 29204
rect 21551 29173 21563 29176
rect 21505 29167 21563 29173
rect 22698 29164 22704 29176
rect 22756 29164 22762 29216
rect 23342 29204 23348 29216
rect 23303 29176 23348 29204
rect 23342 29164 23348 29176
rect 23400 29164 23406 29216
rect 24265 29207 24323 29213
rect 24265 29204 24277 29207
rect 23636 29176 24277 29204
rect 22146 29096 22152 29148
rect 22204 29136 22210 29148
rect 23636 29145 23664 29176
rect 24265 29173 24277 29176
rect 24311 29204 24323 29207
rect 24446 29204 24452 29216
rect 24311 29176 24452 29204
rect 24311 29173 24323 29176
rect 24265 29167 24323 29173
rect 24446 29164 24452 29176
rect 24504 29164 24510 29216
rect 25458 29204 25464 29216
rect 25419 29176 25464 29204
rect 25458 29164 25464 29176
rect 25516 29164 25522 29216
rect 26197 29207 26255 29213
rect 26197 29173 26209 29207
rect 26243 29204 26255 29207
rect 27390 29204 27396 29216
rect 26243 29176 27396 29204
rect 26243 29173 26255 29176
rect 26197 29167 26255 29173
rect 23621 29139 23679 29145
rect 23621 29136 23633 29139
rect 22204 29108 23633 29136
rect 22204 29096 22210 29108
rect 23621 29105 23633 29108
rect 23667 29105 23679 29139
rect 23621 29099 23679 29105
rect 24817 29139 24875 29145
rect 24817 29105 24829 29139
rect 24863 29136 24875 29139
rect 26212 29136 26240 29167
rect 27390 29164 27396 29176
rect 27448 29164 27454 29216
rect 29233 29207 29291 29213
rect 29233 29173 29245 29207
rect 29279 29204 29291 29207
rect 29506 29204 29512 29216
rect 29279 29176 29512 29204
rect 29279 29173 29291 29176
rect 29233 29167 29291 29173
rect 29506 29164 29512 29176
rect 29564 29164 29570 29216
rect 26378 29136 26384 29148
rect 24863 29108 26240 29136
rect 26339 29108 26384 29136
rect 24863 29105 24875 29108
rect 24817 29099 24875 29105
rect 26378 29096 26384 29108
rect 26436 29096 26442 29148
rect 18576 29040 20812 29068
rect 23710 29028 23716 29080
rect 23768 29068 23774 29080
rect 24081 29071 24139 29077
rect 24081 29068 24093 29071
rect 23768 29040 24093 29068
rect 23768 29028 23774 29040
rect 24081 29037 24093 29040
rect 24127 29037 24139 29071
rect 24081 29031 24139 29037
rect 24909 29071 24967 29077
rect 24909 29037 24921 29071
rect 24955 29068 24967 29071
rect 26286 29068 26292 29080
rect 24955 29040 26292 29068
rect 24955 29037 24967 29040
rect 24909 29031 24967 29037
rect 26286 29028 26292 29040
rect 26344 29028 26350 29080
rect 27114 29068 27120 29080
rect 27075 29040 27120 29068
rect 27114 29028 27120 29040
rect 27172 29028 27178 29080
rect 27206 29028 27212 29080
rect 27264 29068 27270 29080
rect 27264 29040 27309 29068
rect 27264 29028 27270 29040
rect 28770 29028 28776 29080
rect 28828 29068 28834 29080
rect 29049 29071 29107 29077
rect 29049 29068 29061 29071
rect 28828 29040 29061 29068
rect 28828 29028 28834 29040
rect 29049 29037 29061 29040
rect 29095 29037 29107 29071
rect 29049 29031 29107 29037
rect 11000 28978 30136 29000
rect 11000 28926 19142 28978
rect 19194 28926 19206 28978
rect 19258 28926 19270 28978
rect 19322 28926 19334 28978
rect 19386 28926 29142 28978
rect 29194 28926 29206 28978
rect 29258 28926 29270 28978
rect 29322 28926 29334 28978
rect 29386 28926 30136 28978
rect 11000 28904 30136 28926
rect 14510 28824 14516 28876
rect 14568 28864 14574 28876
rect 20674 28864 20680 28876
rect 14568 28836 18144 28864
rect 14568 28824 14574 28836
rect 14789 28799 14847 28805
rect 14789 28765 14801 28799
rect 14835 28796 14847 28799
rect 15062 28796 15068 28808
rect 14835 28768 15068 28796
rect 14835 28765 14847 28768
rect 14789 28759 14847 28765
rect 15062 28756 15068 28768
rect 15120 28756 15126 28808
rect 10646 28688 10652 28740
rect 10704 28728 10710 28740
rect 11661 28731 11719 28737
rect 11661 28728 11673 28731
rect 10704 28700 11673 28728
rect 10704 28688 10710 28700
rect 11661 28697 11673 28700
rect 11707 28697 11719 28731
rect 14050 28728 14056 28740
rect 14011 28700 14056 28728
rect 11661 28691 11719 28697
rect 14050 28688 14056 28700
rect 14108 28688 14114 28740
rect 14970 28728 14976 28740
rect 14883 28700 14976 28728
rect 14970 28688 14976 28700
rect 15028 28688 15034 28740
rect 15430 28728 15436 28740
rect 15391 28700 15436 28728
rect 15430 28688 15436 28700
rect 15488 28688 15494 28740
rect 16718 28728 16724 28740
rect 16679 28700 16724 28728
rect 16718 28688 16724 28700
rect 16776 28688 16782 28740
rect 14988 28660 15016 28688
rect 16736 28660 16764 28688
rect 14988 28632 16764 28660
rect 17638 28620 17644 28672
rect 17696 28660 17702 28672
rect 17917 28663 17975 28669
rect 17917 28660 17929 28663
rect 17696 28632 17929 28660
rect 17696 28620 17702 28632
rect 17917 28629 17929 28632
rect 17963 28629 17975 28663
rect 18116 28660 18144 28836
rect 19680 28836 20680 28864
rect 18469 28799 18527 28805
rect 18469 28765 18481 28799
rect 18515 28796 18527 28799
rect 19018 28796 19024 28808
rect 18515 28768 19024 28796
rect 18515 28765 18527 28768
rect 18469 28759 18527 28765
rect 19018 28756 19024 28768
rect 19076 28756 19082 28808
rect 19680 28805 19708 28836
rect 20674 28824 20680 28836
rect 20732 28824 20738 28876
rect 24446 28864 24452 28876
rect 24407 28836 24452 28864
rect 24446 28824 24452 28836
rect 24504 28824 24510 28876
rect 27758 28824 27764 28876
rect 27816 28864 27822 28876
rect 28129 28867 28187 28873
rect 28129 28864 28141 28867
rect 27816 28836 28141 28864
rect 27816 28824 27822 28836
rect 28129 28833 28141 28836
rect 28175 28833 28187 28867
rect 28129 28827 28187 28833
rect 19665 28799 19723 28805
rect 19665 28765 19677 28799
rect 19711 28765 19723 28799
rect 19665 28759 19723 28765
rect 22698 28756 22704 28808
rect 22756 28796 22762 28808
rect 22885 28799 22943 28805
rect 22885 28796 22897 28799
rect 22756 28768 22897 28796
rect 22756 28756 22762 28768
rect 22885 28765 22897 28768
rect 22931 28765 22943 28799
rect 22885 28759 22943 28765
rect 25458 28756 25464 28808
rect 25516 28796 25522 28808
rect 25553 28799 25611 28805
rect 25553 28796 25565 28799
rect 25516 28768 25565 28796
rect 25516 28756 25522 28768
rect 25553 28765 25565 28768
rect 25599 28796 25611 28799
rect 27482 28796 27488 28808
rect 25599 28768 26976 28796
rect 27443 28768 27488 28796
rect 25599 28765 25611 28768
rect 25553 28759 25611 28765
rect 18190 28688 18196 28740
rect 18248 28728 18254 28740
rect 19573 28731 19631 28737
rect 19573 28728 19585 28731
rect 18248 28700 19585 28728
rect 18248 28688 18254 28700
rect 19573 28697 19585 28700
rect 19619 28697 19631 28731
rect 19573 28691 19631 28697
rect 19849 28731 19907 28737
rect 19849 28697 19861 28731
rect 19895 28728 19907 28731
rect 20306 28728 20312 28740
rect 19895 28700 20312 28728
rect 19895 28697 19907 28700
rect 19849 28691 19907 28697
rect 20306 28688 20312 28700
rect 20364 28688 20370 28740
rect 20677 28731 20735 28737
rect 20677 28697 20689 28731
rect 20723 28728 20735 28731
rect 21134 28728 21140 28740
rect 20723 28700 21140 28728
rect 20723 28697 20735 28700
rect 20677 28691 20735 28697
rect 21134 28688 21140 28700
rect 21192 28688 21198 28740
rect 22146 28728 22152 28740
rect 22107 28700 22152 28728
rect 22146 28688 22152 28700
rect 22204 28688 22210 28740
rect 23618 28728 23624 28740
rect 23579 28700 23624 28728
rect 23618 28688 23624 28700
rect 23676 28688 23682 28740
rect 24357 28731 24415 28737
rect 24357 28697 24369 28731
rect 24403 28728 24415 28731
rect 24722 28728 24728 28740
rect 24403 28700 24728 28728
rect 24403 28697 24415 28700
rect 24357 28691 24415 28697
rect 24722 28688 24728 28700
rect 24780 28688 24786 28740
rect 25274 28688 25280 28740
rect 25332 28728 25338 28740
rect 26948 28737 26976 28768
rect 27482 28756 27488 28768
rect 27540 28756 27546 28808
rect 26289 28731 26347 28737
rect 26289 28728 26301 28731
rect 25332 28700 26301 28728
rect 25332 28688 25338 28700
rect 26289 28697 26301 28700
rect 26335 28697 26347 28731
rect 26289 28691 26347 28697
rect 26933 28731 26991 28737
rect 26933 28697 26945 28731
rect 26979 28697 26991 28731
rect 27390 28728 27396 28740
rect 27351 28700 27396 28728
rect 26933 28691 26991 28697
rect 27390 28688 27396 28700
rect 27448 28688 27454 28740
rect 27850 28688 27856 28740
rect 27908 28728 27914 28740
rect 27945 28731 28003 28737
rect 27945 28728 27957 28731
rect 27908 28700 27957 28728
rect 27908 28688 27914 28700
rect 27945 28697 27957 28700
rect 27991 28697 28003 28731
rect 27945 28691 28003 28697
rect 28954 28688 28960 28740
rect 29012 28728 29018 28740
rect 29141 28731 29199 28737
rect 29141 28728 29153 28731
rect 29012 28700 29153 28728
rect 29012 28688 29018 28700
rect 29141 28697 29153 28700
rect 29187 28697 29199 28731
rect 29141 28691 29199 28697
rect 22606 28660 22612 28672
rect 18116 28632 22612 28660
rect 17917 28623 17975 28629
rect 22606 28620 22612 28632
rect 22664 28620 22670 28672
rect 22790 28660 22796 28672
rect 22751 28632 22796 28660
rect 22790 28620 22796 28632
rect 22848 28620 22854 28672
rect 23713 28663 23771 28669
rect 23713 28629 23725 28663
rect 23759 28629 23771 28663
rect 25458 28660 25464 28672
rect 25419 28632 25464 28660
rect 23713 28623 23771 28629
rect 16626 28552 16632 28604
rect 16684 28592 16690 28604
rect 16721 28595 16779 28601
rect 16721 28592 16733 28595
rect 16684 28564 16733 28592
rect 16684 28552 16690 28564
rect 16721 28561 16733 28564
rect 16767 28561 16779 28595
rect 18374 28592 18380 28604
rect 18335 28564 18380 28592
rect 16721 28555 16779 28561
rect 18374 28552 18380 28564
rect 18432 28552 18438 28604
rect 19573 28595 19631 28601
rect 19573 28561 19585 28595
rect 19619 28592 19631 28595
rect 21962 28592 21968 28604
rect 19619 28564 20904 28592
rect 21923 28564 21968 28592
rect 19619 28561 19631 28564
rect 19573 28555 19631 28561
rect 11753 28527 11811 28533
rect 11753 28493 11765 28527
rect 11799 28524 11811 28527
rect 18282 28524 18288 28536
rect 11799 28496 18288 28524
rect 11799 28493 11811 28496
rect 11753 28487 11811 28493
rect 18282 28484 18288 28496
rect 18340 28484 18346 28536
rect 19662 28484 19668 28536
rect 19720 28524 19726 28536
rect 19941 28527 19999 28533
rect 19941 28524 19953 28527
rect 19720 28496 19953 28524
rect 19720 28484 19726 28496
rect 19941 28493 19953 28496
rect 19987 28493 19999 28527
rect 19941 28487 19999 28493
rect 20214 28484 20220 28536
rect 20272 28524 20278 28536
rect 20766 28524 20772 28536
rect 20272 28496 20772 28524
rect 20272 28484 20278 28496
rect 20766 28484 20772 28496
rect 20824 28484 20830 28536
rect 20876 28524 20904 28564
rect 21962 28552 21968 28564
rect 22020 28552 22026 28604
rect 23728 28524 23756 28623
rect 25458 28620 25464 28632
rect 25516 28620 25522 28672
rect 26381 28663 26439 28669
rect 26381 28629 26393 28663
rect 26427 28660 26439 28663
rect 29598 28660 29604 28672
rect 26427 28632 29604 28660
rect 26427 28629 26439 28632
rect 26381 28623 26439 28629
rect 29598 28620 29604 28632
rect 29656 28620 29662 28672
rect 20876 28496 23756 28524
rect 28586 28484 28592 28536
rect 28644 28524 28650 28536
rect 29233 28527 29291 28533
rect 29233 28524 29245 28527
rect 28644 28496 29245 28524
rect 28644 28484 28650 28496
rect 29233 28493 29245 28496
rect 29279 28493 29291 28527
rect 29233 28487 29291 28493
rect 11000 28434 30136 28456
rect 11000 28382 14142 28434
rect 14194 28382 14206 28434
rect 14258 28382 14270 28434
rect 14322 28382 14334 28434
rect 14386 28382 24142 28434
rect 24194 28382 24206 28434
rect 24258 28382 24270 28434
rect 24322 28382 24334 28434
rect 24386 28382 30136 28434
rect 11000 28360 30136 28382
rect 15154 28280 15160 28332
rect 15212 28320 15218 28332
rect 15212 28292 18788 28320
rect 15212 28280 15218 28292
rect 12486 28212 12492 28264
rect 12544 28252 12550 28264
rect 18760 28252 18788 28292
rect 20674 28280 20680 28332
rect 20732 28320 20738 28332
rect 20861 28323 20919 28329
rect 20861 28320 20873 28323
rect 20732 28292 20873 28320
rect 20732 28280 20738 28292
rect 20861 28289 20873 28292
rect 20907 28289 20919 28323
rect 20861 28283 20919 28289
rect 22514 28252 22520 28264
rect 12544 28224 18696 28252
rect 18760 28224 22520 28252
rect 12544 28212 12550 28224
rect 13958 28144 13964 28196
rect 14016 28184 14022 28196
rect 14145 28187 14203 28193
rect 14145 28184 14157 28187
rect 14016 28156 14157 28184
rect 14016 28144 14022 28156
rect 14145 28153 14157 28156
rect 14191 28153 14203 28187
rect 14145 28147 14203 28153
rect 14605 28187 14663 28193
rect 14605 28153 14617 28187
rect 14651 28184 14663 28187
rect 15062 28184 15068 28196
rect 14651 28156 15068 28184
rect 14651 28153 14663 28156
rect 14605 28147 14663 28153
rect 15062 28144 15068 28156
rect 15120 28144 15126 28196
rect 15430 28184 15436 28196
rect 15391 28156 15436 28184
rect 15430 28144 15436 28156
rect 15488 28144 15494 28196
rect 15893 28187 15951 28193
rect 15893 28153 15905 28187
rect 15939 28184 15951 28187
rect 16626 28184 16632 28196
rect 15939 28156 16632 28184
rect 15939 28153 15951 28156
rect 15893 28147 15951 28153
rect 16626 28144 16632 28156
rect 16684 28184 16690 28196
rect 18668 28193 18696 28224
rect 22514 28212 22520 28224
rect 22572 28212 22578 28264
rect 23253 28255 23311 28261
rect 23253 28221 23265 28255
rect 23299 28252 23311 28255
rect 23342 28252 23348 28264
rect 23299 28224 23348 28252
rect 23299 28221 23311 28224
rect 23253 28215 23311 28221
rect 23342 28212 23348 28224
rect 23400 28212 23406 28264
rect 24722 28212 24728 28264
rect 24780 28252 24786 28264
rect 25737 28255 25795 28261
rect 25737 28252 25749 28255
rect 24780 28224 25749 28252
rect 24780 28212 24786 28224
rect 25737 28221 25749 28224
rect 25783 28252 25795 28255
rect 26933 28255 26991 28261
rect 26933 28252 26945 28255
rect 25783 28224 26945 28252
rect 25783 28221 25795 28224
rect 25737 28215 25795 28221
rect 26933 28221 26945 28224
rect 26979 28221 26991 28255
rect 26933 28215 26991 28221
rect 18653 28187 18711 28193
rect 16684 28156 18144 28184
rect 16684 28144 16690 28156
rect 14694 28116 14700 28128
rect 14655 28088 14700 28116
rect 14694 28076 14700 28088
rect 14752 28076 14758 28128
rect 15982 28116 15988 28128
rect 15943 28088 15988 28116
rect 15982 28076 15988 28088
rect 16040 28076 16046 28128
rect 16718 28076 16724 28128
rect 16776 28116 16782 28128
rect 17181 28119 17239 28125
rect 17181 28116 17193 28119
rect 16776 28088 17193 28116
rect 16776 28076 16782 28088
rect 17181 28085 17193 28088
rect 17227 28085 17239 28119
rect 17181 28079 17239 28085
rect 17733 28119 17791 28125
rect 17733 28085 17745 28119
rect 17779 28116 17791 28119
rect 18006 28116 18012 28128
rect 17779 28088 18012 28116
rect 17779 28085 17791 28088
rect 17733 28079 17791 28085
rect 18006 28076 18012 28088
rect 18064 28076 18070 28128
rect 16997 28051 17055 28057
rect 16997 28017 17009 28051
rect 17043 28048 17055 28051
rect 17822 28048 17828 28060
rect 17043 28020 17684 28048
rect 17783 28020 17828 28048
rect 17043 28017 17055 28020
rect 16997 28011 17055 28017
rect 17656 27980 17684 28020
rect 17822 28008 17828 28020
rect 17880 28008 17886 28060
rect 18116 28048 18144 28156
rect 18653 28153 18665 28187
rect 18699 28153 18711 28187
rect 18653 28147 18711 28153
rect 19754 28144 19760 28196
rect 19812 28184 19818 28196
rect 19812 28156 19892 28184
rect 19812 28144 19818 28156
rect 18558 28116 18564 28128
rect 18519 28088 18564 28116
rect 18558 28076 18564 28088
rect 18616 28076 18622 28128
rect 19864 28125 19892 28156
rect 22698 28144 22704 28196
rect 22756 28184 22762 28196
rect 22793 28187 22851 28193
rect 22793 28184 22805 28187
rect 22756 28156 22805 28184
rect 22756 28144 22762 28156
rect 22793 28153 22805 28156
rect 22839 28153 22851 28187
rect 22793 28147 22851 28153
rect 19205 28119 19263 28125
rect 19205 28085 19217 28119
rect 19251 28085 19263 28119
rect 19205 28079 19263 28085
rect 19849 28119 19907 28125
rect 19849 28085 19861 28119
rect 19895 28085 19907 28119
rect 19849 28079 19907 28085
rect 19220 28048 19248 28079
rect 19938 28076 19944 28128
rect 19996 28116 20002 28128
rect 20125 28119 20183 28125
rect 20125 28116 20137 28119
rect 19996 28088 20137 28116
rect 19996 28076 20002 28088
rect 20125 28085 20137 28088
rect 20171 28085 20183 28119
rect 20125 28079 20183 28085
rect 20769 28119 20827 28125
rect 20769 28085 20781 28119
rect 20815 28116 20827 28119
rect 21778 28116 21784 28128
rect 20815 28088 21784 28116
rect 20815 28085 20827 28088
rect 20769 28079 20827 28085
rect 21778 28076 21784 28088
rect 21836 28076 21842 28128
rect 23345 28119 23403 28125
rect 23345 28085 23357 28119
rect 23391 28116 23403 28119
rect 23710 28116 23716 28128
rect 23391 28088 23716 28116
rect 23391 28085 23403 28088
rect 23345 28079 23403 28085
rect 23710 28076 23716 28088
rect 23768 28076 23774 28128
rect 24449 28119 24507 28125
rect 24449 28085 24461 28119
rect 24495 28085 24507 28119
rect 25366 28116 25372 28128
rect 25327 28088 25372 28116
rect 24449 28079 24507 28085
rect 20030 28048 20036 28060
rect 18116 28020 18512 28048
rect 19220 28020 20036 28048
rect 18374 27980 18380 27992
rect 17656 27952 18380 27980
rect 18374 27940 18380 27952
rect 18432 27940 18438 27992
rect 18484 27980 18512 28020
rect 20030 28008 20036 28020
rect 20088 28008 20094 28060
rect 20582 28048 20588 28060
rect 20543 28020 20588 28048
rect 20582 28008 20588 28020
rect 20640 28008 20646 28060
rect 23802 28008 23808 28060
rect 23860 28048 23866 28060
rect 24464 28048 24492 28079
rect 25366 28076 25372 28088
rect 25424 28076 25430 28128
rect 26473 28119 26531 28125
rect 26473 28116 26485 28119
rect 25476 28088 26485 28116
rect 25476 28048 25504 28088
rect 26473 28085 26485 28088
rect 26519 28085 26531 28119
rect 27025 28119 27083 28125
rect 27025 28116 27037 28119
rect 26473 28079 26531 28085
rect 26580 28088 27037 28116
rect 23860 28020 25504 28048
rect 23860 28008 23866 28020
rect 26286 28008 26292 28060
rect 26344 28048 26350 28060
rect 26580 28048 26608 28088
rect 27025 28085 27037 28088
rect 27071 28085 27083 28119
rect 27025 28079 27083 28085
rect 26344 28020 26608 28048
rect 26344 28008 26350 28020
rect 27390 28008 27396 28060
rect 27448 28048 27454 28060
rect 28037 28051 28095 28057
rect 28037 28048 28049 28051
rect 27448 28020 28049 28048
rect 27448 28008 27454 28020
rect 28037 28017 28049 28020
rect 28083 28017 28095 28051
rect 28037 28011 28095 28017
rect 28218 28008 28224 28060
rect 28276 28048 28282 28060
rect 28773 28051 28831 28057
rect 28773 28048 28785 28051
rect 28276 28020 28785 28048
rect 28276 28008 28282 28020
rect 28773 28017 28785 28020
rect 28819 28017 28831 28051
rect 28773 28011 28831 28017
rect 20490 27980 20496 27992
rect 18484 27952 20496 27980
rect 20490 27940 20496 27952
rect 20548 27940 20554 27992
rect 25366 27940 25372 27992
rect 25424 27980 25430 27992
rect 26378 27980 26384 27992
rect 25424 27952 26384 27980
rect 25424 27940 25430 27952
rect 26378 27940 26384 27952
rect 26436 27980 26442 27992
rect 28129 27983 28187 27989
rect 28129 27980 28141 27983
rect 26436 27952 28141 27980
rect 26436 27940 26442 27952
rect 28129 27949 28141 27952
rect 28175 27949 28187 27983
rect 28129 27943 28187 27949
rect 28310 27940 28316 27992
rect 28368 27980 28374 27992
rect 28865 27983 28923 27989
rect 28865 27980 28877 27983
rect 28368 27952 28877 27980
rect 28368 27940 28374 27952
rect 28865 27949 28877 27952
rect 28911 27949 28923 27983
rect 28865 27943 28923 27949
rect 11000 27890 30136 27912
rect 11000 27838 19142 27890
rect 19194 27838 19206 27890
rect 19258 27838 19270 27890
rect 19322 27838 19334 27890
rect 19386 27838 29142 27890
rect 29194 27838 29206 27890
rect 29258 27838 29270 27890
rect 29322 27838 29334 27890
rect 29386 27838 30136 27890
rect 11000 27816 30136 27838
rect 16721 27779 16779 27785
rect 16721 27745 16733 27779
rect 16767 27776 16779 27779
rect 17638 27776 17644 27788
rect 16767 27748 17644 27776
rect 16767 27745 16779 27748
rect 16721 27739 16779 27745
rect 17638 27736 17644 27748
rect 17696 27736 17702 27788
rect 17822 27736 17828 27788
rect 17880 27776 17886 27788
rect 17880 27748 20444 27776
rect 17880 27736 17886 27748
rect 18834 27708 18840 27720
rect 17932 27680 18840 27708
rect 11934 27600 11940 27652
rect 11992 27640 11998 27652
rect 17932 27649 17960 27680
rect 18834 27668 18840 27680
rect 18892 27668 18898 27720
rect 19478 27668 19484 27720
rect 19536 27708 19542 27720
rect 19573 27711 19631 27717
rect 19573 27708 19585 27711
rect 19536 27680 19585 27708
rect 19536 27668 19542 27680
rect 19573 27677 19585 27680
rect 19619 27677 19631 27711
rect 19573 27671 19631 27677
rect 19849 27711 19907 27717
rect 19849 27677 19861 27711
rect 19895 27677 19907 27711
rect 19849 27671 19907 27677
rect 19941 27711 19999 27717
rect 19941 27677 19953 27711
rect 19987 27677 19999 27711
rect 20306 27708 20312 27720
rect 20267 27680 20312 27708
rect 19941 27671 19999 27677
rect 12213 27643 12271 27649
rect 12213 27640 12225 27643
rect 11992 27612 12225 27640
rect 11992 27600 11998 27612
rect 12213 27609 12225 27612
rect 12259 27640 12271 27643
rect 14697 27643 14755 27649
rect 14697 27640 14709 27643
rect 12259 27612 14709 27640
rect 12259 27609 12271 27612
rect 12213 27603 12271 27609
rect 14697 27609 14709 27612
rect 14743 27609 14755 27643
rect 14697 27603 14755 27609
rect 16629 27643 16687 27649
rect 16629 27609 16641 27643
rect 16675 27640 16687 27643
rect 17273 27643 17331 27649
rect 17273 27640 17285 27643
rect 16675 27612 17285 27640
rect 16675 27609 16687 27612
rect 16629 27603 16687 27609
rect 17273 27609 17285 27612
rect 17319 27609 17331 27643
rect 17273 27603 17331 27609
rect 17917 27643 17975 27649
rect 17917 27609 17929 27643
rect 17963 27609 17975 27643
rect 18282 27640 18288 27652
rect 18243 27612 18288 27640
rect 17917 27603 17975 27609
rect 18282 27600 18288 27612
rect 18340 27600 18346 27652
rect 18469 27643 18527 27649
rect 18469 27609 18481 27643
rect 18515 27609 18527 27643
rect 18469 27603 18527 27609
rect 18006 27572 18012 27584
rect 17967 27544 18012 27572
rect 18006 27532 18012 27544
rect 18064 27532 18070 27584
rect 18484 27572 18512 27603
rect 19018 27600 19024 27652
rect 19076 27640 19082 27652
rect 19754 27640 19760 27652
rect 19076 27612 19760 27640
rect 19076 27600 19082 27612
rect 19754 27600 19760 27612
rect 19812 27600 19818 27652
rect 19386 27572 19392 27584
rect 18484 27544 19392 27572
rect 19386 27532 19392 27544
rect 19444 27532 19450 27584
rect 19864 27572 19892 27671
rect 19588 27544 19892 27572
rect 19956 27572 19984 27671
rect 20306 27668 20312 27680
rect 20364 27668 20370 27720
rect 20416 27708 20444 27748
rect 20490 27736 20496 27788
rect 20548 27776 20554 27788
rect 28218 27776 28224 27788
rect 20548 27748 28224 27776
rect 20548 27736 20554 27748
rect 28218 27736 28224 27748
rect 28276 27736 28282 27788
rect 27390 27708 27396 27720
rect 20416 27680 26884 27708
rect 27351 27680 27396 27708
rect 21778 27640 21784 27652
rect 21739 27612 21784 27640
rect 21778 27600 21784 27612
rect 21836 27600 21842 27652
rect 22606 27640 22612 27652
rect 22567 27612 22612 27640
rect 22606 27600 22612 27612
rect 22664 27600 22670 27652
rect 23066 27600 23072 27652
rect 23124 27640 23130 27652
rect 23437 27643 23495 27649
rect 23437 27640 23449 27643
rect 23124 27612 23449 27640
rect 23124 27600 23130 27612
rect 23437 27609 23449 27612
rect 23483 27609 23495 27643
rect 23437 27603 23495 27609
rect 23526 27600 23532 27652
rect 23584 27640 23590 27652
rect 24173 27643 24231 27649
rect 24173 27640 24185 27643
rect 23584 27612 24185 27640
rect 23584 27600 23590 27612
rect 24173 27609 24185 27612
rect 24219 27640 24231 27643
rect 24906 27640 24912 27652
rect 24219 27612 24912 27640
rect 24219 27609 24231 27612
rect 24173 27603 24231 27609
rect 24906 27600 24912 27612
rect 24964 27640 24970 27652
rect 25274 27640 25280 27652
rect 24964 27612 25280 27640
rect 24964 27600 24970 27612
rect 25274 27600 25280 27612
rect 25332 27600 25338 27652
rect 25369 27643 25427 27649
rect 25369 27609 25381 27643
rect 25415 27609 25427 27643
rect 25826 27640 25832 27652
rect 25787 27612 25832 27640
rect 25369 27603 25427 27609
rect 20674 27572 20680 27584
rect 19956 27544 20680 27572
rect 19588 27448 19616 27544
rect 20674 27532 20680 27544
rect 20732 27532 20738 27584
rect 21873 27575 21931 27581
rect 21873 27541 21885 27575
rect 21919 27541 21931 27575
rect 21873 27535 21931 27541
rect 22701 27575 22759 27581
rect 22701 27541 22713 27575
rect 22747 27572 22759 27575
rect 23250 27572 23256 27584
rect 22747 27544 23256 27572
rect 22747 27541 22759 27544
rect 22701 27535 22759 27541
rect 21888 27504 21916 27535
rect 23250 27532 23256 27544
rect 23308 27532 23314 27584
rect 23342 27532 23348 27584
rect 23400 27572 23406 27584
rect 23400 27544 23445 27572
rect 23400 27532 23406 27544
rect 23894 27532 23900 27584
rect 23952 27572 23958 27584
rect 24265 27575 24323 27581
rect 24265 27572 24277 27575
rect 23952 27544 24277 27572
rect 23952 27532 23958 27544
rect 24265 27541 24277 27544
rect 24311 27541 24323 27575
rect 25384 27572 25412 27603
rect 25826 27600 25832 27612
rect 25884 27600 25890 27652
rect 26749 27643 26807 27649
rect 26749 27609 26761 27643
rect 26795 27609 26807 27643
rect 26856 27640 26884 27680
rect 27390 27668 27396 27680
rect 27448 27668 27454 27720
rect 27853 27643 27911 27649
rect 27853 27640 27865 27643
rect 26856 27612 27865 27640
rect 26749 27603 26807 27609
rect 27853 27609 27865 27612
rect 27899 27640 27911 27643
rect 28402 27640 28408 27652
rect 27899 27612 28408 27640
rect 27899 27609 27911 27612
rect 27853 27603 27911 27609
rect 26764 27572 26792 27603
rect 28402 27600 28408 27612
rect 28460 27600 28466 27652
rect 29141 27643 29199 27649
rect 29141 27609 29153 27643
rect 29187 27640 29199 27643
rect 29506 27640 29512 27652
rect 29187 27612 29512 27640
rect 29187 27609 29199 27612
rect 29141 27603 29199 27609
rect 29506 27600 29512 27612
rect 29564 27600 29570 27652
rect 27758 27572 27764 27584
rect 25384 27544 27764 27572
rect 24265 27535 24323 27541
rect 27758 27532 27764 27544
rect 27816 27532 27822 27584
rect 25090 27504 25096 27516
rect 21888 27476 25096 27504
rect 25090 27464 25096 27476
rect 25148 27464 25154 27516
rect 29138 27504 29144 27516
rect 29099 27476 29144 27504
rect 29138 27464 29144 27476
rect 29196 27464 29202 27516
rect 12302 27396 12308 27448
rect 12360 27436 12366 27448
rect 12397 27439 12455 27445
rect 12397 27436 12409 27439
rect 12360 27408 12409 27436
rect 12360 27396 12366 27408
rect 12397 27405 12409 27408
rect 12443 27405 12455 27439
rect 12397 27399 12455 27405
rect 14786 27396 14792 27448
rect 14844 27436 14850 27448
rect 14881 27439 14939 27445
rect 14881 27436 14893 27439
rect 14844 27408 14893 27436
rect 14844 27396 14850 27408
rect 14881 27405 14893 27408
rect 14927 27405 14939 27439
rect 14881 27399 14939 27405
rect 19570 27396 19576 27448
rect 19628 27396 19634 27448
rect 19662 27396 19668 27448
rect 19720 27436 19726 27448
rect 23342 27436 23348 27448
rect 19720 27408 23348 27436
rect 19720 27396 19726 27408
rect 23342 27396 23348 27408
rect 23400 27396 23406 27448
rect 25185 27439 25243 27445
rect 25185 27405 25197 27439
rect 25231 27436 25243 27439
rect 27022 27436 27028 27448
rect 25231 27408 27028 27436
rect 25231 27405 25243 27408
rect 25185 27399 25243 27405
rect 27022 27396 27028 27408
rect 27080 27396 27086 27448
rect 11000 27346 30136 27368
rect 11000 27294 14142 27346
rect 14194 27294 14206 27346
rect 14258 27294 14270 27346
rect 14322 27294 14334 27346
rect 14386 27294 24142 27346
rect 24194 27294 24206 27346
rect 24258 27294 24270 27346
rect 24322 27294 24334 27346
rect 24386 27294 30136 27346
rect 11000 27272 30136 27294
rect 18006 27192 18012 27244
rect 18064 27232 18070 27244
rect 18193 27235 18251 27241
rect 18193 27232 18205 27235
rect 18064 27204 18205 27232
rect 18064 27192 18070 27204
rect 18193 27201 18205 27204
rect 18239 27201 18251 27235
rect 18193 27195 18251 27201
rect 18742 27192 18748 27244
rect 18800 27232 18806 27244
rect 19662 27232 19668 27244
rect 18800 27204 19668 27232
rect 18800 27192 18806 27204
rect 19662 27192 19668 27204
rect 19720 27192 19726 27244
rect 22146 27232 22152 27244
rect 19956 27204 22152 27232
rect 19386 27124 19392 27176
rect 19444 27164 19450 27176
rect 19956 27164 19984 27204
rect 22146 27192 22152 27204
rect 22204 27232 22210 27244
rect 25734 27232 25740 27244
rect 22204 27204 25740 27232
rect 22204 27192 22210 27204
rect 25734 27192 25740 27204
rect 25792 27192 25798 27244
rect 19444 27136 19984 27164
rect 19444 27124 19450 27136
rect 20030 27124 20036 27176
rect 20088 27164 20094 27176
rect 23986 27164 23992 27176
rect 20088 27136 23992 27164
rect 20088 27124 20094 27136
rect 23986 27124 23992 27136
rect 24044 27124 24050 27176
rect 27117 27167 27175 27173
rect 27117 27133 27129 27167
rect 27163 27164 27175 27167
rect 27390 27164 27396 27176
rect 27163 27136 27396 27164
rect 27163 27133 27175 27136
rect 27117 27127 27175 27133
rect 27390 27124 27396 27136
rect 27448 27124 27454 27176
rect 13777 27099 13835 27105
rect 13777 27096 13789 27099
rect 11308 27068 13789 27096
rect 11308 27040 11336 27068
rect 13777 27065 13789 27068
rect 13823 27065 13835 27099
rect 13777 27059 13835 27065
rect 16902 27056 16908 27108
rect 16960 27096 16966 27108
rect 19018 27096 19024 27108
rect 16960 27068 19024 27096
rect 16960 27056 16966 27068
rect 19018 27056 19024 27068
rect 19076 27056 19082 27108
rect 19665 27099 19723 27105
rect 19665 27065 19677 27099
rect 19711 27096 19723 27099
rect 20582 27096 20588 27108
rect 19711 27068 20588 27096
rect 19711 27065 19723 27068
rect 19665 27059 19723 27065
rect 20582 27056 20588 27068
rect 20640 27056 20646 27108
rect 23802 27096 23808 27108
rect 23763 27068 23808 27096
rect 23802 27056 23808 27068
rect 23860 27056 23866 27108
rect 24446 27056 24452 27108
rect 24504 27096 24510 27108
rect 24633 27099 24691 27105
rect 24633 27096 24645 27099
rect 24504 27068 24645 27096
rect 24504 27056 24510 27068
rect 24633 27065 24645 27068
rect 24679 27065 24691 27099
rect 24633 27059 24691 27065
rect 25826 27056 25832 27108
rect 25884 27096 25890 27108
rect 26378 27096 26384 27108
rect 25884 27068 26384 27096
rect 25884 27056 25890 27068
rect 26378 27056 26384 27068
rect 26436 27096 26442 27108
rect 26657 27099 26715 27105
rect 26657 27096 26669 27099
rect 26436 27068 26669 27096
rect 26436 27056 26442 27068
rect 26657 27065 26669 27068
rect 26703 27065 26715 27099
rect 27206 27096 27212 27108
rect 27167 27068 27212 27096
rect 26657 27059 26715 27065
rect 27206 27056 27212 27068
rect 27264 27056 27270 27108
rect 28402 27096 28408 27108
rect 28363 27068 28408 27096
rect 28402 27056 28408 27068
rect 28460 27056 28466 27108
rect 28862 27056 28868 27108
rect 28920 27096 28926 27108
rect 28957 27099 29015 27105
rect 28957 27096 28969 27099
rect 28920 27068 28969 27096
rect 28920 27056 28926 27068
rect 28957 27065 28969 27068
rect 29003 27065 29015 27099
rect 28957 27059 29015 27065
rect 11290 27028 11296 27040
rect 11251 27000 11296 27028
rect 11290 26988 11296 27000
rect 11348 26988 11354 27040
rect 16997 27031 17055 27037
rect 16997 26997 17009 27031
rect 17043 27028 17055 27031
rect 17730 27028 17736 27040
rect 17043 27000 17736 27028
rect 17043 26997 17055 27000
rect 16997 26991 17055 26997
rect 17730 26988 17736 27000
rect 17788 27028 17794 27040
rect 18101 27031 18159 27037
rect 17788 27000 18052 27028
rect 17788 26988 17794 27000
rect 11566 26960 11572 26972
rect 11527 26932 11572 26960
rect 11566 26920 11572 26932
rect 11624 26920 11630 26972
rect 12302 26920 12308 26972
rect 12360 26920 12366 26972
rect 13222 26920 13228 26972
rect 13280 26960 13286 26972
rect 13317 26963 13375 26969
rect 13317 26960 13329 26963
rect 13280 26932 13329 26960
rect 13280 26920 13286 26932
rect 13317 26929 13329 26932
rect 13363 26929 13375 26963
rect 14050 26960 14056 26972
rect 14011 26932 14056 26960
rect 13317 26923 13375 26929
rect 14050 26920 14056 26932
rect 14108 26920 14114 26972
rect 14786 26920 14792 26972
rect 14844 26920 14850 26972
rect 15798 26960 15804 26972
rect 15759 26932 15804 26960
rect 15798 26920 15804 26932
rect 15856 26920 15862 26972
rect 16718 26960 16724 26972
rect 16679 26932 16724 26960
rect 16718 26920 16724 26932
rect 16776 26920 16782 26972
rect 17089 26963 17147 26969
rect 17089 26929 17101 26963
rect 17135 26929 17147 26963
rect 17089 26923 17147 26929
rect 17457 26963 17515 26969
rect 17457 26929 17469 26963
rect 17503 26960 17515 26963
rect 17917 26963 17975 26969
rect 17917 26960 17929 26963
rect 17503 26932 17929 26960
rect 17503 26929 17515 26932
rect 17457 26923 17515 26929
rect 17917 26929 17929 26932
rect 17963 26929 17975 26963
rect 17917 26923 17975 26929
rect 16902 26892 16908 26904
rect 16863 26864 16908 26892
rect 16902 26852 16908 26864
rect 16960 26852 16966 26904
rect 17104 26892 17132 26923
rect 17822 26892 17828 26904
rect 17104 26864 17828 26892
rect 17822 26852 17828 26864
rect 17880 26852 17886 26904
rect 18024 26892 18052 27000
rect 18101 26997 18113 27031
rect 18147 27028 18159 27031
rect 18742 27028 18748 27040
rect 18147 27000 18748 27028
rect 18147 26997 18159 27000
rect 18101 26991 18159 26997
rect 18742 26988 18748 27000
rect 18800 26988 18806 27040
rect 19570 27028 19576 27040
rect 19220 27000 19576 27028
rect 18926 26960 18932 26972
rect 18887 26932 18932 26960
rect 18926 26920 18932 26932
rect 18984 26920 18990 26972
rect 19018 26920 19024 26972
rect 19076 26960 19082 26972
rect 19113 26963 19171 26969
rect 19113 26960 19125 26963
rect 19076 26932 19125 26960
rect 19076 26920 19082 26932
rect 19113 26929 19125 26932
rect 19159 26929 19171 26963
rect 19113 26923 19171 26929
rect 19220 26901 19248 27000
rect 19570 26988 19576 27000
rect 19628 27028 19634 27040
rect 19938 27028 19944 27040
rect 19628 27000 19944 27028
rect 19628 26988 19634 27000
rect 19938 26988 19944 27000
rect 19996 26988 20002 27040
rect 20214 27028 20220 27040
rect 20048 27000 20220 27028
rect 19297 26963 19355 26969
rect 19297 26929 19309 26963
rect 19343 26960 19355 26963
rect 20048 26960 20076 27000
rect 20214 26988 20220 27000
rect 20272 27028 20278 27040
rect 20272 27000 20536 27028
rect 20272 26988 20278 27000
rect 20508 26969 20536 27000
rect 22054 26988 22060 27040
rect 22112 27028 22118 27040
rect 22701 27031 22759 27037
rect 22701 27028 22713 27031
rect 22112 27000 22713 27028
rect 22112 26988 22118 27000
rect 22701 26997 22713 27000
rect 22747 26997 22759 27031
rect 22701 26991 22759 26997
rect 23069 27031 23127 27037
rect 23069 26997 23081 27031
rect 23115 27028 23127 27031
rect 23710 27028 23716 27040
rect 23115 27000 23716 27028
rect 23115 26997 23127 27000
rect 23069 26991 23127 26997
rect 23710 26988 23716 27000
rect 23768 26988 23774 27040
rect 24541 27031 24599 27037
rect 24541 26997 24553 27031
rect 24587 27028 24599 27031
rect 24906 27028 24912 27040
rect 24587 27000 24912 27028
rect 24587 26997 24599 27000
rect 24541 26991 24599 26997
rect 24906 26988 24912 27000
rect 24964 26988 24970 27040
rect 25550 27028 25556 27040
rect 25511 27000 25556 27028
rect 25550 26988 25556 27000
rect 25608 26988 25614 27040
rect 19343 26932 20076 26960
rect 20125 26963 20183 26969
rect 19343 26929 19355 26932
rect 19297 26923 19355 26929
rect 20125 26929 20137 26963
rect 20171 26929 20183 26963
rect 20125 26923 20183 26929
rect 20493 26963 20551 26969
rect 20493 26929 20505 26963
rect 20539 26929 20551 26963
rect 20493 26923 20551 26929
rect 20861 26963 20919 26969
rect 20861 26929 20873 26963
rect 20907 26960 20919 26963
rect 21594 26960 21600 26972
rect 20907 26932 21600 26960
rect 20907 26929 20919 26932
rect 20861 26923 20919 26929
rect 19205 26895 19263 26901
rect 19205 26892 19217 26895
rect 18024 26864 19217 26892
rect 19205 26861 19217 26864
rect 19251 26861 19263 26895
rect 19205 26855 19263 26861
rect 19478 26852 19484 26904
rect 19536 26892 19542 26904
rect 20140 26892 20168 26923
rect 21594 26920 21600 26932
rect 21652 26920 21658 26972
rect 22514 26960 22520 26972
rect 22475 26932 22520 26960
rect 22514 26920 22520 26932
rect 22572 26920 22578 26972
rect 28494 26920 28500 26972
rect 28552 26960 28558 26972
rect 28865 26963 28923 26969
rect 28865 26960 28877 26963
rect 28552 26932 28877 26960
rect 28552 26920 28558 26932
rect 28865 26929 28877 26932
rect 28911 26960 28923 26963
rect 29138 26960 29144 26972
rect 28911 26932 29144 26960
rect 28911 26929 28923 26932
rect 28865 26923 28923 26929
rect 29138 26920 29144 26932
rect 29196 26920 29202 26972
rect 20306 26892 20312 26904
rect 19536 26864 20168 26892
rect 20267 26864 20312 26892
rect 19536 26852 19542 26864
rect 20306 26852 20312 26864
rect 20364 26852 20370 26904
rect 20398 26852 20404 26904
rect 20456 26892 20462 26904
rect 25645 26895 25703 26901
rect 20456 26864 20501 26892
rect 20456 26852 20462 26864
rect 25645 26861 25657 26895
rect 25691 26892 25703 26895
rect 26470 26892 26476 26904
rect 25691 26864 26476 26892
rect 25691 26861 25703 26864
rect 25645 26855 25703 26861
rect 26470 26852 26476 26864
rect 26528 26852 26534 26904
rect 11000 26802 30136 26824
rect 11000 26750 19142 26802
rect 19194 26750 19206 26802
rect 19258 26750 19270 26802
rect 19322 26750 19334 26802
rect 19386 26750 29142 26802
rect 29194 26750 29206 26802
rect 29258 26750 29270 26802
rect 29322 26750 29334 26802
rect 29386 26750 30136 26802
rect 11000 26728 30136 26750
rect 15798 26648 15804 26700
rect 15856 26688 15862 26700
rect 20306 26688 20312 26700
rect 15856 26660 20312 26688
rect 15856 26648 15862 26660
rect 11566 26580 11572 26632
rect 11624 26620 11630 26632
rect 11937 26623 11995 26629
rect 11937 26620 11949 26623
rect 11624 26592 11949 26620
rect 11624 26580 11630 26592
rect 11937 26589 11949 26592
rect 11983 26589 11995 26623
rect 11937 26583 11995 26589
rect 12489 26555 12547 26561
rect 12489 26521 12501 26555
rect 12535 26552 12547 26555
rect 12578 26552 12584 26564
rect 12535 26524 12584 26552
rect 12535 26521 12547 26524
rect 12489 26515 12547 26521
rect 12578 26512 12584 26524
rect 12636 26512 12642 26564
rect 12670 26512 12676 26564
rect 12728 26552 12734 26564
rect 12854 26552 12860 26564
rect 12728 26524 12773 26552
rect 12815 26524 12860 26552
rect 12728 26512 12734 26524
rect 12854 26512 12860 26524
rect 12912 26512 12918 26564
rect 13222 26552 13228 26564
rect 13183 26524 13228 26552
rect 13222 26512 13228 26524
rect 13280 26512 13286 26564
rect 15246 26552 15252 26564
rect 15159 26524 15252 26552
rect 15246 26512 15252 26524
rect 15304 26552 15310 26564
rect 15816 26552 15844 26648
rect 15304 26524 15844 26552
rect 15893 26555 15951 26561
rect 15304 26512 15310 26524
rect 15893 26521 15905 26555
rect 15939 26521 15951 26555
rect 15893 26515 15951 26521
rect 13130 26444 13136 26496
rect 13188 26484 13194 26496
rect 13317 26487 13375 26493
rect 13317 26484 13329 26487
rect 13188 26456 13329 26484
rect 13188 26444 13194 26456
rect 13317 26453 13329 26456
rect 13363 26484 13375 26487
rect 15338 26484 15344 26496
rect 13363 26456 15344 26484
rect 13363 26453 13375 26456
rect 13317 26447 13375 26453
rect 15338 26444 15344 26456
rect 15396 26444 15402 26496
rect 13222 26376 13228 26428
rect 13280 26416 13286 26428
rect 15908 26416 15936 26515
rect 17546 26512 17552 26564
rect 17604 26552 17610 26564
rect 17656 26561 17684 26660
rect 20306 26648 20312 26660
rect 20364 26648 20370 26700
rect 22514 26648 22520 26700
rect 22572 26688 22578 26700
rect 22793 26691 22851 26697
rect 22793 26688 22805 26691
rect 22572 26660 22805 26688
rect 22572 26648 22578 26660
rect 22793 26657 22805 26660
rect 22839 26657 22851 26691
rect 22793 26651 22851 26657
rect 23618 26648 23624 26700
rect 23676 26688 23682 26700
rect 26378 26688 26384 26700
rect 23676 26660 25964 26688
rect 26339 26660 26384 26688
rect 23676 26648 23682 26660
rect 17822 26620 17828 26632
rect 17735 26592 17828 26620
rect 17822 26580 17828 26592
rect 17880 26620 17886 26632
rect 18006 26620 18012 26632
rect 17880 26592 18012 26620
rect 17880 26580 17886 26592
rect 18006 26580 18012 26592
rect 18064 26580 18070 26632
rect 19938 26580 19944 26632
rect 19996 26620 20002 26632
rect 20398 26620 20404 26632
rect 19996 26592 20404 26620
rect 19996 26580 20002 26592
rect 20398 26580 20404 26592
rect 20456 26580 20462 26632
rect 20493 26623 20551 26629
rect 20493 26589 20505 26623
rect 20539 26620 20551 26623
rect 20674 26620 20680 26632
rect 20539 26592 20680 26620
rect 20539 26589 20551 26592
rect 20493 26583 20551 26589
rect 20674 26580 20680 26592
rect 20732 26580 20738 26632
rect 21505 26623 21563 26629
rect 21505 26589 21517 26623
rect 21551 26620 21563 26623
rect 21594 26620 21600 26632
rect 21551 26592 21600 26620
rect 21551 26589 21563 26592
rect 21505 26583 21563 26589
rect 21594 26580 21600 26592
rect 21652 26580 21658 26632
rect 22054 26620 22060 26632
rect 22015 26592 22060 26620
rect 22054 26580 22060 26592
rect 22112 26580 22118 26632
rect 23710 26620 23716 26632
rect 23671 26592 23716 26620
rect 23710 26580 23716 26592
rect 23768 26580 23774 26632
rect 17641 26555 17699 26561
rect 17641 26552 17653 26555
rect 17604 26524 17653 26552
rect 17604 26512 17610 26524
rect 17641 26521 17653 26524
rect 17687 26521 17699 26555
rect 17641 26515 17699 26521
rect 17730 26512 17736 26564
rect 17788 26552 17794 26564
rect 18926 26552 18932 26564
rect 17788 26524 17833 26552
rect 18116 26524 18932 26552
rect 17788 26512 17794 26524
rect 16718 26444 16724 26496
rect 16776 26484 16782 26496
rect 17457 26487 17515 26493
rect 17457 26484 17469 26487
rect 16776 26456 17469 26484
rect 16776 26444 16782 26456
rect 17457 26453 17469 26456
rect 17503 26484 17515 26487
rect 18116 26484 18144 26524
rect 18926 26512 18932 26524
rect 18984 26552 18990 26564
rect 19478 26552 19484 26564
rect 18984 26524 19484 26552
rect 18984 26512 18990 26524
rect 19478 26512 19484 26524
rect 19536 26552 19542 26564
rect 20125 26555 20183 26561
rect 20125 26552 20137 26555
rect 19536 26524 20137 26552
rect 19536 26512 19542 26524
rect 20125 26521 20137 26524
rect 20171 26521 20183 26555
rect 21686 26552 21692 26564
rect 21647 26524 21692 26552
rect 20125 26515 20183 26521
rect 21686 26512 21692 26524
rect 21744 26512 21750 26564
rect 21870 26512 21876 26564
rect 21928 26552 21934 26564
rect 22517 26555 22575 26561
rect 22517 26552 22529 26555
rect 21928 26524 22529 26552
rect 21928 26512 21934 26524
rect 22517 26521 22529 26524
rect 22563 26521 22575 26555
rect 22517 26515 22575 26521
rect 22701 26555 22759 26561
rect 22701 26521 22713 26555
rect 22747 26521 22759 26555
rect 22701 26515 22759 26521
rect 17503 26456 18144 26484
rect 18193 26487 18251 26493
rect 17503 26453 17515 26456
rect 17457 26447 17515 26453
rect 18193 26453 18205 26487
rect 18239 26484 18251 26487
rect 18466 26484 18472 26496
rect 18239 26456 18472 26484
rect 18239 26453 18251 26456
rect 18193 26447 18251 26453
rect 18466 26444 18472 26456
rect 18524 26484 18530 26496
rect 19938 26484 19944 26496
rect 18524 26456 19944 26484
rect 18524 26444 18530 26456
rect 19938 26444 19944 26456
rect 19996 26444 20002 26496
rect 20861 26487 20919 26493
rect 20861 26453 20873 26487
rect 20907 26484 20919 26487
rect 21704 26484 21732 26512
rect 20907 26456 21732 26484
rect 20907 26453 20919 26456
rect 20861 26447 20919 26453
rect 21778 26444 21784 26496
rect 21836 26484 21842 26496
rect 22716 26484 22744 26515
rect 22882 26512 22888 26564
rect 22940 26552 22946 26564
rect 23897 26555 23955 26561
rect 23897 26552 23909 26555
rect 22940 26524 23909 26552
rect 22940 26512 22946 26524
rect 23897 26521 23909 26524
rect 23943 26521 23955 26555
rect 23897 26515 23955 26521
rect 25369 26555 25427 26561
rect 25369 26521 25381 26555
rect 25415 26552 25427 26555
rect 25826 26552 25832 26564
rect 25415 26524 25832 26552
rect 25415 26521 25427 26524
rect 25369 26515 25427 26521
rect 25826 26512 25832 26524
rect 25884 26512 25890 26564
rect 25936 26561 25964 26660
rect 26378 26648 26384 26660
rect 26436 26648 26442 26700
rect 28589 26691 28647 26697
rect 28589 26688 28601 26691
rect 27960 26660 28601 26688
rect 27114 26580 27120 26632
rect 27172 26620 27178 26632
rect 27669 26623 27727 26629
rect 27669 26620 27681 26623
rect 27172 26592 27681 26620
rect 27172 26580 27178 26592
rect 27669 26589 27681 26592
rect 27715 26589 27727 26623
rect 27669 26583 27727 26589
rect 27758 26580 27764 26632
rect 27816 26620 27822 26632
rect 27960 26629 27988 26660
rect 28589 26657 28601 26660
rect 28635 26657 28647 26691
rect 28589 26651 28647 26657
rect 27945 26623 28003 26629
rect 27945 26620 27957 26623
rect 27816 26592 27957 26620
rect 27816 26580 27822 26592
rect 27945 26589 27957 26592
rect 27991 26589 28003 26623
rect 28494 26620 28500 26632
rect 28455 26592 28500 26620
rect 27945 26583 28003 26589
rect 28494 26580 28500 26592
rect 28552 26580 28558 26632
rect 25921 26555 25979 26561
rect 25921 26521 25933 26555
rect 25967 26521 25979 26555
rect 25921 26515 25979 26521
rect 26105 26555 26163 26561
rect 26105 26521 26117 26555
rect 26151 26552 26163 26555
rect 26151 26524 26332 26552
rect 26151 26521 26163 26524
rect 26105 26515 26163 26521
rect 21836 26456 22744 26484
rect 24265 26487 24323 26493
rect 21836 26444 21842 26456
rect 24265 26453 24277 26487
rect 24311 26453 24323 26487
rect 24265 26447 24323 26453
rect 18282 26416 18288 26428
rect 13280 26388 18288 26416
rect 13280 26376 13286 26388
rect 18282 26376 18288 26388
rect 18340 26376 18346 26428
rect 24280 26416 24308 26447
rect 24906 26444 24912 26496
rect 24964 26484 24970 26496
rect 25185 26487 25243 26493
rect 25185 26484 25197 26487
rect 24964 26456 25197 26484
rect 24964 26444 24970 26456
rect 25185 26453 25197 26456
rect 25231 26453 25243 26487
rect 25185 26447 25243 26453
rect 26304 26416 26332 26524
rect 26470 26512 26476 26564
rect 26528 26552 26534 26564
rect 27025 26555 27083 26561
rect 27025 26552 27037 26555
rect 26528 26524 27037 26552
rect 26528 26512 26534 26524
rect 27025 26521 27037 26524
rect 27071 26521 27083 26555
rect 27025 26515 27083 26521
rect 28954 26512 28960 26564
rect 29012 26552 29018 26564
rect 29141 26555 29199 26561
rect 29141 26552 29153 26555
rect 29012 26524 29153 26552
rect 29012 26512 29018 26524
rect 29141 26521 29153 26524
rect 29187 26521 29199 26555
rect 29141 26515 29199 26521
rect 26378 26416 26384 26428
rect 24280 26388 26384 26416
rect 26378 26376 26384 26388
rect 26436 26376 26442 26428
rect 27574 26376 27580 26428
rect 27632 26416 27638 26428
rect 29233 26419 29291 26425
rect 29233 26416 29245 26419
rect 27632 26388 29245 26416
rect 27632 26376 27638 26388
rect 29233 26385 29245 26388
rect 29279 26385 29291 26419
rect 29233 26379 29291 26385
rect 14970 26308 14976 26360
rect 15028 26348 15034 26360
rect 15341 26351 15399 26357
rect 15341 26348 15353 26351
rect 15028 26320 15353 26348
rect 15028 26308 15034 26320
rect 15341 26317 15353 26320
rect 15387 26317 15399 26351
rect 15341 26311 15399 26317
rect 15985 26351 16043 26357
rect 15985 26317 15997 26351
rect 16031 26348 16043 26351
rect 16718 26348 16724 26360
rect 16031 26320 16724 26348
rect 16031 26317 16043 26320
rect 15985 26311 16043 26317
rect 16718 26308 16724 26320
rect 16776 26308 16782 26360
rect 11000 26258 30136 26280
rect 11000 26206 14142 26258
rect 14194 26206 14206 26258
rect 14258 26206 14270 26258
rect 14322 26206 14334 26258
rect 14386 26206 24142 26258
rect 24194 26206 24206 26258
rect 24258 26206 24270 26258
rect 24322 26206 24334 26258
rect 24386 26206 30136 26258
rect 11000 26184 30136 26206
rect 12578 26144 12584 26156
rect 12539 26116 12584 26144
rect 12578 26104 12584 26116
rect 12636 26104 12642 26156
rect 24909 26147 24967 26153
rect 19480 26116 22652 26144
rect 12854 26036 12860 26088
rect 12912 26076 12918 26088
rect 15985 26079 16043 26085
rect 15985 26076 15997 26079
rect 12912 26048 15997 26076
rect 12912 26036 12918 26048
rect 13961 26011 14019 26017
rect 13961 25977 13973 26011
rect 14007 26008 14019 26011
rect 14050 26008 14056 26020
rect 14007 25980 14056 26008
rect 14007 25977 14019 25980
rect 13961 25971 14019 25977
rect 14050 25968 14056 25980
rect 14108 25968 14114 26020
rect 11658 25940 11664 25952
rect 11619 25912 11664 25940
rect 11658 25900 11664 25912
rect 11716 25900 11722 25952
rect 12762 25940 12768 25952
rect 12723 25912 12768 25940
rect 12762 25900 12768 25912
rect 12820 25900 12826 25952
rect 13225 25943 13283 25949
rect 13225 25909 13237 25943
rect 13271 25940 13283 25943
rect 13498 25940 13504 25952
rect 13271 25912 13504 25940
rect 13271 25909 13283 25912
rect 13225 25903 13283 25909
rect 13498 25900 13504 25912
rect 13556 25900 13562 25952
rect 14421 25943 14479 25949
rect 14421 25909 14433 25943
rect 14467 25909 14479 25943
rect 14421 25903 14479 25909
rect 14436 25872 14464 25903
rect 14510 25900 14516 25952
rect 14568 25940 14574 25952
rect 14804 25949 14832 26048
rect 15985 26045 15997 26048
rect 16031 26045 16043 26079
rect 19480 26076 19508 26116
rect 15985 26039 16043 26045
rect 16092 26048 19508 26076
rect 22624 26076 22652 26116
rect 24909 26113 24921 26147
rect 24955 26144 24967 26147
rect 25550 26144 25556 26156
rect 24955 26116 25556 26144
rect 24955 26113 24967 26116
rect 24909 26107 24967 26113
rect 25550 26104 25556 26116
rect 25608 26104 25614 26156
rect 26933 26079 26991 26085
rect 22624 26048 25688 26076
rect 15246 26008 15252 26020
rect 15207 25980 15252 26008
rect 15246 25968 15252 25980
rect 15304 25968 15310 26020
rect 15338 25968 15344 26020
rect 15396 26008 15402 26020
rect 15396 25980 15936 26008
rect 15396 25968 15402 25980
rect 14605 25943 14663 25949
rect 14605 25940 14617 25943
rect 14568 25912 14617 25940
rect 14568 25900 14574 25912
rect 14605 25909 14617 25912
rect 14651 25909 14663 25943
rect 14605 25903 14663 25909
rect 14789 25943 14847 25949
rect 14789 25909 14801 25943
rect 14835 25909 14847 25943
rect 14789 25903 14847 25909
rect 14878 25900 14884 25952
rect 14936 25940 14942 25952
rect 15908 25949 15936 25980
rect 15893 25943 15951 25949
rect 14936 25912 15844 25940
rect 14936 25900 14942 25912
rect 15706 25872 15712 25884
rect 14436 25844 15712 25872
rect 15706 25832 15712 25844
rect 15764 25832 15770 25884
rect 15816 25872 15844 25912
rect 15893 25909 15905 25943
rect 15939 25909 15951 25943
rect 15893 25903 15951 25909
rect 16092 25872 16120 26048
rect 18006 25968 18012 26020
rect 18064 26008 18070 26020
rect 18558 26008 18564 26020
rect 18064 25980 18564 26008
rect 18064 25968 18070 25980
rect 16902 25940 16908 25952
rect 16815 25912 16908 25940
rect 16718 25872 16724 25884
rect 15816 25844 16120 25872
rect 16679 25844 16724 25872
rect 16718 25832 16724 25844
rect 16776 25832 16782 25884
rect 11753 25807 11811 25813
rect 11753 25773 11765 25807
rect 11799 25804 11811 25807
rect 14878 25804 14884 25816
rect 11799 25776 14884 25804
rect 11799 25773 11811 25776
rect 11753 25767 11811 25773
rect 14878 25764 14884 25776
rect 14936 25764 14942 25816
rect 14970 25764 14976 25816
rect 15028 25804 15034 25816
rect 16828 25804 16856 25912
rect 16902 25900 16908 25912
rect 16960 25900 16966 25952
rect 17178 25900 17184 25952
rect 17236 25940 17242 25952
rect 17730 25940 17736 25952
rect 17236 25912 17736 25940
rect 17236 25900 17242 25912
rect 17730 25900 17736 25912
rect 17788 25940 17794 25952
rect 18116 25949 18144 25980
rect 18558 25968 18564 25980
rect 18616 25968 18622 26020
rect 21778 26008 21784 26020
rect 21428 25980 21784 26008
rect 21428 25952 21456 25980
rect 21778 25968 21784 25980
rect 21836 25968 21842 26020
rect 25366 26008 25372 26020
rect 25327 25980 25372 26008
rect 25366 25968 25372 25980
rect 25424 25968 25430 26020
rect 17917 25943 17975 25949
rect 17917 25940 17929 25943
rect 17788 25912 17929 25940
rect 17788 25900 17794 25912
rect 17917 25909 17929 25912
rect 17963 25909 17975 25943
rect 17917 25903 17975 25909
rect 18101 25943 18159 25949
rect 18101 25909 18113 25943
rect 18147 25909 18159 25943
rect 18101 25903 18159 25909
rect 18190 25900 18196 25952
rect 18248 25940 18254 25952
rect 18653 25943 18711 25949
rect 18653 25940 18665 25943
rect 18248 25912 18665 25940
rect 18248 25900 18254 25912
rect 18653 25909 18665 25912
rect 18699 25909 18711 25943
rect 18653 25903 18711 25909
rect 18926 25900 18932 25952
rect 18984 25940 18990 25952
rect 19297 25943 19355 25949
rect 19297 25940 19309 25943
rect 18984 25912 19309 25940
rect 18984 25900 18990 25912
rect 19297 25909 19309 25912
rect 19343 25940 19355 25943
rect 20309 25943 20367 25949
rect 20309 25940 20321 25943
rect 19343 25912 20321 25940
rect 19343 25909 19355 25912
rect 19297 25903 19355 25909
rect 20309 25909 20321 25912
rect 20355 25909 20367 25943
rect 21410 25940 21416 25952
rect 21323 25912 21416 25940
rect 20309 25903 20367 25909
rect 21410 25900 21416 25912
rect 21468 25900 21474 25952
rect 21686 25900 21692 25952
rect 21744 25940 21750 25952
rect 23161 25943 23219 25949
rect 23161 25940 23173 25943
rect 21744 25912 23173 25940
rect 21744 25900 21750 25912
rect 23161 25909 23173 25912
rect 23207 25909 23219 25943
rect 23161 25903 23219 25909
rect 23345 25943 23403 25949
rect 23345 25909 23357 25943
rect 23391 25909 23403 25943
rect 25274 25940 25280 25952
rect 25235 25912 25280 25940
rect 23345 25903 23403 25909
rect 17089 25875 17147 25881
rect 17089 25872 17101 25875
rect 16920 25844 17101 25872
rect 16920 25816 16948 25844
rect 17089 25841 17101 25844
rect 17135 25841 17147 25875
rect 17089 25835 17147 25841
rect 17270 25832 17276 25884
rect 17328 25872 17334 25884
rect 17457 25875 17515 25881
rect 17457 25872 17469 25875
rect 17328 25844 17469 25872
rect 17328 25832 17334 25844
rect 17457 25841 17469 25844
rect 17503 25841 17515 25875
rect 17457 25835 17515 25841
rect 17546 25832 17552 25884
rect 17604 25872 17610 25884
rect 18285 25875 18343 25881
rect 18285 25872 18297 25875
rect 17604 25844 18297 25872
rect 17604 25832 17610 25844
rect 18285 25841 18297 25844
rect 18331 25841 18343 25875
rect 18285 25835 18343 25841
rect 19018 25832 19024 25884
rect 19076 25872 19082 25884
rect 19113 25875 19171 25881
rect 19113 25872 19125 25875
rect 19076 25844 19125 25872
rect 19076 25832 19082 25844
rect 19113 25841 19125 25844
rect 19159 25841 19171 25875
rect 19113 25835 19171 25841
rect 20125 25875 20183 25881
rect 20125 25841 20137 25875
rect 20171 25841 20183 25875
rect 20125 25835 20183 25841
rect 15028 25776 16856 25804
rect 15028 25764 15034 25776
rect 16902 25764 16908 25816
rect 16960 25764 16966 25816
rect 16994 25764 17000 25816
rect 17052 25804 17058 25816
rect 17052 25776 17097 25804
rect 17052 25764 17058 25776
rect 18098 25764 18104 25816
rect 18156 25804 18162 25816
rect 18193 25807 18251 25813
rect 18193 25804 18205 25807
rect 18156 25776 18205 25804
rect 18156 25764 18162 25776
rect 18193 25773 18205 25776
rect 18239 25773 18251 25807
rect 18193 25767 18251 25773
rect 18374 25764 18380 25816
rect 18432 25804 18438 25816
rect 19389 25807 19447 25813
rect 19389 25804 19401 25807
rect 18432 25776 19401 25804
rect 18432 25764 18438 25776
rect 19389 25773 19401 25776
rect 19435 25773 19447 25807
rect 20140 25804 20168 25835
rect 20582 25832 20588 25884
rect 20640 25872 20646 25884
rect 20677 25875 20735 25881
rect 20677 25872 20689 25875
rect 20640 25844 20689 25872
rect 20640 25832 20646 25844
rect 20677 25841 20689 25844
rect 20723 25841 20735 25875
rect 21226 25872 21232 25884
rect 21187 25844 21232 25872
rect 20677 25835 20735 25841
rect 21226 25832 21232 25844
rect 21284 25832 21290 25884
rect 21781 25875 21839 25881
rect 21781 25841 21793 25875
rect 21827 25872 21839 25875
rect 22514 25872 22520 25884
rect 21827 25844 22520 25872
rect 21827 25841 21839 25844
rect 21781 25835 21839 25841
rect 22514 25832 22520 25844
rect 22572 25832 22578 25884
rect 22882 25832 22888 25884
rect 22940 25872 22946 25884
rect 23360 25872 23388 25903
rect 25274 25900 25280 25912
rect 25332 25900 25338 25952
rect 25660 25949 25688 26048
rect 26933 26045 26945 26079
rect 26979 26076 26991 26079
rect 27114 26076 27120 26088
rect 26979 26048 27120 26076
rect 26979 26045 26991 26048
rect 26933 26039 26991 26045
rect 27114 26036 27120 26048
rect 27172 26036 27178 26088
rect 28678 26036 28684 26088
rect 28736 26076 28742 26088
rect 28865 26079 28923 26085
rect 28865 26076 28877 26079
rect 28736 26048 28877 26076
rect 28736 26036 28742 26048
rect 28865 26045 28877 26048
rect 28911 26045 28923 26079
rect 28865 26039 28923 26045
rect 26470 26008 26476 26020
rect 26431 25980 26476 26008
rect 26470 25968 26476 25980
rect 26528 25968 26534 26020
rect 27022 26008 27028 26020
rect 26983 25980 27028 26008
rect 27022 25968 27028 25980
rect 27080 25968 27086 26020
rect 28770 25968 28776 26020
rect 28828 26008 28834 26020
rect 28957 26011 29015 26017
rect 28957 26008 28969 26011
rect 28828 25980 28969 26008
rect 28828 25968 28834 25980
rect 28957 25977 28969 25980
rect 29003 25977 29015 26011
rect 28957 25971 29015 25977
rect 25645 25943 25703 25949
rect 25645 25909 25657 25943
rect 25691 25909 25703 25943
rect 25645 25903 25703 25909
rect 25734 25900 25740 25952
rect 25792 25940 25798 25952
rect 25792 25912 25837 25940
rect 25792 25900 25798 25912
rect 28034 25900 28040 25952
rect 28092 25940 28098 25952
rect 28405 25943 28463 25949
rect 28405 25940 28417 25943
rect 28092 25912 28417 25940
rect 28092 25900 28098 25912
rect 28405 25909 28417 25912
rect 28451 25909 28463 25943
rect 28405 25903 28463 25909
rect 22940 25844 23388 25872
rect 23713 25875 23771 25881
rect 22940 25832 22946 25844
rect 23713 25841 23725 25875
rect 23759 25872 23771 25875
rect 24170 25872 24176 25884
rect 23759 25844 24176 25872
rect 23759 25841 23771 25844
rect 23713 25835 23771 25841
rect 24170 25832 24176 25844
rect 24228 25832 24234 25884
rect 21686 25804 21692 25816
rect 20140 25776 21692 25804
rect 19389 25767 19447 25773
rect 21686 25764 21692 25776
rect 21744 25804 21750 25816
rect 23434 25804 23440 25816
rect 21744 25776 23440 25804
rect 21744 25764 21750 25776
rect 23434 25764 23440 25776
rect 23492 25764 23498 25816
rect 11000 25714 30136 25736
rect 11000 25662 19142 25714
rect 19194 25662 19206 25714
rect 19258 25662 19270 25714
rect 19322 25662 19334 25714
rect 19386 25662 29142 25714
rect 29194 25662 29206 25714
rect 29258 25662 29270 25714
rect 29322 25662 29334 25714
rect 29386 25662 30136 25714
rect 11000 25640 30136 25662
rect 12670 25560 12676 25612
rect 12728 25600 12734 25612
rect 13041 25603 13099 25609
rect 13041 25600 13053 25603
rect 12728 25572 13053 25600
rect 12728 25560 12734 25572
rect 13041 25569 13053 25572
rect 13087 25569 13099 25603
rect 15706 25600 15712 25612
rect 15667 25572 15712 25600
rect 13041 25563 13099 25569
rect 15706 25560 15712 25572
rect 15764 25560 15770 25612
rect 17178 25560 17184 25612
rect 17236 25600 17242 25612
rect 18834 25600 18840 25612
rect 17236 25572 17408 25600
rect 18795 25572 18840 25600
rect 17236 25560 17242 25572
rect 12762 25532 12768 25544
rect 12675 25504 12768 25532
rect 12762 25492 12768 25504
rect 12820 25532 12826 25544
rect 13961 25535 14019 25541
rect 13961 25532 13973 25535
rect 12820 25504 13973 25532
rect 12820 25492 12826 25504
rect 13961 25501 13973 25504
rect 14007 25501 14019 25535
rect 13961 25495 14019 25501
rect 14602 25492 14608 25544
rect 14660 25532 14666 25544
rect 14660 25504 15660 25532
rect 14660 25492 14666 25504
rect 11934 25464 11940 25476
rect 11895 25436 11940 25464
rect 11934 25424 11940 25436
rect 11992 25424 11998 25476
rect 12949 25467 13007 25473
rect 12949 25433 12961 25467
rect 12995 25464 13007 25467
rect 13498 25464 13504 25476
rect 12995 25436 13504 25464
rect 12995 25433 13007 25436
rect 12949 25427 13007 25433
rect 13498 25424 13504 25436
rect 13556 25424 13562 25476
rect 14786 25464 14792 25476
rect 14747 25436 14792 25464
rect 14786 25424 14792 25436
rect 14844 25424 14850 25476
rect 14878 25424 14884 25476
rect 14936 25464 14942 25476
rect 15632 25473 15660 25504
rect 16994 25492 17000 25544
rect 17052 25532 17058 25544
rect 17380 25541 17408 25572
rect 18834 25560 18840 25572
rect 18892 25560 18898 25612
rect 19754 25560 19760 25612
rect 19812 25600 19818 25612
rect 19849 25603 19907 25609
rect 19849 25600 19861 25603
rect 19812 25572 19861 25600
rect 19812 25560 19818 25572
rect 19849 25569 19861 25572
rect 19895 25569 19907 25603
rect 21502 25600 21508 25612
rect 19849 25563 19907 25569
rect 19956 25572 21508 25600
rect 17365 25535 17423 25541
rect 17052 25504 17316 25532
rect 17052 25492 17058 25504
rect 17288 25473 17316 25504
rect 17365 25501 17377 25535
rect 17411 25501 17423 25535
rect 17365 25495 17423 25501
rect 18193 25535 18251 25541
rect 18193 25501 18205 25535
rect 18239 25532 18251 25535
rect 19956 25532 19984 25572
rect 21502 25560 21508 25572
rect 21560 25560 21566 25612
rect 24449 25603 24507 25609
rect 24449 25569 24461 25603
rect 24495 25600 24507 25603
rect 25274 25600 25280 25612
rect 24495 25572 25280 25600
rect 24495 25569 24507 25572
rect 24449 25563 24507 25569
rect 25274 25560 25280 25572
rect 25332 25560 25338 25612
rect 25458 25560 25464 25612
rect 25516 25600 25522 25612
rect 25829 25603 25887 25609
rect 25829 25600 25841 25603
rect 25516 25572 25841 25600
rect 25516 25560 25522 25572
rect 25829 25569 25841 25572
rect 25875 25569 25887 25603
rect 25829 25563 25887 25569
rect 26841 25603 26899 25609
rect 26841 25569 26853 25603
rect 26887 25600 26899 25603
rect 27942 25600 27948 25612
rect 26887 25572 27948 25600
rect 26887 25569 26899 25572
rect 26841 25563 26899 25569
rect 27942 25560 27948 25572
rect 28000 25560 28006 25612
rect 18239 25504 19984 25532
rect 20033 25535 20091 25541
rect 18239 25501 18251 25504
rect 18193 25495 18251 25501
rect 20033 25501 20045 25535
rect 20079 25532 20091 25535
rect 20214 25532 20220 25544
rect 20079 25504 20220 25532
rect 20079 25501 20091 25504
rect 20033 25495 20091 25501
rect 20214 25492 20220 25504
rect 20272 25492 20278 25544
rect 21244 25504 21548 25532
rect 18374 25473 18380 25476
rect 15433 25467 15491 25473
rect 15433 25464 15445 25467
rect 14936 25436 15445 25464
rect 14936 25424 14942 25436
rect 15433 25433 15445 25436
rect 15479 25433 15491 25467
rect 15433 25427 15491 25433
rect 15617 25467 15675 25473
rect 15617 25433 15629 25467
rect 15663 25433 15675 25467
rect 15617 25427 15675 25433
rect 17181 25467 17239 25473
rect 17181 25433 17193 25467
rect 17227 25433 17239 25467
rect 17181 25427 17239 25433
rect 17273 25467 17331 25473
rect 17273 25433 17285 25467
rect 17319 25464 17331 25467
rect 18340 25467 18380 25473
rect 17319 25436 17684 25464
rect 17319 25433 17331 25436
rect 17273 25427 17331 25433
rect 14510 25396 14516 25408
rect 14471 25368 14516 25396
rect 14510 25356 14516 25368
rect 14568 25356 14574 25408
rect 14970 25396 14976 25408
rect 14931 25368 14976 25396
rect 14970 25356 14976 25368
rect 15028 25356 15034 25408
rect 16258 25356 16264 25408
rect 16316 25396 16322 25408
rect 16718 25396 16724 25408
rect 16316 25368 16724 25396
rect 16316 25356 16322 25368
rect 16718 25356 16724 25368
rect 16776 25396 16782 25408
rect 16997 25399 17055 25405
rect 16997 25396 17009 25399
rect 16776 25368 17009 25396
rect 16776 25356 16782 25368
rect 16997 25365 17009 25368
rect 17043 25365 17055 25399
rect 17196 25396 17224 25427
rect 17546 25396 17552 25408
rect 17196 25368 17552 25396
rect 16997 25359 17055 25365
rect 17546 25356 17552 25368
rect 17604 25356 17610 25408
rect 12118 25260 12124 25272
rect 12079 25232 12124 25260
rect 12118 25220 12124 25232
rect 12176 25220 12182 25272
rect 17656 25260 17684 25436
rect 18340 25433 18352 25467
rect 18340 25427 18380 25433
rect 18374 25424 18380 25427
rect 18432 25424 18438 25476
rect 18466 25424 18472 25476
rect 18524 25464 18530 25476
rect 18524 25436 19800 25464
rect 18524 25424 18530 25436
rect 17733 25399 17791 25405
rect 17733 25365 17745 25399
rect 17779 25396 17791 25399
rect 17779 25368 18512 25396
rect 17779 25365 17791 25368
rect 17733 25359 17791 25365
rect 18484 25337 18512 25368
rect 18558 25356 18564 25408
rect 18616 25396 18622 25408
rect 18616 25368 18661 25396
rect 18616 25356 18622 25368
rect 19478 25356 19484 25408
rect 19536 25396 19542 25408
rect 19665 25399 19723 25405
rect 19665 25396 19677 25399
rect 19536 25368 19677 25396
rect 19536 25356 19542 25368
rect 19665 25365 19677 25368
rect 19711 25365 19723 25399
rect 19772 25396 19800 25436
rect 19846 25424 19852 25476
rect 19904 25464 19910 25476
rect 19941 25467 19999 25473
rect 19941 25464 19953 25467
rect 19904 25436 19953 25464
rect 19904 25424 19910 25436
rect 19941 25433 19953 25436
rect 19987 25433 19999 25467
rect 21244 25464 21272 25504
rect 21520 25473 21548 25504
rect 21594 25492 21600 25544
rect 21652 25532 21658 25544
rect 21652 25504 22560 25532
rect 21652 25492 21658 25504
rect 22532 25473 22560 25504
rect 23158 25492 23164 25544
rect 23216 25532 23222 25544
rect 23216 25504 25375 25532
rect 23216 25492 23222 25504
rect 19941 25427 19999 25433
rect 20048 25436 21272 25464
rect 21321 25467 21379 25473
rect 20048 25396 20076 25436
rect 21321 25433 21333 25467
rect 21367 25433 21379 25467
rect 21321 25427 21379 25433
rect 21505 25467 21563 25473
rect 21505 25433 21517 25467
rect 21551 25464 21563 25467
rect 22333 25467 22391 25473
rect 22333 25464 22345 25467
rect 21551 25436 22345 25464
rect 21551 25433 21563 25436
rect 21505 25427 21563 25433
rect 22333 25433 22345 25436
rect 22379 25433 22391 25467
rect 22333 25427 22391 25433
rect 22517 25467 22575 25473
rect 22517 25433 22529 25467
rect 22563 25433 22575 25467
rect 23805 25467 23863 25473
rect 23805 25464 23817 25467
rect 22517 25427 22575 25433
rect 22624 25436 23817 25464
rect 20398 25396 20404 25408
rect 19772 25368 20076 25396
rect 20359 25368 20404 25396
rect 19665 25359 19723 25365
rect 20398 25356 20404 25368
rect 20456 25356 20462 25408
rect 21042 25356 21048 25408
rect 21100 25396 21106 25408
rect 21336 25396 21364 25427
rect 21870 25396 21876 25408
rect 21100 25368 21364 25396
rect 21831 25368 21876 25396
rect 21100 25356 21106 25368
rect 21870 25356 21876 25368
rect 21928 25356 21934 25408
rect 22422 25356 22428 25408
rect 22480 25396 22486 25408
rect 22624 25396 22652 25436
rect 23805 25433 23817 25436
rect 23851 25433 23863 25467
rect 23805 25427 23863 25433
rect 23894 25424 23900 25476
rect 23952 25464 23958 25476
rect 24814 25464 24820 25476
rect 23952 25436 24820 25464
rect 23952 25424 23958 25436
rect 24814 25424 24820 25436
rect 24872 25464 24878 25476
rect 25347 25473 25375 25504
rect 25734 25492 25740 25544
rect 25792 25532 25798 25544
rect 26930 25532 26936 25544
rect 25792 25504 26936 25532
rect 25792 25492 25798 25504
rect 26930 25492 26936 25504
rect 26988 25532 26994 25544
rect 26988 25504 27712 25532
rect 26988 25492 26994 25504
rect 25185 25467 25243 25473
rect 25185 25464 25197 25467
rect 24872 25436 25197 25464
rect 24872 25424 24878 25436
rect 25185 25433 25197 25436
rect 25231 25433 25243 25467
rect 25185 25427 25243 25433
rect 25332 25467 25390 25473
rect 25332 25433 25344 25467
rect 25378 25433 25390 25467
rect 25332 25427 25390 25433
rect 25458 25424 25464 25476
rect 25516 25464 25522 25476
rect 27209 25467 27267 25473
rect 27209 25464 27221 25467
rect 25516 25436 27221 25464
rect 25516 25424 25522 25436
rect 27209 25433 27221 25436
rect 27255 25433 27267 25467
rect 27574 25464 27580 25476
rect 27535 25436 27580 25464
rect 27209 25427 27267 25433
rect 27574 25424 27580 25436
rect 27632 25424 27638 25476
rect 27684 25473 27712 25504
rect 28678 25492 28684 25544
rect 28736 25532 28742 25544
rect 28957 25535 29015 25541
rect 28957 25532 28969 25535
rect 28736 25504 28969 25532
rect 28736 25492 28742 25504
rect 28957 25501 28969 25504
rect 29003 25501 29015 25535
rect 28957 25495 29015 25501
rect 29233 25535 29291 25541
rect 29233 25501 29245 25535
rect 29279 25532 29291 25535
rect 29506 25532 29512 25544
rect 29279 25504 29512 25532
rect 29279 25501 29291 25504
rect 29233 25495 29291 25501
rect 29506 25492 29512 25504
rect 29564 25492 29570 25544
rect 27669 25467 27727 25473
rect 27669 25433 27681 25467
rect 27715 25433 27727 25467
rect 27669 25427 27727 25433
rect 28034 25424 28040 25476
rect 28092 25464 28098 25476
rect 28313 25467 28371 25473
rect 28313 25464 28325 25467
rect 28092 25436 28325 25464
rect 28092 25424 28098 25436
rect 28313 25433 28325 25436
rect 28359 25433 28371 25467
rect 28313 25427 28371 25433
rect 22480 25368 22652 25396
rect 22885 25399 22943 25405
rect 22480 25356 22486 25368
rect 22885 25365 22897 25399
rect 22931 25396 22943 25399
rect 23526 25396 23532 25408
rect 22931 25368 23532 25396
rect 22931 25365 22943 25368
rect 22885 25359 22943 25365
rect 23526 25356 23532 25368
rect 23584 25356 23590 25408
rect 24170 25396 24176 25408
rect 24083 25368 24176 25396
rect 24170 25356 24176 25368
rect 24228 25396 24234 25408
rect 24998 25396 25004 25408
rect 24228 25368 25004 25396
rect 24228 25356 24234 25368
rect 24998 25356 25004 25368
rect 25056 25396 25062 25408
rect 25553 25399 25611 25405
rect 25553 25396 25565 25399
rect 25056 25368 25565 25396
rect 25056 25356 25062 25368
rect 25553 25365 25565 25368
rect 25599 25365 25611 25399
rect 27022 25396 27028 25408
rect 26983 25368 27028 25396
rect 25553 25359 25611 25365
rect 27022 25356 27028 25368
rect 27080 25356 27086 25408
rect 18469 25331 18527 25337
rect 18469 25297 18481 25331
rect 18515 25297 18527 25331
rect 18469 25291 18527 25297
rect 18834 25288 18840 25340
rect 18892 25328 18898 25340
rect 25918 25328 25924 25340
rect 18892 25300 25924 25328
rect 18892 25288 18898 25300
rect 25918 25288 25924 25300
rect 25976 25288 25982 25340
rect 18852 25260 18880 25288
rect 17656 25232 18880 25260
rect 23802 25220 23808 25272
rect 23860 25260 23866 25272
rect 23943 25263 24001 25269
rect 23943 25260 23955 25263
rect 23860 25232 23955 25260
rect 23860 25220 23866 25232
rect 23943 25229 23955 25232
rect 23989 25229 24001 25263
rect 23943 25223 24001 25229
rect 24081 25263 24139 25269
rect 24081 25229 24093 25263
rect 24127 25260 24139 25263
rect 24630 25260 24636 25272
rect 24127 25232 24636 25260
rect 24127 25229 24139 25232
rect 24081 25223 24139 25229
rect 24630 25220 24636 25232
rect 24688 25260 24694 25272
rect 25461 25263 25519 25269
rect 25461 25260 25473 25263
rect 24688 25232 25473 25260
rect 24688 25220 24694 25232
rect 25461 25229 25473 25232
rect 25507 25229 25519 25263
rect 25461 25223 25519 25229
rect 11000 25170 30136 25192
rect 11000 25118 14142 25170
rect 14194 25118 14206 25170
rect 14258 25118 14270 25170
rect 14322 25118 14334 25170
rect 14386 25118 24142 25170
rect 24194 25118 24206 25170
rect 24258 25118 24270 25170
rect 24322 25118 24334 25170
rect 24386 25118 30136 25170
rect 11000 25096 30136 25118
rect 18558 25016 18564 25068
rect 18616 25056 18622 25068
rect 21229 25059 21287 25065
rect 18616 25028 20996 25056
rect 18616 25016 18622 25028
rect 14510 24988 14516 25000
rect 14344 24960 14516 24988
rect 14344 24929 14372 24960
rect 14510 24948 14516 24960
rect 14568 24948 14574 25000
rect 16997 24991 17055 24997
rect 16997 24957 17009 24991
rect 17043 24988 17055 24991
rect 17546 24988 17552 25000
rect 17043 24960 17552 24988
rect 17043 24957 17055 24960
rect 16997 24951 17055 24957
rect 17546 24948 17552 24960
rect 17604 24948 17610 25000
rect 20398 24948 20404 25000
rect 20456 24988 20462 25000
rect 20861 24991 20919 24997
rect 20861 24988 20873 24991
rect 20456 24960 20873 24988
rect 20456 24948 20462 24960
rect 20861 24957 20873 24960
rect 20907 24957 20919 24991
rect 20861 24951 20919 24957
rect 14329 24923 14387 24929
rect 14329 24889 14341 24923
rect 14375 24889 14387 24923
rect 14878 24920 14884 24932
rect 14329 24883 14387 24889
rect 14436 24892 14884 24920
rect 11290 24852 11296 24864
rect 11251 24824 11296 24852
rect 11290 24812 11296 24824
rect 11348 24812 11354 24864
rect 14237 24855 14295 24861
rect 14237 24821 14249 24855
rect 14283 24852 14295 24855
rect 14436 24852 14464 24892
rect 14878 24880 14884 24892
rect 14936 24880 14942 24932
rect 16718 24880 16724 24932
rect 16776 24920 16782 24932
rect 16868 24923 16926 24929
rect 16868 24920 16880 24923
rect 16776 24892 16880 24920
rect 16776 24880 16782 24892
rect 16868 24889 16880 24892
rect 16914 24889 16926 24923
rect 16868 24883 16926 24889
rect 17089 24923 17147 24929
rect 17089 24889 17101 24923
rect 17135 24920 17147 24923
rect 18193 24923 18251 24929
rect 18193 24920 18205 24923
rect 17135 24892 18205 24920
rect 17135 24889 17147 24892
rect 17089 24883 17147 24889
rect 18193 24889 18205 24892
rect 18239 24920 18251 24923
rect 18282 24920 18288 24932
rect 18239 24892 18288 24920
rect 18239 24889 18251 24892
rect 18193 24883 18251 24889
rect 18282 24880 18288 24892
rect 18340 24880 18346 24932
rect 18926 24920 18932 24932
rect 18887 24892 18932 24920
rect 18926 24880 18932 24892
rect 18984 24880 18990 24932
rect 19389 24923 19447 24929
rect 19389 24889 19401 24923
rect 19435 24920 19447 24923
rect 19478 24920 19484 24932
rect 19435 24892 19484 24920
rect 19435 24889 19447 24892
rect 19389 24883 19447 24889
rect 19478 24880 19484 24892
rect 19536 24880 19542 24932
rect 14283 24824 14464 24852
rect 14283 24821 14295 24824
rect 14237 24815 14295 24821
rect 14510 24812 14516 24864
rect 14568 24852 14574 24864
rect 15798 24852 15804 24864
rect 14568 24824 14613 24852
rect 15759 24824 15804 24852
rect 14568 24812 14574 24824
rect 15798 24812 15804 24824
rect 15856 24812 15862 24864
rect 20125 24855 20183 24861
rect 20125 24821 20137 24855
rect 20171 24852 20183 24855
rect 20732 24855 20790 24861
rect 20732 24852 20744 24855
rect 20171 24824 20744 24852
rect 20171 24821 20183 24824
rect 20125 24815 20183 24821
rect 20732 24821 20744 24824
rect 20778 24821 20790 24855
rect 20876 24852 20904 24951
rect 20968 24929 20996 25028
rect 21229 25025 21241 25059
rect 21275 25056 21287 25059
rect 22330 25056 22336 25068
rect 21275 25028 22336 25056
rect 21275 25025 21287 25028
rect 21229 25019 21287 25025
rect 22330 25016 22336 25028
rect 22388 25016 22394 25068
rect 22609 25059 22667 25065
rect 22609 25056 22621 25059
rect 22440 25028 22621 25056
rect 21042 24948 21048 25000
rect 21100 24988 21106 25000
rect 22440 24988 22468 25028
rect 22609 25025 22621 25028
rect 22655 25025 22667 25059
rect 22609 25019 22667 25025
rect 23434 25016 23440 25068
rect 23492 25056 23498 25068
rect 23989 25059 24047 25065
rect 23989 25056 24001 25059
rect 23492 25028 24001 25056
rect 23492 25016 23498 25028
rect 23989 25025 24001 25028
rect 24035 25025 24047 25059
rect 23989 25019 24047 25025
rect 24357 25059 24415 25065
rect 24357 25025 24369 25059
rect 24403 25056 24415 25059
rect 25458 25056 25464 25068
rect 24403 25028 25464 25056
rect 24403 25025 24415 25028
rect 24357 25019 24415 25025
rect 25458 25016 25464 25028
rect 25516 25016 25522 25068
rect 28034 25056 28040 25068
rect 27995 25028 28040 25056
rect 28034 25016 28040 25028
rect 28092 25016 28098 25068
rect 21100 24960 22468 24988
rect 22498 24991 22556 24997
rect 21100 24948 21106 24960
rect 22498 24957 22510 24991
rect 22544 24988 22556 24991
rect 22544 24960 23296 24988
rect 22544 24957 22556 24960
rect 22498 24951 22556 24957
rect 20953 24923 21011 24929
rect 20953 24889 20965 24923
rect 20999 24889 21011 24923
rect 22513 24920 22541 24951
rect 20953 24883 21011 24889
rect 22256 24892 22541 24920
rect 22701 24923 22759 24929
rect 22256 24852 22284 24892
rect 22701 24889 22713 24923
rect 22747 24889 22759 24923
rect 22701 24883 22759 24889
rect 23069 24923 23127 24929
rect 23069 24889 23081 24923
rect 23115 24920 23127 24923
rect 23158 24920 23164 24932
rect 23115 24892 23164 24920
rect 23115 24889 23127 24892
rect 23069 24883 23127 24889
rect 20876 24824 22284 24852
rect 22333 24855 22391 24861
rect 20732 24815 20790 24821
rect 22333 24821 22345 24855
rect 22379 24852 22391 24855
rect 22422 24852 22428 24864
rect 22379 24824 22428 24852
rect 22379 24821 22391 24824
rect 22333 24815 22391 24821
rect 22422 24812 22428 24824
rect 22480 24812 22486 24864
rect 22716 24852 22744 24883
rect 23158 24880 23164 24892
rect 23216 24880 23222 24932
rect 23268 24920 23296 24960
rect 23526 24948 23532 25000
rect 23584 24988 23590 25000
rect 23584 24960 25136 24988
rect 23584 24948 23590 24960
rect 24081 24923 24139 24929
rect 23268 24892 23986 24920
rect 23434 24852 23440 24864
rect 22716 24824 23440 24852
rect 23434 24812 23440 24824
rect 23492 24812 23498 24864
rect 23802 24812 23808 24864
rect 23860 24861 23866 24864
rect 23860 24855 23918 24861
rect 23860 24821 23872 24855
rect 23906 24821 23918 24855
rect 23958 24852 23986 24892
rect 24081 24889 24093 24923
rect 24127 24920 24139 24923
rect 24998 24920 25004 24932
rect 24127 24892 25004 24920
rect 24127 24889 24139 24892
rect 24081 24883 24139 24889
rect 24998 24880 25004 24892
rect 25056 24880 25062 24932
rect 24538 24852 24544 24864
rect 23958 24824 24544 24852
rect 23860 24815 23918 24821
rect 23860 24812 23866 24815
rect 24538 24812 24544 24824
rect 24596 24812 24602 24864
rect 25108 24861 25136 24960
rect 25550 24948 25556 25000
rect 25608 24988 25614 25000
rect 28310 24988 28316 25000
rect 25608 24960 28316 24988
rect 25608 24948 25614 24960
rect 28310 24948 28316 24960
rect 28368 24948 28374 25000
rect 25918 24920 25924 24932
rect 25879 24892 25924 24920
rect 25918 24880 25924 24892
rect 25976 24880 25982 24932
rect 26746 24880 26752 24932
rect 26804 24920 26810 24932
rect 28954 24920 28960 24932
rect 26804 24892 28960 24920
rect 26804 24880 26810 24892
rect 28954 24880 28960 24892
rect 29012 24920 29018 24932
rect 29049 24923 29107 24929
rect 29049 24920 29061 24923
rect 29012 24892 29061 24920
rect 29012 24880 29018 24892
rect 29049 24889 29061 24892
rect 29095 24889 29107 24923
rect 29049 24883 29107 24889
rect 25093 24855 25151 24861
rect 25093 24821 25105 24855
rect 25139 24821 25151 24855
rect 26010 24852 26016 24864
rect 25971 24824 26016 24852
rect 25093 24815 25151 24821
rect 26010 24812 26016 24824
rect 26068 24812 26074 24864
rect 27942 24852 27948 24864
rect 27903 24824 27948 24852
rect 27942 24812 27948 24824
rect 28000 24812 28006 24864
rect 28586 24852 28592 24864
rect 28547 24824 28592 24852
rect 28586 24812 28592 24824
rect 28644 24812 28650 24864
rect 11566 24784 11572 24796
rect 11527 24756 11572 24784
rect 11566 24744 11572 24756
rect 11624 24744 11630 24796
rect 12118 24744 12124 24796
rect 12176 24744 12182 24796
rect 13317 24787 13375 24793
rect 13317 24753 13329 24787
rect 13363 24784 13375 24787
rect 13406 24784 13412 24796
rect 13363 24756 13412 24784
rect 13363 24753 13375 24756
rect 13317 24747 13375 24753
rect 13406 24744 13412 24756
rect 13464 24744 13470 24796
rect 15614 24784 15620 24796
rect 15575 24756 15620 24784
rect 15614 24744 15620 24756
rect 15672 24744 15678 24796
rect 16169 24787 16227 24793
rect 16169 24753 16181 24787
rect 16215 24753 16227 24787
rect 16169 24747 16227 24753
rect 16721 24787 16779 24793
rect 16721 24753 16733 24787
rect 16767 24784 16779 24787
rect 16810 24784 16816 24796
rect 16767 24756 16816 24784
rect 16767 24753 16779 24756
rect 16721 24747 16779 24753
rect 16184 24716 16212 24747
rect 16810 24744 16816 24756
rect 16868 24744 16874 24796
rect 17178 24744 17184 24796
rect 17236 24784 17242 24796
rect 18098 24784 18104 24796
rect 17236 24756 18104 24784
rect 17236 24744 17242 24756
rect 18098 24744 18104 24756
rect 18156 24784 18162 24796
rect 18469 24787 18527 24793
rect 18469 24784 18481 24787
rect 18156 24756 18481 24784
rect 18156 24744 18162 24756
rect 18469 24753 18481 24756
rect 18515 24753 18527 24787
rect 18469 24747 18527 24753
rect 18561 24787 18619 24793
rect 18561 24753 18573 24787
rect 18607 24784 18619 24787
rect 18834 24784 18840 24796
rect 18607 24756 18840 24784
rect 18607 24753 18619 24756
rect 18561 24747 18619 24753
rect 18834 24744 18840 24756
rect 18892 24744 18898 24796
rect 19754 24784 19760 24796
rect 19715 24756 19760 24784
rect 19754 24744 19760 24756
rect 19812 24744 19818 24796
rect 20582 24784 20588 24796
rect 20543 24756 20588 24784
rect 20582 24744 20588 24756
rect 20640 24744 20646 24796
rect 23342 24744 23348 24796
rect 23400 24784 23406 24796
rect 23713 24787 23771 24793
rect 23713 24784 23725 24787
rect 23400 24756 23725 24784
rect 23400 24744 23406 24756
rect 23713 24753 23725 24756
rect 23759 24784 23771 24787
rect 24909 24787 24967 24793
rect 24909 24784 24921 24787
rect 23759 24756 24921 24784
rect 23759 24753 23771 24756
rect 23713 24747 23771 24753
rect 24909 24753 24921 24756
rect 24955 24753 24967 24787
rect 24909 24747 24967 24753
rect 25366 24744 25372 24796
rect 25424 24784 25430 24796
rect 25461 24787 25519 24793
rect 25461 24784 25473 24787
rect 25424 24756 25473 24784
rect 25424 24744 25430 24756
rect 25461 24753 25473 24756
rect 25507 24753 25519 24787
rect 25461 24747 25519 24753
rect 26473 24787 26531 24793
rect 26473 24753 26485 24787
rect 26519 24784 26531 24787
rect 28126 24784 28132 24796
rect 26519 24756 28132 24784
rect 26519 24753 26531 24756
rect 26473 24747 26531 24753
rect 28126 24744 28132 24756
rect 28184 24744 28190 24796
rect 29141 24787 29199 24793
rect 29141 24753 29153 24787
rect 29187 24753 29199 24787
rect 29141 24747 29199 24753
rect 16994 24716 17000 24728
rect 16184 24688 17000 24716
rect 16994 24676 17000 24688
rect 17052 24676 17058 24728
rect 17362 24716 17368 24728
rect 17323 24688 17368 24716
rect 17362 24676 17368 24688
rect 17420 24676 17426 24728
rect 17546 24676 17552 24728
rect 17604 24716 17610 24728
rect 18377 24719 18435 24725
rect 18377 24716 18389 24719
rect 17604 24688 18389 24716
rect 17604 24676 17610 24688
rect 18377 24685 18389 24688
rect 18423 24716 18435 24719
rect 19573 24719 19631 24725
rect 19573 24716 19585 24719
rect 18423 24688 19585 24716
rect 18423 24685 18435 24688
rect 18377 24679 18435 24685
rect 19573 24685 19585 24688
rect 19619 24685 19631 24719
rect 19573 24679 19631 24685
rect 19662 24676 19668 24728
rect 19720 24716 19726 24728
rect 19846 24716 19852 24728
rect 19720 24688 19852 24716
rect 19720 24676 19726 24688
rect 19846 24676 19852 24688
rect 19904 24676 19910 24728
rect 26562 24676 26568 24728
rect 26620 24716 26626 24728
rect 26933 24719 26991 24725
rect 26933 24716 26945 24719
rect 26620 24688 26945 24716
rect 26620 24676 26626 24688
rect 26933 24685 26945 24688
rect 26979 24685 26991 24719
rect 26933 24679 26991 24685
rect 27022 24676 27028 24728
rect 27080 24716 27086 24728
rect 27080 24688 27125 24716
rect 27080 24676 27086 24688
rect 27206 24676 27212 24728
rect 27264 24716 27270 24728
rect 29156 24716 29184 24747
rect 27264 24688 29184 24716
rect 27264 24676 27270 24688
rect 11000 24626 30136 24648
rect 11000 24574 19142 24626
rect 19194 24574 19206 24626
rect 19258 24574 19270 24626
rect 19322 24574 19334 24626
rect 19386 24574 29142 24626
rect 29194 24574 29206 24626
rect 29258 24574 29270 24626
rect 29322 24574 29334 24626
rect 29386 24574 30136 24626
rect 11000 24552 30136 24574
rect 15982 24512 15988 24524
rect 13976 24484 15988 24512
rect 12029 24379 12087 24385
rect 12029 24345 12041 24379
rect 12075 24376 12087 24379
rect 12118 24376 12124 24388
rect 12075 24348 12124 24376
rect 12075 24345 12087 24348
rect 12029 24339 12087 24345
rect 12118 24336 12124 24348
rect 12176 24336 12182 24388
rect 12213 24379 12271 24385
rect 12213 24345 12225 24379
rect 12259 24376 12271 24379
rect 12394 24376 12400 24388
rect 12259 24348 12400 24376
rect 12259 24345 12271 24348
rect 12213 24339 12271 24345
rect 12394 24336 12400 24348
rect 12452 24336 12458 24388
rect 13406 24336 13412 24388
rect 13464 24376 13470 24388
rect 13976 24385 14004 24484
rect 15982 24472 15988 24484
rect 16040 24512 16046 24524
rect 16718 24512 16724 24524
rect 16040 24484 16724 24512
rect 16040 24472 16046 24484
rect 16718 24472 16724 24484
rect 16776 24512 16782 24524
rect 18006 24512 18012 24524
rect 16776 24484 18012 24512
rect 16776 24472 16782 24484
rect 18006 24472 18012 24484
rect 18064 24512 18070 24524
rect 19662 24512 19668 24524
rect 18064 24484 19668 24512
rect 18064 24472 18070 24484
rect 19662 24472 19668 24484
rect 19720 24472 19726 24524
rect 21502 24512 21508 24524
rect 21463 24484 21508 24512
rect 21502 24472 21508 24484
rect 21560 24472 21566 24524
rect 25185 24515 25243 24521
rect 25185 24481 25197 24515
rect 25231 24512 25243 24515
rect 27206 24512 27212 24524
rect 25231 24484 27212 24512
rect 25231 24481 25243 24484
rect 25185 24475 25243 24481
rect 27206 24472 27212 24484
rect 27264 24472 27270 24524
rect 27758 24512 27764 24524
rect 27719 24484 27764 24512
rect 27758 24472 27764 24484
rect 27816 24472 27822 24524
rect 29506 24512 29512 24524
rect 29432 24484 29512 24512
rect 15249 24447 15307 24453
rect 15249 24413 15261 24447
rect 15295 24444 15307 24447
rect 17089 24447 17147 24453
rect 15295 24416 17040 24444
rect 15295 24413 15307 24416
rect 15249 24407 15307 24413
rect 13961 24379 14019 24385
rect 13961 24376 13973 24379
rect 13464 24348 13973 24376
rect 13464 24336 13470 24348
rect 13961 24345 13973 24348
rect 14007 24345 14019 24379
rect 13961 24339 14019 24345
rect 15157 24379 15215 24385
rect 15157 24345 15169 24379
rect 15203 24345 15215 24379
rect 15157 24339 15215 24345
rect 15801 24379 15859 24385
rect 15801 24345 15813 24379
rect 15847 24376 15859 24379
rect 16810 24376 16816 24388
rect 15847 24348 16816 24376
rect 15847 24345 15859 24348
rect 15801 24339 15859 24345
rect 15172 24240 15200 24339
rect 16810 24336 16816 24348
rect 16868 24336 16874 24388
rect 15982 24317 15988 24320
rect 15948 24311 15988 24317
rect 15948 24277 15960 24311
rect 15948 24271 15988 24277
rect 15982 24268 15988 24271
rect 16040 24268 16046 24320
rect 16166 24308 16172 24320
rect 16127 24280 16172 24308
rect 16166 24268 16172 24280
rect 16224 24268 16230 24320
rect 16261 24243 16319 24249
rect 16261 24240 16273 24243
rect 15172 24212 16273 24240
rect 16261 24209 16273 24212
rect 16307 24209 16319 24243
rect 17012 24240 17040 24416
rect 17089 24413 17101 24447
rect 17135 24444 17147 24447
rect 18190 24444 18196 24456
rect 17135 24416 18196 24444
rect 17135 24413 17147 24416
rect 17089 24407 17147 24413
rect 18190 24404 18196 24416
rect 18248 24404 18254 24456
rect 18285 24447 18343 24453
rect 18285 24413 18297 24447
rect 18331 24444 18343 24447
rect 18374 24444 18380 24456
rect 18331 24416 18380 24444
rect 18331 24413 18343 24416
rect 18285 24407 18343 24413
rect 18374 24404 18380 24416
rect 18432 24404 18438 24456
rect 19021 24447 19079 24453
rect 19021 24413 19033 24447
rect 19067 24444 19079 24447
rect 20769 24447 20827 24453
rect 19067 24416 20536 24444
rect 19067 24413 19079 24416
rect 19021 24407 19079 24413
rect 17270 24376 17276 24388
rect 17231 24348 17276 24376
rect 17270 24336 17276 24348
rect 17328 24336 17334 24388
rect 18624 24379 18682 24385
rect 18624 24345 18636 24379
rect 18670 24376 18682 24379
rect 19573 24379 19631 24385
rect 18670 24348 19524 24376
rect 18670 24345 18682 24348
rect 18624 24339 18682 24345
rect 17641 24311 17699 24317
rect 17641 24277 17653 24311
rect 17687 24308 17699 24311
rect 19496 24308 19524 24348
rect 19573 24345 19585 24379
rect 19619 24376 19631 24379
rect 19754 24376 19760 24388
rect 19619 24348 19760 24376
rect 19619 24345 19631 24348
rect 19573 24339 19631 24345
rect 19754 24336 19760 24348
rect 19812 24376 19818 24388
rect 20122 24376 20128 24388
rect 19812 24348 20128 24376
rect 19812 24336 19818 24348
rect 20122 24336 20128 24348
rect 20180 24336 20186 24388
rect 20217 24379 20275 24385
rect 20217 24345 20229 24379
rect 20263 24345 20275 24379
rect 20217 24339 20275 24345
rect 20401 24379 20459 24385
rect 20401 24345 20413 24379
rect 20447 24345 20459 24379
rect 20401 24339 20459 24345
rect 19662 24308 19668 24320
rect 17687 24280 19432 24308
rect 19496 24280 19668 24308
rect 17687 24277 17699 24280
rect 17641 24271 17699 24277
rect 18558 24240 18564 24252
rect 17012 24212 18564 24240
rect 16261 24203 16319 24209
rect 18558 24200 18564 24212
rect 18616 24200 18622 24252
rect 19404 24240 19432 24280
rect 19662 24268 19668 24280
rect 19720 24268 19726 24320
rect 20232 24240 20260 24339
rect 19404 24212 20260 24240
rect 20416 24240 20444 24339
rect 20508 24308 20536 24416
rect 20769 24413 20781 24447
rect 20815 24444 20827 24447
rect 23802 24444 23808 24456
rect 20815 24416 23808 24444
rect 20815 24413 20827 24416
rect 20769 24407 20827 24413
rect 20950 24336 20956 24388
rect 21008 24376 21014 24388
rect 21229 24379 21287 24385
rect 21229 24376 21241 24379
rect 21008 24348 21241 24376
rect 21008 24336 21014 24348
rect 21229 24345 21241 24348
rect 21275 24345 21287 24379
rect 21229 24339 21287 24345
rect 21413 24379 21471 24385
rect 21413 24345 21425 24379
rect 21459 24376 21471 24379
rect 22054 24376 22060 24388
rect 21459 24348 22060 24376
rect 21459 24345 21471 24348
rect 21413 24339 21471 24345
rect 22054 24336 22060 24348
rect 22112 24336 22118 24388
rect 23158 24376 23164 24388
rect 23119 24348 23164 24376
rect 23158 24336 23164 24348
rect 23216 24336 23222 24388
rect 23544 24317 23572 24416
rect 23802 24404 23808 24416
rect 23860 24404 23866 24456
rect 24449 24447 24507 24453
rect 24449 24413 24461 24447
rect 24495 24444 24507 24447
rect 26746 24444 26752 24456
rect 24495 24416 26752 24444
rect 24495 24413 24507 24416
rect 24449 24407 24507 24413
rect 26746 24404 26752 24416
rect 26804 24404 26810 24456
rect 29322 24444 29328 24456
rect 26948 24416 28264 24444
rect 26948 24388 26976 24416
rect 25369 24379 25427 24385
rect 25369 24345 25381 24379
rect 25415 24376 25427 24379
rect 25550 24376 25556 24388
rect 25415 24348 25556 24376
rect 25415 24345 25427 24348
rect 25369 24339 25427 24345
rect 25550 24336 25556 24348
rect 25608 24336 25614 24388
rect 26010 24336 26016 24388
rect 26068 24376 26074 24388
rect 26289 24379 26347 24385
rect 26289 24376 26301 24379
rect 26068 24348 26301 24376
rect 26068 24336 26074 24348
rect 26289 24345 26301 24348
rect 26335 24345 26347 24379
rect 26470 24376 26476 24388
rect 26431 24348 26476 24376
rect 26289 24339 26347 24345
rect 26470 24336 26476 24348
rect 26528 24336 26534 24388
rect 26838 24376 26844 24388
rect 26799 24348 26844 24376
rect 26838 24336 26844 24348
rect 26896 24336 26902 24388
rect 26930 24336 26936 24388
rect 26988 24376 26994 24388
rect 27945 24379 28003 24385
rect 27945 24376 27957 24379
rect 26988 24348 27033 24376
rect 27408 24348 27957 24376
rect 26988 24336 26994 24348
rect 23308 24311 23366 24317
rect 23308 24308 23320 24311
rect 20508 24280 23320 24308
rect 23308 24277 23320 24280
rect 23354 24277 23366 24311
rect 23308 24271 23366 24277
rect 23529 24311 23587 24317
rect 23529 24277 23541 24311
rect 23575 24277 23587 24311
rect 26488 24308 26516 24336
rect 27408 24308 27436 24348
rect 27945 24345 27957 24348
rect 27991 24345 28003 24379
rect 28126 24376 28132 24388
rect 28087 24348 28132 24376
rect 27945 24339 28003 24345
rect 28126 24336 28132 24348
rect 28184 24336 28190 24388
rect 26488 24280 27436 24308
rect 28236 24308 28264 24416
rect 28604 24416 29328 24444
rect 28494 24376 28500 24388
rect 28455 24348 28500 24376
rect 28494 24336 28500 24348
rect 28552 24336 28558 24388
rect 28405 24311 28463 24317
rect 28405 24308 28417 24311
rect 28236 24280 28417 24308
rect 23529 24271 23587 24277
rect 28405 24277 28417 24280
rect 28451 24277 28463 24311
rect 28405 24271 28463 24277
rect 23158 24240 23164 24252
rect 20416 24212 23164 24240
rect 12026 24132 12032 24184
rect 12084 24172 12090 24184
rect 12305 24175 12363 24181
rect 12305 24172 12317 24175
rect 12084 24144 12317 24172
rect 12084 24132 12090 24144
rect 12305 24141 12317 24144
rect 12351 24141 12363 24175
rect 12305 24135 12363 24141
rect 12946 24132 12952 24184
rect 13004 24172 13010 24184
rect 14053 24175 14111 24181
rect 14053 24172 14065 24175
rect 13004 24144 14065 24172
rect 13004 24132 13010 24144
rect 14053 24141 14065 24144
rect 14099 24172 14111 24175
rect 15982 24172 15988 24184
rect 14099 24144 15988 24172
rect 14099 24141 14111 24144
rect 14053 24135 14111 24141
rect 15982 24132 15988 24144
rect 16040 24132 16046 24184
rect 16077 24175 16135 24181
rect 16077 24141 16089 24175
rect 16123 24172 16135 24175
rect 16166 24172 16172 24184
rect 16123 24144 16172 24172
rect 16123 24141 16135 24144
rect 16077 24135 16135 24141
rect 16166 24132 16172 24144
rect 16224 24132 16230 24184
rect 18190 24132 18196 24184
rect 18248 24172 18254 24184
rect 18466 24181 18472 24184
rect 18423 24175 18472 24181
rect 18423 24172 18435 24175
rect 18248 24144 18435 24172
rect 18248 24132 18254 24144
rect 18423 24141 18435 24144
rect 18469 24141 18472 24175
rect 18423 24135 18472 24141
rect 18466 24132 18472 24135
rect 18524 24172 18530 24184
rect 18524 24144 18571 24172
rect 18524 24132 18530 24144
rect 18650 24132 18656 24184
rect 18708 24172 18714 24184
rect 19665 24175 19723 24181
rect 19665 24172 19677 24175
rect 18708 24144 19677 24172
rect 18708 24132 18714 24144
rect 19665 24141 19677 24144
rect 19711 24141 19723 24175
rect 20232 24172 20260 24212
rect 23158 24200 23164 24212
rect 23216 24240 23222 24252
rect 23618 24240 23624 24252
rect 23216 24212 23624 24240
rect 23216 24200 23222 24212
rect 23618 24200 23624 24212
rect 23676 24200 23682 24252
rect 24541 24243 24599 24249
rect 24541 24209 24553 24243
rect 24587 24240 24599 24243
rect 24587 24212 26240 24240
rect 24587 24209 24599 24212
rect 24541 24203 24599 24209
rect 21226 24172 21232 24184
rect 20232 24144 21232 24172
rect 19665 24135 19723 24141
rect 21226 24132 21232 24144
rect 21284 24132 21290 24184
rect 23434 24172 23440 24184
rect 23395 24144 23440 24172
rect 23434 24132 23440 24144
rect 23492 24132 23498 24184
rect 23802 24172 23808 24184
rect 23763 24144 23808 24172
rect 23802 24132 23808 24144
rect 23860 24132 23866 24184
rect 26102 24172 26108 24184
rect 26063 24144 26108 24172
rect 26102 24132 26108 24144
rect 26160 24132 26166 24184
rect 26212 24172 26240 24212
rect 26838 24200 26844 24252
rect 26896 24240 26902 24252
rect 28604 24240 28632 24416
rect 29322 24404 29328 24416
rect 29380 24404 29386 24456
rect 29432 24453 29460 24484
rect 29506 24472 29512 24484
rect 29564 24472 29570 24524
rect 29417 24447 29475 24453
rect 29417 24413 29429 24447
rect 29463 24413 29475 24447
rect 29417 24407 29475 24413
rect 29233 24379 29291 24385
rect 29233 24345 29245 24379
rect 29279 24376 29291 24379
rect 29506 24376 29512 24388
rect 29279 24348 29512 24376
rect 29279 24345 29291 24348
rect 29233 24339 29291 24345
rect 29506 24336 29512 24348
rect 29564 24336 29570 24388
rect 26896 24212 28632 24240
rect 26896 24200 26902 24212
rect 28494 24172 28500 24184
rect 26212 24144 28500 24172
rect 28494 24132 28500 24144
rect 28552 24132 28558 24184
rect 11000 24082 30136 24104
rect 11000 24030 14142 24082
rect 14194 24030 14206 24082
rect 14258 24030 14270 24082
rect 14322 24030 14334 24082
rect 14386 24030 24142 24082
rect 24194 24030 24206 24082
rect 24258 24030 24270 24082
rect 24322 24030 24334 24082
rect 24386 24030 30136 24082
rect 11000 24008 30136 24030
rect 14421 23971 14479 23977
rect 14421 23937 14433 23971
rect 14467 23968 14479 23971
rect 14878 23968 14884 23980
rect 14467 23940 14884 23968
rect 14467 23937 14479 23940
rect 14421 23931 14479 23937
rect 14878 23928 14884 23940
rect 14936 23928 14942 23980
rect 16077 23971 16135 23977
rect 16077 23937 16089 23971
rect 16123 23968 16135 23971
rect 21042 23968 21048 23980
rect 16123 23940 21048 23968
rect 16123 23937 16135 23940
rect 16077 23931 16135 23937
rect 21042 23928 21048 23940
rect 21100 23928 21106 23980
rect 21210 23971 21268 23977
rect 21210 23937 21222 23971
rect 21256 23968 21268 23971
rect 21502 23968 21508 23980
rect 21256 23940 21508 23968
rect 21256 23937 21268 23940
rect 21210 23931 21268 23937
rect 21502 23928 21508 23940
rect 21560 23928 21566 23980
rect 29233 23971 29291 23977
rect 29233 23937 29245 23971
rect 29279 23968 29291 23971
rect 29322 23968 29328 23980
rect 29279 23940 29328 23968
rect 29279 23937 29291 23940
rect 29233 23931 29291 23937
rect 29322 23928 29328 23940
rect 29380 23928 29386 23980
rect 14786 23860 14792 23912
rect 14844 23860 14850 23912
rect 15982 23860 15988 23912
rect 16040 23900 16046 23912
rect 17178 23900 17184 23912
rect 16040 23872 17184 23900
rect 16040 23860 16046 23872
rect 17178 23860 17184 23872
rect 17236 23909 17242 23912
rect 17236 23903 17285 23909
rect 17236 23869 17239 23903
rect 17273 23869 17285 23903
rect 17236 23863 17285 23869
rect 17365 23903 17423 23909
rect 17365 23869 17377 23903
rect 17411 23900 17423 23903
rect 17546 23900 17552 23912
rect 17411 23872 17552 23900
rect 17411 23869 17423 23872
rect 17365 23863 17423 23869
rect 17236 23860 17242 23863
rect 17546 23860 17552 23872
rect 17604 23860 17610 23912
rect 18742 23900 18748 23912
rect 18300 23872 18748 23900
rect 11566 23832 11572 23844
rect 11527 23804 11572 23832
rect 11566 23792 11572 23804
rect 11624 23792 11630 23844
rect 12857 23835 12915 23841
rect 12857 23801 12869 23835
rect 12903 23832 12915 23835
rect 13406 23832 13412 23844
rect 12903 23804 13412 23832
rect 12903 23801 12915 23804
rect 12857 23795 12915 23801
rect 13406 23792 13412 23804
rect 13464 23792 13470 23844
rect 14694 23832 14700 23844
rect 14655 23804 14700 23832
rect 14694 23792 14700 23804
rect 14752 23792 14758 23844
rect 14804 23832 14832 23860
rect 18300 23844 18328 23872
rect 18742 23860 18748 23872
rect 18800 23860 18806 23912
rect 21321 23903 21379 23909
rect 21321 23869 21333 23903
rect 21367 23900 21379 23903
rect 23618 23900 23624 23912
rect 21367 23872 23624 23900
rect 21367 23869 21379 23872
rect 21321 23863 21379 23869
rect 23618 23860 23624 23872
rect 23676 23860 23682 23912
rect 23710 23860 23716 23912
rect 23768 23900 23774 23912
rect 26010 23900 26016 23912
rect 23768 23872 24676 23900
rect 23768 23860 23774 23872
rect 14804 23804 15200 23832
rect 12026 23764 12032 23776
rect 11987 23736 12032 23764
rect 12026 23724 12032 23736
rect 12084 23724 12090 23776
rect 12210 23764 12216 23776
rect 12171 23736 12216 23764
rect 12210 23724 12216 23736
rect 12268 23724 12274 23776
rect 12397 23767 12455 23773
rect 12397 23733 12409 23767
rect 12443 23733 12455 23767
rect 13038 23764 13044 23776
rect 12999 23736 13044 23764
rect 12397 23727 12455 23733
rect 12412 23696 12440 23727
rect 13038 23724 13044 23736
rect 13096 23724 13102 23776
rect 13498 23764 13504 23776
rect 13411 23736 13504 23764
rect 13498 23724 13504 23736
rect 13556 23764 13562 23776
rect 13958 23764 13964 23776
rect 13556 23736 13964 23764
rect 13556 23724 13562 23736
rect 13958 23724 13964 23736
rect 14016 23724 14022 23776
rect 14789 23767 14847 23773
rect 14789 23733 14801 23767
rect 14835 23764 14847 23767
rect 15062 23764 15068 23776
rect 14835 23736 15068 23764
rect 14835 23733 14847 23736
rect 14789 23727 14847 23733
rect 15062 23724 15068 23736
rect 15120 23724 15126 23776
rect 15172 23773 15200 23804
rect 15246 23792 15252 23844
rect 15304 23832 15310 23844
rect 17457 23835 17515 23841
rect 17457 23832 17469 23835
rect 15304 23804 17469 23832
rect 15304 23792 15310 23804
rect 17457 23801 17469 23804
rect 17503 23832 17515 23835
rect 18282 23832 18288 23844
rect 17503 23804 18288 23832
rect 17503 23801 17515 23804
rect 17457 23795 17515 23801
rect 18282 23792 18288 23804
rect 18340 23792 18346 23844
rect 18377 23835 18435 23841
rect 18377 23801 18389 23835
rect 18423 23832 18435 23835
rect 18929 23835 18987 23841
rect 18423 23804 18880 23832
rect 18423 23801 18435 23804
rect 18377 23795 18435 23801
rect 15157 23767 15215 23773
rect 15157 23733 15169 23767
rect 15203 23733 15215 23767
rect 15157 23727 15215 23733
rect 15341 23767 15399 23773
rect 15341 23733 15353 23767
rect 15387 23733 15399 23767
rect 15341 23727 15399 23733
rect 15985 23767 16043 23773
rect 15985 23733 15997 23767
rect 16031 23764 16043 23767
rect 17362 23764 17368 23776
rect 16031 23736 17368 23764
rect 16031 23733 16043 23736
rect 15985 23727 16043 23733
rect 12578 23696 12584 23708
rect 12412 23668 12584 23696
rect 12578 23656 12584 23668
rect 12636 23656 12642 23708
rect 14970 23656 14976 23708
rect 15028 23696 15034 23708
rect 15356 23696 15384 23727
rect 17362 23724 17368 23736
rect 17420 23724 17426 23776
rect 18469 23767 18527 23773
rect 18469 23733 18481 23767
rect 18515 23764 18527 23767
rect 18650 23764 18656 23776
rect 18515 23736 18656 23764
rect 18515 23733 18527 23736
rect 18469 23727 18527 23733
rect 18650 23724 18656 23736
rect 18708 23724 18714 23776
rect 18852 23764 18880 23804
rect 18929 23801 18941 23835
rect 18975 23832 18987 23835
rect 19018 23832 19024 23844
rect 18975 23804 19024 23832
rect 18975 23801 18987 23804
rect 18929 23795 18987 23801
rect 19018 23792 19024 23804
rect 19076 23792 19082 23844
rect 20033 23835 20091 23841
rect 20033 23832 20045 23835
rect 19956 23804 20045 23832
rect 19956 23764 19984 23804
rect 20033 23801 20045 23804
rect 20079 23832 20091 23835
rect 21042 23832 21048 23844
rect 20079 23804 21048 23832
rect 20079 23801 20091 23804
rect 20033 23795 20091 23801
rect 21042 23792 21048 23804
rect 21100 23792 21106 23844
rect 21413 23835 21471 23841
rect 21413 23801 21425 23835
rect 21459 23832 21471 23835
rect 21870 23832 21876 23844
rect 21459 23804 21876 23832
rect 21459 23801 21471 23804
rect 21413 23795 21471 23801
rect 21870 23792 21876 23804
rect 21928 23792 21934 23844
rect 23342 23792 23348 23844
rect 23400 23832 23406 23844
rect 23894 23832 23900 23844
rect 23400 23804 23756 23832
rect 23855 23804 23900 23832
rect 23400 23792 23406 23804
rect 23728 23776 23756 23804
rect 23894 23792 23900 23804
rect 23952 23792 23958 23844
rect 24648 23841 24676 23872
rect 25200 23872 26016 23900
rect 25200 23841 25228 23872
rect 26010 23860 26016 23872
rect 26068 23860 26074 23912
rect 24633 23835 24691 23841
rect 24633 23801 24645 23835
rect 24679 23801 24691 23835
rect 24633 23795 24691 23801
rect 25185 23835 25243 23841
rect 25185 23801 25197 23835
rect 25231 23801 25243 23835
rect 25185 23795 25243 23801
rect 25645 23835 25703 23841
rect 25645 23801 25657 23835
rect 25691 23832 25703 23835
rect 25918 23832 25924 23844
rect 25691 23804 25924 23832
rect 25691 23801 25703 23804
rect 25645 23795 25703 23801
rect 20122 23764 20128 23776
rect 18852 23736 19984 23764
rect 20083 23736 20128 23764
rect 20122 23724 20128 23736
rect 20180 23724 20186 23776
rect 20585 23767 20643 23773
rect 20585 23733 20597 23767
rect 20631 23764 20643 23767
rect 20950 23764 20956 23776
rect 20631 23736 20956 23764
rect 20631 23733 20643 23736
rect 20585 23727 20643 23733
rect 20950 23724 20956 23736
rect 21008 23724 21014 23776
rect 21318 23724 21324 23776
rect 21376 23764 21382 23776
rect 21781 23767 21839 23773
rect 21781 23764 21793 23767
rect 21376 23736 21793 23764
rect 21376 23724 21382 23736
rect 21781 23733 21793 23736
rect 21827 23733 21839 23767
rect 21781 23727 21839 23733
rect 22054 23724 22060 23776
rect 22112 23764 22118 23776
rect 22517 23767 22575 23773
rect 22517 23764 22529 23767
rect 22112 23736 22529 23764
rect 22112 23724 22118 23736
rect 22517 23733 22529 23736
rect 22563 23733 22575 23767
rect 22517 23727 22575 23733
rect 22885 23767 22943 23773
rect 22885 23733 22897 23767
rect 22931 23764 22943 23767
rect 22974 23764 22980 23776
rect 22931 23736 22980 23764
rect 22931 23733 22943 23736
rect 22885 23727 22943 23733
rect 22974 23724 22980 23736
rect 23032 23724 23038 23776
rect 23526 23764 23532 23776
rect 23487 23736 23532 23764
rect 23526 23724 23532 23736
rect 23584 23724 23590 23776
rect 23710 23724 23716 23776
rect 23768 23764 23774 23776
rect 25200 23764 25228 23795
rect 25918 23792 25924 23804
rect 25976 23792 25982 23844
rect 27758 23832 27764 23844
rect 26948 23804 27764 23832
rect 23768 23736 25228 23764
rect 25461 23767 25519 23773
rect 23768 23724 23774 23736
rect 25461 23733 25473 23767
rect 25507 23733 25519 23767
rect 26102 23764 26108 23776
rect 26063 23736 26108 23764
rect 25461 23727 25519 23733
rect 16166 23696 16172 23708
rect 15028 23668 16172 23696
rect 15028 23656 15034 23668
rect 16166 23656 16172 23668
rect 16224 23656 16230 23708
rect 16810 23656 16816 23708
rect 16868 23696 16874 23708
rect 17089 23699 17147 23705
rect 17089 23696 17101 23699
rect 16868 23668 17101 23696
rect 16868 23656 16874 23668
rect 17089 23665 17101 23668
rect 17135 23665 17147 23699
rect 19478 23696 19484 23708
rect 17089 23659 17147 23665
rect 17656 23668 19484 23696
rect 13590 23628 13596 23640
rect 13551 23600 13596 23628
rect 13590 23588 13596 23600
rect 13648 23588 13654 23640
rect 15614 23588 15620 23640
rect 15672 23628 15678 23640
rect 17656 23628 17684 23668
rect 19478 23656 19484 23668
rect 19536 23696 19542 23708
rect 19536 23668 20812 23696
rect 19536 23656 19542 23668
rect 15672 23600 17684 23628
rect 17733 23631 17791 23637
rect 15672 23588 15678 23600
rect 17733 23597 17745 23631
rect 17779 23628 17791 23631
rect 19570 23628 19576 23640
rect 17779 23600 19576 23628
rect 17779 23597 17791 23600
rect 17733 23591 17791 23597
rect 19570 23588 19576 23600
rect 19628 23588 19634 23640
rect 20784 23628 20812 23668
rect 20858 23656 20864 23708
rect 20916 23696 20922 23708
rect 21045 23699 21103 23705
rect 21045 23696 21057 23699
rect 20916 23668 21057 23696
rect 20916 23656 20922 23668
rect 21045 23665 21057 23668
rect 21091 23665 21103 23699
rect 21045 23659 21103 23665
rect 22333 23699 22391 23705
rect 22333 23665 22345 23699
rect 22379 23696 22391 23699
rect 23345 23699 23403 23705
rect 23345 23696 23357 23699
rect 22379 23668 23357 23696
rect 22379 23665 22391 23668
rect 22333 23659 22391 23665
rect 23345 23665 23357 23668
rect 23391 23665 23403 23699
rect 23345 23659 23403 23665
rect 22348 23628 22376 23659
rect 20784 23600 22376 23628
rect 22422 23588 22428 23640
rect 22480 23628 22486 23640
rect 25476 23628 25504 23727
rect 26102 23724 26108 23736
rect 26160 23724 26166 23776
rect 26948 23773 26976 23804
rect 27758 23792 27764 23804
rect 27816 23792 27822 23844
rect 28494 23832 28500 23844
rect 28455 23804 28500 23832
rect 28494 23792 28500 23804
rect 28552 23792 28558 23844
rect 26933 23767 26991 23773
rect 26933 23733 26945 23767
rect 26979 23733 26991 23767
rect 26933 23727 26991 23733
rect 27025 23767 27083 23773
rect 27025 23733 27037 23767
rect 27071 23764 27083 23767
rect 27390 23764 27396 23776
rect 27071 23736 27396 23764
rect 27071 23733 27083 23736
rect 27025 23727 27083 23733
rect 27390 23724 27396 23736
rect 27448 23764 27454 23776
rect 27945 23767 28003 23773
rect 27945 23764 27957 23767
rect 27448 23736 27957 23764
rect 27448 23724 27454 23736
rect 27945 23733 27957 23736
rect 27991 23733 28003 23767
rect 29138 23764 29144 23776
rect 29099 23736 29144 23764
rect 27945 23727 28003 23733
rect 29138 23724 29144 23736
rect 29196 23724 29202 23776
rect 28402 23696 28408 23708
rect 28363 23668 28408 23696
rect 28402 23656 28408 23668
rect 28460 23656 28466 23708
rect 26194 23628 26200 23640
rect 22480 23600 25504 23628
rect 26155 23600 26200 23628
rect 22480 23588 22486 23600
rect 26194 23588 26200 23600
rect 26252 23588 26258 23640
rect 11000 23538 30136 23560
rect 11000 23486 19142 23538
rect 19194 23486 19206 23538
rect 19258 23486 19270 23538
rect 19322 23486 19334 23538
rect 19386 23486 29142 23538
rect 29194 23486 29206 23538
rect 29258 23486 29270 23538
rect 29322 23486 29334 23538
rect 29386 23486 30136 23538
rect 11000 23464 30136 23486
rect 14786 23424 14792 23436
rect 12872 23396 14792 23424
rect 12118 23316 12124 23368
rect 12176 23356 12182 23368
rect 12213 23359 12271 23365
rect 12213 23356 12225 23359
rect 12176 23328 12225 23356
rect 12176 23316 12182 23328
rect 12213 23325 12225 23328
rect 12259 23325 12271 23359
rect 12213 23319 12271 23325
rect 12872 23297 12900 23396
rect 14786 23384 14792 23396
rect 14844 23384 14850 23436
rect 16261 23427 16319 23433
rect 16261 23393 16273 23427
rect 16307 23424 16319 23427
rect 17086 23424 17092 23436
rect 16307 23396 17092 23424
rect 16307 23393 16319 23396
rect 16261 23387 16319 23393
rect 17086 23384 17092 23396
rect 17144 23424 17150 23436
rect 17273 23427 17331 23433
rect 17273 23424 17285 23427
rect 17144 23396 17285 23424
rect 17144 23384 17150 23396
rect 17273 23393 17285 23396
rect 17319 23393 17331 23427
rect 18190 23424 18196 23436
rect 18151 23396 18196 23424
rect 17273 23387 17331 23393
rect 18190 23384 18196 23396
rect 18248 23384 18254 23436
rect 19662 23424 19668 23436
rect 19623 23396 19668 23424
rect 19662 23384 19668 23396
rect 19720 23384 19726 23436
rect 20858 23424 20864 23436
rect 20819 23396 20864 23424
rect 20858 23384 20864 23396
rect 20916 23384 20922 23436
rect 20950 23384 20956 23436
rect 21008 23424 21014 23436
rect 25461 23427 25519 23433
rect 25461 23424 25473 23427
rect 21008 23396 24032 23424
rect 21008 23384 21014 23396
rect 13590 23316 13596 23368
rect 13648 23356 13654 23368
rect 13648 23328 14648 23356
rect 13648 23316 13654 23328
rect 12857 23291 12915 23297
rect 12857 23257 12869 23291
rect 12903 23257 12915 23291
rect 13222 23288 13228 23300
rect 13183 23260 13228 23288
rect 12857 23251 12915 23257
rect 13222 23248 13228 23260
rect 13280 23248 13286 23300
rect 13406 23288 13412 23300
rect 13367 23260 13412 23288
rect 13406 23248 13412 23260
rect 13464 23248 13470 23300
rect 13866 23248 13872 23300
rect 13924 23288 13930 23300
rect 14510 23288 14516 23300
rect 13924 23260 14096 23288
rect 14471 23260 14516 23288
rect 13924 23248 13930 23260
rect 12946 23220 12952 23232
rect 12907 23192 12952 23220
rect 12946 23180 12952 23192
rect 13004 23180 13010 23232
rect 13961 23223 14019 23229
rect 13961 23189 13973 23223
rect 14007 23189 14019 23223
rect 13961 23183 14019 23189
rect 12394 23112 12400 23164
rect 12452 23152 12458 23164
rect 13976 23152 14004 23183
rect 12452 23124 14004 23152
rect 14068 23152 14096 23260
rect 14510 23248 14516 23260
rect 14568 23248 14574 23300
rect 14620 23297 14648 23328
rect 15982 23316 15988 23368
rect 16040 23356 16046 23368
rect 16353 23359 16411 23365
rect 16353 23356 16365 23359
rect 16040 23328 16365 23356
rect 16040 23316 16046 23328
rect 16353 23325 16365 23328
rect 16399 23325 16411 23359
rect 16353 23319 16411 23325
rect 16994 23316 17000 23368
rect 17052 23356 17058 23368
rect 20217 23359 20275 23365
rect 20217 23356 20229 23359
rect 17052 23328 20229 23356
rect 17052 23316 17058 23328
rect 20217 23325 20229 23328
rect 20263 23356 20275 23359
rect 22238 23356 22244 23368
rect 20263 23328 22244 23356
rect 20263 23325 20275 23328
rect 20217 23319 20275 23325
rect 22238 23316 22244 23328
rect 22296 23316 22302 23368
rect 22333 23359 22391 23365
rect 22333 23325 22345 23359
rect 22379 23356 22391 23359
rect 22514 23356 22520 23368
rect 22379 23328 22520 23356
rect 22379 23325 22391 23328
rect 22333 23319 22391 23325
rect 22514 23316 22520 23328
rect 22572 23356 22578 23368
rect 23434 23356 23440 23368
rect 22572 23328 23440 23356
rect 22572 23316 22578 23328
rect 23434 23316 23440 23328
rect 23492 23316 23498 23368
rect 23710 23356 23716 23368
rect 23544 23328 23716 23356
rect 14605 23291 14663 23297
rect 14605 23257 14617 23291
rect 14651 23257 14663 23291
rect 14878 23288 14884 23300
rect 14839 23260 14884 23288
rect 14605 23251 14663 23257
rect 14878 23248 14884 23260
rect 14936 23248 14942 23300
rect 15430 23288 15436 23300
rect 15391 23260 15436 23288
rect 15430 23248 15436 23260
rect 15488 23248 15494 23300
rect 16166 23288 16172 23300
rect 16127 23260 16172 23288
rect 16166 23248 16172 23260
rect 16224 23248 16230 23300
rect 17086 23248 17092 23300
rect 17144 23288 17150 23300
rect 17181 23291 17239 23297
rect 17181 23288 17193 23291
rect 17144 23260 17193 23288
rect 17144 23248 17150 23260
rect 17181 23257 17193 23260
rect 17227 23257 17239 23291
rect 18006 23288 18012 23300
rect 17967 23260 18012 23288
rect 17181 23251 17239 23257
rect 18006 23248 18012 23260
rect 18064 23248 18070 23300
rect 18374 23288 18380 23300
rect 18335 23260 18380 23288
rect 18374 23248 18380 23260
rect 18432 23248 18438 23300
rect 19570 23288 19576 23300
rect 18484 23260 19432 23288
rect 19531 23260 19576 23288
rect 15062 23220 15068 23232
rect 15023 23192 15068 23220
rect 15062 23180 15068 23192
rect 15120 23180 15126 23232
rect 15985 23223 16043 23229
rect 15985 23189 15997 23223
rect 16031 23220 16043 23223
rect 16258 23220 16264 23232
rect 16031 23192 16264 23220
rect 16031 23189 16043 23192
rect 15985 23183 16043 23189
rect 16258 23180 16264 23192
rect 16316 23180 16322 23232
rect 16534 23180 16540 23232
rect 16592 23220 16598 23232
rect 16721 23223 16779 23229
rect 16721 23220 16733 23223
rect 16592 23192 16733 23220
rect 16592 23180 16598 23192
rect 16721 23189 16733 23192
rect 16767 23220 16779 23223
rect 18484 23220 18512 23260
rect 16767 23192 18512 23220
rect 19404 23220 19432 23260
rect 19570 23248 19576 23260
rect 19628 23248 19634 23300
rect 20030 23248 20036 23300
rect 20088 23288 20094 23300
rect 20858 23288 20864 23300
rect 20088 23260 20864 23288
rect 20088 23248 20094 23260
rect 20858 23248 20864 23260
rect 20916 23248 20922 23300
rect 22054 23248 22060 23300
rect 22112 23288 22118 23300
rect 23544 23297 23572 23328
rect 23710 23316 23716 23328
rect 23768 23316 23774 23368
rect 24004 23365 24032 23396
rect 24096 23396 25473 23424
rect 23989 23359 24047 23365
rect 23989 23325 24001 23359
rect 24035 23325 24047 23359
rect 23989 23319 24047 23325
rect 22977 23291 23035 23297
rect 22977 23288 22989 23291
rect 22112 23260 22989 23288
rect 22112 23248 22118 23260
rect 22977 23257 22989 23260
rect 23023 23257 23035 23291
rect 22977 23251 23035 23257
rect 23345 23291 23403 23297
rect 23345 23257 23357 23291
rect 23391 23257 23403 23291
rect 23529 23291 23587 23297
rect 23529 23288 23541 23291
rect 23345 23251 23403 23257
rect 23452 23260 23541 23288
rect 19754 23220 19760 23232
rect 19404 23192 19760 23220
rect 16767 23189 16779 23192
rect 16721 23183 16779 23189
rect 19754 23180 19760 23192
rect 19812 23180 19818 23232
rect 19938 23180 19944 23232
rect 19996 23220 20002 23232
rect 20398 23229 20404 23232
rect 20364 23223 20404 23229
rect 20364 23220 20376 23223
rect 19996 23192 20376 23220
rect 19996 23180 20002 23192
rect 20364 23189 20376 23192
rect 20364 23183 20404 23189
rect 20398 23180 20404 23183
rect 20456 23180 20462 23232
rect 20490 23180 20496 23232
rect 20548 23220 20554 23232
rect 20585 23223 20643 23229
rect 20585 23220 20597 23223
rect 20548 23192 20597 23220
rect 20548 23180 20554 23192
rect 20585 23189 20597 23192
rect 20631 23189 20643 23223
rect 20585 23183 20643 23189
rect 20674 23180 20680 23232
rect 20732 23220 20738 23232
rect 20732 23192 22836 23220
rect 20732 23180 20738 23192
rect 22808 23152 22836 23192
rect 22882 23180 22888 23232
rect 22940 23220 22946 23232
rect 22940 23192 22985 23220
rect 22940 23180 22946 23192
rect 23360 23152 23388 23251
rect 23452 23232 23480 23260
rect 23529 23257 23541 23260
rect 23575 23257 23587 23291
rect 23529 23251 23587 23257
rect 23618 23248 23624 23300
rect 23676 23288 23682 23300
rect 24096 23288 24124 23396
rect 25461 23393 25473 23396
rect 25507 23393 25519 23427
rect 25461 23387 25519 23393
rect 24538 23316 24544 23368
rect 24596 23356 24602 23368
rect 25185 23359 25243 23365
rect 25185 23356 25197 23359
rect 24596 23328 25197 23356
rect 24596 23316 24602 23328
rect 25185 23325 25197 23328
rect 25231 23325 25243 23359
rect 25185 23319 25243 23325
rect 26749 23359 26807 23365
rect 26749 23325 26761 23359
rect 26795 23356 26807 23359
rect 28402 23356 28408 23368
rect 26795 23328 28408 23356
rect 26795 23325 26807 23328
rect 26749 23319 26807 23325
rect 28402 23316 28408 23328
rect 28460 23356 28466 23368
rect 28957 23359 29015 23365
rect 28957 23356 28969 23359
rect 28460 23328 28969 23356
rect 28460 23316 28466 23328
rect 28957 23325 28969 23328
rect 29003 23325 29015 23359
rect 28957 23319 29015 23325
rect 23676 23260 24124 23288
rect 24173 23291 24231 23297
rect 23676 23248 23682 23260
rect 24173 23257 24185 23291
rect 24219 23288 24231 23291
rect 25090 23288 25096 23300
rect 24219 23260 25096 23288
rect 24219 23257 24231 23260
rect 24173 23251 24231 23257
rect 25090 23248 25096 23260
rect 25148 23248 25154 23300
rect 25369 23291 25427 23297
rect 25369 23257 25381 23291
rect 25415 23257 25427 23291
rect 27390 23288 27396 23300
rect 27351 23260 27396 23288
rect 25369 23251 25427 23257
rect 23434 23180 23440 23232
rect 23492 23180 23498 23232
rect 24538 23180 24544 23232
rect 24596 23220 24602 23232
rect 25384 23220 25412 23251
rect 27390 23248 27396 23260
rect 27448 23248 27454 23300
rect 28218 23248 28224 23300
rect 28276 23288 28282 23300
rect 28313 23291 28371 23297
rect 28313 23288 28325 23291
rect 28276 23260 28325 23288
rect 28276 23248 28282 23260
rect 28313 23257 28325 23260
rect 28359 23257 28371 23291
rect 28313 23251 28371 23257
rect 24596 23192 25412 23220
rect 24596 23180 24602 23192
rect 14068 23124 22560 23152
rect 22808 23124 23388 23152
rect 12452 23112 12458 23124
rect 17546 23044 17552 23096
rect 17604 23084 17610 23096
rect 18190 23084 18196 23096
rect 17604 23056 18196 23084
rect 17604 23044 17610 23056
rect 18190 23044 18196 23056
rect 18248 23084 18254 23096
rect 19294 23084 19300 23096
rect 18248 23056 19300 23084
rect 18248 23044 18254 23056
rect 19294 23044 19300 23056
rect 19352 23044 19358 23096
rect 19754 23044 19760 23096
rect 19812 23084 19818 23096
rect 20493 23087 20551 23093
rect 20493 23084 20505 23087
rect 19812 23056 20505 23084
rect 19812 23044 19818 23056
rect 20493 23053 20505 23056
rect 20539 23053 20551 23087
rect 20493 23047 20551 23053
rect 20858 23044 20864 23096
rect 20916 23084 20922 23096
rect 22422 23084 22428 23096
rect 20916 23056 22428 23084
rect 20916 23044 20922 23056
rect 22422 23044 22428 23056
rect 22480 23044 22486 23096
rect 22532 23084 22560 23124
rect 23802 23112 23808 23164
rect 23860 23152 23866 23164
rect 28310 23152 28316 23164
rect 23860 23124 28316 23152
rect 23860 23112 23866 23124
rect 28310 23112 28316 23124
rect 28368 23112 28374 23164
rect 23526 23084 23532 23096
rect 22532 23056 23532 23084
rect 23526 23044 23532 23056
rect 23584 23044 23590 23096
rect 23894 23044 23900 23096
rect 23952 23084 23958 23096
rect 24265 23087 24323 23093
rect 24265 23084 24277 23087
rect 23952 23056 24277 23084
rect 23952 23044 23958 23056
rect 24265 23053 24277 23056
rect 24311 23053 24323 23087
rect 24265 23047 24323 23053
rect 26654 23044 26660 23096
rect 26712 23084 26718 23096
rect 26841 23087 26899 23093
rect 26841 23084 26853 23087
rect 26712 23056 26853 23084
rect 26712 23044 26718 23056
rect 26841 23053 26853 23056
rect 26887 23053 26899 23087
rect 26841 23047 26899 23053
rect 11000 22994 30136 23016
rect 11000 22942 14142 22994
rect 14194 22942 14206 22994
rect 14258 22942 14270 22994
rect 14322 22942 14334 22994
rect 14386 22942 24142 22994
rect 24194 22942 24206 22994
rect 24258 22942 24270 22994
rect 24322 22942 24334 22994
rect 24386 22942 30136 22994
rect 11000 22920 30136 22942
rect 13222 22840 13228 22892
rect 13280 22880 13286 22892
rect 13961 22883 14019 22889
rect 13961 22880 13973 22883
rect 13280 22852 13973 22880
rect 13280 22840 13286 22852
rect 13961 22849 13973 22852
rect 14007 22880 14019 22883
rect 15062 22880 15068 22892
rect 14007 22852 15068 22880
rect 14007 22849 14019 22852
rect 13961 22843 14019 22849
rect 15062 22840 15068 22852
rect 15120 22840 15126 22892
rect 15246 22840 15252 22892
rect 15304 22880 15310 22892
rect 16626 22880 16632 22892
rect 15304 22852 16632 22880
rect 15304 22840 15310 22852
rect 16626 22840 16632 22852
rect 16684 22840 16690 22892
rect 19662 22840 19668 22892
rect 19720 22880 19726 22892
rect 20447 22883 20505 22889
rect 20447 22880 20459 22883
rect 19720 22852 20459 22880
rect 19720 22840 19726 22852
rect 20447 22849 20459 22852
rect 20493 22849 20505 22883
rect 22790 22880 22796 22892
rect 20447 22843 20505 22849
rect 20600 22852 22796 22880
rect 20122 22812 20128 22824
rect 18024 22784 20128 22812
rect 12210 22744 12216 22756
rect 12171 22716 12216 22744
rect 12210 22704 12216 22716
rect 12268 22704 12274 22756
rect 15430 22704 15436 22756
rect 15488 22744 15494 22756
rect 15617 22747 15675 22753
rect 15617 22744 15629 22747
rect 15488 22716 15629 22744
rect 15488 22704 15494 22716
rect 15617 22713 15629 22716
rect 15663 22744 15675 22747
rect 16994 22744 17000 22756
rect 15663 22716 17000 22744
rect 15663 22713 15675 22716
rect 15617 22707 15675 22713
rect 16994 22704 17000 22716
rect 17052 22744 17058 22756
rect 17052 22716 17500 22744
rect 17052 22704 17058 22716
rect 12118 22676 12124 22688
rect 12079 22648 12124 22676
rect 12118 22636 12124 22648
rect 12176 22636 12182 22688
rect 12394 22676 12400 22688
rect 12355 22648 12400 22676
rect 12394 22636 12400 22648
rect 12452 22636 12458 22688
rect 13869 22679 13927 22685
rect 13869 22676 13881 22679
rect 13700 22648 13881 22676
rect 13700 22620 13728 22648
rect 13869 22645 13881 22648
rect 13915 22676 13927 22679
rect 14786 22676 14792 22688
rect 13915 22648 14792 22676
rect 13915 22645 13927 22648
rect 13869 22639 13927 22645
rect 14786 22636 14792 22648
rect 14844 22636 14850 22688
rect 15246 22676 15252 22688
rect 15207 22648 15252 22676
rect 15246 22636 15252 22648
rect 15304 22636 15310 22688
rect 16626 22636 16632 22688
rect 16684 22676 16690 22688
rect 16721 22679 16779 22685
rect 16721 22676 16733 22679
rect 16684 22648 16733 22676
rect 16684 22636 16690 22648
rect 16721 22645 16733 22648
rect 16767 22645 16779 22679
rect 16721 22639 16779 22645
rect 16905 22679 16963 22685
rect 16905 22645 16917 22679
rect 16951 22645 16963 22679
rect 17086 22676 17092 22688
rect 17047 22648 17092 22676
rect 16905 22639 16963 22645
rect 13682 22568 13688 22620
rect 13740 22568 13746 22620
rect 14694 22568 14700 22620
rect 14752 22608 14758 22620
rect 15065 22611 15123 22617
rect 15065 22608 15077 22611
rect 14752 22580 15077 22608
rect 14752 22568 14758 22580
rect 15065 22577 15077 22580
rect 15111 22577 15123 22611
rect 15065 22571 15123 22577
rect 15080 22540 15108 22571
rect 16166 22568 16172 22620
rect 16224 22608 16230 22620
rect 16920 22608 16948 22639
rect 17086 22636 17092 22648
rect 17144 22636 17150 22688
rect 17472 22685 17500 22716
rect 18024 22688 18052 22784
rect 18285 22747 18343 22753
rect 18285 22713 18297 22747
rect 18331 22744 18343 22747
rect 18374 22744 18380 22756
rect 18331 22716 18380 22744
rect 18331 22713 18343 22716
rect 18285 22707 18343 22713
rect 18374 22704 18380 22716
rect 18432 22704 18438 22756
rect 18742 22704 18748 22756
rect 18800 22744 18806 22756
rect 19113 22747 19171 22753
rect 19113 22744 19125 22747
rect 18800 22716 19125 22744
rect 18800 22704 18806 22716
rect 19113 22713 19125 22716
rect 19159 22713 19171 22747
rect 19113 22707 19171 22713
rect 17457 22679 17515 22685
rect 17457 22645 17469 22679
rect 17503 22645 17515 22679
rect 17457 22639 17515 22645
rect 17710 22679 17768 22685
rect 17710 22645 17722 22679
rect 17756 22676 17768 22679
rect 18006 22676 18012 22688
rect 17756 22648 18012 22676
rect 17756 22645 17768 22648
rect 17710 22639 17768 22645
rect 18006 22636 18012 22648
rect 18064 22636 18070 22688
rect 19294 22676 19300 22688
rect 19255 22648 19300 22676
rect 19294 22636 19300 22648
rect 19352 22636 19358 22688
rect 17270 22608 17276 22620
rect 16224 22580 17276 22608
rect 16224 22568 16230 22580
rect 17270 22568 17276 22580
rect 17328 22568 17334 22620
rect 18098 22568 18104 22620
rect 18156 22608 18162 22620
rect 19404 22608 19432 22784
rect 20122 22772 20128 22784
rect 20180 22772 20186 22824
rect 20600 22821 20628 22852
rect 22790 22840 22796 22852
rect 22848 22840 22854 22892
rect 22885 22883 22943 22889
rect 22885 22849 22897 22883
rect 22931 22880 22943 22883
rect 23342 22880 23348 22892
rect 22931 22852 23348 22880
rect 22931 22849 22943 22852
rect 22885 22843 22943 22849
rect 23342 22840 23348 22852
rect 23400 22840 23406 22892
rect 23526 22840 23532 22892
rect 23584 22880 23590 22892
rect 23584 22852 24860 22880
rect 23584 22840 23590 22852
rect 20585 22815 20643 22821
rect 20585 22812 20597 22815
rect 20416 22784 20597 22812
rect 20416 22756 20444 22784
rect 20585 22781 20597 22784
rect 20631 22781 20643 22815
rect 21042 22812 21048 22824
rect 20585 22775 20643 22781
rect 20692 22784 21048 22812
rect 19478 22704 19484 22756
rect 19536 22744 19542 22756
rect 19849 22747 19907 22753
rect 19849 22744 19861 22747
rect 19536 22716 19861 22744
rect 19536 22704 19542 22716
rect 19849 22713 19861 22716
rect 19895 22713 19907 22747
rect 19849 22707 19907 22713
rect 20398 22704 20404 22756
rect 20456 22704 20462 22756
rect 20692 22753 20720 22784
rect 21042 22772 21048 22784
rect 21100 22812 21106 22824
rect 23434 22812 23440 22824
rect 21100 22784 23440 22812
rect 21100 22772 21106 22784
rect 21520 22756 21548 22784
rect 23434 22772 23440 22784
rect 23492 22772 23498 22824
rect 23710 22772 23716 22824
rect 23768 22812 23774 22824
rect 23768 22784 24032 22812
rect 23768 22772 23774 22784
rect 20677 22747 20735 22753
rect 20677 22713 20689 22747
rect 20723 22713 20735 22747
rect 20677 22707 20735 22713
rect 21502 22704 21508 22756
rect 21560 22704 21566 22756
rect 22977 22747 23035 22753
rect 22977 22713 22989 22747
rect 23023 22744 23035 22747
rect 23158 22744 23164 22756
rect 23023 22716 23164 22744
rect 23023 22713 23035 22716
rect 22977 22707 23035 22713
rect 23158 22704 23164 22716
rect 23216 22704 23222 22756
rect 23894 22744 23900 22756
rect 23855 22716 23900 22744
rect 23894 22704 23900 22716
rect 23952 22704 23958 22756
rect 24004 22753 24032 22784
rect 24832 22753 24860 22852
rect 25090 22840 25096 22892
rect 25148 22880 25154 22892
rect 25645 22883 25703 22889
rect 25645 22880 25657 22883
rect 25148 22852 25657 22880
rect 25148 22840 25154 22852
rect 25645 22849 25657 22852
rect 25691 22849 25703 22883
rect 25645 22843 25703 22849
rect 23989 22747 24047 22753
rect 23989 22713 24001 22747
rect 24035 22713 24047 22747
rect 23989 22707 24047 22713
rect 24817 22747 24875 22753
rect 24817 22713 24829 22747
rect 24863 22713 24875 22747
rect 24817 22707 24875 22713
rect 24998 22704 25004 22756
rect 25056 22744 25062 22756
rect 25056 22716 25596 22744
rect 25056 22704 25062 22716
rect 20214 22636 20220 22688
rect 20272 22676 20278 22688
rect 20309 22679 20367 22685
rect 20309 22676 20321 22679
rect 20272 22648 20321 22676
rect 20272 22636 20278 22648
rect 20309 22645 20321 22648
rect 20355 22645 20367 22679
rect 21042 22676 21048 22688
rect 21003 22648 21048 22676
rect 20309 22639 20367 22645
rect 21042 22636 21048 22648
rect 21100 22636 21106 22688
rect 22514 22636 22520 22688
rect 22572 22676 22578 22688
rect 22609 22679 22667 22685
rect 22609 22676 22621 22679
rect 22572 22648 22621 22676
rect 22572 22636 22578 22648
rect 22609 22645 22621 22648
rect 22655 22645 22667 22679
rect 22609 22639 22667 22645
rect 22756 22679 22814 22685
rect 22756 22645 22768 22679
rect 22802 22676 22814 22679
rect 23250 22676 23256 22688
rect 22802 22648 23256 22676
rect 22802 22645 22814 22648
rect 22756 22639 22814 22645
rect 23250 22636 23256 22648
rect 23308 22636 23314 22688
rect 23345 22679 23403 22685
rect 23345 22645 23357 22679
rect 23391 22676 23403 22679
rect 23802 22676 23808 22688
rect 23391 22648 23808 22676
rect 23391 22645 23403 22648
rect 23345 22639 23403 22645
rect 23802 22636 23808 22648
rect 23860 22636 23866 22688
rect 24538 22676 24544 22688
rect 23912 22648 24544 22676
rect 19465 22611 19523 22617
rect 19465 22608 19477 22611
rect 18156 22580 19156 22608
rect 19404 22580 19477 22608
rect 18156 22568 18162 22580
rect 16442 22540 16448 22552
rect 15080 22512 16448 22540
rect 16442 22500 16448 22512
rect 16500 22500 16506 22552
rect 19128 22540 19156 22580
rect 19465 22577 19477 22580
rect 19511 22577 19523 22611
rect 19465 22571 19523 22577
rect 21226 22568 21232 22620
rect 21284 22608 21290 22620
rect 23912 22608 23940 22648
rect 24538 22636 24544 22648
rect 24596 22636 24602 22688
rect 24725 22679 24783 22685
rect 24725 22645 24737 22679
rect 24771 22676 24783 22679
rect 24906 22676 24912 22688
rect 24771 22648 24912 22676
rect 24771 22645 24783 22648
rect 24725 22639 24783 22645
rect 24906 22636 24912 22648
rect 24964 22636 24970 22688
rect 25366 22676 25372 22688
rect 25327 22648 25372 22676
rect 25366 22636 25372 22648
rect 25424 22636 25430 22688
rect 25568 22685 25596 22716
rect 26194 22704 26200 22756
rect 26252 22744 26258 22756
rect 26381 22747 26439 22753
rect 26381 22744 26393 22747
rect 26252 22716 26393 22744
rect 26252 22704 26258 22716
rect 26381 22713 26393 22716
rect 26427 22713 26439 22747
rect 26381 22707 26439 22713
rect 26933 22747 26991 22753
rect 26933 22713 26945 22747
rect 26979 22744 26991 22747
rect 27022 22744 27028 22756
rect 26979 22716 27028 22744
rect 26979 22713 26991 22716
rect 26933 22707 26991 22713
rect 27022 22704 27028 22716
rect 27080 22704 27086 22756
rect 25553 22679 25611 22685
rect 25553 22645 25565 22679
rect 25599 22645 25611 22679
rect 25553 22639 25611 22645
rect 28405 22679 28463 22685
rect 28405 22645 28417 22679
rect 28451 22676 28463 22679
rect 28586 22676 28592 22688
rect 28451 22648 28592 22676
rect 28451 22645 28463 22648
rect 28405 22639 28463 22645
rect 28586 22636 28592 22648
rect 28644 22636 28650 22688
rect 28954 22636 28960 22688
rect 29012 22676 29018 22688
rect 29049 22679 29107 22685
rect 29049 22676 29061 22679
rect 29012 22648 29061 22676
rect 29012 22636 29018 22648
rect 29049 22645 29061 22648
rect 29095 22645 29107 22679
rect 29049 22639 29107 22645
rect 21284 22580 23940 22608
rect 26841 22611 26899 22617
rect 21284 22568 21290 22580
rect 26841 22577 26853 22611
rect 26887 22608 26899 22611
rect 27390 22608 27396 22620
rect 26887 22580 27396 22608
rect 26887 22577 26899 22580
rect 26841 22571 26899 22577
rect 27390 22568 27396 22580
rect 27448 22568 27454 22620
rect 28218 22568 28224 22620
rect 28276 22608 28282 22620
rect 29325 22611 29383 22617
rect 29325 22608 29337 22611
rect 28276 22580 29337 22608
rect 28276 22568 28282 22580
rect 29325 22577 29337 22580
rect 29371 22577 29383 22611
rect 29325 22571 29383 22577
rect 19389 22543 19447 22549
rect 19389 22540 19401 22543
rect 19128 22512 19401 22540
rect 19389 22509 19401 22512
rect 19435 22509 19447 22543
rect 19389 22503 19447 22509
rect 22330 22500 22336 22552
rect 22388 22540 22394 22552
rect 23250 22540 23256 22552
rect 22388 22512 23256 22540
rect 22388 22500 22394 22512
rect 23250 22500 23256 22512
rect 23308 22500 23314 22552
rect 11000 22450 30136 22472
rect 11000 22398 19142 22450
rect 19194 22398 19206 22450
rect 19258 22398 19270 22450
rect 19322 22398 19334 22450
rect 19386 22398 29142 22450
rect 29194 22398 29206 22450
rect 29258 22398 29270 22450
rect 29322 22398 29334 22450
rect 29386 22398 30136 22450
rect 11000 22376 30136 22398
rect 19665 22339 19723 22345
rect 19665 22305 19677 22339
rect 19711 22336 19723 22339
rect 20674 22336 20680 22348
rect 19711 22308 20680 22336
rect 19711 22305 19723 22308
rect 19665 22299 19723 22305
rect 20674 22296 20680 22308
rect 20732 22296 20738 22348
rect 21962 22336 21968 22348
rect 21428 22308 21968 22336
rect 21428 22280 21456 22308
rect 21962 22296 21968 22308
rect 22020 22296 22026 22348
rect 22606 22296 22612 22348
rect 22664 22336 22670 22348
rect 24265 22339 24323 22345
rect 24265 22336 24277 22339
rect 22664 22308 24277 22336
rect 22664 22296 22670 22308
rect 24265 22305 24277 22308
rect 24311 22305 24323 22339
rect 24265 22299 24323 22305
rect 13958 22268 13964 22280
rect 13919 22240 13964 22268
rect 13958 22228 13964 22240
rect 14016 22228 14022 22280
rect 15062 22228 15068 22280
rect 15120 22268 15126 22280
rect 15433 22271 15491 22277
rect 15433 22268 15445 22271
rect 15120 22240 15445 22268
rect 15120 22228 15126 22240
rect 15433 22237 15445 22240
rect 15479 22237 15491 22271
rect 16994 22268 17000 22280
rect 15433 22231 15491 22237
rect 16828 22240 17000 22268
rect 11845 22203 11903 22209
rect 11845 22169 11857 22203
rect 11891 22200 11903 22203
rect 11934 22200 11940 22212
rect 11891 22172 11940 22200
rect 11891 22169 11903 22172
rect 11845 22163 11903 22169
rect 11934 22160 11940 22172
rect 11992 22160 11998 22212
rect 14786 22200 14792 22212
rect 14747 22172 14792 22200
rect 14786 22160 14792 22172
rect 14844 22160 14850 22212
rect 14973 22203 15031 22209
rect 14973 22169 14985 22203
rect 15019 22200 15031 22203
rect 15246 22200 15252 22212
rect 15019 22172 15252 22200
rect 15019 22169 15031 22172
rect 14973 22163 15031 22169
rect 15246 22160 15252 22172
rect 15304 22160 15310 22212
rect 15617 22203 15675 22209
rect 15617 22169 15629 22203
rect 15663 22200 15675 22203
rect 16258 22200 16264 22212
rect 15663 22172 16264 22200
rect 15663 22169 15675 22172
rect 15617 22163 15675 22169
rect 16258 22160 16264 22172
rect 16316 22160 16322 22212
rect 16828 22209 16856 22240
rect 16994 22228 17000 22240
rect 17052 22268 17058 22280
rect 18561 22271 18619 22277
rect 17052 22240 18512 22268
rect 17052 22228 17058 22240
rect 16813 22203 16871 22209
rect 16813 22169 16825 22203
rect 16859 22169 16871 22203
rect 18098 22200 18104 22212
rect 18059 22172 18104 22200
rect 16813 22163 16871 22169
rect 18098 22160 18104 22172
rect 18156 22160 18162 22212
rect 18374 22200 18380 22212
rect 18335 22172 18380 22200
rect 18374 22160 18380 22172
rect 18432 22160 18438 22212
rect 18484 22200 18512 22240
rect 18561 22237 18573 22271
rect 18607 22268 18619 22271
rect 20214 22268 20220 22280
rect 18607 22240 20220 22268
rect 18607 22237 18619 22240
rect 18561 22231 18619 22237
rect 20214 22228 20220 22240
rect 20272 22228 20278 22280
rect 20861 22271 20919 22277
rect 20861 22237 20873 22271
rect 20907 22268 20919 22271
rect 21410 22268 21416 22280
rect 20907 22240 21416 22268
rect 20907 22237 20919 22240
rect 20861 22231 20919 22237
rect 21410 22228 21416 22240
rect 21468 22228 21474 22280
rect 21597 22271 21655 22277
rect 21597 22237 21609 22271
rect 21643 22268 21655 22271
rect 21643 22240 22983 22268
rect 21643 22237 21655 22240
rect 21597 22231 21655 22237
rect 22955 22212 22983 22240
rect 23894 22228 23900 22280
rect 23952 22268 23958 22280
rect 28497 22271 28555 22277
rect 23952 22240 24216 22268
rect 23952 22228 23958 22240
rect 19573 22203 19631 22209
rect 19573 22200 19585 22203
rect 18484 22172 19585 22200
rect 19573 22169 19585 22172
rect 19619 22169 19631 22203
rect 19573 22163 19631 22169
rect 19754 22160 19760 22212
rect 19812 22200 19818 22212
rect 20309 22203 20367 22209
rect 20309 22200 20321 22203
rect 19812 22172 20321 22200
rect 19812 22160 19818 22172
rect 20309 22169 20321 22172
rect 20355 22169 20367 22203
rect 20490 22200 20496 22212
rect 20451 22172 20496 22200
rect 20309 22163 20367 22169
rect 20490 22160 20496 22172
rect 20548 22160 20554 22212
rect 21686 22160 21692 22212
rect 21744 22200 21750 22212
rect 22955 22209 22980 22212
rect 22793 22203 22851 22209
rect 22793 22200 22805 22203
rect 21744 22172 22805 22200
rect 21744 22160 21750 22172
rect 22793 22169 22805 22172
rect 22839 22169 22851 22203
rect 22793 22163 22851 22169
rect 22940 22203 22980 22209
rect 22940 22169 22952 22203
rect 22940 22163 22980 22169
rect 22974 22160 22980 22163
rect 23032 22160 23038 22212
rect 23250 22160 23256 22212
rect 23308 22200 23314 22212
rect 24188 22209 24216 22240
rect 28497 22237 28509 22271
rect 28543 22268 28555 22271
rect 28586 22268 28592 22280
rect 28543 22240 28592 22268
rect 28543 22237 28555 22240
rect 28497 22231 28555 22237
rect 28586 22228 28592 22240
rect 28644 22228 28650 22280
rect 23989 22203 24047 22209
rect 23989 22200 24001 22203
rect 23308 22172 24001 22200
rect 23308 22160 23314 22172
rect 23989 22169 24001 22172
rect 24035 22169 24047 22203
rect 23989 22163 24047 22169
rect 24173 22203 24231 22209
rect 24173 22169 24185 22203
rect 24219 22169 24231 22203
rect 24173 22163 24231 22169
rect 25090 22160 25096 22212
rect 25148 22200 25154 22212
rect 25185 22203 25243 22209
rect 25185 22200 25197 22203
rect 25148 22172 25197 22200
rect 25148 22160 25154 22172
rect 25185 22169 25197 22172
rect 25231 22169 25243 22203
rect 25185 22163 25243 22169
rect 25921 22203 25979 22209
rect 25921 22169 25933 22203
rect 25967 22200 25979 22203
rect 26194 22200 26200 22212
rect 25967 22172 26200 22200
rect 25967 22169 25979 22172
rect 25921 22163 25979 22169
rect 26194 22160 26200 22172
rect 26252 22160 26258 22212
rect 26378 22160 26384 22212
rect 26436 22200 26442 22212
rect 26841 22203 26899 22209
rect 26841 22200 26853 22203
rect 26436 22172 26853 22200
rect 26436 22160 26442 22172
rect 26841 22169 26853 22172
rect 26887 22169 26899 22203
rect 26841 22163 26899 22169
rect 29233 22203 29291 22209
rect 29233 22169 29245 22203
rect 29279 22200 29291 22203
rect 29874 22200 29880 22212
rect 29279 22172 29880 22200
rect 29279 22169 29291 22172
rect 29233 22163 29291 22169
rect 29874 22160 29880 22172
rect 29932 22160 29938 22212
rect 14513 22135 14571 22141
rect 14513 22101 14525 22135
rect 14559 22101 14571 22135
rect 14513 22095 14571 22101
rect 16721 22135 16779 22141
rect 16721 22101 16733 22135
rect 16767 22132 16779 22135
rect 17178 22132 17184 22144
rect 16767 22104 17184 22132
rect 16767 22101 16779 22104
rect 16721 22095 16779 22101
rect 12026 21996 12032 22008
rect 11987 21968 12032 21996
rect 12026 21956 12032 21968
rect 12084 21956 12090 22008
rect 14528 21996 14556 22095
rect 17178 22092 17184 22104
rect 17236 22092 17242 22144
rect 20398 22092 20404 22144
rect 20456 22132 20462 22144
rect 20582 22132 20588 22144
rect 20456 22104 20588 22132
rect 20456 22092 20462 22104
rect 20582 22092 20588 22104
rect 20640 22092 20646 22144
rect 21870 22092 21876 22144
rect 21928 22092 21934 22144
rect 21962 22092 21968 22144
rect 22020 22132 22026 22144
rect 23158 22132 23164 22144
rect 22020 22104 22065 22132
rect 22440 22104 23164 22132
rect 22020 22092 22026 22104
rect 21762 22067 21820 22073
rect 21762 22033 21774 22067
rect 21808 22064 21820 22067
rect 21888 22064 21916 22092
rect 22440 22064 22468 22104
rect 23158 22092 23164 22104
rect 23216 22092 23222 22144
rect 23529 22135 23587 22141
rect 23529 22101 23541 22135
rect 23575 22132 23587 22135
rect 28405 22135 28463 22141
rect 28405 22132 28417 22135
rect 23575 22104 28417 22132
rect 23575 22101 23587 22104
rect 23529 22095 23587 22101
rect 28405 22101 28417 22104
rect 28451 22101 28463 22135
rect 29322 22132 29328 22144
rect 29283 22104 29328 22132
rect 28405 22095 28463 22101
rect 29322 22092 29328 22104
rect 29380 22092 29386 22144
rect 21808 22036 22468 22064
rect 23069 22067 23127 22073
rect 21808 22033 21820 22036
rect 21762 22027 21820 22033
rect 23069 22033 23081 22067
rect 23115 22064 23127 22067
rect 23618 22064 23624 22076
rect 23115 22036 23624 22064
rect 23115 22033 23127 22036
rect 23069 22027 23127 22033
rect 15709 21999 15767 22005
rect 15709 21996 15721 21999
rect 14528 21968 15721 21996
rect 15709 21965 15721 21968
rect 15755 21996 15767 21999
rect 15798 21996 15804 22008
rect 15755 21968 15804 21996
rect 15755 21965 15767 21968
rect 15709 21959 15767 21965
rect 15798 21956 15804 21968
rect 15856 21956 15862 22008
rect 16810 21956 16816 22008
rect 16868 21996 16874 22008
rect 16997 21999 17055 22005
rect 16997 21996 17009 21999
rect 16868 21968 17009 21996
rect 16868 21956 16874 21968
rect 16997 21965 17009 21968
rect 17043 21965 17055 21999
rect 16997 21959 17055 21965
rect 21226 21956 21232 22008
rect 21284 21996 21290 22008
rect 21873 21999 21931 22005
rect 21873 21996 21885 21999
rect 21284 21968 21885 21996
rect 21284 21956 21290 21968
rect 21873 21965 21885 21968
rect 21919 21965 21931 21999
rect 21873 21959 21931 21965
rect 21962 21956 21968 22008
rect 22020 21996 22026 22008
rect 22057 21999 22115 22005
rect 22057 21996 22069 21999
rect 22020 21968 22069 21996
rect 22020 21956 22026 21968
rect 22057 21965 22069 21968
rect 22103 21965 22115 21999
rect 22057 21959 22115 21965
rect 22330 21956 22336 22008
rect 22388 21996 22394 22008
rect 23084 21996 23112 22027
rect 23618 22024 23624 22036
rect 23676 22024 23682 22076
rect 27390 22064 27396 22076
rect 27351 22036 27396 22064
rect 27390 22024 27396 22036
rect 27448 22024 27454 22076
rect 25274 21996 25280 22008
rect 22388 21968 23112 21996
rect 25235 21968 25280 21996
rect 22388 21956 22394 21968
rect 25274 21956 25280 21968
rect 25332 21956 25338 22008
rect 11000 21906 30136 21928
rect 11000 21854 14142 21906
rect 14194 21854 14206 21906
rect 14258 21854 14270 21906
rect 14322 21854 14334 21906
rect 14386 21854 24142 21906
rect 24194 21854 24206 21906
rect 24258 21854 24270 21906
rect 24322 21854 24334 21906
rect 24386 21854 30136 21906
rect 11000 21832 30136 21854
rect 16994 21792 17000 21804
rect 16955 21764 17000 21792
rect 16994 21752 17000 21764
rect 17052 21752 17058 21804
rect 18006 21792 18012 21804
rect 17967 21764 18012 21792
rect 18006 21752 18012 21764
rect 18064 21752 18070 21804
rect 19570 21752 19576 21804
rect 19628 21792 19634 21804
rect 21686 21792 21692 21804
rect 19628 21764 21456 21792
rect 21647 21764 21692 21792
rect 19628 21752 19634 21764
rect 14510 21724 14516 21736
rect 14068 21696 14516 21724
rect 13038 21616 13044 21668
rect 13096 21656 13102 21668
rect 14068 21665 14096 21696
rect 14510 21684 14516 21696
rect 14568 21684 14574 21736
rect 16810 21724 16816 21736
rect 14804 21696 16816 21724
rect 13225 21659 13283 21665
rect 13225 21656 13237 21659
rect 13096 21628 13237 21656
rect 13096 21616 13102 21628
rect 13225 21625 13237 21628
rect 13271 21625 13283 21659
rect 13225 21619 13283 21625
rect 14053 21659 14111 21665
rect 14053 21625 14065 21659
rect 14099 21625 14111 21659
rect 14053 21619 14111 21625
rect 12210 21548 12216 21600
rect 12268 21588 12274 21600
rect 12305 21591 12363 21597
rect 12305 21588 12317 21591
rect 12268 21560 12317 21588
rect 12268 21548 12274 21560
rect 12305 21557 12317 21560
rect 12351 21557 12363 21591
rect 12305 21551 12363 21557
rect 12581 21591 12639 21597
rect 12581 21557 12593 21591
rect 12627 21557 12639 21591
rect 12581 21551 12639 21557
rect 11842 21520 11848 21532
rect 11803 21492 11848 21520
rect 11842 21480 11848 21492
rect 11900 21480 11906 21532
rect 12596 21520 12624 21551
rect 12670 21548 12676 21600
rect 12728 21588 12734 21600
rect 13130 21588 13136 21600
rect 12728 21560 12773 21588
rect 13091 21560 13136 21588
rect 12728 21548 12734 21560
rect 13130 21548 13136 21560
rect 13188 21548 13194 21600
rect 14510 21588 14516 21600
rect 14471 21560 14516 21588
rect 14510 21548 14516 21560
rect 14568 21548 14574 21600
rect 14804 21597 14832 21696
rect 16810 21684 16816 21696
rect 16868 21684 16874 21736
rect 20030 21684 20036 21736
rect 20088 21724 20094 21736
rect 20493 21727 20551 21733
rect 20493 21724 20505 21727
rect 20088 21696 20505 21724
rect 20088 21684 20094 21696
rect 20493 21693 20505 21696
rect 20539 21693 20551 21727
rect 20493 21687 20551 21693
rect 20582 21684 20588 21736
rect 20640 21724 20646 21736
rect 21321 21727 21379 21733
rect 21321 21724 21333 21727
rect 20640 21696 21333 21724
rect 20640 21684 20646 21696
rect 21321 21693 21333 21696
rect 21367 21693 21379 21727
rect 21428 21724 21456 21764
rect 21686 21752 21692 21764
rect 21744 21752 21750 21804
rect 23802 21752 23808 21804
rect 23860 21792 23866 21804
rect 23943 21795 24001 21801
rect 23943 21792 23955 21795
rect 23860 21764 23955 21792
rect 23860 21752 23866 21764
rect 23943 21761 23955 21764
rect 23989 21761 24001 21795
rect 23943 21755 24001 21761
rect 22885 21727 22943 21733
rect 22885 21724 22897 21727
rect 21428 21696 22897 21724
rect 21321 21687 21379 21693
rect 22885 21693 22897 21696
rect 22931 21693 22943 21727
rect 22885 21687 22943 21693
rect 23158 21684 23164 21736
rect 23216 21724 23222 21736
rect 24081 21727 24139 21733
rect 24081 21724 24093 21727
rect 23216 21696 24093 21724
rect 23216 21684 23222 21696
rect 24081 21693 24093 21696
rect 24127 21693 24139 21727
rect 24081 21687 24139 21693
rect 15062 21616 15068 21668
rect 15120 21656 15126 21668
rect 15157 21659 15215 21665
rect 15157 21656 15169 21659
rect 15120 21628 15169 21656
rect 15120 21616 15126 21628
rect 15157 21625 15169 21628
rect 15203 21625 15215 21659
rect 15157 21619 15215 21625
rect 18742 21616 18748 21668
rect 18800 21656 18806 21668
rect 19018 21656 19024 21668
rect 18800 21628 19024 21656
rect 18800 21616 18806 21628
rect 19018 21616 19024 21628
rect 19076 21656 19082 21668
rect 19205 21659 19263 21665
rect 19205 21656 19217 21659
rect 19076 21628 19217 21656
rect 19076 21616 19082 21628
rect 19205 21625 19217 21628
rect 19251 21625 19263 21659
rect 19205 21619 19263 21625
rect 14789 21591 14847 21597
rect 14789 21557 14801 21591
rect 14835 21557 14847 21591
rect 14789 21551 14847 21557
rect 14973 21591 15031 21597
rect 14973 21557 14985 21591
rect 15019 21557 15031 21591
rect 15522 21588 15528 21600
rect 15483 21560 15528 21588
rect 14973 21551 15031 21557
rect 12762 21520 12768 21532
rect 12596 21492 12768 21520
rect 12762 21480 12768 21492
rect 12820 21480 12826 21532
rect 14988 21520 15016 21551
rect 15522 21548 15528 21560
rect 15580 21548 15586 21600
rect 16905 21591 16963 21597
rect 16905 21557 16917 21591
rect 16951 21588 16963 21591
rect 17822 21588 17828 21600
rect 16951 21560 17828 21588
rect 16951 21557 16963 21560
rect 16905 21551 16963 21557
rect 17822 21548 17828 21560
rect 17880 21588 17886 21600
rect 17917 21591 17975 21597
rect 17917 21588 17929 21591
rect 17880 21560 17929 21588
rect 17880 21548 17886 21560
rect 17917 21557 17929 21560
rect 17963 21557 17975 21591
rect 17917 21551 17975 21557
rect 18098 21548 18104 21600
rect 18156 21588 18162 21600
rect 19481 21591 19539 21597
rect 19481 21588 19493 21591
rect 18156 21560 19493 21588
rect 18156 21548 18162 21560
rect 19481 21557 19493 21560
rect 19527 21557 19539 21591
rect 20048 21588 20076 21684
rect 21413 21659 21471 21665
rect 21413 21625 21425 21659
rect 21459 21656 21471 21659
rect 21502 21656 21508 21668
rect 21459 21628 21508 21656
rect 21459 21625 21471 21628
rect 21413 21619 21471 21625
rect 21502 21616 21508 21628
rect 21560 21616 21566 21668
rect 22698 21616 22704 21668
rect 22756 21665 22762 21668
rect 22756 21659 22814 21665
rect 22756 21625 22768 21659
rect 22802 21625 22814 21659
rect 22756 21619 22814 21625
rect 22977 21659 23035 21665
rect 22977 21625 22989 21659
rect 23023 21656 23035 21659
rect 23434 21656 23440 21668
rect 23023 21628 23440 21656
rect 23023 21625 23035 21628
rect 22977 21619 23035 21625
rect 22756 21616 22762 21619
rect 23434 21616 23440 21628
rect 23492 21616 23498 21668
rect 24173 21659 24231 21665
rect 24173 21625 24185 21659
rect 24219 21625 24231 21659
rect 24173 21619 24231 21625
rect 28497 21659 28555 21665
rect 28497 21625 28509 21659
rect 28543 21656 28555 21659
rect 29690 21656 29696 21668
rect 28543 21628 29696 21656
rect 28543 21625 28555 21628
rect 28497 21619 28555 21625
rect 20398 21588 20404 21600
rect 19481 21551 19539 21557
rect 19588 21560 20076 21588
rect 20359 21560 20404 21588
rect 15430 21520 15436 21532
rect 14988 21492 15436 21520
rect 15430 21480 15436 21492
rect 15488 21480 15494 21532
rect 16721 21523 16779 21529
rect 16721 21489 16733 21523
rect 16767 21489 16779 21523
rect 17730 21520 17736 21532
rect 17691 21492 17736 21520
rect 16721 21483 16779 21489
rect 15246 21412 15252 21464
rect 15304 21452 15310 21464
rect 16736 21452 16764 21483
rect 17730 21480 17736 21492
rect 17788 21480 17794 21532
rect 19588 21529 19616 21560
rect 20398 21548 20404 21560
rect 20456 21548 20462 21600
rect 21134 21548 21140 21600
rect 21192 21597 21198 21600
rect 21192 21591 21250 21597
rect 21192 21557 21204 21591
rect 21238 21557 21250 21591
rect 22606 21588 22612 21600
rect 22567 21560 22612 21588
rect 21192 21551 21250 21557
rect 21192 21548 21198 21551
rect 22606 21548 22612 21560
rect 22664 21548 22670 21600
rect 24188 21588 24216 21619
rect 29690 21616 29696 21628
rect 29748 21616 29754 21668
rect 25550 21588 25556 21600
rect 22716 21560 24216 21588
rect 25511 21560 25556 21588
rect 19573 21523 19631 21529
rect 19573 21489 19585 21523
rect 19619 21489 19631 21523
rect 19573 21483 19631 21489
rect 19941 21523 19999 21529
rect 19941 21489 19953 21523
rect 19987 21520 19999 21523
rect 20214 21520 20220 21532
rect 19987 21492 20220 21520
rect 19987 21489 19999 21492
rect 19941 21483 19999 21489
rect 20214 21480 20220 21492
rect 20272 21480 20278 21532
rect 21045 21523 21103 21529
rect 21045 21489 21057 21523
rect 21091 21520 21103 21523
rect 21410 21520 21416 21532
rect 21091 21492 21416 21520
rect 21091 21489 21103 21492
rect 21045 21483 21103 21489
rect 21410 21480 21416 21492
rect 21468 21520 21474 21532
rect 22716 21520 22744 21560
rect 25550 21548 25556 21560
rect 25608 21548 25614 21600
rect 25642 21548 25648 21600
rect 25700 21588 25706 21600
rect 26378 21588 26384 21600
rect 25700 21560 26384 21588
rect 25700 21548 25706 21560
rect 26378 21548 26384 21560
rect 26436 21588 26442 21600
rect 26473 21591 26531 21597
rect 26473 21588 26485 21591
rect 26436 21560 26485 21588
rect 26436 21548 26442 21560
rect 26473 21557 26485 21560
rect 26519 21588 26531 21591
rect 27209 21591 27267 21597
rect 27209 21588 27221 21591
rect 26519 21560 27221 21588
rect 26519 21557 26531 21560
rect 26473 21551 26531 21557
rect 27209 21557 27221 21560
rect 27255 21557 27267 21591
rect 27942 21588 27948 21600
rect 27903 21560 27948 21588
rect 27209 21551 27267 21557
rect 27942 21548 27948 21560
rect 28000 21548 28006 21600
rect 28405 21591 28463 21597
rect 28405 21557 28417 21591
rect 28451 21588 28463 21591
rect 28770 21588 28776 21600
rect 28451 21560 28776 21588
rect 28451 21557 28463 21560
rect 28405 21551 28463 21557
rect 28770 21548 28776 21560
rect 28828 21548 28834 21600
rect 23342 21520 23348 21532
rect 21468 21492 22744 21520
rect 23303 21492 23348 21520
rect 21468 21480 21474 21492
rect 23342 21480 23348 21492
rect 23400 21480 23406 21532
rect 23805 21523 23863 21529
rect 23805 21489 23817 21523
rect 23851 21489 23863 21523
rect 23805 21483 23863 21489
rect 26289 21523 26347 21529
rect 26289 21489 26301 21523
rect 26335 21520 26347 21523
rect 26562 21520 26568 21532
rect 26335 21492 26568 21520
rect 26335 21489 26347 21492
rect 26289 21483 26347 21489
rect 15304 21424 16764 21452
rect 15304 21412 15310 21424
rect 17270 21412 17276 21464
rect 17328 21452 17334 21464
rect 18558 21452 18564 21464
rect 17328 21424 18564 21452
rect 17328 21412 17334 21424
rect 18558 21412 18564 21424
rect 18616 21452 18622 21464
rect 19389 21455 19447 21461
rect 19389 21452 19401 21455
rect 18616 21424 19401 21452
rect 18616 21412 18622 21424
rect 19389 21421 19401 21424
rect 19435 21421 19447 21455
rect 19389 21415 19447 21421
rect 22698 21412 22704 21464
rect 22756 21452 22762 21464
rect 23820 21452 23848 21483
rect 26562 21480 26568 21492
rect 26620 21520 26626 21532
rect 26746 21520 26752 21532
rect 26620 21492 26752 21520
rect 26620 21480 26626 21492
rect 26746 21480 26752 21492
rect 26804 21480 26810 21532
rect 26838 21480 26844 21532
rect 26896 21520 26902 21532
rect 27025 21523 27083 21529
rect 27025 21520 27037 21523
rect 26896 21492 27037 21520
rect 26896 21480 26902 21492
rect 27025 21489 27037 21492
rect 27071 21489 27083 21523
rect 27025 21483 27083 21489
rect 27390 21480 27396 21532
rect 27448 21520 27454 21532
rect 29049 21523 29107 21529
rect 29049 21520 29061 21523
rect 27448 21492 29061 21520
rect 27448 21480 27454 21492
rect 29049 21489 29061 21492
rect 29095 21489 29107 21523
rect 29049 21483 29107 21489
rect 29233 21523 29291 21529
rect 29233 21489 29245 21523
rect 29279 21520 29291 21523
rect 29598 21520 29604 21532
rect 29279 21492 29604 21520
rect 29279 21489 29291 21492
rect 29233 21483 29291 21489
rect 29598 21480 29604 21492
rect 29656 21480 29662 21532
rect 22756 21424 23848 21452
rect 22756 21412 22762 21424
rect 23894 21412 23900 21464
rect 23952 21452 23958 21464
rect 24449 21455 24507 21461
rect 24449 21452 24461 21455
rect 23952 21424 24461 21452
rect 23952 21412 23958 21424
rect 24449 21421 24461 21424
rect 24495 21421 24507 21455
rect 24449 21415 24507 21421
rect 11000 21362 30136 21384
rect 11000 21310 19142 21362
rect 19194 21310 19206 21362
rect 19258 21310 19270 21362
rect 19322 21310 19334 21362
rect 19386 21310 29142 21362
rect 29194 21310 29206 21362
rect 29258 21310 29270 21362
rect 29322 21310 29334 21362
rect 29386 21310 30136 21362
rect 11000 21288 30136 21310
rect 17086 21208 17092 21260
rect 17144 21208 17150 21260
rect 18561 21251 18619 21257
rect 18561 21217 18573 21251
rect 18607 21248 18619 21251
rect 19846 21248 19852 21260
rect 18607 21220 19852 21248
rect 18607 21217 18619 21220
rect 18561 21211 18619 21217
rect 19846 21208 19852 21220
rect 19904 21208 19910 21260
rect 24906 21248 24912 21260
rect 24464 21220 24912 21248
rect 11569 21183 11627 21189
rect 11569 21149 11581 21183
rect 11615 21180 11627 21183
rect 11842 21180 11848 21192
rect 11615 21152 11848 21180
rect 11615 21149 11627 21152
rect 11569 21143 11627 21149
rect 11842 21140 11848 21152
rect 11900 21140 11906 21192
rect 12026 21140 12032 21192
rect 12084 21140 12090 21192
rect 15157 21183 15215 21189
rect 15157 21180 15169 21183
rect 14436 21152 15169 21180
rect 11290 21112 11296 21124
rect 11251 21084 11296 21112
rect 11290 21072 11296 21084
rect 11348 21072 11354 21124
rect 13130 21072 13136 21124
rect 13188 21112 13194 21124
rect 14436 21121 14464 21152
rect 15157 21149 15169 21152
rect 15203 21180 15215 21183
rect 15246 21180 15252 21192
rect 15203 21152 15252 21180
rect 15203 21149 15215 21152
rect 15157 21143 15215 21149
rect 15246 21140 15252 21152
rect 15304 21140 15310 21192
rect 15522 21140 15528 21192
rect 15580 21180 15586 21192
rect 15709 21183 15767 21189
rect 15709 21180 15721 21183
rect 15580 21152 15721 21180
rect 15580 21140 15586 21152
rect 15709 21149 15721 21152
rect 15755 21180 15767 21183
rect 17104 21180 17132 21208
rect 15755 21152 17132 21180
rect 15755 21149 15767 21152
rect 15709 21143 15767 21149
rect 13317 21115 13375 21121
rect 13317 21112 13329 21115
rect 13188 21084 13329 21112
rect 13188 21072 13194 21084
rect 13317 21081 13329 21084
rect 13363 21112 13375 21115
rect 14421 21115 14479 21121
rect 14421 21112 14433 21115
rect 13363 21084 14433 21112
rect 13363 21081 13375 21084
rect 13317 21075 13375 21081
rect 14421 21081 14433 21084
rect 14467 21081 14479 21115
rect 15341 21115 15399 21121
rect 15341 21112 15353 21115
rect 14421 21075 14479 21081
rect 15264 21084 15353 21112
rect 15264 21056 15292 21084
rect 15341 21081 15353 21084
rect 15387 21081 15399 21115
rect 16258 21112 16264 21124
rect 16219 21084 16264 21112
rect 15341 21075 15399 21081
rect 16258 21072 16264 21084
rect 16316 21072 16322 21124
rect 16442 21112 16448 21124
rect 16403 21084 16448 21112
rect 16442 21072 16448 21084
rect 16500 21072 16506 21124
rect 16644 21121 16672 21152
rect 17822 21140 17828 21192
rect 17880 21180 17886 21192
rect 18653 21183 18711 21189
rect 18653 21180 18665 21183
rect 17880 21152 18665 21180
rect 17880 21140 17886 21152
rect 18653 21149 18665 21152
rect 18699 21149 18711 21183
rect 18653 21143 18711 21149
rect 19021 21183 19079 21189
rect 19021 21149 19033 21183
rect 19067 21180 19079 21183
rect 19570 21180 19576 21192
rect 19067 21152 19576 21180
rect 19067 21149 19079 21152
rect 19021 21143 19079 21149
rect 19570 21140 19576 21152
rect 19628 21140 19634 21192
rect 19662 21140 19668 21192
rect 19720 21180 19726 21192
rect 23713 21183 23771 21189
rect 19720 21152 22284 21180
rect 19720 21140 19726 21152
rect 16629 21115 16687 21121
rect 16629 21081 16641 21115
rect 16675 21081 16687 21115
rect 16902 21112 16908 21124
rect 16863 21084 16908 21112
rect 16629 21075 16687 21081
rect 16902 21072 16908 21084
rect 16960 21072 16966 21124
rect 17178 21121 17184 21124
rect 17158 21115 17184 21121
rect 17158 21081 17170 21115
rect 17158 21075 17184 21081
rect 17178 21072 17184 21075
rect 17236 21072 17242 21124
rect 18469 21115 18527 21121
rect 18469 21081 18481 21115
rect 18515 21112 18527 21115
rect 18558 21112 18564 21124
rect 18515 21084 18564 21112
rect 18515 21081 18527 21084
rect 18469 21075 18527 21081
rect 18558 21072 18564 21084
rect 18616 21072 18622 21124
rect 20214 21112 20220 21124
rect 20175 21084 20220 21112
rect 20214 21072 20220 21084
rect 20272 21072 20278 21124
rect 20398 21072 20404 21124
rect 20456 21112 20462 21124
rect 20585 21115 20643 21121
rect 20585 21112 20597 21115
rect 20456 21084 20597 21112
rect 20456 21072 20462 21084
rect 20585 21081 20597 21084
rect 20631 21081 20643 21115
rect 20585 21075 20643 21081
rect 20769 21115 20827 21121
rect 20769 21081 20781 21115
rect 20815 21112 20827 21115
rect 21502 21112 21508 21124
rect 20815 21084 21508 21112
rect 20815 21081 20827 21084
rect 20769 21075 20827 21081
rect 21502 21072 21508 21084
rect 21560 21072 21566 21124
rect 21870 21112 21876 21124
rect 21831 21084 21876 21112
rect 21870 21072 21876 21084
rect 21928 21072 21934 21124
rect 22256 21121 22284 21152
rect 23713 21149 23725 21183
rect 23759 21180 23771 21183
rect 23986 21180 23992 21192
rect 23759 21152 23992 21180
rect 23759 21149 23771 21152
rect 23713 21143 23771 21149
rect 23986 21140 23992 21152
rect 24044 21140 24050 21192
rect 22241 21115 22299 21121
rect 22241 21081 22253 21115
rect 22287 21081 22299 21115
rect 22241 21075 22299 21081
rect 23342 21072 23348 21124
rect 23400 21112 23406 21124
rect 24464 21121 24492 21220
rect 24906 21208 24912 21220
rect 24964 21208 24970 21260
rect 25458 21180 25464 21192
rect 24556 21152 25464 21180
rect 24556 21121 24584 21152
rect 25458 21140 25464 21152
rect 25516 21140 25522 21192
rect 25550 21140 25556 21192
rect 25608 21180 25614 21192
rect 25608 21152 26700 21180
rect 25608 21140 25614 21152
rect 23621 21115 23679 21121
rect 23621 21112 23633 21115
rect 23400 21084 23633 21112
rect 23400 21072 23406 21084
rect 23621 21081 23633 21084
rect 23667 21081 23679 21115
rect 23621 21075 23679 21081
rect 24449 21115 24507 21121
rect 24449 21081 24461 21115
rect 24495 21081 24507 21115
rect 24449 21075 24507 21081
rect 24541 21115 24599 21121
rect 24541 21081 24553 21115
rect 24587 21081 24599 21115
rect 24541 21075 24599 21081
rect 25182 21072 25188 21124
rect 25240 21112 25246 21124
rect 26672 21121 26700 21152
rect 26746 21140 26752 21192
rect 26804 21180 26810 21192
rect 27117 21183 27175 21189
rect 27117 21180 27129 21183
rect 26804 21152 27129 21180
rect 26804 21140 26810 21152
rect 27117 21149 27129 21152
rect 27163 21149 27175 21183
rect 27117 21143 27175 21149
rect 29417 21183 29475 21189
rect 29417 21149 29429 21183
rect 29463 21180 29475 21183
rect 29506 21180 29512 21192
rect 29463 21152 29512 21180
rect 29463 21149 29475 21152
rect 29417 21143 29475 21149
rect 29506 21140 29512 21152
rect 29564 21140 29570 21192
rect 25645 21115 25703 21121
rect 25645 21112 25657 21115
rect 25240 21084 25657 21112
rect 25240 21072 25246 21084
rect 25645 21081 25657 21084
rect 25691 21081 25703 21115
rect 25645 21075 25703 21081
rect 26657 21115 26715 21121
rect 26657 21081 26669 21115
rect 26703 21081 26715 21115
rect 26657 21075 26715 21081
rect 27853 21115 27911 21121
rect 27853 21081 27865 21115
rect 27899 21112 27911 21115
rect 28586 21112 28592 21124
rect 27899 21084 28592 21112
rect 27899 21081 27911 21084
rect 27853 21075 27911 21081
rect 28586 21072 28592 21084
rect 28644 21072 28650 21124
rect 29141 21115 29199 21121
rect 29141 21081 29153 21115
rect 29187 21112 29199 21115
rect 29598 21112 29604 21124
rect 29187 21084 29604 21112
rect 29187 21081 29199 21084
rect 29141 21075 29199 21081
rect 29598 21072 29604 21084
rect 29656 21072 29662 21124
rect 15246 21004 15252 21056
rect 15304 21004 15310 21056
rect 17733 21047 17791 21053
rect 17733 21013 17745 21047
rect 17779 21044 17791 21047
rect 18098 21044 18104 21056
rect 17779 21016 18104 21044
rect 17779 21013 17791 21016
rect 17733 21007 17791 21013
rect 18098 21004 18104 21016
rect 18156 21004 18162 21056
rect 18285 21047 18343 21053
rect 18285 21013 18297 21047
rect 18331 21044 18343 21047
rect 19018 21044 19024 21056
rect 18331 21016 19024 21044
rect 18331 21013 18343 21016
rect 18285 21007 18343 21013
rect 19018 21004 19024 21016
rect 19076 21004 19082 21056
rect 20122 21044 20128 21056
rect 20083 21016 20128 21044
rect 20122 21004 20128 21016
rect 20180 21044 20186 21056
rect 21134 21044 21140 21056
rect 20180 21016 21140 21044
rect 20180 21004 20186 21016
rect 21134 21004 21140 21016
rect 21192 21004 21198 21056
rect 21686 21044 21692 21056
rect 21647 21016 21692 21044
rect 21686 21004 21692 21016
rect 21744 21044 21750 21056
rect 21962 21044 21968 21056
rect 21744 21016 21968 21044
rect 21744 21004 21750 21016
rect 21962 21004 21968 21016
rect 22020 21004 22026 21056
rect 22146 21044 22152 21056
rect 22107 21016 22152 21044
rect 22146 21004 22152 21016
rect 22204 21004 22210 21056
rect 26197 21047 26255 21053
rect 26197 21044 26209 21047
rect 24648 21016 26209 21044
rect 17178 20936 17184 20988
rect 17236 20976 17242 20988
rect 17546 20976 17552 20988
rect 17236 20948 17552 20976
rect 17236 20936 17242 20948
rect 17546 20936 17552 20948
rect 17604 20976 17610 20988
rect 20398 20976 20404 20988
rect 17604 20948 20404 20976
rect 17604 20936 17610 20948
rect 20398 20936 20404 20948
rect 20456 20936 20462 20988
rect 21152 20976 21180 21004
rect 21778 20976 21784 20988
rect 21152 20948 21784 20976
rect 21778 20936 21784 20948
rect 21836 20936 21842 20988
rect 23526 20936 23532 20988
rect 23584 20976 23590 20988
rect 24648 20976 24676 21016
rect 26197 21013 26209 21016
rect 26243 21013 26255 21047
rect 27206 21044 27212 21056
rect 27167 21016 27212 21044
rect 26197 21007 26255 21013
rect 27206 21004 27212 21016
rect 27264 21004 27270 21056
rect 23584 20948 24676 20976
rect 26105 20979 26163 20985
rect 23584 20936 23590 20948
rect 26105 20945 26117 20979
rect 26151 20976 26163 20979
rect 26838 20976 26844 20988
rect 26151 20948 26844 20976
rect 26151 20945 26163 20948
rect 26105 20939 26163 20945
rect 26838 20936 26844 20948
rect 26896 20936 26902 20988
rect 13866 20868 13872 20920
rect 13924 20908 13930 20920
rect 14513 20911 14571 20917
rect 14513 20908 14525 20911
rect 13924 20880 14525 20908
rect 13924 20868 13930 20880
rect 14513 20877 14525 20880
rect 14559 20908 14571 20911
rect 17730 20908 17736 20920
rect 14559 20880 17736 20908
rect 14559 20877 14571 20880
rect 14513 20871 14571 20877
rect 17730 20868 17736 20880
rect 17788 20868 17794 20920
rect 19665 20911 19723 20917
rect 19665 20877 19677 20911
rect 19711 20908 19723 20911
rect 19938 20908 19944 20920
rect 19711 20880 19944 20908
rect 19711 20877 19723 20880
rect 19665 20871 19723 20877
rect 19938 20868 19944 20880
rect 19996 20868 20002 20920
rect 21505 20911 21563 20917
rect 21505 20877 21517 20911
rect 21551 20908 21563 20911
rect 24630 20908 24636 20920
rect 21551 20880 24636 20908
rect 21551 20877 21563 20880
rect 21505 20871 21563 20877
rect 24630 20868 24636 20880
rect 24688 20868 24694 20920
rect 11000 20818 30136 20840
rect 11000 20766 14142 20818
rect 14194 20766 14206 20818
rect 14258 20766 14270 20818
rect 14322 20766 14334 20818
rect 14386 20766 24142 20818
rect 24194 20766 24206 20818
rect 24258 20766 24270 20818
rect 24322 20766 24334 20818
rect 24386 20766 30136 20818
rect 11000 20744 30136 20766
rect 15430 20704 15436 20716
rect 15391 20676 15436 20704
rect 15430 20664 15436 20676
rect 15488 20664 15494 20716
rect 19205 20707 19263 20713
rect 19205 20673 19217 20707
rect 19251 20704 19263 20707
rect 20122 20704 20128 20716
rect 19251 20676 20128 20704
rect 19251 20673 19263 20676
rect 19205 20667 19263 20673
rect 20122 20664 20128 20676
rect 20180 20664 20186 20716
rect 20585 20707 20643 20713
rect 20585 20673 20597 20707
rect 20631 20704 20643 20707
rect 21870 20704 21876 20716
rect 20631 20676 21876 20704
rect 20631 20673 20643 20676
rect 20585 20667 20643 20673
rect 21870 20664 21876 20676
rect 21928 20664 21934 20716
rect 22609 20707 22667 20713
rect 22609 20673 22621 20707
rect 22655 20704 22667 20707
rect 22698 20704 22704 20716
rect 22655 20676 22704 20704
rect 22655 20673 22667 20676
rect 22609 20667 22667 20673
rect 22698 20664 22704 20676
rect 22756 20664 22762 20716
rect 23989 20707 24047 20713
rect 23989 20673 24001 20707
rect 24035 20704 24047 20707
rect 27206 20704 27212 20716
rect 24035 20676 27212 20704
rect 24035 20673 24047 20676
rect 23989 20667 24047 20673
rect 27206 20664 27212 20676
rect 27264 20664 27270 20716
rect 14510 20636 14516 20648
rect 13240 20608 14516 20636
rect 12210 20568 12216 20580
rect 12171 20540 12216 20568
rect 12210 20528 12216 20540
rect 12268 20528 12274 20580
rect 13130 20568 13136 20580
rect 13091 20540 13136 20568
rect 13130 20528 13136 20540
rect 13188 20528 13194 20580
rect 11845 20503 11903 20509
rect 11845 20469 11857 20503
rect 11891 20500 11903 20503
rect 12946 20500 12952 20512
rect 11891 20472 12952 20500
rect 11891 20469 11903 20472
rect 11845 20463 11903 20469
rect 12946 20460 12952 20472
rect 13004 20500 13010 20512
rect 13240 20500 13268 20608
rect 14510 20596 14516 20608
rect 14568 20596 14574 20648
rect 15706 20596 15712 20648
rect 15764 20636 15770 20648
rect 19662 20636 19668 20648
rect 15764 20608 19668 20636
rect 15764 20596 15770 20608
rect 19662 20596 19668 20608
rect 19720 20596 19726 20648
rect 20217 20639 20275 20645
rect 20217 20605 20229 20639
rect 20263 20636 20275 20639
rect 20398 20636 20404 20648
rect 20263 20608 20404 20636
rect 20263 20605 20275 20608
rect 20217 20599 20275 20605
rect 20398 20596 20404 20608
rect 20456 20636 20462 20648
rect 23434 20636 23440 20648
rect 20456 20608 23440 20636
rect 20456 20596 20462 20608
rect 23434 20596 23440 20608
rect 23492 20596 23498 20648
rect 24725 20639 24783 20645
rect 24725 20605 24737 20639
rect 24771 20636 24783 20639
rect 25550 20636 25556 20648
rect 24771 20608 25556 20636
rect 24771 20605 24783 20608
rect 24725 20599 24783 20605
rect 25550 20596 25556 20608
rect 25608 20596 25614 20648
rect 15062 20568 15068 20580
rect 13332 20540 15068 20568
rect 13332 20509 13360 20540
rect 15062 20528 15068 20540
rect 15120 20528 15126 20580
rect 18006 20568 18012 20580
rect 17932 20540 18012 20568
rect 13004 20472 13268 20500
rect 13317 20503 13375 20509
rect 13004 20460 13010 20472
rect 13317 20469 13329 20503
rect 13363 20469 13375 20503
rect 13682 20500 13688 20512
rect 13643 20472 13688 20500
rect 13317 20463 13375 20469
rect 13682 20460 13688 20472
rect 13740 20460 13746 20512
rect 13866 20500 13872 20512
rect 13827 20472 13872 20500
rect 13866 20460 13872 20472
rect 13924 20460 13930 20512
rect 14513 20503 14571 20509
rect 14513 20469 14525 20503
rect 14559 20500 14571 20503
rect 14602 20500 14608 20512
rect 14559 20472 14608 20500
rect 14559 20469 14571 20472
rect 14513 20463 14571 20469
rect 14602 20460 14608 20472
rect 14660 20500 14666 20512
rect 17932 20509 17960 20540
rect 18006 20528 18012 20540
rect 18064 20528 18070 20580
rect 18377 20571 18435 20577
rect 18377 20537 18389 20571
rect 18423 20568 18435 20571
rect 20088 20571 20146 20577
rect 20088 20568 20100 20571
rect 18423 20540 20100 20568
rect 18423 20537 18435 20540
rect 18377 20531 18435 20537
rect 20088 20537 20100 20540
rect 20134 20537 20146 20571
rect 20088 20531 20146 20537
rect 20309 20571 20367 20577
rect 20309 20537 20321 20571
rect 20355 20568 20367 20571
rect 20582 20568 20588 20580
rect 20355 20540 20588 20568
rect 20355 20537 20367 20540
rect 20309 20531 20367 20537
rect 20582 20528 20588 20540
rect 20640 20528 20646 20580
rect 21594 20528 21600 20580
rect 21652 20568 21658 20580
rect 21689 20571 21747 20577
rect 21689 20568 21701 20571
rect 21652 20540 21701 20568
rect 21652 20528 21658 20540
rect 21689 20537 21701 20540
rect 21735 20537 21747 20571
rect 25642 20568 25648 20580
rect 21689 20531 21747 20537
rect 22256 20540 22560 20568
rect 15341 20503 15399 20509
rect 15341 20500 15353 20503
rect 14660 20472 15353 20500
rect 14660 20460 14666 20472
rect 15341 20469 15353 20472
rect 15387 20469 15399 20503
rect 15341 20463 15399 20469
rect 17917 20503 17975 20509
rect 17917 20469 17929 20503
rect 17963 20469 17975 20503
rect 18098 20500 18104 20512
rect 18059 20472 18104 20500
rect 17917 20463 17975 20469
rect 18098 20460 18104 20472
rect 18156 20460 18162 20512
rect 19113 20503 19171 20509
rect 19113 20469 19125 20503
rect 19159 20469 19171 20503
rect 19938 20500 19944 20512
rect 19899 20472 19944 20500
rect 19113 20463 19171 20469
rect 11661 20435 11719 20441
rect 11661 20401 11673 20435
rect 11707 20401 11719 20435
rect 11661 20395 11719 20401
rect 14329 20435 14387 20441
rect 14329 20401 14341 20435
rect 14375 20432 14387 20435
rect 14418 20432 14424 20444
rect 14375 20404 14424 20432
rect 14375 20401 14387 20404
rect 14329 20395 14387 20401
rect 11676 20364 11704 20395
rect 14418 20392 14424 20404
rect 14476 20392 14482 20444
rect 14878 20432 14884 20444
rect 14839 20404 14884 20432
rect 14878 20392 14884 20404
rect 14936 20392 14942 20444
rect 18926 20432 18932 20444
rect 18887 20404 18932 20432
rect 18926 20392 18932 20404
rect 18984 20392 18990 20444
rect 19128 20432 19156 20463
rect 19938 20460 19944 20472
rect 19996 20460 20002 20512
rect 20214 20460 20220 20512
rect 20272 20500 20278 20512
rect 21137 20503 21195 20509
rect 21137 20500 21149 20503
rect 20272 20472 21149 20500
rect 20272 20460 20278 20472
rect 21137 20469 21149 20472
rect 21183 20469 21195 20503
rect 21137 20463 21195 20469
rect 21229 20503 21287 20509
rect 21229 20469 21241 20503
rect 21275 20500 21287 20503
rect 21502 20500 21508 20512
rect 21275 20472 21508 20500
rect 21275 20469 21287 20472
rect 21229 20463 21287 20469
rect 21502 20460 21508 20472
rect 21560 20460 21566 20512
rect 21778 20460 21784 20512
rect 21836 20500 21842 20512
rect 22256 20500 22284 20540
rect 21836 20472 22284 20500
rect 21836 20460 21842 20472
rect 22330 20460 22336 20512
rect 22388 20500 22394 20512
rect 22532 20509 22560 20540
rect 24188 20540 25648 20568
rect 24188 20509 24216 20540
rect 25642 20528 25648 20540
rect 25700 20528 25706 20580
rect 26838 20568 26844 20580
rect 26799 20540 26844 20568
rect 26838 20528 26844 20540
rect 26896 20528 26902 20580
rect 22517 20503 22575 20509
rect 22388 20472 22433 20500
rect 22388 20460 22394 20472
rect 22517 20469 22529 20503
rect 22563 20469 22575 20503
rect 22517 20463 22575 20469
rect 24173 20503 24231 20509
rect 24173 20469 24185 20503
rect 24219 20469 24231 20503
rect 24630 20500 24636 20512
rect 24591 20472 24636 20500
rect 24173 20463 24231 20469
rect 24630 20460 24636 20472
rect 24688 20460 24694 20512
rect 25182 20460 25188 20512
rect 25240 20500 25246 20512
rect 25277 20503 25335 20509
rect 25277 20500 25289 20503
rect 25240 20472 25289 20500
rect 25240 20460 25246 20472
rect 25277 20469 25289 20472
rect 25323 20469 25335 20503
rect 26470 20500 26476 20512
rect 26431 20472 26476 20500
rect 25277 20463 25335 20469
rect 26470 20460 26476 20472
rect 26528 20460 26534 20512
rect 27942 20500 27948 20512
rect 27903 20472 27948 20500
rect 27942 20460 27948 20472
rect 28000 20460 28006 20512
rect 19662 20432 19668 20444
rect 19128 20404 19668 20432
rect 19662 20392 19668 20404
rect 19720 20432 19726 20444
rect 24538 20432 24544 20444
rect 19720 20404 24544 20432
rect 19720 20392 19726 20404
rect 24538 20392 24544 20404
rect 24596 20392 24602 20444
rect 28681 20435 28739 20441
rect 28681 20401 28693 20435
rect 28727 20432 28739 20435
rect 28770 20432 28776 20444
rect 28727 20404 28776 20432
rect 28727 20401 28739 20404
rect 28681 20395 28739 20401
rect 28770 20392 28776 20404
rect 28828 20392 28834 20444
rect 28865 20435 28923 20441
rect 28865 20401 28877 20435
rect 28911 20432 28923 20435
rect 29598 20432 29604 20444
rect 28911 20404 29604 20432
rect 28911 20401 28923 20404
rect 28865 20395 28923 20401
rect 29598 20392 29604 20404
rect 29656 20392 29662 20444
rect 12670 20364 12676 20376
rect 11676 20336 12676 20364
rect 12670 20324 12676 20336
rect 12728 20364 12734 20376
rect 12765 20367 12823 20373
rect 12765 20364 12777 20367
rect 12728 20336 12777 20364
rect 12728 20324 12734 20336
rect 12765 20333 12777 20336
rect 12811 20333 12823 20367
rect 12765 20327 12823 20333
rect 19754 20324 19760 20376
rect 19812 20364 19818 20376
rect 20214 20364 20220 20376
rect 19812 20336 20220 20364
rect 19812 20324 19818 20336
rect 20214 20324 20220 20336
rect 20272 20324 20278 20376
rect 11000 20274 30136 20296
rect 11000 20222 19142 20274
rect 19194 20222 19206 20274
rect 19258 20222 19270 20274
rect 19322 20222 19334 20274
rect 19386 20222 29142 20274
rect 29194 20222 29206 20274
rect 29258 20222 29270 20274
rect 29322 20222 29334 20274
rect 29386 20222 30136 20274
rect 11000 20200 30136 20222
rect 16442 20120 16448 20172
rect 16500 20160 16506 20172
rect 18190 20160 18196 20172
rect 16500 20132 18196 20160
rect 16500 20120 16506 20132
rect 18190 20120 18196 20132
rect 18248 20160 18254 20172
rect 18377 20163 18435 20169
rect 18377 20160 18389 20163
rect 18248 20132 18389 20160
rect 18248 20120 18254 20132
rect 18377 20129 18389 20132
rect 18423 20129 18435 20163
rect 18377 20123 18435 20129
rect 18469 20163 18527 20169
rect 18469 20129 18481 20163
rect 18515 20160 18527 20163
rect 19846 20160 19852 20172
rect 18515 20132 19852 20160
rect 18515 20129 18527 20132
rect 18469 20123 18527 20129
rect 19220 20104 19248 20132
rect 15798 20092 15804 20104
rect 15759 20064 15804 20092
rect 15798 20052 15804 20064
rect 15856 20052 15862 20104
rect 16994 20092 17000 20104
rect 16907 20064 17000 20092
rect 16994 20052 17000 20064
rect 17052 20092 17058 20104
rect 17546 20092 17552 20104
rect 17052 20064 17316 20092
rect 17507 20064 17552 20092
rect 17052 20052 17058 20064
rect 11658 20024 11664 20036
rect 11619 19996 11664 20024
rect 11658 19984 11664 19996
rect 11716 19984 11722 20036
rect 12670 19984 12676 20036
rect 12728 20024 12734 20036
rect 12946 20024 12952 20036
rect 12728 19996 12773 20024
rect 12907 19996 12952 20024
rect 12728 19984 12734 19996
rect 12946 19984 12952 19996
rect 13004 19984 13010 20036
rect 14237 20027 14295 20033
rect 14237 19993 14249 20027
rect 14283 20024 14295 20027
rect 14418 20024 14424 20036
rect 14283 19996 14424 20024
rect 14283 19993 14295 19996
rect 14237 19987 14295 19993
rect 14418 19984 14424 19996
rect 14476 19984 14482 20036
rect 14602 20024 14608 20036
rect 14563 19996 14608 20024
rect 14602 19984 14608 19996
rect 14660 19984 14666 20036
rect 17178 20024 17184 20036
rect 17139 19996 17184 20024
rect 17178 19984 17184 19996
rect 17236 19984 17242 20036
rect 17288 20024 17316 20064
rect 17546 20052 17552 20064
rect 17604 20052 17610 20104
rect 17822 20052 17828 20104
rect 17880 20092 17886 20104
rect 18561 20095 18619 20101
rect 18561 20092 18573 20095
rect 17880 20064 18573 20092
rect 17880 20052 17886 20064
rect 18561 20061 18573 20064
rect 18607 20061 18619 20095
rect 18926 20092 18932 20104
rect 18887 20064 18932 20092
rect 18561 20055 18619 20061
rect 18926 20052 18932 20064
rect 18984 20052 18990 20104
rect 19202 20052 19208 20104
rect 19260 20052 19266 20104
rect 19588 20101 19616 20132
rect 19846 20120 19852 20132
rect 19904 20120 19910 20172
rect 21413 20163 21471 20169
rect 21413 20129 21425 20163
rect 21459 20160 21471 20163
rect 27209 20163 27267 20169
rect 21459 20132 27160 20160
rect 21459 20129 21471 20132
rect 21413 20123 21471 20129
rect 19573 20095 19631 20101
rect 19573 20061 19585 20095
rect 19619 20061 19631 20095
rect 19754 20092 19760 20104
rect 19715 20064 19760 20092
rect 19573 20055 19631 20061
rect 19754 20052 19760 20064
rect 19812 20052 19818 20104
rect 19938 20092 19944 20104
rect 19899 20064 19944 20092
rect 19938 20052 19944 20064
rect 19996 20052 20002 20104
rect 21502 20052 21508 20104
rect 21560 20092 21566 20104
rect 24081 20095 24139 20101
rect 24081 20092 24093 20095
rect 21560 20064 24093 20092
rect 21560 20052 21566 20064
rect 24081 20061 24093 20064
rect 24127 20061 24139 20095
rect 24081 20055 24139 20061
rect 26381 20095 26439 20101
rect 26381 20061 26393 20095
rect 26427 20092 26439 20095
rect 26470 20092 26476 20104
rect 26427 20064 26476 20092
rect 26427 20061 26439 20064
rect 26381 20055 26439 20061
rect 26470 20052 26476 20064
rect 26528 20052 26534 20104
rect 17730 20024 17736 20036
rect 17288 19996 17736 20024
rect 17730 19984 17736 19996
rect 17788 19984 17794 20036
rect 19849 20027 19907 20033
rect 19849 19993 19861 20027
rect 19895 19993 19907 20027
rect 19849 19987 19907 19993
rect 12762 19956 12768 19968
rect 12723 19928 12768 19956
rect 12762 19916 12768 19928
rect 12820 19916 12826 19968
rect 14329 19959 14387 19965
rect 14329 19925 14341 19959
rect 14375 19956 14387 19959
rect 14694 19956 14700 19968
rect 14375 19928 14700 19956
rect 14375 19925 14387 19928
rect 14329 19919 14387 19925
rect 14694 19916 14700 19928
rect 14752 19916 14758 19968
rect 16169 19959 16227 19965
rect 16169 19925 16181 19959
rect 16215 19956 16227 19959
rect 18006 19956 18012 19968
rect 16215 19928 18012 19956
rect 16215 19925 16227 19928
rect 16169 19919 16227 19925
rect 18006 19916 18012 19928
rect 18064 19916 18070 19968
rect 18193 19959 18251 19965
rect 18193 19925 18205 19959
rect 18239 19925 18251 19959
rect 19864 19956 19892 19987
rect 21042 19984 21048 20036
rect 21100 20024 21106 20036
rect 21781 20027 21839 20033
rect 21781 20024 21793 20027
rect 21100 19996 21793 20024
rect 21100 19984 21106 19996
rect 21781 19993 21793 19996
rect 21827 19993 21839 20027
rect 22146 20024 22152 20036
rect 22107 19996 22152 20024
rect 21781 19987 21839 19993
rect 22146 19984 22152 19996
rect 22204 19984 22210 20036
rect 22238 19984 22244 20036
rect 22296 20024 22302 20036
rect 23345 20027 23403 20033
rect 22296 19996 22341 20024
rect 22296 19984 22302 19996
rect 23345 19993 23357 20027
rect 23391 19993 23403 20027
rect 23526 20024 23532 20036
rect 23487 19996 23532 20024
rect 23345 19987 23403 19993
rect 20214 19956 20220 19968
rect 18193 19919 18251 19925
rect 18944 19928 20220 19956
rect 11753 19891 11811 19897
rect 11753 19857 11765 19891
rect 11799 19888 11811 19891
rect 15706 19888 15712 19900
rect 11799 19860 15712 19888
rect 11799 19857 11811 19860
rect 11753 19851 11811 19857
rect 15706 19848 15712 19860
rect 15764 19848 15770 19900
rect 15890 19848 15896 19900
rect 15948 19897 15954 19900
rect 15948 19891 15997 19897
rect 15948 19857 15951 19891
rect 15985 19857 15997 19891
rect 15948 19851 15997 19857
rect 15948 19848 15954 19851
rect 16258 19848 16264 19900
rect 16316 19888 16322 19900
rect 18208 19888 18236 19919
rect 18944 19900 18972 19928
rect 20214 19916 20220 19928
rect 20272 19916 20278 19968
rect 20309 19959 20367 19965
rect 20309 19925 20321 19959
rect 20355 19956 20367 19959
rect 20398 19956 20404 19968
rect 20355 19928 20404 19956
rect 20355 19925 20367 19928
rect 20309 19919 20367 19925
rect 20398 19916 20404 19928
rect 20456 19916 20462 19968
rect 21686 19956 21692 19968
rect 21647 19928 21692 19956
rect 21686 19916 21692 19928
rect 21744 19916 21750 19968
rect 23360 19956 23388 19987
rect 23526 19984 23532 19996
rect 23584 19984 23590 20036
rect 23986 20024 23992 20036
rect 23899 19996 23992 20024
rect 23986 19984 23992 19996
rect 24044 20024 24050 20036
rect 24630 20024 24636 20036
rect 24044 19996 24636 20024
rect 24044 19984 24050 19996
rect 24630 19984 24636 19996
rect 24688 19984 24694 20036
rect 25461 20027 25519 20033
rect 25461 19993 25473 20027
rect 25507 20024 25519 20027
rect 25550 20024 25556 20036
rect 25507 19996 25556 20024
rect 25507 19993 25519 19996
rect 25461 19987 25519 19993
rect 25550 19984 25556 19996
rect 25608 19984 25614 20036
rect 27132 20033 27160 20132
rect 27209 20129 27221 20163
rect 27255 20160 27267 20163
rect 27942 20160 27948 20172
rect 27255 20132 27948 20160
rect 27255 20129 27267 20132
rect 27209 20123 27267 20129
rect 27942 20120 27948 20132
rect 28000 20120 28006 20172
rect 29049 20095 29107 20101
rect 29049 20061 29061 20095
rect 29095 20092 29107 20095
rect 29506 20092 29512 20104
rect 29095 20064 29512 20092
rect 29095 20061 29107 20064
rect 29049 20055 29107 20061
rect 29506 20052 29512 20064
rect 29564 20052 29570 20104
rect 26105 20027 26163 20033
rect 26105 19993 26117 20027
rect 26151 19993 26163 20027
rect 26105 19987 26163 19993
rect 27117 20027 27175 20033
rect 27117 19993 27129 20027
rect 27163 19993 27175 20027
rect 27117 19987 27175 19993
rect 26010 19956 26016 19968
rect 23360 19928 26016 19956
rect 26010 19916 26016 19928
rect 26068 19956 26074 19968
rect 26120 19956 26148 19987
rect 27298 19984 27304 20036
rect 27356 20024 27362 20036
rect 27945 20027 28003 20033
rect 27945 20024 27957 20027
rect 27356 19996 27957 20024
rect 27356 19984 27362 19996
rect 27945 19993 27957 19996
rect 27991 19993 28003 20027
rect 28586 20024 28592 20036
rect 28547 19996 28592 20024
rect 27945 19987 28003 19993
rect 28586 19984 28592 19996
rect 28644 19984 28650 20036
rect 26068 19928 26148 19956
rect 26068 19916 26074 19928
rect 28862 19916 28868 19968
rect 28920 19956 28926 19968
rect 29141 19959 29199 19965
rect 29141 19956 29153 19959
rect 28920 19928 29153 19956
rect 28920 19916 28926 19928
rect 29141 19925 29153 19928
rect 29187 19925 29199 19959
rect 29141 19919 29199 19925
rect 18926 19888 18932 19900
rect 16316 19860 18932 19888
rect 16316 19848 16322 19860
rect 18926 19848 18932 19860
rect 18984 19848 18990 19900
rect 24906 19848 24912 19900
rect 24964 19888 24970 19900
rect 26194 19888 26200 19900
rect 24964 19860 26200 19888
rect 24964 19848 24970 19860
rect 26194 19848 26200 19860
rect 26252 19848 26258 19900
rect 16074 19820 16080 19832
rect 16035 19792 16080 19820
rect 16074 19780 16080 19792
rect 16132 19780 16138 19832
rect 16445 19823 16503 19829
rect 16445 19789 16457 19823
rect 16491 19820 16503 19823
rect 16718 19820 16724 19832
rect 16491 19792 16724 19820
rect 16491 19789 16503 19792
rect 16445 19783 16503 19789
rect 16718 19780 16724 19792
rect 16776 19780 16782 19832
rect 27758 19820 27764 19832
rect 27719 19792 27764 19820
rect 27758 19780 27764 19792
rect 27816 19780 27822 19832
rect 11000 19730 30136 19752
rect 11000 19678 14142 19730
rect 14194 19678 14206 19730
rect 14258 19678 14270 19730
rect 14322 19678 14334 19730
rect 14386 19678 24142 19730
rect 24194 19678 24206 19730
rect 24258 19678 24270 19730
rect 24322 19678 24334 19730
rect 24386 19678 30136 19730
rect 11000 19656 30136 19678
rect 24556 19588 26056 19616
rect 17178 19548 17184 19560
rect 15448 19520 17184 19548
rect 12762 19440 12768 19492
rect 12820 19480 12826 19492
rect 13317 19483 13375 19489
rect 13317 19480 13329 19483
rect 12820 19452 13329 19480
rect 12820 19440 12826 19452
rect 13317 19449 13329 19452
rect 13363 19449 13375 19483
rect 13317 19443 13375 19449
rect 13777 19483 13835 19489
rect 13777 19449 13789 19483
rect 13823 19480 13835 19483
rect 13866 19480 13872 19492
rect 13823 19452 13872 19480
rect 13823 19449 13835 19452
rect 13777 19443 13835 19449
rect 13866 19440 13872 19452
rect 13924 19440 13930 19492
rect 14602 19440 14608 19492
rect 14660 19480 14666 19492
rect 14697 19483 14755 19489
rect 14697 19480 14709 19483
rect 14660 19452 14709 19480
rect 14660 19440 14666 19452
rect 14697 19449 14709 19452
rect 14743 19449 14755 19483
rect 14697 19443 14755 19449
rect 15246 19440 15252 19492
rect 15304 19480 15310 19492
rect 15448 19489 15476 19520
rect 17178 19508 17184 19520
rect 17236 19508 17242 19560
rect 19938 19508 19944 19560
rect 19996 19548 20002 19560
rect 20217 19551 20275 19557
rect 20217 19548 20229 19551
rect 19996 19520 20229 19548
rect 19996 19508 20002 19520
rect 20217 19517 20229 19520
rect 20263 19517 20275 19551
rect 24262 19548 24268 19560
rect 24223 19520 24268 19548
rect 20217 19511 20275 19517
rect 24262 19508 24268 19520
rect 24320 19508 24326 19560
rect 15433 19483 15491 19489
rect 15433 19480 15445 19483
rect 15304 19452 15445 19480
rect 15304 19440 15310 19452
rect 15433 19449 15445 19452
rect 15479 19449 15491 19483
rect 17822 19480 17828 19492
rect 15433 19443 15491 19449
rect 16092 19452 17828 19480
rect 16092 19424 16120 19452
rect 17822 19440 17828 19452
rect 17880 19440 17886 19492
rect 18926 19480 18932 19492
rect 18887 19452 18932 19480
rect 18926 19440 18932 19452
rect 18984 19440 18990 19492
rect 19662 19480 19668 19492
rect 19623 19452 19668 19480
rect 19662 19440 19668 19452
rect 19720 19440 19726 19492
rect 20861 19483 20919 19489
rect 20861 19449 20873 19483
rect 20907 19480 20919 19483
rect 23986 19480 23992 19492
rect 20907 19452 23992 19480
rect 20907 19449 20919 19452
rect 20861 19443 20919 19449
rect 23986 19440 23992 19452
rect 24044 19440 24050 19492
rect 13593 19415 13651 19421
rect 13593 19381 13605 19415
rect 13639 19412 13651 19415
rect 13682 19412 13688 19424
rect 13639 19384 13688 19412
rect 13639 19381 13651 19384
rect 13593 19375 13651 19381
rect 13682 19372 13688 19384
rect 13740 19412 13746 19424
rect 13958 19412 13964 19424
rect 13740 19384 13964 19412
rect 13740 19372 13746 19384
rect 13958 19372 13964 19384
rect 14016 19412 14022 19424
rect 15341 19415 15399 19421
rect 15341 19412 15353 19415
rect 14016 19384 15353 19412
rect 14016 19372 14022 19384
rect 15341 19381 15353 19384
rect 15387 19381 15399 19415
rect 15341 19375 15399 19381
rect 15709 19415 15767 19421
rect 15709 19381 15721 19415
rect 15755 19381 15767 19415
rect 15709 19375 15767 19381
rect 15893 19415 15951 19421
rect 15893 19381 15905 19415
rect 15939 19412 15951 19415
rect 16074 19412 16080 19424
rect 15939 19384 16080 19412
rect 15939 19381 15951 19384
rect 15893 19375 15951 19381
rect 12765 19347 12823 19353
rect 12765 19313 12777 19347
rect 12811 19344 12823 19347
rect 14510 19344 14516 19356
rect 12811 19316 14516 19344
rect 12811 19313 12823 19316
rect 12765 19307 12823 19313
rect 14510 19304 14516 19316
rect 14568 19304 14574 19356
rect 15062 19236 15068 19288
rect 15120 19276 15126 19288
rect 15338 19276 15344 19288
rect 15120 19248 15344 19276
rect 15120 19236 15126 19248
rect 15338 19236 15344 19248
rect 15396 19276 15402 19288
rect 15724 19276 15752 19375
rect 16074 19372 16080 19384
rect 16132 19372 16138 19424
rect 16718 19412 16724 19424
rect 16679 19384 16724 19412
rect 16718 19372 16724 19384
rect 16776 19372 16782 19424
rect 17178 19372 17184 19424
rect 17236 19412 17242 19424
rect 17733 19415 17791 19421
rect 17733 19412 17745 19415
rect 17236 19384 17745 19412
rect 17236 19372 17242 19384
rect 17733 19381 17745 19384
rect 17779 19381 17791 19415
rect 19202 19412 19208 19424
rect 19163 19384 19208 19412
rect 17733 19375 17791 19381
rect 17748 19344 17776 19375
rect 19202 19372 19208 19384
rect 19260 19412 19266 19424
rect 19478 19412 19484 19424
rect 19260 19384 19484 19412
rect 19260 19372 19266 19384
rect 19478 19372 19484 19384
rect 19536 19412 19542 19424
rect 20125 19415 20183 19421
rect 20125 19412 20137 19415
rect 19536 19384 20137 19412
rect 19536 19372 19542 19384
rect 20125 19381 20137 19384
rect 20171 19381 20183 19415
rect 20125 19375 20183 19381
rect 20214 19372 20220 19424
rect 20272 19412 20278 19424
rect 20401 19415 20459 19421
rect 20401 19412 20413 19415
rect 20272 19384 20413 19412
rect 20272 19372 20278 19384
rect 20401 19381 20413 19384
rect 20447 19381 20459 19415
rect 22974 19412 22980 19424
rect 22935 19384 22980 19412
rect 20401 19375 20459 19381
rect 22974 19372 22980 19384
rect 23032 19372 23038 19424
rect 23066 19372 23072 19424
rect 23124 19412 23130 19424
rect 24449 19415 24507 19421
rect 24449 19412 24461 19415
rect 23124 19384 24461 19412
rect 23124 19372 23130 19384
rect 24449 19381 24461 19384
rect 24495 19412 24507 19415
rect 24556 19412 24584 19588
rect 25274 19508 25280 19560
rect 25332 19548 25338 19560
rect 25458 19548 25464 19560
rect 25332 19520 25464 19548
rect 25332 19508 25338 19520
rect 25458 19508 25464 19520
rect 25516 19548 25522 19560
rect 26028 19548 26056 19588
rect 26470 19576 26476 19628
rect 26528 19616 26534 19628
rect 27117 19619 27175 19625
rect 27117 19616 27129 19619
rect 26528 19588 27129 19616
rect 26528 19576 26534 19588
rect 27117 19585 27129 19588
rect 27163 19616 27175 19619
rect 27298 19616 27304 19628
rect 27163 19588 27304 19616
rect 27163 19585 27175 19588
rect 27117 19579 27175 19585
rect 27298 19576 27304 19588
rect 27356 19576 27362 19628
rect 26654 19548 26660 19560
rect 25516 19520 25964 19548
rect 26028 19520 26660 19548
rect 25516 19508 25522 19520
rect 24630 19440 24636 19492
rect 24688 19480 24694 19492
rect 25936 19480 25964 19520
rect 26654 19508 26660 19520
rect 26712 19508 26718 19560
rect 28586 19508 28592 19560
rect 28644 19548 28650 19560
rect 28681 19551 28739 19557
rect 28681 19548 28693 19551
rect 28644 19520 28693 19548
rect 28644 19508 28650 19520
rect 28681 19517 28693 19520
rect 28727 19517 28739 19551
rect 28681 19511 28739 19517
rect 29874 19480 29880 19492
rect 24688 19452 25872 19480
rect 25936 19452 28908 19480
rect 24688 19440 24694 19452
rect 25458 19412 25464 19424
rect 24495 19384 24584 19412
rect 25419 19384 25464 19412
rect 24495 19381 24507 19384
rect 24449 19375 24507 19381
rect 25458 19372 25464 19384
rect 25516 19372 25522 19424
rect 25844 19421 25872 19452
rect 25645 19415 25703 19421
rect 25645 19381 25657 19415
rect 25691 19381 25703 19415
rect 25645 19375 25703 19381
rect 25829 19415 25887 19421
rect 25829 19381 25841 19415
rect 25875 19381 25887 19415
rect 26194 19412 26200 19424
rect 26155 19384 26200 19412
rect 25829 19375 25887 19381
rect 19297 19347 19355 19353
rect 19297 19344 19309 19347
rect 17748 19316 19309 19344
rect 19297 19313 19309 19316
rect 19343 19344 19355 19347
rect 19754 19344 19760 19356
rect 19343 19316 19760 19344
rect 19343 19313 19355 19316
rect 19297 19307 19355 19313
rect 19754 19304 19760 19316
rect 19812 19304 19818 19356
rect 25001 19347 25059 19353
rect 25001 19313 25013 19347
rect 25047 19344 25059 19347
rect 25550 19344 25556 19356
rect 25047 19316 25556 19344
rect 25047 19313 25059 19316
rect 25001 19307 25059 19313
rect 25550 19304 25556 19316
rect 25608 19304 25614 19356
rect 16810 19276 16816 19288
rect 15396 19248 15752 19276
rect 16771 19248 16816 19276
rect 15396 19236 15402 19248
rect 16810 19236 16816 19248
rect 16868 19236 16874 19288
rect 19018 19236 19024 19288
rect 19076 19276 19082 19288
rect 19113 19279 19171 19285
rect 19113 19276 19125 19279
rect 19076 19248 19125 19276
rect 19076 19236 19082 19248
rect 19113 19245 19125 19248
rect 19159 19245 19171 19279
rect 19113 19239 19171 19245
rect 20306 19236 20312 19288
rect 20364 19276 20370 19288
rect 25660 19276 25688 19375
rect 26194 19372 26200 19384
rect 26252 19372 26258 19424
rect 28880 19421 28908 19452
rect 29248 19452 29880 19480
rect 29248 19421 29276 19452
rect 29874 19440 29880 19452
rect 29932 19440 29938 19492
rect 26473 19415 26531 19421
rect 26473 19381 26485 19415
rect 26519 19412 26531 19415
rect 28865 19415 28923 19421
rect 26519 19384 28816 19412
rect 26519 19381 26531 19384
rect 26473 19375 26531 19381
rect 27022 19344 27028 19356
rect 26983 19316 27028 19344
rect 27022 19304 27028 19316
rect 27080 19304 27086 19356
rect 28788 19344 28816 19384
rect 28865 19381 28877 19415
rect 28911 19381 28923 19415
rect 28865 19375 28923 19381
rect 29233 19415 29291 19421
rect 29233 19381 29245 19415
rect 29279 19381 29291 19415
rect 29233 19375 29291 19381
rect 29325 19415 29383 19421
rect 29325 19381 29337 19415
rect 29371 19412 29383 19415
rect 29506 19412 29512 19424
rect 29371 19384 29512 19412
rect 29371 19381 29383 19384
rect 29325 19375 29383 19381
rect 29506 19372 29512 19384
rect 29564 19372 29570 19424
rect 29966 19344 29972 19356
rect 28788 19316 29972 19344
rect 29966 19304 29972 19316
rect 30024 19304 30030 19356
rect 20364 19248 25688 19276
rect 20364 19236 20370 19248
rect 11000 19186 30136 19208
rect 11000 19134 19142 19186
rect 19194 19134 19206 19186
rect 19258 19134 19270 19186
rect 19322 19134 19334 19186
rect 19386 19134 29142 19186
rect 29194 19134 29206 19186
rect 29258 19134 29270 19186
rect 29322 19134 29334 19186
rect 29386 19134 30136 19186
rect 11000 19112 30136 19134
rect 13866 19072 13872 19084
rect 12688 19044 13872 19072
rect 12688 18945 12716 19044
rect 13866 19032 13872 19044
rect 13924 19032 13930 19084
rect 20306 19072 20312 19084
rect 20267 19044 20312 19072
rect 20306 19032 20312 19044
rect 20364 19032 20370 19084
rect 21413 19075 21471 19081
rect 21413 19041 21425 19075
rect 21459 19072 21471 19075
rect 22146 19072 22152 19084
rect 21459 19044 22152 19072
rect 21459 19041 21471 19044
rect 21413 19035 21471 19041
rect 22146 19032 22152 19044
rect 22204 19032 22210 19084
rect 22790 19072 22796 19084
rect 22703 19044 22796 19072
rect 12854 18964 12860 19016
rect 12912 19004 12918 19016
rect 13225 19007 13283 19013
rect 13225 19004 13237 19007
rect 12912 18976 13237 19004
rect 12912 18964 12918 18976
rect 13225 18973 13237 18976
rect 13271 18973 13283 19007
rect 13225 18967 13283 18973
rect 14237 19007 14295 19013
rect 14237 18973 14249 19007
rect 14283 19004 14295 19007
rect 16813 19007 16871 19013
rect 16813 19004 16825 19007
rect 14283 18976 16825 19004
rect 14283 18973 14295 18976
rect 14237 18967 14295 18973
rect 16813 18973 16825 18976
rect 16859 18973 16871 19007
rect 16813 18967 16871 18973
rect 17454 18964 17460 19016
rect 17512 18964 17518 19016
rect 18561 19007 18619 19013
rect 18561 18973 18573 19007
rect 18607 19004 18619 19007
rect 19665 19007 19723 19013
rect 19665 19004 19677 19007
rect 18607 18976 19677 19004
rect 18607 18973 18619 18976
rect 18561 18967 18619 18973
rect 19665 18973 19677 18976
rect 19711 19004 19723 19007
rect 19754 19004 19760 19016
rect 19711 18976 19760 19004
rect 19711 18973 19723 18976
rect 19665 18967 19723 18973
rect 19754 18964 19760 18976
rect 19812 18964 19818 19016
rect 22716 19013 22744 19044
rect 22790 19032 22796 19044
rect 22848 19072 22854 19084
rect 24357 19075 24415 19081
rect 24357 19072 24369 19075
rect 22848 19044 24369 19072
rect 22848 19032 22854 19044
rect 24357 19041 24369 19044
rect 24403 19041 24415 19075
rect 24357 19035 24415 19041
rect 26933 19075 26991 19081
rect 26933 19041 26945 19075
rect 26979 19072 26991 19075
rect 27022 19072 27028 19084
rect 26979 19044 27028 19072
rect 26979 19041 26991 19044
rect 26933 19035 26991 19041
rect 27022 19032 27028 19044
rect 27080 19032 27086 19084
rect 29233 19075 29291 19081
rect 29233 19041 29245 19075
rect 29279 19072 29291 19075
rect 29690 19072 29696 19084
rect 29279 19044 29696 19072
rect 29279 19041 29291 19044
rect 29233 19035 29291 19041
rect 29690 19032 29696 19044
rect 29748 19032 29754 19084
rect 22701 19007 22759 19013
rect 22701 18973 22713 19007
rect 22747 18973 22759 19007
rect 22701 18967 22759 18973
rect 22885 19007 22943 19013
rect 22885 18973 22897 19007
rect 22931 19004 22943 19007
rect 23066 19004 23072 19016
rect 22931 18976 23072 19004
rect 22931 18973 22943 18976
rect 22885 18967 22943 18973
rect 23066 18964 23072 18976
rect 23124 18964 23130 19016
rect 23805 19007 23863 19013
rect 23805 18973 23817 19007
rect 23851 19004 23863 19007
rect 23986 19004 23992 19016
rect 23851 18976 23992 19004
rect 23851 18973 23863 18976
rect 23805 18967 23863 18973
rect 23986 18964 23992 18976
rect 24044 19004 24050 19016
rect 24262 19004 24268 19016
rect 24044 18976 24268 19004
rect 24044 18964 24050 18976
rect 24262 18964 24268 18976
rect 24320 18964 24326 19016
rect 26010 19004 26016 19016
rect 25971 18976 26016 19004
rect 26010 18964 26016 18976
rect 26068 18964 26074 19016
rect 26105 19007 26163 19013
rect 26105 18973 26117 19007
rect 26151 19004 26163 19007
rect 27758 19004 27764 19016
rect 26151 18976 27764 19004
rect 26151 18973 26163 18976
rect 26105 18967 26163 18973
rect 27758 18964 27764 18976
rect 27816 18964 27822 19016
rect 12673 18939 12731 18945
rect 12673 18905 12685 18939
rect 12719 18905 12731 18939
rect 12946 18936 12952 18948
rect 12907 18908 12952 18936
rect 12673 18899 12731 18905
rect 12946 18896 12952 18908
rect 13004 18896 13010 18948
rect 14694 18936 14700 18948
rect 14655 18908 14700 18936
rect 14694 18896 14700 18908
rect 14752 18896 14758 18948
rect 14878 18936 14884 18948
rect 14839 18908 14884 18936
rect 14878 18896 14884 18908
rect 14936 18896 14942 18948
rect 15062 18936 15068 18948
rect 15023 18908 15068 18936
rect 15062 18896 15068 18908
rect 15120 18896 15126 18948
rect 15246 18896 15252 18948
rect 15304 18936 15310 18948
rect 15341 18939 15399 18945
rect 15341 18936 15353 18939
rect 15304 18908 15353 18936
rect 15304 18896 15310 18908
rect 15341 18905 15353 18908
rect 15387 18905 15399 18939
rect 15341 18899 15399 18905
rect 20950 18896 20956 18948
rect 21008 18936 21014 18948
rect 21321 18939 21379 18945
rect 21321 18936 21333 18939
rect 21008 18908 21333 18936
rect 21008 18896 21014 18908
rect 21321 18905 21333 18908
rect 21367 18905 21379 18939
rect 21962 18936 21968 18948
rect 21923 18908 21968 18936
rect 21321 18899 21379 18905
rect 21962 18896 21968 18908
rect 22020 18896 22026 18948
rect 22974 18896 22980 18948
rect 23032 18936 23038 18948
rect 23345 18939 23403 18945
rect 23345 18936 23357 18939
rect 23032 18908 23357 18936
rect 23032 18896 23038 18908
rect 23345 18905 23357 18908
rect 23391 18905 23403 18939
rect 25550 18936 25556 18948
rect 25511 18908 25556 18936
rect 23345 18899 23403 18905
rect 25550 18896 25556 18908
rect 25608 18896 25614 18948
rect 27942 18936 27948 18948
rect 27903 18908 27948 18936
rect 27942 18896 27948 18908
rect 28000 18896 28006 18948
rect 29417 18939 29475 18945
rect 29417 18905 29429 18939
rect 29463 18936 29475 18939
rect 29598 18936 29604 18948
rect 29463 18908 29604 18936
rect 29463 18905 29475 18908
rect 29417 18899 29475 18905
rect 29598 18896 29604 18908
rect 29656 18896 29662 18948
rect 12305 18871 12363 18877
rect 12305 18837 12317 18871
rect 12351 18868 12363 18871
rect 13314 18868 13320 18880
rect 12351 18840 13320 18868
rect 12351 18837 12363 18840
rect 12305 18831 12363 18837
rect 13314 18828 13320 18840
rect 13372 18828 13378 18880
rect 15617 18871 15675 18877
rect 15617 18837 15629 18871
rect 15663 18837 15675 18871
rect 15617 18831 15675 18837
rect 13038 18760 13044 18812
rect 13096 18800 13102 18812
rect 15632 18800 15660 18831
rect 16442 18828 16448 18880
rect 16500 18868 16506 18880
rect 16537 18871 16595 18877
rect 16537 18868 16549 18871
rect 16500 18840 16549 18868
rect 16500 18828 16506 18840
rect 16537 18837 16549 18840
rect 16583 18837 16595 18871
rect 16537 18831 16595 18837
rect 19478 18828 19484 18880
rect 19536 18868 19542 18880
rect 19812 18871 19870 18877
rect 19812 18868 19824 18871
rect 19536 18840 19824 18868
rect 19536 18828 19542 18840
rect 19812 18837 19824 18840
rect 19858 18837 19870 18871
rect 19812 18831 19870 18837
rect 20033 18871 20091 18877
rect 20033 18837 20045 18871
rect 20079 18868 20091 18871
rect 20214 18868 20220 18880
rect 20079 18840 20220 18868
rect 20079 18837 20091 18840
rect 20033 18831 20091 18837
rect 20214 18828 20220 18840
rect 20272 18828 20278 18880
rect 23897 18871 23955 18877
rect 23897 18837 23909 18871
rect 23943 18868 23955 18871
rect 24449 18871 24507 18877
rect 24449 18868 24461 18871
rect 23943 18840 24461 18868
rect 23943 18837 23955 18840
rect 23897 18831 23955 18837
rect 24449 18837 24461 18840
rect 24495 18837 24507 18871
rect 26562 18868 26568 18880
rect 26523 18840 26568 18868
rect 24449 18831 24507 18837
rect 26562 18828 26568 18840
rect 26620 18828 26626 18880
rect 26930 18800 26936 18812
rect 13096 18772 15660 18800
rect 26891 18772 26936 18800
rect 13096 18760 13102 18772
rect 15632 18732 15660 18772
rect 26930 18760 26936 18772
rect 26988 18760 26994 18812
rect 27761 18803 27819 18809
rect 27761 18769 27773 18803
rect 27807 18800 27819 18803
rect 27850 18800 27856 18812
rect 27807 18772 27856 18800
rect 27807 18769 27819 18772
rect 27761 18763 27819 18769
rect 27850 18760 27856 18772
rect 27908 18760 27914 18812
rect 16902 18732 16908 18744
rect 15632 18704 16908 18732
rect 16902 18692 16908 18704
rect 16960 18692 16966 18744
rect 18558 18692 18564 18744
rect 18616 18732 18622 18744
rect 19018 18732 19024 18744
rect 18616 18704 19024 18732
rect 18616 18692 18622 18704
rect 19018 18692 19024 18704
rect 19076 18732 19082 18744
rect 19941 18735 19999 18741
rect 19941 18732 19953 18735
rect 19076 18704 19953 18732
rect 19076 18692 19082 18704
rect 19941 18701 19953 18704
rect 19987 18701 19999 18735
rect 19941 18695 19999 18701
rect 11000 18642 30136 18664
rect 11000 18590 14142 18642
rect 14194 18590 14206 18642
rect 14258 18590 14270 18642
rect 14322 18590 14334 18642
rect 14386 18590 24142 18642
rect 24194 18590 24206 18642
rect 24258 18590 24270 18642
rect 24322 18590 24334 18642
rect 24386 18590 30136 18642
rect 11000 18568 30136 18590
rect 27942 18528 27948 18540
rect 27903 18500 27948 18528
rect 27942 18488 27948 18500
rect 28000 18488 28006 18540
rect 29690 18488 29696 18540
rect 29748 18528 29754 18540
rect 29966 18528 29972 18540
rect 29748 18500 29972 18528
rect 29748 18488 29754 18500
rect 29966 18488 29972 18500
rect 30024 18488 30030 18540
rect 12578 18420 12584 18472
rect 12636 18460 12642 18472
rect 15062 18460 15068 18472
rect 12636 18432 15068 18460
rect 12636 18420 12642 18432
rect 15062 18420 15068 18432
rect 15120 18420 15126 18472
rect 15709 18463 15767 18469
rect 15709 18429 15721 18463
rect 15755 18429 15767 18463
rect 15890 18460 15896 18472
rect 15851 18432 15896 18460
rect 15709 18423 15767 18429
rect 13314 18392 13320 18404
rect 13275 18364 13320 18392
rect 13314 18352 13320 18364
rect 13372 18392 13378 18404
rect 15580 18395 15638 18401
rect 15580 18392 15592 18395
rect 13372 18364 15592 18392
rect 13372 18352 13378 18364
rect 15580 18361 15592 18364
rect 15626 18361 15638 18395
rect 15580 18355 15638 18361
rect 12854 18324 12860 18336
rect 12815 18296 12860 18324
rect 12854 18284 12860 18296
rect 12912 18284 12918 18336
rect 13041 18327 13099 18333
rect 13041 18293 13053 18327
rect 13087 18293 13099 18327
rect 13041 18287 13099 18293
rect 13409 18327 13467 18333
rect 13409 18293 13421 18327
rect 13455 18324 13467 18327
rect 13866 18324 13872 18336
rect 13455 18296 13872 18324
rect 13455 18293 13467 18296
rect 13409 18287 13467 18293
rect 13056 18256 13084 18287
rect 13866 18284 13872 18296
rect 13924 18284 13930 18336
rect 14145 18327 14203 18333
rect 14145 18293 14157 18327
rect 14191 18324 14203 18327
rect 14602 18324 14608 18336
rect 14191 18296 14608 18324
rect 14191 18293 14203 18296
rect 14145 18287 14203 18293
rect 14602 18284 14608 18296
rect 14660 18284 14666 18336
rect 15724 18324 15752 18423
rect 15890 18420 15896 18432
rect 15948 18420 15954 18472
rect 17454 18460 17460 18472
rect 17415 18432 17460 18460
rect 17454 18420 17460 18432
rect 17512 18420 17518 18472
rect 18285 18463 18343 18469
rect 18285 18429 18297 18463
rect 18331 18460 18343 18463
rect 21962 18460 21968 18472
rect 18331 18432 21968 18460
rect 18331 18429 18343 18432
rect 18285 18423 18343 18429
rect 21962 18420 21968 18432
rect 22020 18420 22026 18472
rect 22238 18420 22244 18472
rect 22296 18460 22302 18472
rect 22790 18460 22796 18472
rect 22296 18432 22468 18460
rect 22751 18432 22796 18460
rect 22296 18420 22302 18432
rect 15801 18395 15859 18401
rect 15801 18361 15813 18395
rect 15847 18392 15859 18395
rect 18558 18392 18564 18404
rect 15847 18364 18564 18392
rect 15847 18361 15859 18364
rect 15801 18355 15859 18361
rect 18558 18352 18564 18364
rect 18616 18352 18622 18404
rect 18745 18395 18803 18401
rect 18745 18361 18757 18395
rect 18791 18392 18803 18395
rect 21980 18392 22008 18420
rect 22333 18395 22391 18401
rect 22333 18392 22345 18395
rect 18791 18364 20260 18392
rect 21980 18364 22345 18392
rect 18791 18361 18803 18364
rect 18745 18355 18803 18361
rect 16994 18324 17000 18336
rect 15724 18296 17000 18324
rect 16994 18284 17000 18296
rect 17052 18284 17058 18336
rect 17273 18327 17331 18333
rect 17273 18293 17285 18327
rect 17319 18324 17331 18327
rect 17914 18324 17920 18336
rect 17319 18296 17920 18324
rect 17319 18293 17331 18296
rect 17273 18287 17331 18293
rect 17914 18284 17920 18296
rect 17972 18284 17978 18336
rect 18650 18324 18656 18336
rect 18611 18296 18656 18324
rect 18650 18284 18656 18296
rect 18708 18284 18714 18336
rect 18834 18284 18840 18336
rect 18892 18324 18898 18336
rect 19021 18327 19079 18333
rect 19021 18324 19033 18327
rect 18892 18296 19033 18324
rect 18892 18284 18898 18296
rect 19021 18293 19033 18296
rect 19067 18293 19079 18327
rect 19021 18287 19079 18293
rect 19205 18327 19263 18333
rect 19205 18293 19217 18327
rect 19251 18324 19263 18327
rect 19478 18324 19484 18336
rect 19251 18296 19484 18324
rect 19251 18293 19263 18296
rect 19205 18287 19263 18293
rect 19478 18284 19484 18296
rect 19536 18284 19542 18336
rect 20232 18333 20260 18364
rect 22333 18361 22345 18364
rect 22379 18361 22391 18395
rect 22333 18355 22391 18361
rect 20033 18327 20091 18333
rect 20033 18293 20045 18327
rect 20079 18293 20091 18327
rect 20033 18287 20091 18293
rect 20217 18327 20275 18333
rect 20217 18293 20229 18327
rect 20263 18324 20275 18327
rect 22440 18324 22468 18432
rect 22790 18420 22796 18432
rect 22848 18420 22854 18472
rect 27301 18463 27359 18469
rect 27301 18460 27313 18463
rect 23452 18432 27313 18460
rect 23452 18324 23480 18432
rect 27301 18429 27313 18432
rect 27347 18429 27359 18463
rect 28862 18460 28868 18472
rect 28823 18432 28868 18460
rect 27301 18423 27359 18429
rect 28862 18420 28868 18432
rect 28920 18420 28926 18472
rect 25645 18395 25703 18401
rect 25645 18361 25657 18395
rect 25691 18392 25703 18395
rect 26930 18392 26936 18404
rect 25691 18364 26936 18392
rect 25691 18361 25703 18364
rect 25645 18355 25703 18361
rect 26930 18352 26936 18364
rect 26988 18352 26994 18404
rect 27022 18352 27028 18404
rect 27080 18392 27086 18404
rect 27758 18392 27764 18404
rect 27080 18364 27764 18392
rect 27080 18352 27086 18364
rect 27758 18352 27764 18364
rect 27816 18392 27822 18404
rect 27816 18364 27988 18392
rect 27816 18352 27822 18364
rect 20263 18296 23480 18324
rect 23529 18327 23587 18333
rect 20263 18293 20275 18296
rect 20217 18287 20275 18293
rect 23529 18293 23541 18327
rect 23575 18293 23587 18327
rect 23529 18287 23587 18293
rect 15430 18256 15436 18268
rect 13056 18228 14648 18256
rect 15391 18228 15436 18256
rect 12486 18148 12492 18200
rect 12544 18188 12550 18200
rect 12673 18191 12731 18197
rect 12673 18188 12685 18191
rect 12544 18160 12685 18188
rect 12544 18148 12550 18160
rect 12673 18157 12685 18160
rect 12719 18188 12731 18191
rect 13958 18188 13964 18200
rect 12719 18160 13964 18188
rect 12719 18157 12731 18160
rect 12673 18151 12731 18157
rect 13958 18148 13964 18160
rect 14016 18148 14022 18200
rect 14237 18191 14295 18197
rect 14237 18157 14249 18191
rect 14283 18188 14295 18191
rect 14510 18188 14516 18200
rect 14283 18160 14516 18188
rect 14283 18157 14295 18160
rect 14237 18151 14295 18157
rect 14510 18148 14516 18160
rect 14568 18148 14574 18200
rect 14620 18188 14648 18228
rect 15430 18216 15436 18228
rect 15488 18216 15494 18268
rect 15338 18188 15344 18200
rect 14620 18160 15344 18188
rect 15338 18148 15344 18160
rect 15396 18148 15402 18200
rect 20048 18188 20076 18287
rect 20122 18216 20128 18268
rect 20180 18256 20186 18268
rect 20677 18259 20735 18265
rect 20180 18228 20225 18256
rect 20180 18216 20186 18228
rect 20677 18225 20689 18259
rect 20723 18256 20735 18259
rect 21134 18256 21140 18268
rect 20723 18228 21140 18256
rect 20723 18225 20735 18228
rect 20677 18219 20735 18225
rect 21134 18216 21140 18228
rect 21192 18216 21198 18268
rect 22885 18259 22943 18265
rect 22885 18225 22897 18259
rect 22931 18225 22943 18259
rect 22885 18219 22943 18225
rect 20766 18188 20772 18200
rect 20048 18160 20772 18188
rect 20766 18148 20772 18160
rect 20824 18148 20830 18200
rect 22900 18188 22928 18219
rect 23066 18216 23072 18268
rect 23124 18256 23130 18268
rect 23544 18256 23572 18287
rect 23986 18284 23992 18336
rect 24044 18324 24050 18336
rect 24173 18327 24231 18333
rect 24173 18324 24185 18327
rect 24044 18296 24185 18324
rect 24044 18284 24050 18296
rect 24173 18293 24185 18296
rect 24219 18293 24231 18327
rect 24173 18287 24231 18293
rect 24357 18327 24415 18333
rect 24357 18293 24369 18327
rect 24403 18324 24415 18327
rect 24998 18324 25004 18336
rect 24403 18296 25004 18324
rect 24403 18293 24415 18296
rect 24357 18287 24415 18293
rect 24998 18284 25004 18296
rect 25056 18284 25062 18336
rect 26473 18327 26531 18333
rect 26473 18293 26485 18327
rect 26519 18324 26531 18327
rect 26562 18324 26568 18336
rect 26519 18296 26568 18324
rect 26519 18293 26531 18296
rect 26473 18287 26531 18293
rect 26562 18284 26568 18296
rect 26620 18284 26626 18336
rect 27960 18333 27988 18364
rect 27209 18327 27267 18333
rect 27209 18293 27221 18327
rect 27255 18293 27267 18327
rect 27209 18287 27267 18293
rect 27945 18327 28003 18333
rect 27945 18293 27957 18327
rect 27991 18293 28003 18327
rect 28770 18324 28776 18336
rect 28731 18296 28776 18324
rect 27945 18287 28003 18293
rect 23124 18228 23572 18256
rect 26289 18259 26347 18265
rect 23124 18216 23130 18228
rect 26289 18225 26301 18259
rect 26335 18256 26347 18259
rect 26378 18256 26384 18268
rect 26335 18228 26384 18256
rect 26335 18225 26347 18228
rect 26289 18219 26347 18225
rect 26378 18216 26384 18228
rect 26436 18216 26442 18268
rect 26654 18256 26660 18268
rect 26615 18228 26660 18256
rect 26654 18216 26660 18228
rect 26712 18216 26718 18268
rect 27224 18256 27252 18287
rect 28770 18284 28776 18296
rect 28828 18284 28834 18336
rect 29874 18256 29880 18268
rect 27224 18228 29880 18256
rect 23345 18191 23403 18197
rect 23345 18188 23357 18191
rect 22900 18160 23357 18188
rect 23345 18157 23357 18160
rect 23391 18157 23403 18191
rect 24814 18188 24820 18200
rect 24775 18160 24820 18188
rect 23345 18151 23403 18157
rect 24814 18148 24820 18160
rect 24872 18148 24878 18200
rect 26194 18148 26200 18200
rect 26252 18188 26258 18200
rect 27224 18188 27252 18228
rect 29874 18216 29880 18228
rect 29932 18216 29938 18268
rect 26252 18160 27252 18188
rect 26252 18148 26258 18160
rect 11000 18098 30136 18120
rect 11000 18046 19142 18098
rect 19194 18046 19206 18098
rect 19258 18046 19270 18098
rect 19322 18046 19334 18098
rect 19386 18046 29142 18098
rect 29194 18046 29206 18098
rect 29258 18046 29270 18098
rect 29322 18046 29334 18098
rect 29386 18046 30136 18098
rect 11000 18024 30136 18046
rect 14237 17987 14295 17993
rect 14237 17984 14249 17987
rect 13424 17956 14249 17984
rect 13424 17916 13452 17956
rect 14237 17953 14249 17956
rect 14283 17953 14295 17987
rect 14237 17947 14295 17953
rect 15709 17987 15767 17993
rect 15709 17953 15721 17987
rect 15755 17984 15767 17987
rect 16534 17984 16540 17996
rect 15755 17956 16540 17984
rect 15755 17953 15767 17956
rect 15709 17947 15767 17953
rect 16534 17944 16540 17956
rect 16592 17944 16598 17996
rect 16810 17984 16816 17996
rect 16644 17956 16816 17984
rect 13958 17916 13964 17928
rect 12228 17888 13452 17916
rect 13919 17888 13964 17916
rect 12228 17857 12256 17888
rect 13958 17876 13964 17888
rect 14016 17876 14022 17928
rect 15430 17876 15436 17928
rect 15488 17916 15494 17928
rect 16644 17925 16672 17956
rect 16810 17944 16816 17956
rect 16868 17944 16874 17996
rect 16902 17944 16908 17996
rect 16960 17984 16966 17996
rect 16960 17956 17005 17984
rect 16960 17944 16966 17956
rect 18834 17944 18840 17996
rect 18892 17984 18898 17996
rect 20490 17984 20496 17996
rect 18892 17956 20496 17984
rect 18892 17944 18898 17956
rect 20490 17944 20496 17956
rect 20548 17984 20554 17996
rect 23342 17984 23348 17996
rect 20548 17956 23348 17984
rect 20548 17944 20554 17956
rect 23342 17944 23348 17956
rect 23400 17944 23406 17996
rect 15617 17919 15675 17925
rect 15617 17916 15629 17919
rect 15488 17888 15629 17916
rect 15488 17876 15494 17888
rect 15617 17885 15629 17888
rect 15663 17885 15675 17919
rect 15617 17879 15675 17885
rect 15801 17919 15859 17925
rect 15801 17885 15813 17919
rect 15847 17885 15859 17919
rect 15801 17879 15859 17885
rect 16629 17919 16687 17925
rect 16629 17885 16641 17919
rect 16675 17885 16687 17919
rect 16629 17879 16687 17885
rect 12213 17851 12271 17857
rect 12213 17817 12225 17851
rect 12259 17817 12271 17851
rect 12213 17811 12271 17817
rect 12397 17851 12455 17857
rect 12397 17817 12409 17851
rect 12443 17817 12455 17851
rect 12578 17848 12584 17860
rect 12539 17820 12584 17848
rect 12397 17811 12455 17817
rect 11658 17780 11664 17792
rect 11619 17752 11664 17780
rect 11658 17740 11664 17752
rect 11716 17740 11722 17792
rect 12412 17780 12440 17811
rect 12578 17808 12584 17820
rect 12636 17808 12642 17860
rect 12854 17848 12860 17860
rect 12815 17820 12860 17848
rect 12854 17808 12860 17820
rect 12912 17808 12918 17860
rect 13038 17848 13044 17860
rect 12999 17820 13044 17848
rect 13038 17808 13044 17820
rect 13096 17808 13102 17860
rect 14145 17851 14203 17857
rect 14145 17817 14157 17851
rect 14191 17817 14203 17851
rect 14145 17811 14203 17817
rect 12946 17780 12952 17792
rect 12412 17752 12952 17780
rect 12946 17740 12952 17752
rect 13004 17740 13010 17792
rect 12762 17672 12768 17724
rect 12820 17712 12826 17724
rect 14160 17712 14188 17811
rect 15338 17808 15344 17860
rect 15396 17848 15402 17860
rect 15816 17848 15844 17879
rect 17914 17876 17920 17928
rect 17972 17916 17978 17928
rect 24357 17919 24415 17925
rect 17972 17888 21180 17916
rect 17972 17876 17978 17888
rect 21152 17860 21180 17888
rect 24357 17885 24369 17919
rect 24403 17916 24415 17919
rect 24998 17916 25004 17928
rect 24403 17888 25004 17916
rect 24403 17885 24415 17888
rect 24357 17879 24415 17885
rect 24998 17876 25004 17888
rect 25056 17876 25062 17928
rect 26562 17916 26568 17928
rect 25108 17888 26568 17916
rect 16810 17848 16816 17860
rect 15396 17820 15844 17848
rect 16771 17820 16816 17848
rect 15396 17808 15402 17820
rect 16810 17808 16816 17820
rect 16868 17808 16874 17860
rect 19938 17848 19944 17860
rect 19899 17820 19944 17848
rect 19938 17808 19944 17820
rect 19996 17808 20002 17860
rect 20677 17851 20735 17857
rect 20677 17817 20689 17851
rect 20723 17848 20735 17851
rect 20766 17848 20772 17860
rect 20723 17820 20772 17848
rect 20723 17817 20735 17820
rect 20677 17811 20735 17817
rect 20766 17808 20772 17820
rect 20824 17808 20830 17860
rect 21134 17848 21140 17860
rect 21047 17820 21140 17848
rect 21134 17808 21140 17820
rect 21192 17848 21198 17860
rect 22330 17848 22336 17860
rect 21192 17820 22336 17848
rect 21192 17808 21198 17820
rect 22330 17808 22336 17820
rect 22388 17808 22394 17860
rect 23434 17848 23440 17860
rect 23395 17820 23440 17848
rect 23434 17808 23440 17820
rect 23492 17808 23498 17860
rect 23986 17808 23992 17860
rect 24044 17848 24050 17860
rect 24081 17851 24139 17857
rect 24081 17848 24093 17851
rect 24044 17820 24093 17848
rect 24044 17808 24050 17820
rect 24081 17817 24093 17820
rect 24127 17817 24139 17851
rect 24081 17811 24139 17817
rect 15433 17783 15491 17789
rect 15433 17780 15445 17783
rect 15080 17752 15445 17780
rect 14970 17712 14976 17724
rect 12820 17684 14976 17712
rect 12820 17672 12826 17684
rect 14970 17672 14976 17684
rect 15028 17672 15034 17724
rect 13314 17604 13320 17656
rect 13372 17644 13378 17656
rect 15080 17644 15108 17752
rect 15433 17749 15445 17752
rect 15479 17749 15491 17783
rect 15433 17743 15491 17749
rect 16169 17783 16227 17789
rect 16169 17749 16181 17783
rect 16215 17780 16227 17783
rect 16718 17780 16724 17792
rect 16215 17752 16724 17780
rect 16215 17749 16227 17752
rect 16169 17743 16227 17749
rect 16718 17740 16724 17752
rect 16776 17740 16782 17792
rect 20309 17783 20367 17789
rect 20309 17749 20321 17783
rect 20355 17780 20367 17783
rect 25108 17780 25136 17888
rect 26562 17876 26568 17888
rect 26620 17876 26626 17928
rect 29233 17919 29291 17925
rect 27776 17888 28632 17916
rect 26473 17851 26531 17857
rect 26473 17817 26485 17851
rect 26519 17848 26531 17851
rect 26654 17848 26660 17860
rect 26519 17820 26660 17848
rect 26519 17817 26531 17820
rect 26473 17811 26531 17817
rect 26654 17808 26660 17820
rect 26712 17808 26718 17860
rect 27776 17857 27804 17888
rect 28604 17860 28632 17888
rect 29233 17885 29245 17919
rect 29279 17916 29291 17919
rect 29598 17916 29604 17928
rect 29279 17888 29604 17916
rect 29279 17885 29291 17888
rect 29233 17879 29291 17885
rect 29598 17876 29604 17888
rect 29656 17876 29662 17928
rect 27761 17851 27819 17857
rect 27761 17817 27773 17851
rect 27807 17817 27819 17851
rect 28494 17848 28500 17860
rect 28455 17820 28500 17848
rect 27761 17811 27819 17817
rect 20355 17752 25136 17780
rect 25185 17783 25243 17789
rect 20355 17749 20367 17752
rect 20309 17743 20367 17749
rect 25185 17749 25197 17783
rect 25231 17749 25243 17783
rect 25734 17780 25740 17792
rect 25695 17752 25740 17780
rect 25185 17743 25243 17749
rect 23710 17672 23716 17724
rect 23768 17712 23774 17724
rect 25200 17712 25228 17743
rect 25734 17740 25740 17752
rect 25792 17740 25798 17792
rect 27776 17780 27804 17811
rect 28494 17808 28500 17820
rect 28552 17808 28558 17860
rect 28586 17808 28592 17860
rect 28644 17848 28650 17860
rect 29417 17851 29475 17857
rect 29417 17848 29429 17851
rect 28644 17820 29429 17848
rect 28644 17808 28650 17820
rect 29417 17817 29429 17820
rect 29463 17817 29475 17851
rect 29417 17811 29475 17817
rect 25844 17752 27804 17780
rect 23768 17684 25228 17712
rect 23768 17672 23774 17684
rect 25550 17672 25556 17724
rect 25608 17712 25614 17724
rect 25645 17715 25703 17721
rect 25645 17712 25657 17715
rect 25608 17684 25657 17712
rect 25608 17672 25614 17684
rect 25645 17681 25657 17684
rect 25691 17712 25703 17715
rect 25844 17712 25872 17752
rect 27758 17712 27764 17724
rect 25691 17684 25872 17712
rect 27719 17684 27764 17712
rect 25691 17681 25703 17684
rect 25645 17675 25703 17681
rect 27758 17672 27764 17684
rect 27816 17672 27822 17724
rect 13372 17616 15108 17644
rect 13372 17604 13378 17616
rect 20674 17604 20680 17656
rect 20732 17644 20738 17656
rect 21321 17647 21379 17653
rect 21321 17644 21333 17647
rect 20732 17616 21333 17644
rect 20732 17604 20738 17616
rect 21321 17613 21333 17616
rect 21367 17613 21379 17647
rect 21321 17607 21379 17613
rect 11000 17554 30136 17576
rect 11000 17502 14142 17554
rect 14194 17502 14206 17554
rect 14258 17502 14270 17554
rect 14322 17502 14334 17554
rect 14386 17502 24142 17554
rect 24194 17502 24206 17554
rect 24258 17502 24270 17554
rect 24322 17502 24334 17554
rect 24386 17502 30136 17554
rect 11000 17480 30136 17502
rect 13314 17400 13320 17452
rect 13372 17440 13378 17452
rect 13501 17443 13559 17449
rect 13501 17440 13513 17443
rect 13372 17412 13513 17440
rect 13372 17400 13378 17412
rect 13501 17409 13513 17412
rect 13547 17409 13559 17443
rect 27114 17440 27120 17452
rect 13501 17403 13559 17409
rect 16828 17412 27120 17440
rect 16828 17381 16856 17412
rect 27114 17400 27120 17412
rect 27172 17400 27178 17452
rect 16813 17375 16871 17381
rect 16813 17341 16825 17375
rect 16859 17341 16871 17375
rect 23894 17372 23900 17384
rect 16813 17335 16871 17341
rect 22532 17344 23900 17372
rect 12581 17307 12639 17313
rect 12581 17273 12593 17307
rect 12627 17304 12639 17307
rect 12946 17304 12952 17316
rect 12627 17276 12952 17304
rect 12627 17273 12639 17276
rect 12581 17267 12639 17273
rect 12946 17264 12952 17276
rect 13004 17264 13010 17316
rect 14602 17304 14608 17316
rect 14563 17276 14608 17304
rect 14602 17264 14608 17276
rect 14660 17264 14666 17316
rect 14970 17304 14976 17316
rect 14931 17276 14976 17304
rect 14970 17264 14976 17276
rect 15028 17264 15034 17316
rect 15062 17264 15068 17316
rect 15120 17304 15126 17316
rect 15430 17304 15436 17316
rect 15120 17276 15292 17304
rect 15391 17276 15436 17304
rect 15120 17264 15126 17276
rect 12486 17236 12492 17248
rect 12447 17208 12492 17236
rect 12486 17196 12492 17208
rect 12544 17196 12550 17248
rect 12762 17236 12768 17248
rect 12723 17208 12768 17236
rect 12762 17196 12768 17208
rect 12820 17196 12826 17248
rect 12854 17196 12860 17248
rect 12912 17236 12918 17248
rect 13314 17236 13320 17248
rect 12912 17208 13320 17236
rect 12912 17196 12918 17208
rect 13314 17196 13320 17208
rect 13372 17236 13378 17248
rect 13409 17239 13467 17245
rect 13409 17236 13421 17239
rect 13372 17208 13421 17236
rect 13372 17196 13378 17208
rect 13409 17205 13421 17208
rect 13455 17205 13467 17239
rect 13409 17199 13467 17205
rect 15157 17239 15215 17245
rect 15157 17205 15169 17239
rect 15203 17205 15215 17239
rect 15264 17236 15292 17276
rect 15430 17264 15436 17276
rect 15488 17264 15494 17316
rect 22532 17313 22560 17344
rect 23894 17332 23900 17344
rect 23952 17332 23958 17384
rect 25550 17372 25556 17384
rect 25511 17344 25556 17372
rect 25550 17332 25556 17344
rect 25608 17332 25614 17384
rect 22517 17307 22575 17313
rect 22517 17273 22529 17307
rect 22563 17273 22575 17307
rect 22517 17267 22575 17273
rect 23437 17307 23495 17313
rect 23437 17273 23449 17307
rect 23483 17304 23495 17307
rect 23526 17304 23532 17316
rect 23483 17276 23532 17304
rect 23483 17273 23495 17276
rect 23437 17267 23495 17273
rect 23526 17264 23532 17276
rect 23584 17264 23590 17316
rect 25366 17264 25372 17316
rect 25424 17304 25430 17316
rect 26197 17307 26255 17313
rect 26197 17304 26209 17307
rect 25424 17276 26209 17304
rect 25424 17264 25430 17276
rect 26197 17273 26209 17276
rect 26243 17273 26255 17307
rect 28494 17304 28500 17316
rect 28455 17276 28500 17304
rect 26197 17267 26255 17273
rect 28494 17264 28500 17276
rect 28552 17264 28558 17316
rect 28954 17264 28960 17316
rect 29012 17304 29018 17316
rect 29325 17307 29383 17313
rect 29325 17304 29337 17307
rect 29012 17276 29337 17304
rect 29012 17264 29018 17276
rect 29325 17273 29337 17276
rect 29371 17273 29383 17307
rect 29325 17267 29383 17273
rect 15525 17239 15583 17245
rect 15525 17236 15537 17239
rect 15264 17208 15537 17236
rect 15157 17199 15215 17205
rect 15525 17205 15537 17208
rect 15571 17205 15583 17239
rect 16718 17236 16724 17248
rect 16679 17208 16724 17236
rect 15525 17199 15583 17205
rect 15172 17168 15200 17199
rect 16718 17196 16724 17208
rect 16776 17196 16782 17248
rect 16994 17236 17000 17248
rect 16955 17208 17000 17236
rect 16994 17196 17000 17208
rect 17052 17196 17058 17248
rect 17914 17236 17920 17248
rect 17875 17208 17920 17236
rect 17914 17196 17920 17208
rect 17972 17196 17978 17248
rect 19297 17239 19355 17245
rect 19297 17205 19309 17239
rect 19343 17205 19355 17239
rect 19297 17199 19355 17205
rect 16810 17168 16816 17180
rect 15172 17140 16816 17168
rect 16810 17128 16816 17140
rect 16868 17168 16874 17180
rect 17457 17171 17515 17177
rect 17457 17168 17469 17171
rect 16868 17140 17469 17168
rect 16868 17128 16874 17140
rect 17457 17137 17469 17140
rect 17503 17137 17515 17171
rect 17457 17131 17515 17137
rect 18098 17100 18104 17112
rect 18059 17072 18104 17100
rect 18098 17060 18104 17072
rect 18156 17060 18162 17112
rect 19312 17100 19340 17199
rect 20674 17196 20680 17248
rect 20732 17196 20738 17248
rect 23342 17236 23348 17248
rect 23255 17208 23348 17236
rect 23342 17196 23348 17208
rect 23400 17236 23406 17248
rect 23400 17208 23664 17236
rect 23400 17196 23406 17208
rect 19570 17168 19576 17180
rect 19531 17140 19576 17168
rect 19570 17128 19576 17140
rect 19628 17128 19634 17180
rect 21318 17168 21324 17180
rect 21279 17140 21324 17168
rect 21318 17128 21324 17140
rect 21376 17128 21382 17180
rect 22609 17171 22667 17177
rect 22609 17137 22621 17171
rect 22655 17137 22667 17171
rect 23636 17168 23664 17208
rect 23710 17196 23716 17248
rect 23768 17236 23774 17248
rect 24081 17239 24139 17245
rect 24081 17236 24093 17239
rect 23768 17208 24093 17236
rect 23768 17196 23774 17208
rect 24081 17205 24093 17208
rect 24127 17205 24139 17239
rect 24998 17236 25004 17248
rect 24959 17208 25004 17236
rect 24081 17199 24139 17205
rect 24998 17196 25004 17208
rect 25056 17196 25062 17248
rect 27025 17239 27083 17245
rect 27025 17236 27037 17239
rect 25108 17208 27037 17236
rect 25108 17168 25136 17208
rect 27025 17205 27037 17208
rect 27071 17205 27083 17239
rect 27025 17199 27083 17205
rect 27117 17239 27175 17245
rect 27117 17205 27129 17239
rect 27163 17236 27175 17239
rect 27206 17236 27212 17248
rect 27163 17208 27212 17236
rect 27163 17205 27175 17208
rect 27117 17199 27175 17205
rect 23636 17140 25136 17168
rect 26289 17171 26347 17177
rect 22609 17131 22667 17137
rect 26289 17137 26301 17171
rect 26335 17168 26347 17171
rect 26470 17168 26476 17180
rect 26335 17140 26476 17168
rect 26335 17137 26347 17140
rect 26289 17131 26347 17137
rect 19478 17100 19484 17112
rect 19312 17072 19484 17100
rect 19478 17060 19484 17072
rect 19536 17060 19542 17112
rect 22624 17100 22652 17131
rect 26470 17128 26476 17140
rect 26528 17128 26534 17180
rect 27040 17168 27068 17199
rect 27206 17196 27212 17208
rect 27264 17196 27270 17248
rect 28310 17196 28316 17248
rect 28368 17236 28374 17248
rect 28405 17239 28463 17245
rect 28405 17236 28417 17239
rect 28368 17208 28417 17236
rect 28368 17196 28374 17208
rect 28405 17205 28417 17208
rect 28451 17205 28463 17239
rect 28405 17199 28463 17205
rect 29233 17239 29291 17245
rect 29233 17205 29245 17239
rect 29279 17236 29291 17239
rect 29874 17236 29880 17248
rect 29279 17208 29880 17236
rect 29279 17205 29291 17208
rect 29233 17199 29291 17205
rect 29248 17168 29276 17199
rect 29874 17196 29880 17208
rect 29932 17196 29938 17248
rect 27040 17140 29276 17168
rect 23434 17100 23440 17112
rect 22624 17072 23440 17100
rect 23434 17060 23440 17072
rect 23492 17060 23498 17112
rect 11000 17010 30136 17032
rect 11000 16958 19142 17010
rect 19194 16958 19206 17010
rect 19258 16958 19270 17010
rect 19322 16958 19334 17010
rect 19386 16958 29142 17010
rect 29194 16958 29206 17010
rect 29258 16958 29270 17010
rect 29322 16958 29334 17010
rect 29386 16958 30136 17010
rect 11000 16936 30136 16958
rect 16442 16896 16448 16908
rect 13976 16868 16448 16896
rect 11569 16831 11627 16837
rect 11569 16797 11581 16831
rect 11615 16828 11627 16831
rect 11658 16828 11664 16840
rect 11615 16800 11664 16828
rect 11615 16797 11627 16800
rect 11569 16791 11627 16797
rect 11658 16788 11664 16800
rect 11716 16788 11722 16840
rect 12118 16788 12124 16840
rect 12176 16788 12182 16840
rect 13314 16828 13320 16840
rect 13275 16800 13320 16828
rect 13314 16788 13320 16800
rect 13372 16788 13378 16840
rect 11290 16760 11296 16772
rect 11251 16732 11296 16760
rect 11290 16720 11296 16732
rect 11348 16720 11354 16772
rect 12946 16720 12952 16772
rect 13004 16760 13010 16772
rect 13976 16769 14004 16868
rect 16442 16856 16448 16868
rect 16500 16896 16506 16908
rect 17638 16896 17644 16908
rect 16500 16868 17644 16896
rect 16500 16856 16506 16868
rect 14237 16831 14295 16837
rect 14237 16797 14249 16831
rect 14283 16828 14295 16831
rect 14510 16828 14516 16840
rect 14283 16800 14516 16828
rect 14283 16797 14295 16800
rect 14237 16791 14295 16797
rect 14510 16788 14516 16800
rect 14568 16788 14574 16840
rect 14694 16788 14700 16840
rect 14752 16788 14758 16840
rect 16736 16769 16764 16868
rect 17638 16856 17644 16868
rect 17696 16896 17702 16908
rect 19478 16896 19484 16908
rect 17696 16868 19484 16896
rect 17696 16856 17702 16868
rect 19478 16856 19484 16868
rect 19536 16856 19542 16908
rect 19570 16856 19576 16908
rect 19628 16896 19634 16908
rect 19941 16899 19999 16905
rect 19941 16896 19953 16899
rect 19628 16868 19953 16896
rect 19628 16856 19634 16868
rect 19941 16865 19953 16868
rect 19987 16865 19999 16899
rect 19941 16859 19999 16865
rect 25734 16856 25740 16908
rect 25792 16896 25798 16908
rect 26013 16899 26071 16905
rect 26013 16896 26025 16899
rect 25792 16868 26025 16896
rect 25792 16856 25798 16868
rect 26013 16865 26025 16868
rect 26059 16865 26071 16899
rect 26013 16859 26071 16865
rect 24081 16831 24139 16837
rect 24081 16797 24093 16831
rect 24127 16828 24139 16831
rect 24814 16828 24820 16840
rect 24127 16800 24820 16828
rect 24127 16797 24139 16800
rect 24081 16791 24139 16797
rect 24814 16788 24820 16800
rect 24872 16788 24878 16840
rect 27577 16831 27635 16837
rect 27577 16797 27589 16831
rect 27623 16828 27635 16831
rect 27758 16828 27764 16840
rect 27623 16800 27764 16828
rect 27623 16797 27635 16800
rect 27577 16791 27635 16797
rect 27758 16788 27764 16800
rect 27816 16788 27822 16840
rect 13961 16763 14019 16769
rect 13961 16760 13973 16763
rect 13004 16732 13973 16760
rect 13004 16720 13010 16732
rect 13961 16729 13973 16732
rect 14007 16729 14019 16763
rect 13961 16723 14019 16729
rect 16721 16763 16779 16769
rect 16721 16729 16733 16763
rect 16767 16729 16779 16763
rect 16721 16723 16779 16729
rect 18098 16720 18104 16772
rect 18156 16720 18162 16772
rect 19570 16720 19576 16772
rect 19628 16760 19634 16772
rect 19665 16763 19723 16769
rect 19665 16760 19677 16763
rect 19628 16732 19677 16760
rect 19628 16720 19634 16732
rect 19665 16729 19677 16732
rect 19711 16729 19723 16763
rect 19665 16723 19723 16729
rect 19849 16763 19907 16769
rect 19849 16729 19861 16763
rect 19895 16760 19907 16763
rect 20766 16760 20772 16772
rect 19895 16732 20772 16760
rect 19895 16729 19907 16732
rect 19849 16723 19907 16729
rect 20766 16720 20772 16732
rect 20824 16720 20830 16772
rect 22514 16760 22520 16772
rect 22270 16732 22520 16760
rect 22514 16720 22520 16732
rect 22572 16720 22578 16772
rect 23434 16720 23440 16772
rect 23492 16760 23498 16772
rect 23529 16763 23587 16769
rect 23529 16760 23541 16763
rect 23492 16732 23541 16760
rect 23492 16720 23498 16732
rect 23529 16729 23541 16732
rect 23575 16729 23587 16763
rect 25185 16763 25243 16769
rect 25185 16760 25197 16763
rect 23529 16723 23587 16729
rect 23820 16732 25197 16760
rect 11308 16692 11336 16720
rect 12964 16692 12992 16720
rect 11308 16664 12992 16692
rect 14970 16652 14976 16704
rect 15028 16692 15034 16704
rect 15985 16695 16043 16701
rect 15985 16692 15997 16695
rect 15028 16664 15997 16692
rect 15028 16652 15034 16664
rect 15985 16661 15997 16664
rect 16031 16661 16043 16695
rect 15985 16655 16043 16661
rect 16997 16695 17055 16701
rect 16997 16661 17009 16695
rect 17043 16692 17055 16695
rect 18006 16692 18012 16704
rect 17043 16664 18012 16692
rect 17043 16661 17055 16664
rect 16997 16655 17055 16661
rect 18006 16652 18012 16664
rect 18064 16652 18070 16704
rect 18745 16695 18803 16701
rect 18745 16661 18757 16695
rect 18791 16661 18803 16695
rect 18745 16655 18803 16661
rect 17178 16516 17184 16568
rect 17236 16556 17242 16568
rect 18760 16556 18788 16655
rect 19478 16652 19484 16704
rect 19536 16692 19542 16704
rect 20858 16692 20864 16704
rect 19536 16664 20864 16692
rect 19536 16652 19542 16664
rect 20858 16652 20864 16664
rect 20916 16652 20922 16704
rect 21134 16692 21140 16704
rect 21095 16664 21140 16692
rect 21134 16652 21140 16664
rect 21192 16652 21198 16704
rect 22885 16695 22943 16701
rect 22885 16692 22897 16695
rect 22256 16664 22897 16692
rect 22256 16636 22284 16664
rect 22885 16661 22897 16664
rect 22931 16661 22943 16695
rect 22885 16655 22943 16661
rect 22238 16584 22244 16636
rect 22296 16584 22302 16636
rect 22330 16584 22336 16636
rect 22388 16624 22394 16636
rect 23820 16624 23848 16732
rect 25185 16729 25197 16732
rect 25231 16760 25243 16763
rect 25826 16760 25832 16772
rect 25231 16732 25832 16760
rect 25231 16729 25243 16732
rect 25185 16723 25243 16729
rect 25826 16720 25832 16732
rect 25884 16720 25890 16772
rect 25921 16763 25979 16769
rect 25921 16729 25933 16763
rect 25967 16729 25979 16763
rect 25921 16723 25979 16729
rect 23986 16692 23992 16704
rect 23899 16664 23992 16692
rect 23986 16652 23992 16664
rect 24044 16692 24050 16704
rect 25936 16692 25964 16723
rect 26470 16720 26476 16772
rect 26528 16760 26534 16772
rect 27117 16763 27175 16769
rect 27117 16760 27129 16763
rect 26528 16732 27129 16760
rect 26528 16720 26534 16732
rect 27117 16729 27129 16732
rect 27163 16729 27175 16763
rect 27117 16723 27175 16729
rect 28494 16720 28500 16772
rect 28552 16760 28558 16772
rect 28589 16763 28647 16769
rect 28589 16760 28601 16763
rect 28552 16732 28601 16760
rect 28552 16720 28558 16732
rect 28589 16729 28601 16732
rect 28635 16729 28647 16763
rect 28589 16723 28647 16729
rect 24044 16664 25964 16692
rect 27669 16695 27727 16701
rect 24044 16652 24050 16664
rect 27669 16661 27681 16695
rect 27715 16692 27727 16695
rect 28770 16692 28776 16704
rect 27715 16664 28776 16692
rect 27715 16661 27727 16664
rect 27669 16655 27727 16661
rect 28770 16652 28776 16664
rect 28828 16652 28834 16704
rect 28862 16652 28868 16704
rect 28920 16692 28926 16704
rect 29141 16695 29199 16701
rect 29141 16692 29153 16695
rect 28920 16664 29153 16692
rect 28920 16652 28926 16664
rect 29141 16661 29153 16664
rect 29187 16661 29199 16695
rect 29141 16655 29199 16661
rect 22388 16596 23848 16624
rect 29049 16627 29107 16633
rect 22388 16584 22394 16596
rect 29049 16593 29061 16627
rect 29095 16624 29107 16627
rect 29598 16624 29604 16636
rect 29095 16596 29604 16624
rect 29095 16593 29107 16596
rect 29049 16587 29107 16593
rect 29598 16584 29604 16596
rect 29656 16584 29662 16636
rect 25366 16556 25372 16568
rect 17236 16528 18788 16556
rect 25327 16528 25372 16556
rect 17236 16516 17242 16528
rect 25366 16516 25372 16528
rect 25424 16516 25430 16568
rect 11000 16466 30136 16488
rect 11000 16414 14142 16466
rect 14194 16414 14206 16466
rect 14258 16414 14270 16466
rect 14322 16414 14334 16466
rect 14386 16414 24142 16466
rect 24194 16414 24206 16466
rect 24258 16414 24270 16466
rect 24322 16414 24334 16466
rect 24386 16414 30136 16466
rect 11000 16392 30136 16414
rect 12118 16352 12124 16364
rect 12079 16324 12124 16352
rect 12118 16312 12124 16324
rect 12176 16312 12182 16364
rect 14605 16355 14663 16361
rect 14605 16321 14617 16355
rect 14651 16352 14663 16355
rect 14694 16352 14700 16364
rect 14651 16324 14700 16352
rect 14651 16321 14663 16324
rect 14605 16315 14663 16321
rect 14694 16312 14700 16324
rect 14752 16312 14758 16364
rect 15341 16355 15399 16361
rect 15341 16321 15353 16355
rect 15387 16352 15399 16355
rect 15430 16352 15436 16364
rect 15387 16324 15436 16352
rect 15387 16321 15399 16324
rect 15341 16315 15399 16321
rect 15430 16312 15436 16324
rect 15488 16312 15494 16364
rect 15985 16355 16043 16361
rect 15985 16321 15997 16355
rect 16031 16352 16043 16355
rect 16994 16352 17000 16364
rect 16031 16324 17000 16352
rect 16031 16321 16043 16324
rect 15985 16315 16043 16321
rect 16994 16312 17000 16324
rect 17052 16312 17058 16364
rect 17914 16352 17920 16364
rect 17104 16324 17920 16352
rect 17104 16216 17132 16324
rect 17914 16312 17920 16324
rect 17972 16312 17978 16364
rect 19570 16352 19576 16364
rect 19531 16324 19576 16352
rect 19570 16312 19576 16324
rect 19628 16312 19634 16364
rect 22514 16352 22520 16364
rect 22475 16324 22520 16352
rect 22514 16312 22520 16324
rect 22572 16312 22578 16364
rect 27114 16352 27120 16364
rect 27075 16324 27120 16352
rect 27114 16312 27120 16324
rect 27172 16312 27178 16364
rect 18006 16284 18012 16296
rect 17967 16256 18012 16284
rect 18006 16244 18012 16256
rect 18064 16244 18070 16296
rect 20858 16244 20864 16296
rect 20916 16284 20922 16296
rect 20916 16256 23112 16284
rect 20916 16244 20922 16256
rect 14436 16188 17132 16216
rect 20953 16219 21011 16225
rect 11934 16148 11940 16160
rect 11895 16120 11940 16148
rect 11934 16108 11940 16120
rect 11992 16148 11998 16160
rect 13774 16148 13780 16160
rect 11992 16120 13780 16148
rect 11992 16108 11998 16120
rect 13774 16108 13780 16120
rect 13832 16148 13838 16160
rect 14436 16157 14464 16188
rect 20953 16185 20965 16219
rect 20999 16216 21011 16219
rect 21134 16216 21140 16228
rect 20999 16188 21140 16216
rect 20999 16185 21011 16188
rect 20953 16179 21011 16185
rect 21134 16176 21140 16188
rect 21192 16176 21198 16228
rect 14421 16151 14479 16157
rect 14421 16148 14433 16151
rect 13832 16120 14433 16148
rect 13832 16108 13838 16120
rect 14421 16117 14433 16120
rect 14467 16117 14479 16151
rect 14421 16111 14479 16117
rect 14970 16108 14976 16160
rect 15028 16148 15034 16160
rect 15249 16151 15307 16157
rect 15249 16148 15261 16151
rect 15028 16120 15261 16148
rect 15028 16108 15034 16120
rect 15249 16117 15261 16120
rect 15295 16117 15307 16151
rect 15249 16111 15307 16117
rect 15893 16151 15951 16157
rect 15893 16117 15905 16151
rect 15939 16117 15951 16151
rect 15893 16111 15951 16117
rect 17089 16151 17147 16157
rect 17089 16117 17101 16151
rect 17135 16117 17147 16151
rect 17089 16111 17147 16117
rect 14878 16040 14884 16092
rect 14936 16080 14942 16092
rect 15908 16080 15936 16111
rect 14936 16052 15936 16080
rect 17104 16080 17132 16111
rect 17178 16108 17184 16160
rect 17236 16148 17242 16160
rect 17638 16148 17644 16160
rect 17236 16120 17281 16148
rect 17599 16120 17644 16148
rect 17236 16108 17242 16120
rect 17638 16108 17644 16120
rect 17696 16108 17702 16160
rect 17825 16151 17883 16157
rect 17825 16117 17837 16151
rect 17871 16148 17883 16151
rect 18282 16148 18288 16160
rect 17871 16120 18288 16148
rect 17871 16117 17883 16120
rect 17825 16111 17883 16117
rect 18282 16108 18288 16120
rect 18340 16108 18346 16160
rect 18926 16108 18932 16160
rect 18984 16148 18990 16160
rect 19113 16151 19171 16157
rect 19113 16148 19125 16151
rect 18984 16120 19125 16148
rect 18984 16108 18990 16120
rect 19113 16117 19125 16120
rect 19159 16117 19171 16151
rect 19113 16111 19171 16117
rect 19389 16151 19447 16157
rect 19389 16117 19401 16151
rect 19435 16117 19447 16151
rect 19389 16111 19447 16117
rect 20585 16151 20643 16157
rect 20585 16117 20597 16151
rect 20631 16148 20643 16151
rect 20766 16148 20772 16160
rect 20631 16120 20772 16148
rect 20631 16117 20643 16120
rect 20585 16111 20643 16117
rect 17656 16080 17684 16108
rect 17104 16052 17684 16080
rect 14936 16040 14942 16052
rect 17656 16012 17684 16052
rect 19018 16040 19024 16092
rect 19076 16080 19082 16092
rect 19297 16083 19355 16089
rect 19297 16080 19309 16083
rect 19076 16052 19309 16080
rect 19076 16040 19082 16052
rect 19297 16049 19309 16052
rect 19343 16049 19355 16083
rect 19297 16043 19355 16049
rect 19404 16012 19432 16111
rect 20766 16108 20772 16120
rect 20824 16108 20830 16160
rect 21410 16148 21416 16160
rect 21371 16120 21416 16148
rect 21410 16108 21416 16120
rect 21468 16108 21474 16160
rect 22330 16108 22336 16160
rect 22388 16148 22394 16160
rect 23084 16148 23112 16256
rect 23158 16176 23164 16228
rect 23216 16216 23222 16228
rect 25645 16219 25703 16225
rect 25645 16216 25657 16219
rect 23216 16188 25657 16216
rect 23216 16176 23222 16188
rect 25645 16185 25657 16188
rect 25691 16185 25703 16219
rect 25645 16179 25703 16185
rect 26120 16188 28632 16216
rect 23621 16151 23679 16157
rect 23621 16148 23633 16151
rect 22388 16120 22433 16148
rect 23084 16120 23633 16148
rect 22388 16108 22394 16120
rect 23621 16117 23633 16120
rect 23667 16117 23679 16151
rect 25366 16148 25372 16160
rect 25030 16120 25372 16148
rect 23621 16111 23679 16117
rect 20401 16083 20459 16089
rect 20401 16049 20413 16083
rect 20447 16080 20459 16083
rect 21505 16083 21563 16089
rect 21505 16080 21517 16083
rect 20447 16052 21517 16080
rect 20447 16049 20459 16052
rect 20401 16043 20459 16049
rect 21505 16049 21517 16052
rect 21551 16049 21563 16083
rect 21505 16043 21563 16049
rect 17656 15984 19432 16012
rect 23636 16012 23664 16111
rect 25366 16108 25372 16120
rect 25424 16108 25430 16160
rect 25826 16108 25832 16160
rect 25884 16148 25890 16160
rect 26120 16157 26148 16188
rect 26105 16151 26163 16157
rect 26105 16148 26117 16151
rect 25884 16120 26117 16148
rect 25884 16108 25890 16120
rect 26105 16117 26117 16120
rect 26151 16117 26163 16151
rect 27022 16148 27028 16160
rect 26983 16120 27028 16148
rect 26105 16111 26163 16117
rect 27022 16108 27028 16120
rect 27080 16108 27086 16160
rect 27850 16108 27856 16160
rect 27908 16148 27914 16160
rect 28604 16157 28632 16188
rect 27945 16151 28003 16157
rect 27945 16148 27957 16151
rect 27908 16120 27957 16148
rect 27908 16108 27914 16120
rect 27945 16117 27957 16120
rect 27991 16117 28003 16151
rect 27945 16111 28003 16117
rect 28589 16151 28647 16157
rect 28589 16117 28601 16151
rect 28635 16148 28647 16151
rect 28954 16148 28960 16160
rect 28635 16120 28960 16148
rect 28635 16117 28647 16120
rect 28589 16111 28647 16117
rect 28954 16108 28960 16120
rect 29012 16108 29018 16160
rect 23894 16080 23900 16092
rect 23855 16052 23900 16080
rect 23894 16040 23900 16052
rect 23952 16040 23958 16092
rect 25274 16012 25280 16024
rect 23636 15984 25280 16012
rect 25274 15972 25280 15984
rect 25332 15972 25338 16024
rect 26286 16012 26292 16024
rect 26247 15984 26292 16012
rect 26286 15972 26292 15984
rect 26344 15972 26350 16024
rect 27942 15972 27948 16024
rect 28000 16012 28006 16024
rect 28037 16015 28095 16021
rect 28037 16012 28049 16015
rect 28000 15984 28049 16012
rect 28000 15972 28006 15984
rect 28037 15981 28049 15984
rect 28083 16012 28095 16015
rect 28586 16012 28592 16024
rect 28083 15984 28592 16012
rect 28083 15981 28095 15984
rect 28037 15975 28095 15981
rect 28586 15972 28592 15984
rect 28644 15972 28650 16024
rect 28678 15972 28684 16024
rect 28736 16012 28742 16024
rect 28773 16015 28831 16021
rect 28773 16012 28785 16015
rect 28736 15984 28785 16012
rect 28736 15972 28742 15984
rect 28773 15981 28785 15984
rect 28819 15981 28831 16015
rect 28773 15975 28831 15981
rect 11000 15922 30136 15944
rect 11000 15870 19142 15922
rect 19194 15870 19206 15922
rect 19258 15870 19270 15922
rect 19322 15870 19334 15922
rect 19386 15870 29142 15922
rect 29194 15870 29206 15922
rect 29258 15870 29270 15922
rect 29322 15870 29334 15922
rect 29386 15870 30136 15922
rect 11000 15848 30136 15870
rect 23894 15768 23900 15820
rect 23952 15808 23958 15820
rect 24081 15811 24139 15817
rect 24081 15808 24093 15811
rect 23952 15780 24093 15808
rect 23952 15768 23958 15780
rect 24081 15777 24093 15780
rect 24127 15777 24139 15811
rect 24081 15771 24139 15777
rect 27942 15740 27948 15752
rect 22072 15712 22468 15740
rect 11750 15672 11756 15684
rect 11711 15644 11756 15672
rect 11750 15632 11756 15644
rect 11808 15632 11814 15684
rect 13038 15672 13044 15684
rect 12999 15644 13044 15672
rect 13038 15632 13044 15644
rect 13096 15632 13102 15684
rect 14697 15675 14755 15681
rect 14697 15641 14709 15675
rect 14743 15641 14755 15675
rect 14697 15635 14755 15641
rect 11658 15604 11664 15616
rect 11571 15576 11664 15604
rect 11658 15564 11664 15576
rect 11716 15604 11722 15616
rect 12670 15604 12676 15616
rect 11716 15576 12676 15604
rect 11716 15564 11722 15576
rect 12670 15564 12676 15576
rect 12728 15564 12734 15616
rect 14712 15604 14740 15635
rect 14786 15632 14792 15684
rect 14844 15672 14850 15684
rect 15246 15672 15252 15684
rect 14844 15644 14889 15672
rect 15207 15644 15252 15672
rect 14844 15632 14850 15644
rect 15246 15632 15252 15644
rect 15304 15632 15310 15684
rect 15433 15675 15491 15681
rect 15433 15641 15445 15675
rect 15479 15672 15491 15675
rect 16074 15672 16080 15684
rect 15479 15644 16080 15672
rect 15479 15641 15491 15644
rect 15433 15635 15491 15641
rect 16074 15632 16080 15644
rect 16132 15632 16138 15684
rect 17178 15672 17184 15684
rect 17139 15644 17184 15672
rect 17178 15632 17184 15644
rect 17236 15632 17242 15684
rect 17733 15675 17791 15681
rect 17733 15641 17745 15675
rect 17779 15672 17791 15675
rect 18190 15672 18196 15684
rect 17779 15644 18196 15672
rect 17779 15641 17791 15644
rect 17733 15635 17791 15641
rect 18190 15632 18196 15644
rect 18248 15632 18254 15684
rect 18282 15632 18288 15684
rect 18340 15672 18346 15684
rect 18377 15675 18435 15681
rect 18377 15672 18389 15675
rect 18340 15644 18389 15672
rect 18340 15632 18346 15644
rect 18377 15641 18389 15644
rect 18423 15641 18435 15675
rect 18558 15672 18564 15684
rect 18519 15644 18564 15672
rect 18377 15635 18435 15641
rect 18558 15632 18564 15644
rect 18616 15632 18622 15684
rect 20033 15675 20091 15681
rect 20033 15672 20045 15675
rect 18668 15644 20045 15672
rect 18208 15604 18236 15632
rect 18668 15604 18696 15644
rect 20033 15641 20045 15644
rect 20079 15641 20091 15675
rect 20033 15635 20091 15641
rect 20125 15675 20183 15681
rect 20125 15641 20137 15675
rect 20171 15641 20183 15675
rect 20125 15635 20183 15641
rect 21873 15675 21931 15681
rect 21873 15641 21885 15675
rect 21919 15672 21931 15675
rect 22072 15672 22100 15712
rect 22238 15672 22244 15684
rect 21919 15644 22100 15672
rect 22199 15644 22244 15672
rect 21919 15641 21931 15644
rect 21873 15635 21931 15641
rect 18926 15604 18932 15616
rect 14712 15576 14832 15604
rect 18208 15576 18696 15604
rect 18887 15576 18932 15604
rect 13133 15539 13191 15545
rect 13133 15505 13145 15539
rect 13179 15536 13191 15539
rect 14694 15536 14700 15548
rect 13179 15508 14700 15536
rect 13179 15505 13191 15508
rect 13133 15499 13191 15505
rect 14694 15496 14700 15508
rect 14752 15496 14758 15548
rect 14804 15536 14832 15576
rect 18926 15564 18932 15576
rect 18984 15564 18990 15616
rect 20140 15604 20168 15635
rect 22238 15632 22244 15644
rect 22296 15632 22302 15684
rect 22440 15672 22468 15712
rect 23084 15712 23388 15740
rect 22514 15672 22520 15684
rect 22440 15644 22520 15672
rect 22514 15632 22520 15644
rect 22572 15632 22578 15684
rect 23084 15681 23112 15712
rect 23069 15675 23127 15681
rect 23069 15641 23081 15675
rect 23115 15641 23127 15675
rect 23360 15672 23388 15712
rect 23636 15712 23940 15740
rect 23636 15681 23664 15712
rect 23621 15675 23679 15681
rect 23621 15672 23633 15675
rect 23069 15635 23127 15641
rect 23268 15644 23633 15672
rect 22256 15604 22284 15632
rect 20140 15576 22284 15604
rect 22333 15607 22391 15613
rect 22333 15573 22345 15607
rect 22379 15604 22391 15607
rect 22977 15607 23035 15613
rect 22977 15604 22989 15607
rect 22379 15576 22989 15604
rect 22379 15573 22391 15576
rect 22333 15567 22391 15573
rect 22977 15573 22989 15576
rect 23023 15604 23035 15607
rect 23158 15604 23164 15616
rect 23023 15576 23164 15604
rect 23023 15573 23035 15576
rect 22977 15567 23035 15573
rect 23158 15564 23164 15576
rect 23216 15564 23222 15616
rect 15246 15536 15252 15548
rect 14804 15508 15252 15536
rect 15246 15496 15252 15508
rect 15304 15536 15310 15548
rect 17638 15536 17644 15548
rect 15304 15508 17644 15536
rect 15304 15496 15310 15508
rect 17638 15496 17644 15508
rect 17696 15496 17702 15548
rect 19846 15536 19852 15548
rect 19759 15508 19852 15536
rect 19846 15496 19852 15508
rect 19904 15536 19910 15548
rect 21318 15536 21324 15548
rect 19904 15508 21324 15536
rect 19904 15496 19910 15508
rect 21318 15496 21324 15508
rect 21376 15496 21382 15548
rect 21689 15539 21747 15545
rect 21689 15505 21701 15539
rect 21735 15536 21747 15539
rect 22422 15536 22428 15548
rect 21735 15508 22428 15536
rect 21735 15505 21747 15508
rect 21689 15499 21747 15505
rect 22422 15496 22428 15508
rect 22480 15496 22486 15548
rect 11937 15471 11995 15477
rect 11937 15437 11949 15471
rect 11983 15468 11995 15471
rect 12026 15468 12032 15480
rect 11983 15440 12032 15468
rect 11983 15437 11995 15440
rect 11937 15431 11995 15437
rect 12026 15428 12032 15440
rect 12084 15428 12090 15480
rect 13222 15428 13228 15480
rect 13280 15468 13286 15480
rect 15709 15471 15767 15477
rect 15709 15468 15721 15471
rect 13280 15440 15721 15468
rect 13280 15428 13286 15440
rect 15709 15437 15721 15440
rect 15755 15437 15767 15471
rect 15709 15431 15767 15437
rect 17089 15471 17147 15477
rect 17089 15437 17101 15471
rect 17135 15468 17147 15471
rect 17178 15468 17184 15480
rect 17135 15440 17184 15468
rect 17135 15437 17147 15440
rect 17089 15431 17147 15437
rect 17178 15428 17184 15440
rect 17236 15428 17242 15480
rect 20306 15468 20312 15480
rect 20267 15440 20312 15468
rect 20306 15428 20312 15440
rect 20364 15428 20370 15480
rect 20398 15428 20404 15480
rect 20456 15468 20462 15480
rect 23268 15468 23296 15644
rect 23621 15641 23633 15644
rect 23667 15641 23679 15675
rect 23802 15672 23808 15684
rect 23763 15644 23808 15672
rect 23621 15635 23679 15641
rect 23802 15632 23808 15644
rect 23860 15632 23866 15684
rect 23912 15672 23940 15712
rect 27408 15712 27948 15740
rect 25461 15675 25519 15681
rect 25461 15672 25473 15675
rect 23912 15644 25473 15672
rect 25461 15641 25473 15644
rect 25507 15641 25519 15675
rect 25461 15635 25519 15641
rect 25553 15675 25611 15681
rect 25553 15641 25565 15675
rect 25599 15672 25611 15675
rect 25918 15672 25924 15684
rect 25599 15644 25924 15672
rect 25599 15641 25611 15644
rect 25553 15635 25611 15641
rect 25476 15536 25504 15635
rect 25918 15632 25924 15644
rect 25976 15632 25982 15684
rect 26010 15632 26016 15684
rect 26068 15672 26074 15684
rect 26197 15675 26255 15681
rect 26068 15644 26113 15672
rect 26068 15632 26074 15644
rect 26197 15641 26209 15675
rect 26243 15672 26255 15675
rect 27408 15672 27436 15712
rect 27942 15700 27948 15712
rect 28000 15700 28006 15752
rect 28678 15700 28684 15752
rect 28736 15700 28742 15752
rect 26243 15644 27436 15672
rect 26243 15641 26255 15644
rect 26197 15635 26255 15641
rect 27393 15607 27451 15613
rect 27393 15573 27405 15607
rect 27439 15573 27451 15607
rect 27393 15567 27451 15573
rect 27669 15607 27727 15613
rect 27669 15573 27681 15607
rect 27715 15604 27727 15607
rect 29138 15604 29144 15616
rect 27715 15576 29144 15604
rect 27715 15573 27727 15576
rect 27669 15567 27727 15573
rect 26010 15536 26016 15548
rect 25476 15508 26016 15536
rect 26010 15496 26016 15508
rect 26068 15496 26074 15548
rect 27408 15480 27436 15567
rect 29138 15564 29144 15576
rect 29196 15564 29202 15616
rect 29417 15607 29475 15613
rect 29417 15604 29429 15607
rect 29248 15576 29429 15604
rect 20456 15440 23296 15468
rect 20456 15428 20462 15440
rect 25550 15428 25556 15480
rect 25608 15468 25614 15480
rect 26473 15471 26531 15477
rect 26473 15468 26485 15471
rect 25608 15440 26485 15468
rect 25608 15428 25614 15440
rect 26473 15437 26485 15440
rect 26519 15437 26531 15471
rect 27390 15468 27396 15480
rect 27303 15440 27396 15468
rect 26473 15431 26531 15437
rect 27390 15428 27396 15440
rect 27448 15468 27454 15480
rect 27758 15468 27764 15480
rect 27448 15440 27764 15468
rect 27448 15428 27454 15440
rect 27758 15428 27764 15440
rect 27816 15428 27822 15480
rect 27850 15428 27856 15480
rect 27908 15468 27914 15480
rect 29248 15468 29276 15576
rect 29417 15573 29429 15576
rect 29463 15573 29475 15607
rect 29417 15567 29475 15573
rect 27908 15440 29276 15468
rect 27908 15428 27914 15440
rect 11000 15378 30136 15400
rect 11000 15326 14142 15378
rect 14194 15326 14206 15378
rect 14258 15326 14270 15378
rect 14322 15326 14334 15378
rect 14386 15326 24142 15378
rect 24194 15326 24206 15378
rect 24258 15326 24270 15378
rect 24322 15326 24334 15378
rect 24386 15326 30136 15378
rect 11000 15304 30136 15326
rect 13958 15224 13964 15276
rect 14016 15264 14022 15276
rect 18650 15264 18656 15276
rect 14016 15236 18656 15264
rect 14016 15224 14022 15236
rect 18650 15224 18656 15236
rect 18708 15224 18714 15276
rect 19018 15224 19024 15276
rect 19076 15264 19082 15276
rect 19113 15267 19171 15273
rect 19113 15264 19125 15267
rect 19076 15236 19125 15264
rect 19076 15224 19082 15236
rect 19113 15233 19125 15236
rect 19159 15233 19171 15267
rect 19113 15227 19171 15233
rect 19941 15267 19999 15273
rect 19941 15233 19953 15267
rect 19987 15264 19999 15267
rect 21410 15264 21416 15276
rect 19987 15236 21416 15264
rect 19987 15233 19999 15236
rect 19941 15227 19999 15233
rect 21410 15224 21416 15236
rect 21468 15224 21474 15276
rect 22514 15224 22520 15276
rect 22572 15264 22578 15276
rect 24173 15267 24231 15273
rect 24173 15264 24185 15267
rect 22572 15236 24185 15264
rect 22572 15224 22578 15236
rect 24173 15233 24185 15236
rect 24219 15233 24231 15267
rect 29138 15264 29144 15276
rect 29099 15236 29144 15264
rect 24173 15227 24231 15233
rect 29138 15224 29144 15236
rect 29196 15224 29202 15276
rect 21597 15199 21655 15205
rect 21597 15165 21609 15199
rect 21643 15196 21655 15199
rect 22974 15196 22980 15208
rect 21643 15168 22980 15196
rect 21643 15165 21655 15168
rect 21597 15159 21655 15165
rect 11934 15128 11940 15140
rect 11895 15100 11940 15128
rect 11934 15088 11940 15100
rect 11992 15088 11998 15140
rect 12946 15128 12952 15140
rect 12907 15100 12952 15128
rect 12946 15088 12952 15100
rect 13004 15088 13010 15140
rect 13222 15128 13228 15140
rect 13183 15100 13228 15128
rect 13222 15088 13228 15100
rect 13280 15088 13286 15140
rect 14786 15088 14792 15140
rect 14844 15128 14850 15140
rect 14973 15131 15031 15137
rect 14973 15128 14985 15131
rect 14844 15100 14985 15128
rect 14844 15088 14850 15100
rect 14973 15097 14985 15100
rect 15019 15097 15031 15131
rect 14973 15091 15031 15097
rect 11658 15060 11664 15072
rect 11619 15032 11664 15060
rect 11658 15020 11664 15032
rect 11716 15020 11722 15072
rect 11750 15020 11756 15072
rect 11808 15060 11814 15072
rect 11845 15063 11903 15069
rect 11845 15060 11857 15063
rect 11808 15032 11857 15060
rect 11808 15020 11814 15032
rect 11845 15029 11857 15032
rect 11891 15029 11903 15063
rect 14988 15060 15016 15091
rect 16074 15088 16080 15140
rect 16132 15128 16138 15140
rect 18558 15128 18564 15140
rect 16132 15100 18564 15128
rect 16132 15088 16138 15100
rect 18558 15088 18564 15100
rect 18616 15088 18622 15140
rect 21612 15128 21640 15159
rect 22974 15156 22980 15168
rect 23032 15196 23038 15208
rect 23032 15168 23848 15196
rect 23032 15156 23038 15168
rect 23820 15140 23848 15168
rect 20876 15100 21640 15128
rect 15433 15063 15491 15069
rect 15433 15060 15445 15063
rect 14988 15032 15445 15060
rect 11845 15023 11903 15029
rect 15433 15029 15445 15032
rect 15479 15029 15491 15063
rect 15433 15023 15491 15029
rect 11860 14924 11888 15023
rect 17178 15020 17184 15072
rect 17236 15060 17242 15072
rect 17273 15063 17331 15069
rect 17273 15060 17285 15063
rect 17236 15032 17285 15060
rect 17236 15020 17242 15032
rect 17273 15029 17285 15032
rect 17319 15029 17331 15063
rect 17273 15023 17331 15029
rect 17362 15020 17368 15072
rect 17420 15060 17426 15072
rect 17549 15063 17607 15069
rect 17549 15060 17561 15063
rect 17420 15032 17561 15060
rect 17420 15020 17426 15032
rect 17549 15029 17561 15032
rect 17595 15029 17607 15063
rect 17549 15023 17607 15029
rect 17733 15063 17791 15069
rect 17733 15029 17745 15063
rect 17779 15060 17791 15063
rect 18190 15060 18196 15072
rect 17779 15032 18196 15060
rect 17779 15029 17791 15032
rect 17733 15023 17791 15029
rect 18190 15020 18196 15032
rect 18248 15060 18254 15072
rect 19021 15063 19079 15069
rect 18248 15032 18880 15060
rect 18248 15020 18254 15032
rect 14234 14952 14240 15004
rect 14292 14952 14298 15004
rect 14602 14952 14608 15004
rect 14660 14992 14666 15004
rect 18852 15001 18880 15032
rect 19021 15029 19033 15063
rect 19067 15060 19079 15063
rect 19846 15060 19852 15072
rect 19067 15032 19852 15060
rect 19067 15029 19079 15032
rect 19021 15023 19079 15029
rect 19846 15020 19852 15032
rect 19904 15020 19910 15072
rect 20306 15020 20312 15072
rect 20364 15060 20370 15072
rect 20493 15063 20551 15069
rect 20493 15060 20505 15063
rect 20364 15032 20505 15060
rect 20364 15020 20370 15032
rect 20493 15029 20505 15032
rect 20539 15029 20551 15063
rect 20493 15023 20551 15029
rect 20582 15020 20588 15072
rect 20640 15060 20646 15072
rect 20876 15069 20904 15100
rect 22330 15088 22336 15140
rect 22388 15128 22394 15140
rect 23345 15131 23403 15137
rect 23345 15128 23357 15131
rect 22388 15100 23357 15128
rect 22388 15088 22394 15100
rect 23345 15097 23357 15100
rect 23391 15097 23403 15131
rect 23345 15091 23403 15097
rect 23802 15088 23808 15140
rect 23860 15128 23866 15140
rect 23897 15131 23955 15137
rect 23897 15128 23909 15131
rect 23860 15100 23909 15128
rect 23860 15088 23866 15100
rect 23897 15097 23909 15100
rect 23943 15097 23955 15131
rect 25550 15128 25556 15140
rect 25511 15100 25556 15128
rect 23897 15091 23955 15097
rect 25550 15088 25556 15100
rect 25608 15088 25614 15140
rect 25918 15088 25924 15140
rect 25976 15128 25982 15140
rect 27301 15131 27359 15137
rect 27301 15128 27313 15131
rect 25976 15100 27313 15128
rect 25976 15088 25982 15100
rect 27301 15097 27313 15100
rect 27347 15097 27359 15131
rect 27301 15091 27359 15097
rect 20861 15063 20919 15069
rect 20640 15032 20685 15060
rect 20640 15020 20646 15032
rect 20861 15029 20873 15063
rect 20907 15029 20919 15063
rect 20861 15023 20919 15029
rect 20953 15063 21011 15069
rect 20953 15029 20965 15063
rect 20999 15029 21011 15063
rect 20953 15023 21011 15029
rect 21505 15063 21563 15069
rect 21505 15029 21517 15063
rect 21551 15060 21563 15063
rect 22238 15060 22244 15072
rect 21551 15032 22244 15060
rect 21551 15029 21563 15032
rect 21505 15023 21563 15029
rect 16721 14995 16779 15001
rect 16721 14992 16733 14995
rect 14660 14964 16733 14992
rect 14660 14952 14666 14964
rect 16721 14961 16733 14964
rect 16767 14961 16779 14995
rect 16721 14955 16779 14961
rect 18837 14995 18895 15001
rect 18837 14961 18849 14995
rect 18883 14961 18895 14995
rect 18837 14955 18895 14961
rect 15338 14924 15344 14936
rect 11860 14896 15344 14924
rect 15338 14884 15344 14896
rect 15396 14884 15402 14936
rect 15522 14924 15528 14936
rect 15483 14896 15528 14924
rect 15522 14884 15528 14896
rect 15580 14884 15586 14936
rect 18282 14924 18288 14936
rect 18243 14896 18288 14924
rect 18282 14884 18288 14896
rect 18340 14884 18346 14936
rect 18852 14924 18880 14955
rect 18926 14952 18932 15004
rect 18984 14992 18990 15004
rect 20968 14992 20996 15023
rect 22238 15020 22244 15032
rect 22296 15020 22302 15072
rect 22422 15060 22428 15072
rect 22383 15032 22428 15060
rect 22422 15020 22428 15032
rect 22480 15020 22486 15072
rect 22606 15020 22612 15072
rect 22664 15060 22670 15072
rect 23253 15063 23311 15069
rect 23253 15060 23265 15063
rect 22664 15032 23265 15060
rect 22664 15020 22670 15032
rect 23253 15029 23265 15032
rect 23299 15029 23311 15063
rect 23253 15023 23311 15029
rect 23986 15020 23992 15072
rect 24044 15060 24050 15072
rect 25274 15060 25280 15072
rect 24044 15032 24089 15060
rect 25187 15032 25280 15060
rect 24044 15020 24050 15032
rect 25274 15020 25280 15032
rect 25332 15020 25338 15072
rect 27942 15060 27948 15072
rect 27903 15032 27948 15060
rect 27942 15020 27948 15032
rect 28000 15020 28006 15072
rect 28129 15063 28187 15069
rect 28129 15029 28141 15063
rect 28175 15029 28187 15063
rect 28586 15060 28592 15072
rect 28547 15032 28592 15060
rect 28129 15023 28187 15029
rect 18984 14964 20996 14992
rect 22517 14995 22575 15001
rect 18984 14952 18990 14964
rect 22517 14961 22529 14995
rect 22563 14992 22575 14995
rect 23802 14992 23808 15004
rect 22563 14964 23808 14992
rect 22563 14961 22575 14964
rect 22517 14955 22575 14961
rect 23802 14952 23808 14964
rect 23860 14952 23866 15004
rect 19018 14924 19024 14936
rect 18852 14896 19024 14924
rect 19018 14884 19024 14896
rect 19076 14884 19082 14936
rect 25292 14924 25320 15020
rect 26286 14952 26292 15004
rect 26344 14952 26350 15004
rect 27758 14952 27764 15004
rect 27816 14992 27822 15004
rect 28144 14992 28172 15023
rect 28586 15020 28592 15032
rect 28644 15020 28650 15072
rect 28681 15063 28739 15069
rect 28681 15029 28693 15063
rect 28727 15029 28739 15063
rect 28681 15023 28739 15029
rect 28696 14992 28724 15023
rect 27816 14964 28724 14992
rect 27816 14952 27822 14964
rect 26562 14924 26568 14936
rect 25292 14896 26568 14924
rect 26562 14884 26568 14896
rect 26620 14884 26626 14936
rect 11000 14834 30136 14856
rect 11000 14782 19142 14834
rect 19194 14782 19206 14834
rect 19258 14782 19270 14834
rect 19322 14782 19334 14834
rect 19386 14782 29142 14834
rect 29194 14782 29206 14834
rect 29258 14782 29270 14834
rect 29322 14782 29334 14834
rect 29386 14782 30136 14834
rect 11000 14760 30136 14782
rect 14145 14723 14203 14729
rect 14145 14689 14157 14723
rect 14191 14720 14203 14723
rect 14234 14720 14240 14732
rect 14191 14692 14240 14720
rect 14191 14689 14203 14692
rect 14145 14683 14203 14689
rect 14234 14680 14240 14692
rect 14292 14680 14298 14732
rect 15338 14680 15344 14732
rect 15396 14720 15402 14732
rect 18193 14723 18251 14729
rect 18193 14720 18205 14723
rect 15396 14692 18205 14720
rect 15396 14680 15402 14692
rect 18193 14689 18205 14692
rect 18239 14689 18251 14723
rect 18193 14683 18251 14689
rect 18558 14680 18564 14732
rect 18616 14720 18622 14732
rect 18929 14723 18987 14729
rect 18929 14720 18941 14723
rect 18616 14692 18941 14720
rect 18616 14680 18622 14692
rect 18929 14689 18941 14692
rect 18975 14689 18987 14723
rect 18929 14683 18987 14689
rect 23529 14723 23587 14729
rect 23529 14689 23541 14723
rect 23575 14720 23587 14723
rect 23986 14720 23992 14732
rect 23575 14692 23992 14720
rect 23575 14689 23587 14692
rect 23529 14683 23587 14689
rect 19846 14652 19852 14664
rect 15172 14624 16120 14652
rect 11934 14584 11940 14596
rect 11895 14556 11940 14584
rect 11934 14544 11940 14556
rect 11992 14544 11998 14596
rect 12305 14587 12363 14593
rect 12305 14553 12317 14587
rect 12351 14553 12363 14587
rect 12305 14547 12363 14553
rect 12026 14516 12032 14528
rect 11987 14488 12032 14516
rect 12026 14476 12032 14488
rect 12084 14476 12090 14528
rect 11566 14408 11572 14460
rect 11624 14448 11630 14460
rect 12320 14448 12348 14547
rect 12946 14544 12952 14596
rect 13004 14593 13010 14596
rect 13004 14584 13015 14593
rect 13004 14556 13049 14584
rect 13004 14547 13015 14556
rect 13004 14544 13010 14547
rect 13774 14544 13780 14596
rect 13832 14584 13838 14596
rect 15172 14593 15200 14624
rect 16092 14596 16120 14624
rect 17196 14624 17776 14652
rect 17196 14596 17224 14624
rect 13961 14587 14019 14593
rect 13961 14584 13973 14587
rect 13832 14556 13973 14584
rect 13832 14544 13838 14556
rect 13961 14553 13973 14556
rect 14007 14553 14019 14587
rect 13961 14547 14019 14553
rect 15157 14587 15215 14593
rect 15157 14553 15169 14587
rect 15203 14553 15215 14587
rect 15157 14547 15215 14553
rect 15341 14587 15399 14593
rect 15341 14553 15353 14587
rect 15387 14584 15399 14587
rect 15522 14584 15528 14596
rect 15387 14556 15528 14584
rect 15387 14553 15399 14556
rect 15341 14547 15399 14553
rect 15522 14544 15528 14556
rect 15580 14584 15586 14596
rect 15890 14584 15896 14596
rect 15580 14556 15896 14584
rect 15580 14544 15586 14556
rect 15890 14544 15896 14556
rect 15948 14544 15954 14596
rect 16074 14584 16080 14596
rect 16035 14556 16080 14584
rect 16074 14544 16080 14556
rect 16132 14584 16138 14596
rect 16442 14584 16448 14596
rect 16132 14556 16448 14584
rect 16132 14544 16138 14556
rect 16442 14544 16448 14556
rect 16500 14544 16506 14596
rect 17178 14584 17184 14596
rect 17139 14556 17184 14584
rect 17178 14544 17184 14556
rect 17236 14544 17242 14596
rect 17748 14593 17776 14624
rect 18852 14624 19852 14652
rect 18852 14593 18880 14624
rect 19846 14612 19852 14624
rect 19904 14612 19910 14664
rect 23544 14652 23572 14683
rect 23986 14680 23992 14692
rect 24044 14680 24050 14732
rect 25918 14680 25924 14732
rect 25976 14720 25982 14732
rect 26473 14723 26531 14729
rect 26473 14720 26485 14723
rect 25976 14692 26485 14720
rect 25976 14680 25982 14692
rect 26473 14689 26485 14692
rect 26519 14689 26531 14723
rect 27942 14720 27948 14732
rect 26473 14683 26531 14689
rect 26580 14692 27948 14720
rect 26580 14661 26608 14692
rect 27942 14680 27948 14692
rect 28000 14720 28006 14732
rect 28000 14692 29644 14720
rect 28000 14680 28006 14692
rect 22808 14624 23572 14652
rect 26565 14655 26623 14661
rect 17641 14587 17699 14593
rect 17641 14584 17653 14587
rect 17288 14556 17653 14584
rect 12394 14476 12400 14528
rect 12452 14516 12458 14528
rect 14602 14516 14608 14528
rect 12452 14488 14608 14516
rect 12452 14476 12458 14488
rect 14602 14476 14608 14488
rect 14660 14476 14666 14528
rect 16997 14519 17055 14525
rect 16997 14485 17009 14519
rect 17043 14516 17055 14519
rect 17288 14516 17316 14556
rect 17641 14553 17653 14556
rect 17687 14553 17699 14587
rect 17641 14547 17699 14553
rect 17733 14587 17791 14593
rect 17733 14553 17745 14587
rect 17779 14553 17791 14587
rect 17733 14547 17791 14553
rect 18837 14587 18895 14593
rect 18837 14553 18849 14587
rect 18883 14553 18895 14587
rect 18837 14547 18895 14553
rect 19757 14587 19815 14593
rect 19757 14553 19769 14587
rect 19803 14584 19815 14587
rect 20306 14584 20312 14596
rect 19803 14556 20312 14584
rect 19803 14553 19815 14556
rect 19757 14547 19815 14553
rect 20306 14544 20312 14556
rect 20364 14544 20370 14596
rect 22425 14587 22483 14593
rect 22425 14553 22437 14587
rect 22471 14584 22483 14587
rect 22606 14584 22612 14596
rect 22471 14556 22612 14584
rect 22471 14553 22483 14556
rect 22425 14547 22483 14553
rect 22606 14544 22612 14556
rect 22664 14544 22670 14596
rect 22808 14593 22836 14624
rect 26565 14621 26577 14655
rect 26611 14621 26623 14655
rect 26565 14615 26623 14621
rect 26933 14655 26991 14661
rect 26933 14621 26945 14655
rect 26979 14652 26991 14655
rect 27022 14652 27028 14664
rect 26979 14624 27028 14652
rect 26979 14621 26991 14624
rect 26933 14615 26991 14621
rect 27022 14612 27028 14624
rect 27080 14612 27086 14664
rect 27758 14652 27764 14664
rect 27408 14624 27764 14652
rect 22793 14587 22851 14593
rect 22793 14553 22805 14587
rect 22839 14553 22851 14587
rect 22974 14584 22980 14596
rect 22935 14556 22980 14584
rect 22793 14547 22851 14553
rect 22974 14544 22980 14556
rect 23032 14544 23038 14596
rect 23158 14544 23164 14596
rect 23216 14584 23222 14596
rect 23437 14587 23495 14593
rect 23437 14584 23449 14587
rect 23216 14556 23449 14584
rect 23216 14544 23222 14556
rect 23437 14553 23449 14556
rect 23483 14553 23495 14587
rect 25274 14584 25280 14596
rect 25235 14556 25280 14584
rect 23437 14547 23495 14553
rect 25274 14544 25280 14556
rect 25332 14544 25338 14596
rect 26381 14587 26439 14593
rect 26381 14584 26393 14587
rect 26120 14556 26393 14584
rect 17043 14488 17316 14516
rect 19665 14519 19723 14525
rect 17043 14485 17055 14488
rect 16997 14479 17055 14485
rect 19665 14485 19677 14519
rect 19711 14516 19723 14519
rect 20030 14516 20036 14528
rect 19711 14488 20036 14516
rect 19711 14485 19723 14488
rect 19665 14479 19723 14485
rect 12946 14448 12952 14460
rect 11624 14420 12348 14448
rect 12688 14420 12952 14448
rect 11624 14408 11630 14420
rect 11385 14383 11443 14389
rect 11385 14349 11397 14383
rect 11431 14380 11443 14383
rect 12688 14380 12716 14420
rect 12946 14408 12952 14420
rect 13004 14408 13010 14460
rect 16258 14448 16264 14460
rect 16219 14420 16264 14448
rect 16258 14408 16264 14420
rect 16316 14448 16322 14460
rect 17012 14448 17040 14479
rect 20030 14476 20036 14488
rect 20088 14476 20094 14528
rect 22514 14516 22520 14528
rect 22475 14488 22520 14516
rect 22514 14476 22520 14488
rect 22572 14476 22578 14528
rect 23894 14476 23900 14528
rect 23952 14516 23958 14528
rect 25185 14519 25243 14525
rect 25185 14516 25197 14519
rect 23952 14488 25197 14516
rect 23952 14476 23958 14488
rect 25185 14485 25197 14488
rect 25231 14485 25243 14519
rect 25185 14479 25243 14485
rect 16316 14420 17040 14448
rect 16316 14408 16322 14420
rect 20582 14408 20588 14460
rect 20640 14448 20646 14460
rect 25918 14448 25924 14460
rect 20640 14420 25924 14448
rect 20640 14408 20646 14420
rect 25918 14408 25924 14420
rect 25976 14448 25982 14460
rect 26120 14448 26148 14556
rect 26381 14553 26393 14556
rect 26427 14584 26439 14587
rect 27408 14584 27436 14624
rect 27758 14612 27764 14624
rect 27816 14612 27822 14664
rect 29506 14652 29512 14664
rect 28894 14624 29512 14652
rect 29506 14612 29512 14624
rect 29564 14612 29570 14664
rect 26427 14556 27436 14584
rect 29417 14587 29475 14593
rect 26427 14553 26439 14556
rect 26381 14547 26439 14553
rect 29417 14553 29429 14587
rect 29463 14584 29475 14587
rect 29616 14584 29644 14692
rect 29463 14556 29644 14584
rect 29463 14553 29475 14556
rect 29417 14547 29475 14553
rect 26197 14519 26255 14525
rect 26197 14485 26209 14519
rect 26243 14485 26255 14519
rect 26197 14479 26255 14485
rect 25976 14420 26148 14448
rect 25976 14408 25982 14420
rect 11431 14352 12716 14380
rect 11431 14349 11443 14352
rect 11385 14343 11443 14349
rect 12762 14340 12768 14392
rect 12820 14380 12826 14392
rect 13041 14383 13099 14389
rect 13041 14380 13053 14383
rect 12820 14352 13053 14380
rect 12820 14340 12826 14352
rect 13041 14349 13053 14352
rect 13087 14349 13099 14383
rect 13041 14343 13099 14349
rect 18926 14340 18932 14392
rect 18984 14380 18990 14392
rect 19941 14383 19999 14389
rect 19941 14380 19953 14383
rect 18984 14352 19953 14380
rect 18984 14340 18990 14352
rect 19941 14349 19953 14352
rect 19987 14349 19999 14383
rect 22054 14380 22060 14392
rect 22015 14352 22060 14380
rect 19941 14343 19999 14349
rect 22054 14340 22060 14352
rect 22112 14340 22118 14392
rect 25458 14380 25464 14392
rect 25419 14352 25464 14380
rect 25458 14340 25464 14352
rect 25516 14340 25522 14392
rect 26212 14380 26240 14479
rect 26562 14476 26568 14528
rect 26620 14516 26626 14528
rect 27390 14516 27396 14528
rect 26620 14488 27396 14516
rect 26620 14476 26626 14488
rect 27390 14476 27396 14488
rect 27448 14476 27454 14528
rect 27669 14519 27727 14525
rect 27669 14485 27681 14519
rect 27715 14516 27727 14519
rect 28218 14516 28224 14528
rect 27715 14488 28224 14516
rect 27715 14485 27727 14488
rect 27669 14479 27727 14485
rect 28218 14476 28224 14488
rect 28276 14476 28282 14528
rect 27850 14380 27856 14392
rect 26212 14352 27856 14380
rect 27850 14340 27856 14352
rect 27908 14340 27914 14392
rect 11000 14290 30136 14312
rect 11000 14238 14142 14290
rect 14194 14238 14206 14290
rect 14258 14238 14270 14290
rect 14322 14238 14334 14290
rect 14386 14238 24142 14290
rect 24194 14238 24206 14290
rect 24258 14238 24270 14290
rect 24322 14238 24334 14290
rect 24386 14238 30136 14290
rect 11000 14216 30136 14238
rect 13038 14176 13044 14188
rect 12999 14148 13044 14176
rect 13038 14136 13044 14148
rect 13096 14136 13102 14188
rect 13866 14136 13872 14188
rect 13924 14176 13930 14188
rect 14881 14179 14939 14185
rect 14881 14176 14893 14179
rect 13924 14148 14893 14176
rect 13924 14136 13930 14148
rect 14881 14145 14893 14148
rect 14927 14145 14939 14179
rect 14881 14139 14939 14145
rect 16810 14136 16816 14188
rect 16868 14176 16874 14188
rect 17914 14176 17920 14188
rect 16868 14148 17920 14176
rect 16868 14136 16874 14148
rect 17914 14136 17920 14148
rect 17972 14136 17978 14188
rect 22422 14136 22428 14188
rect 22480 14176 22486 14188
rect 22609 14179 22667 14185
rect 22609 14176 22621 14179
rect 22480 14148 22621 14176
rect 22480 14136 22486 14148
rect 22609 14145 22621 14148
rect 22655 14145 22667 14179
rect 28218 14176 28224 14188
rect 28179 14148 28224 14176
rect 22609 14139 22667 14145
rect 28218 14136 28224 14148
rect 28276 14136 28282 14188
rect 28862 14136 28868 14188
rect 28920 14176 28926 14188
rect 28957 14179 29015 14185
rect 28957 14176 28969 14179
rect 28920 14148 28969 14176
rect 28920 14136 28926 14148
rect 28957 14145 28969 14148
rect 29003 14145 29015 14179
rect 28957 14139 29015 14145
rect 25458 14108 25464 14120
rect 18852 14080 25464 14108
rect 12394 14040 12400 14052
rect 11952 14012 12400 14040
rect 11566 13972 11572 13984
rect 11527 13944 11572 13972
rect 11566 13932 11572 13944
rect 11624 13932 11630 13984
rect 11952 13981 11980 14012
rect 12394 14000 12400 14012
rect 12452 14000 12458 14052
rect 18852 14040 18880 14080
rect 25458 14068 25464 14080
rect 25516 14068 25522 14120
rect 13608 14012 18880 14040
rect 24633 14043 24691 14049
rect 11937 13975 11995 13981
rect 11937 13941 11949 13975
rect 11983 13941 11995 13975
rect 11937 13935 11995 13941
rect 12305 13975 12363 13981
rect 12305 13941 12317 13975
rect 12351 13972 12363 13975
rect 12762 13972 12768 13984
rect 12351 13944 12768 13972
rect 12351 13941 12363 13944
rect 12305 13935 12363 13941
rect 12762 13932 12768 13944
rect 12820 13932 12826 13984
rect 13608 13981 13636 14012
rect 24633 14009 24645 14043
rect 24679 14040 24691 14043
rect 24679 14012 25504 14040
rect 24679 14009 24691 14012
rect 24633 14003 24691 14009
rect 25476 13984 25504 14012
rect 27942 14000 27948 14052
rect 28000 14040 28006 14052
rect 28000 14012 28172 14040
rect 28000 14000 28006 14012
rect 13593 13975 13651 13981
rect 13593 13941 13605 13975
rect 13639 13941 13651 13975
rect 13593 13935 13651 13941
rect 13682 13932 13688 13984
rect 13740 13972 13746 13984
rect 13740 13944 13785 13972
rect 13740 13932 13746 13944
rect 13866 13932 13872 13984
rect 13924 13972 13930 13984
rect 13961 13975 14019 13981
rect 13961 13972 13973 13975
rect 13924 13944 13973 13972
rect 13924 13932 13930 13944
rect 13961 13941 13973 13944
rect 14007 13941 14019 13975
rect 13961 13935 14019 13941
rect 14145 13975 14203 13981
rect 14145 13941 14157 13975
rect 14191 13972 14203 13975
rect 14191 13944 14740 13972
rect 14191 13941 14203 13944
rect 14145 13935 14203 13941
rect 12489 13907 12547 13913
rect 12489 13873 12501 13907
rect 12535 13904 12547 13907
rect 14234 13904 14240 13916
rect 12535 13876 14240 13904
rect 12535 13873 12547 13876
rect 12489 13867 12547 13873
rect 14234 13864 14240 13876
rect 14292 13864 14298 13916
rect 14605 13907 14663 13913
rect 14605 13904 14617 13907
rect 14344 13876 14617 13904
rect 13958 13796 13964 13848
rect 14016 13836 14022 13848
rect 14344 13836 14372 13876
rect 14605 13873 14617 13876
rect 14651 13873 14663 13907
rect 14712 13904 14740 13944
rect 14786 13932 14792 13984
rect 14844 13972 14850 13984
rect 15617 13975 15675 13981
rect 14844 13944 14889 13972
rect 14844 13932 14850 13944
rect 15617 13941 15629 13975
rect 15663 13941 15675 13975
rect 16810 13972 16816 13984
rect 16771 13944 16816 13972
rect 15617 13935 15675 13941
rect 15632 13904 15660 13935
rect 16810 13932 16816 13944
rect 16868 13932 16874 13984
rect 16902 13932 16908 13984
rect 16960 13972 16966 13984
rect 17546 13972 17552 13984
rect 16960 13944 17552 13972
rect 16960 13932 16966 13944
rect 17546 13932 17552 13944
rect 17604 13932 17610 13984
rect 19110 13932 19116 13984
rect 19168 13972 19174 13984
rect 19573 13975 19631 13981
rect 19573 13972 19585 13975
rect 19168 13944 19585 13972
rect 19168 13932 19174 13944
rect 19573 13941 19585 13944
rect 19619 13941 19631 13975
rect 20030 13972 20036 13984
rect 19991 13944 20036 13972
rect 19573 13935 19631 13941
rect 20030 13932 20036 13944
rect 20088 13932 20094 13984
rect 20217 13975 20275 13981
rect 20217 13941 20229 13975
rect 20263 13972 20275 13975
rect 20306 13972 20312 13984
rect 20263 13944 20312 13972
rect 20263 13941 20275 13944
rect 20217 13935 20275 13941
rect 20306 13932 20312 13944
rect 20364 13932 20370 13984
rect 20766 13972 20772 13984
rect 20727 13944 20772 13972
rect 20766 13932 20772 13944
rect 20824 13932 20830 13984
rect 22330 13932 22336 13984
rect 22388 13972 22394 13984
rect 22517 13975 22575 13981
rect 22388 13944 22433 13972
rect 22388 13932 22394 13944
rect 22517 13941 22529 13975
rect 22563 13972 22575 13975
rect 22606 13972 22612 13984
rect 22563 13944 22612 13972
rect 22563 13941 22575 13944
rect 22517 13935 22575 13941
rect 22606 13932 22612 13944
rect 22664 13932 22670 13984
rect 23802 13932 23808 13984
rect 23860 13972 23866 13984
rect 24173 13975 24231 13981
rect 24173 13972 24185 13975
rect 23860 13944 24185 13972
rect 23860 13932 23866 13944
rect 24173 13941 24185 13944
rect 24219 13941 24231 13975
rect 24173 13935 24231 13941
rect 24817 13975 24875 13981
rect 24817 13941 24829 13975
rect 24863 13941 24875 13975
rect 25090 13972 25096 13984
rect 25051 13944 25096 13972
rect 24817 13935 24875 13941
rect 17270 13904 17276 13916
rect 14712 13876 17276 13904
rect 14605 13867 14663 13873
rect 17270 13864 17276 13876
rect 17328 13864 17334 13916
rect 17730 13864 17736 13916
rect 17788 13904 17794 13916
rect 17825 13907 17883 13913
rect 17825 13904 17837 13907
rect 17788 13876 17837 13904
rect 17788 13864 17794 13876
rect 17825 13873 17837 13876
rect 17871 13873 17883 13907
rect 20398 13904 20404 13916
rect 17825 13867 17883 13873
rect 14016 13808 14372 13836
rect 14016 13796 14022 13808
rect 14970 13796 14976 13848
rect 15028 13836 15034 13848
rect 15709 13839 15767 13845
rect 15709 13836 15721 13839
rect 15028 13808 15721 13836
rect 15028 13796 15034 13808
rect 15709 13805 15721 13808
rect 15755 13805 15767 13839
rect 15709 13799 15767 13805
rect 16997 13839 17055 13845
rect 16997 13805 17009 13839
rect 17043 13836 17055 13839
rect 18300 13836 18328 13890
rect 20359 13876 20404 13904
rect 20398 13864 20404 13876
rect 20456 13864 20462 13916
rect 17043 13808 18328 13836
rect 17043 13805 17055 13808
rect 16997 13799 17055 13805
rect 18742 13796 18748 13848
rect 18800 13836 18806 13848
rect 20309 13839 20367 13845
rect 20309 13836 20321 13839
rect 18800 13808 20321 13836
rect 18800 13796 18806 13808
rect 20309 13805 20321 13808
rect 20355 13805 20367 13839
rect 20309 13799 20367 13805
rect 24262 13796 24268 13848
rect 24320 13836 24326 13848
rect 24832 13836 24860 13935
rect 25090 13932 25096 13944
rect 25148 13932 25154 13984
rect 25369 13975 25427 13981
rect 25369 13941 25381 13975
rect 25415 13941 25427 13975
rect 25369 13935 25427 13941
rect 24906 13864 24912 13916
rect 24964 13904 24970 13916
rect 25384 13904 25412 13935
rect 25458 13932 25464 13984
rect 25516 13932 25522 13984
rect 28144 13981 28172 14012
rect 28129 13975 28187 13981
rect 28129 13941 28141 13975
rect 28175 13941 28187 13975
rect 28129 13935 28187 13941
rect 28494 13932 28500 13984
rect 28552 13972 28558 13984
rect 29141 13975 29199 13981
rect 29141 13972 29153 13975
rect 28552 13944 29153 13972
rect 28552 13932 28558 13944
rect 29141 13941 29153 13944
rect 29187 13941 29199 13975
rect 29141 13935 29199 13941
rect 24964 13876 25412 13904
rect 24964 13864 24970 13876
rect 27850 13864 27856 13916
rect 27908 13904 27914 13916
rect 27945 13907 28003 13913
rect 27945 13904 27957 13907
rect 27908 13876 27957 13904
rect 27908 13864 27914 13876
rect 27945 13873 27957 13876
rect 27991 13873 28003 13907
rect 27945 13867 28003 13873
rect 25182 13836 25188 13848
rect 24320 13808 25188 13836
rect 24320 13796 24326 13808
rect 25182 13796 25188 13808
rect 25240 13796 25246 13848
rect 11000 13746 30136 13768
rect 11000 13694 19142 13746
rect 19194 13694 19206 13746
rect 19258 13694 19270 13746
rect 19322 13694 19334 13746
rect 19386 13694 29142 13746
rect 29194 13694 29206 13746
rect 29258 13694 29270 13746
rect 29322 13694 29334 13746
rect 29386 13694 30136 13746
rect 11000 13672 30136 13694
rect 15801 13635 15859 13641
rect 15801 13601 15813 13635
rect 15847 13632 15859 13635
rect 15847 13604 19524 13632
rect 15847 13601 15859 13604
rect 15801 13595 15859 13601
rect 12305 13567 12363 13573
rect 12305 13533 12317 13567
rect 12351 13564 12363 13567
rect 12762 13564 12768 13576
rect 12351 13536 12768 13564
rect 12351 13533 12363 13536
rect 12305 13527 12363 13533
rect 12762 13524 12768 13536
rect 12820 13524 12826 13576
rect 12857 13567 12915 13573
rect 12857 13533 12869 13567
rect 12903 13564 12915 13567
rect 13866 13564 13872 13576
rect 12903 13536 13872 13564
rect 12903 13533 12915 13536
rect 12857 13527 12915 13533
rect 13866 13524 13872 13536
rect 13924 13524 13930 13576
rect 14697 13567 14755 13573
rect 14697 13533 14709 13567
rect 14743 13564 14755 13567
rect 14878 13564 14884 13576
rect 14743 13536 14884 13564
rect 14743 13533 14755 13536
rect 14697 13527 14755 13533
rect 14878 13524 14884 13536
rect 14936 13524 14942 13576
rect 15890 13524 15896 13576
rect 15948 13564 15954 13576
rect 17730 13564 17736 13576
rect 15948 13536 16580 13564
rect 17691 13536 17736 13564
rect 15948 13524 15954 13536
rect 12026 13456 12032 13508
rect 12084 13496 12090 13508
rect 12489 13499 12547 13505
rect 12489 13496 12501 13499
rect 12084 13468 12501 13496
rect 12084 13456 12090 13468
rect 12489 13465 12501 13468
rect 12535 13465 12547 13499
rect 12489 13459 12547 13465
rect 13130 13456 13136 13508
rect 13188 13496 13194 13508
rect 13958 13496 13964 13508
rect 13188 13468 13964 13496
rect 13188 13456 13194 13468
rect 13958 13456 13964 13468
rect 14016 13456 14022 13508
rect 16552 13505 16580 13536
rect 17730 13524 17736 13536
rect 17788 13524 17794 13576
rect 19496 13564 19524 13604
rect 19570 13592 19576 13644
rect 19628 13632 19634 13644
rect 19665 13635 19723 13641
rect 19665 13632 19677 13635
rect 19628 13604 19677 13632
rect 19628 13592 19634 13604
rect 19665 13601 19677 13604
rect 19711 13601 19723 13635
rect 22606 13632 22612 13644
rect 19665 13595 19723 13601
rect 19772 13604 22612 13632
rect 19772 13564 19800 13604
rect 22606 13592 22612 13604
rect 22664 13592 22670 13644
rect 23529 13635 23587 13641
rect 23529 13601 23541 13635
rect 23575 13632 23587 13635
rect 23894 13632 23900 13644
rect 23575 13604 23900 13632
rect 23575 13601 23587 13604
rect 23529 13595 23587 13601
rect 23894 13592 23900 13604
rect 23952 13592 23958 13644
rect 29233 13635 29291 13641
rect 29233 13601 29245 13635
rect 29279 13632 29291 13635
rect 29506 13632 29512 13644
rect 29279 13604 29512 13632
rect 29279 13601 29291 13604
rect 29233 13595 29291 13601
rect 29506 13592 29512 13604
rect 29564 13592 29570 13644
rect 28126 13564 28132 13576
rect 19496 13536 19800 13564
rect 21428 13536 22008 13564
rect 16169 13499 16227 13505
rect 16169 13465 16181 13499
rect 16215 13496 16227 13499
rect 16537 13499 16595 13505
rect 16215 13468 16396 13496
rect 16215 13465 16227 13468
rect 16169 13459 16227 13465
rect 14329 13431 14387 13437
rect 14329 13397 14341 13431
rect 14375 13428 14387 13431
rect 14970 13428 14976 13440
rect 14375 13400 14976 13428
rect 14375 13397 14387 13400
rect 14329 13391 14387 13397
rect 14970 13388 14976 13400
rect 15028 13388 15034 13440
rect 16258 13428 16264 13440
rect 16219 13400 16264 13428
rect 16258 13388 16264 13400
rect 16316 13388 16322 13440
rect 14234 13360 14240 13372
rect 14195 13332 14240 13360
rect 14234 13320 14240 13332
rect 14292 13320 14298 13372
rect 16368 13360 16396 13468
rect 16537 13465 16549 13499
rect 16583 13465 16595 13499
rect 18374 13496 18380 13508
rect 18335 13468 18380 13496
rect 16537 13459 16595 13465
rect 18374 13456 18380 13468
rect 18432 13456 18438 13508
rect 18742 13496 18748 13508
rect 18703 13468 18748 13496
rect 18742 13456 18748 13468
rect 18800 13456 18806 13508
rect 18926 13496 18932 13508
rect 18887 13468 18932 13496
rect 18926 13456 18932 13468
rect 18984 13456 18990 13508
rect 19849 13499 19907 13505
rect 19849 13465 19861 13499
rect 19895 13496 19907 13499
rect 20030 13496 20036 13508
rect 19895 13468 20036 13496
rect 19895 13465 19907 13468
rect 19849 13459 19907 13465
rect 20030 13456 20036 13468
rect 20088 13456 20094 13508
rect 20125 13499 20183 13505
rect 20125 13465 20137 13499
rect 20171 13496 20183 13499
rect 20306 13496 20312 13508
rect 20171 13468 20312 13496
rect 20171 13465 20183 13468
rect 20125 13459 20183 13465
rect 20306 13456 20312 13468
rect 20364 13456 20370 13508
rect 21134 13456 21140 13508
rect 21192 13496 21198 13508
rect 21428 13505 21456 13536
rect 21980 13505 22008 13536
rect 23452 13536 25504 13564
rect 28066 13536 28132 13564
rect 21413 13499 21471 13505
rect 21413 13496 21425 13499
rect 21192 13468 21425 13496
rect 21192 13456 21198 13468
rect 21413 13465 21425 13468
rect 21459 13465 21471 13499
rect 21873 13499 21931 13505
rect 21873 13496 21885 13499
rect 21413 13459 21471 13465
rect 21612 13468 21885 13496
rect 16442 13388 16448 13440
rect 16500 13428 16506 13440
rect 18282 13428 18288 13440
rect 16500 13400 16545 13428
rect 18243 13400 18288 13428
rect 16500 13388 16506 13400
rect 18282 13388 18288 13400
rect 18340 13388 18346 13440
rect 21226 13428 21232 13440
rect 21187 13400 21232 13428
rect 21226 13388 21232 13400
rect 21284 13428 21290 13440
rect 21612 13428 21640 13468
rect 21873 13465 21885 13468
rect 21919 13465 21931 13499
rect 21873 13459 21931 13465
rect 21965 13499 22023 13505
rect 21965 13465 21977 13499
rect 22011 13496 22023 13499
rect 22054 13496 22060 13508
rect 22011 13468 22060 13496
rect 22011 13465 22023 13468
rect 21965 13459 22023 13465
rect 22054 13456 22060 13468
rect 22112 13456 22118 13508
rect 23452 13505 23480 13536
rect 25476 13508 25504 13536
rect 28126 13524 28132 13536
rect 28184 13524 28190 13576
rect 23437 13499 23495 13505
rect 23437 13465 23449 13499
rect 23483 13465 23495 13499
rect 23437 13459 23495 13465
rect 23802 13456 23808 13508
rect 23860 13496 23866 13508
rect 24081 13499 24139 13505
rect 24081 13496 24093 13499
rect 23860 13468 24093 13496
rect 23860 13456 23866 13468
rect 24081 13465 24093 13468
rect 24127 13465 24139 13499
rect 24262 13496 24268 13508
rect 24223 13468 24268 13496
rect 24081 13459 24139 13465
rect 24262 13456 24268 13468
rect 24320 13456 24326 13508
rect 24633 13499 24691 13505
rect 24633 13465 24645 13499
rect 24679 13496 24691 13499
rect 25369 13499 25427 13505
rect 25369 13496 25381 13499
rect 24679 13468 25381 13496
rect 24679 13465 24691 13468
rect 24633 13459 24691 13465
rect 25369 13465 25381 13468
rect 25415 13465 25427 13499
rect 25369 13459 25427 13465
rect 25458 13456 25464 13508
rect 25516 13496 25522 13508
rect 26562 13496 26568 13508
rect 25516 13468 25561 13496
rect 26523 13468 26568 13496
rect 25516 13456 25522 13468
rect 26562 13456 26568 13468
rect 26620 13456 26626 13508
rect 28954 13456 28960 13508
rect 29012 13496 29018 13508
rect 29049 13499 29107 13505
rect 29049 13496 29061 13499
rect 29012 13468 29061 13496
rect 29012 13456 29018 13468
rect 29049 13465 29061 13468
rect 29095 13465 29107 13499
rect 29049 13459 29107 13465
rect 21284 13400 21640 13428
rect 25185 13431 25243 13437
rect 21284 13388 21290 13400
rect 25185 13397 25197 13431
rect 25231 13428 25243 13431
rect 25274 13428 25280 13440
rect 25231 13400 25280 13428
rect 25231 13397 25243 13400
rect 25185 13391 25243 13397
rect 25274 13388 25280 13400
rect 25332 13388 25338 13440
rect 26841 13431 26899 13437
rect 26841 13397 26853 13431
rect 26887 13428 26899 13431
rect 27482 13428 27488 13440
rect 26887 13400 27488 13428
rect 26887 13397 26899 13400
rect 26841 13391 26899 13397
rect 27482 13388 27488 13400
rect 27540 13388 27546 13440
rect 28586 13428 28592 13440
rect 28547 13400 28592 13428
rect 28586 13388 28592 13400
rect 28644 13388 28650 13440
rect 17178 13360 17184 13372
rect 16368 13332 17184 13360
rect 17178 13320 17184 13332
rect 17236 13320 17242 13372
rect 17270 13320 17276 13372
rect 17328 13360 17334 13372
rect 17328 13332 25688 13360
rect 17328 13320 17334 13332
rect 12946 13252 12952 13304
rect 13004 13292 13010 13304
rect 13682 13292 13688 13304
rect 13004 13264 13688 13292
rect 13004 13252 13010 13264
rect 13682 13252 13688 13264
rect 13740 13292 13746 13304
rect 14099 13295 14157 13301
rect 14099 13292 14111 13295
rect 13740 13264 14111 13292
rect 13740 13252 13746 13264
rect 14099 13261 14111 13264
rect 14145 13261 14157 13295
rect 14099 13255 14157 13261
rect 22425 13295 22483 13301
rect 22425 13261 22437 13295
rect 22471 13292 22483 13295
rect 24906 13292 24912 13304
rect 22471 13264 24912 13292
rect 22471 13261 22483 13264
rect 22425 13255 22483 13261
rect 24906 13252 24912 13264
rect 24964 13252 24970 13304
rect 25660 13301 25688 13332
rect 25645 13295 25703 13301
rect 25645 13261 25657 13295
rect 25691 13261 25703 13295
rect 25645 13255 25703 13261
rect 11000 13202 30136 13224
rect 11000 13150 14142 13202
rect 14194 13150 14206 13202
rect 14258 13150 14270 13202
rect 14322 13150 14334 13202
rect 14386 13150 24142 13202
rect 24194 13150 24206 13202
rect 24258 13150 24270 13202
rect 24322 13150 24334 13202
rect 24386 13150 30136 13202
rect 11000 13128 30136 13150
rect 18374 13048 18380 13100
rect 18432 13088 18438 13100
rect 20582 13088 20588 13100
rect 18432 13060 20588 13088
rect 18432 13048 18438 13060
rect 14513 13023 14571 13029
rect 14513 13020 14525 13023
rect 13240 12992 14525 13020
rect 12946 12952 12952 12964
rect 12907 12924 12952 12952
rect 12946 12912 12952 12924
rect 13004 12912 13010 12964
rect 12026 12844 12032 12896
rect 12084 12884 12090 12896
rect 12397 12887 12455 12893
rect 12397 12884 12409 12887
rect 12084 12856 12409 12884
rect 12084 12844 12090 12856
rect 12397 12853 12409 12856
rect 12443 12853 12455 12887
rect 12397 12847 12455 12853
rect 12489 12887 12547 12893
rect 12489 12853 12501 12887
rect 12535 12884 12547 12887
rect 12578 12884 12584 12896
rect 12535 12856 12584 12884
rect 12535 12853 12547 12856
rect 12489 12847 12547 12853
rect 12578 12844 12584 12856
rect 12636 12884 12642 12896
rect 13240 12884 13268 12992
rect 14513 12989 14525 12992
rect 14559 12989 14571 13023
rect 14513 12983 14571 12989
rect 13406 12952 13412 12964
rect 13367 12924 13412 12952
rect 13406 12912 13412 12924
rect 13464 12952 13470 12964
rect 18834 12952 18840 12964
rect 13464 12924 13820 12952
rect 13464 12912 13470 12924
rect 12636 12856 13268 12884
rect 13593 12887 13651 12893
rect 12636 12844 12642 12856
rect 13593 12853 13605 12887
rect 13639 12884 13651 12887
rect 13792 12884 13820 12924
rect 14896 12924 18840 12952
rect 14053 12887 14111 12893
rect 14053 12884 14065 12887
rect 13639 12856 13728 12884
rect 13792 12856 14065 12884
rect 13639 12853 13651 12856
rect 13593 12847 13651 12853
rect 13314 12708 13320 12760
rect 13372 12748 13378 12760
rect 13700 12748 13728 12856
rect 14053 12853 14065 12856
rect 14099 12853 14111 12887
rect 14053 12847 14111 12853
rect 14142 12844 14148 12896
rect 14200 12884 14206 12896
rect 14200 12856 14245 12884
rect 14200 12844 14206 12856
rect 14326 12844 14332 12896
rect 14384 12884 14390 12896
rect 14896 12884 14924 12924
rect 18834 12912 18840 12924
rect 18892 12912 18898 12964
rect 18944 12961 18972 13060
rect 20582 13048 20588 13060
rect 20640 13048 20646 13100
rect 25185 13091 25243 13097
rect 25185 13057 25197 13091
rect 25231 13088 25243 13091
rect 25274 13088 25280 13100
rect 25231 13060 25280 13088
rect 25231 13057 25243 13060
rect 25185 13051 25243 13057
rect 25274 13048 25280 13060
rect 25332 13048 25338 13100
rect 28126 13088 28132 13100
rect 28087 13060 28132 13088
rect 28126 13048 28132 13060
rect 28184 13048 28190 13100
rect 19018 12980 19024 13032
rect 19076 13020 19082 13032
rect 21045 13023 21103 13029
rect 19076 12992 19524 13020
rect 19076 12980 19082 12992
rect 18929 12955 18987 12961
rect 18929 12921 18941 12955
rect 18975 12921 18987 12955
rect 19294 12952 19300 12964
rect 18929 12915 18987 12921
rect 19036 12924 19300 12952
rect 14384 12856 14924 12884
rect 14384 12844 14390 12856
rect 14970 12844 14976 12896
rect 15028 12884 15034 12896
rect 19036 12893 19064 12924
rect 19294 12912 19300 12924
rect 19352 12912 19358 12964
rect 19496 12961 19524 12992
rect 21045 12989 21057 13023
rect 21091 13020 21103 13023
rect 21226 13020 21232 13032
rect 21091 12992 21232 13020
rect 21091 12989 21103 12992
rect 21045 12983 21103 12989
rect 21226 12980 21232 12992
rect 21284 12980 21290 13032
rect 19481 12955 19539 12961
rect 19481 12921 19493 12955
rect 19527 12921 19539 12955
rect 19481 12915 19539 12921
rect 20030 12912 20036 12964
rect 20088 12952 20094 12964
rect 20674 12952 20680 12964
rect 20088 12924 20680 12952
rect 20088 12912 20094 12924
rect 20674 12912 20680 12924
rect 20732 12952 20738 12964
rect 20732 12924 22376 12952
rect 20732 12912 20738 12924
rect 15249 12887 15307 12893
rect 15249 12884 15261 12887
rect 15028 12856 15261 12884
rect 15028 12844 15034 12856
rect 15249 12853 15261 12856
rect 15295 12853 15307 12887
rect 15249 12847 15307 12853
rect 19021 12887 19079 12893
rect 19021 12853 19033 12887
rect 19067 12853 19079 12887
rect 19386 12884 19392 12896
rect 19347 12856 19392 12884
rect 19021 12847 19079 12853
rect 19386 12844 19392 12856
rect 19444 12844 19450 12896
rect 21226 12884 21232 12896
rect 21187 12856 21232 12884
rect 21226 12844 21232 12856
rect 21284 12844 21290 12896
rect 21612 12893 21640 12924
rect 21597 12887 21655 12893
rect 21597 12853 21609 12887
rect 21643 12853 21655 12887
rect 21597 12847 21655 12853
rect 21689 12887 21747 12893
rect 21689 12853 21701 12887
rect 21735 12884 21747 12887
rect 22146 12884 22152 12896
rect 21735 12856 22152 12884
rect 21735 12853 21747 12856
rect 21689 12847 21747 12853
rect 22146 12844 22152 12856
rect 22204 12844 22210 12896
rect 22348 12893 22376 12924
rect 25182 12912 25188 12964
rect 25240 12952 25246 12964
rect 27390 12952 27396 12964
rect 25240 12924 27396 12952
rect 25240 12912 25246 12924
rect 27390 12912 27396 12924
rect 27448 12912 27454 12964
rect 28770 12952 28776 12964
rect 28731 12924 28776 12952
rect 28770 12912 28776 12924
rect 28828 12912 28834 12964
rect 22333 12887 22391 12893
rect 22333 12853 22345 12887
rect 22379 12853 22391 12887
rect 22333 12847 22391 12853
rect 23897 12887 23955 12893
rect 23897 12853 23909 12887
rect 23943 12884 23955 12887
rect 24722 12884 24728 12896
rect 23943 12856 24728 12884
rect 23943 12853 23955 12856
rect 23897 12847 23955 12853
rect 24722 12844 24728 12856
rect 24780 12844 24786 12896
rect 24906 12884 24912 12896
rect 24867 12856 24912 12884
rect 24906 12844 24912 12856
rect 24964 12844 24970 12896
rect 25090 12844 25096 12896
rect 25148 12884 25154 12896
rect 25918 12884 25924 12896
rect 25148 12856 25241 12884
rect 25879 12856 25924 12884
rect 25148 12844 25154 12856
rect 25918 12844 25924 12856
rect 25976 12844 25982 12896
rect 26010 12844 26016 12896
rect 26068 12884 26074 12896
rect 27945 12887 28003 12893
rect 26068 12856 26113 12884
rect 26068 12844 26074 12856
rect 27945 12853 27957 12887
rect 27991 12853 28003 12887
rect 27945 12847 28003 12853
rect 28681 12887 28739 12893
rect 28681 12853 28693 12887
rect 28727 12884 28739 12887
rect 29598 12884 29604 12896
rect 28727 12856 29604 12884
rect 28727 12853 28739 12856
rect 28681 12847 28739 12853
rect 18377 12819 18435 12825
rect 18377 12785 18389 12819
rect 18423 12816 18435 12819
rect 19570 12816 19576 12828
rect 18423 12788 19576 12816
rect 18423 12785 18435 12788
rect 18377 12779 18435 12785
rect 19570 12776 19576 12788
rect 19628 12776 19634 12828
rect 25108 12816 25136 12844
rect 27758 12816 27764 12828
rect 25108 12788 27764 12816
rect 27758 12776 27764 12788
rect 27816 12776 27822 12828
rect 27960 12816 27988 12847
rect 29598 12844 29604 12856
rect 29656 12844 29662 12896
rect 28954 12816 28960 12828
rect 27960 12788 28960 12816
rect 14142 12748 14148 12760
rect 13372 12720 14148 12748
rect 13372 12708 13378 12720
rect 14142 12708 14148 12720
rect 14200 12708 14206 12760
rect 14786 12708 14792 12760
rect 14844 12748 14850 12760
rect 15341 12751 15399 12757
rect 15341 12748 15353 12751
rect 14844 12720 15353 12748
rect 14844 12708 14850 12720
rect 15341 12717 15353 12720
rect 15387 12717 15399 12751
rect 15341 12711 15399 12717
rect 15982 12708 15988 12760
rect 16040 12748 16046 12760
rect 19938 12748 19944 12760
rect 16040 12720 19944 12748
rect 16040 12708 16046 12720
rect 19938 12708 19944 12720
rect 19996 12708 20002 12760
rect 21686 12708 21692 12760
rect 21744 12748 21750 12760
rect 22425 12751 22483 12757
rect 22425 12748 22437 12751
rect 21744 12720 22437 12748
rect 21744 12708 21750 12720
rect 22425 12717 22437 12720
rect 22471 12717 22483 12751
rect 23894 12748 23900 12760
rect 23855 12720 23900 12748
rect 22425 12711 22483 12717
rect 23894 12708 23900 12720
rect 23952 12708 23958 12760
rect 25366 12708 25372 12760
rect 25424 12748 25430 12760
rect 26378 12748 26384 12760
rect 25424 12720 26384 12748
rect 25424 12708 25430 12720
rect 26378 12708 26384 12720
rect 26436 12748 26442 12760
rect 27960 12748 27988 12788
rect 28954 12776 28960 12788
rect 29012 12776 29018 12828
rect 26436 12720 27988 12748
rect 26436 12708 26442 12720
rect 11000 12658 30136 12680
rect 11000 12606 19142 12658
rect 19194 12606 19206 12658
rect 19258 12606 19270 12658
rect 19322 12606 19334 12658
rect 19386 12606 29142 12658
rect 29194 12606 29206 12658
rect 29258 12606 29270 12658
rect 29322 12606 29334 12658
rect 29386 12606 30136 12658
rect 11000 12584 30136 12606
rect 12302 12504 12308 12556
rect 12360 12544 12366 12556
rect 12360 12516 13544 12544
rect 12360 12504 12366 12516
rect 13130 12476 13136 12488
rect 13091 12448 13136 12476
rect 13130 12436 13136 12448
rect 13188 12436 13194 12488
rect 12026 12408 12032 12420
rect 11987 12380 12032 12408
rect 12026 12368 12032 12380
rect 12084 12368 12090 12420
rect 12578 12408 12584 12420
rect 12539 12380 12584 12408
rect 12578 12368 12584 12380
rect 12636 12368 12642 12420
rect 12762 12368 12768 12420
rect 12820 12408 12826 12420
rect 12857 12411 12915 12417
rect 12857 12408 12869 12411
rect 12820 12380 12869 12408
rect 12820 12368 12826 12380
rect 12857 12377 12869 12380
rect 12903 12377 12915 12411
rect 12857 12371 12915 12377
rect 13516 12340 13544 12516
rect 14142 12504 14148 12556
rect 14200 12544 14206 12556
rect 14200 12516 18880 12544
rect 14200 12504 14206 12516
rect 16902 12476 16908 12488
rect 13976 12448 14924 12476
rect 13682 12368 13688 12420
rect 13740 12408 13746 12420
rect 13976 12417 14004 12448
rect 13961 12411 14019 12417
rect 13961 12408 13973 12411
rect 13740 12380 13973 12408
rect 13740 12368 13746 12380
rect 13961 12377 13973 12380
rect 14007 12377 14019 12411
rect 13961 12371 14019 12377
rect 14145 12411 14203 12417
rect 14145 12377 14157 12411
rect 14191 12408 14203 12411
rect 14697 12411 14755 12417
rect 14697 12408 14709 12411
rect 14191 12380 14709 12408
rect 14191 12377 14203 12380
rect 14145 12371 14203 12377
rect 14697 12377 14709 12380
rect 14743 12408 14755 12411
rect 14786 12408 14792 12420
rect 14743 12380 14792 12408
rect 14743 12377 14755 12380
rect 14697 12371 14755 12377
rect 14786 12368 14792 12380
rect 14844 12368 14850 12420
rect 14896 12417 14924 12448
rect 16644 12448 16908 12476
rect 14881 12411 14939 12417
rect 14881 12377 14893 12411
rect 14927 12408 14939 12411
rect 15798 12408 15804 12420
rect 14927 12380 15804 12408
rect 14927 12377 14939 12380
rect 14881 12371 14939 12377
rect 15798 12368 15804 12380
rect 15856 12368 15862 12420
rect 15893 12411 15951 12417
rect 15893 12377 15905 12411
rect 15939 12408 15951 12411
rect 16534 12408 16540 12420
rect 15939 12380 16540 12408
rect 15939 12377 15951 12380
rect 15893 12371 15951 12377
rect 16534 12368 16540 12380
rect 16592 12368 16598 12420
rect 16644 12417 16672 12448
rect 16902 12436 16908 12448
rect 16960 12436 16966 12488
rect 17546 12436 17552 12488
rect 17604 12436 17610 12488
rect 18190 12436 18196 12488
rect 18248 12476 18254 12488
rect 18653 12479 18711 12485
rect 18653 12476 18665 12479
rect 18248 12448 18665 12476
rect 18248 12436 18254 12448
rect 18653 12445 18665 12448
rect 18699 12476 18711 12479
rect 18742 12476 18748 12488
rect 18699 12448 18748 12476
rect 18699 12445 18711 12448
rect 18653 12439 18711 12445
rect 18742 12436 18748 12448
rect 18800 12436 18806 12488
rect 18852 12476 18880 12516
rect 19846 12504 19852 12556
rect 19904 12544 19910 12556
rect 23526 12544 23532 12556
rect 19904 12516 23532 12544
rect 19904 12504 19910 12516
rect 23526 12504 23532 12516
rect 23584 12504 23590 12556
rect 26562 12544 26568 12556
rect 25476 12516 26568 12544
rect 20493 12479 20551 12485
rect 20493 12476 20505 12479
rect 18852 12448 20505 12476
rect 20493 12445 20505 12448
rect 20539 12445 20551 12479
rect 25366 12476 25372 12488
rect 23742 12448 25372 12476
rect 20493 12439 20551 12445
rect 25366 12436 25372 12448
rect 25424 12436 25430 12488
rect 25476 12420 25504 12516
rect 26562 12504 26568 12516
rect 26620 12504 26626 12556
rect 27850 12504 27856 12556
rect 27908 12544 27914 12556
rect 29141 12547 29199 12553
rect 29141 12544 29153 12547
rect 27908 12516 29153 12544
rect 27908 12504 27914 12516
rect 29141 12513 29153 12516
rect 29187 12513 29199 12547
rect 29141 12507 29199 12513
rect 26470 12436 26476 12488
rect 26528 12436 26534 12488
rect 27482 12476 27488 12488
rect 27443 12448 27488 12476
rect 27482 12436 27488 12448
rect 27540 12436 27546 12488
rect 28034 12476 28040 12488
rect 27947 12448 28040 12476
rect 16629 12411 16687 12417
rect 16629 12377 16641 12411
rect 16675 12377 16687 12411
rect 19570 12408 19576 12420
rect 19531 12380 19576 12408
rect 16629 12371 16687 12377
rect 14326 12340 14332 12352
rect 13516 12312 14332 12340
rect 14326 12300 14332 12312
rect 14384 12300 14390 12352
rect 13406 12232 13412 12284
rect 13464 12272 13470 12284
rect 15065 12275 15123 12281
rect 15065 12272 15077 12275
rect 13464 12244 15077 12272
rect 13464 12232 13470 12244
rect 15065 12241 15077 12244
rect 15111 12241 15123 12275
rect 16644 12272 16672 12371
rect 19570 12368 19576 12380
rect 19628 12368 19634 12420
rect 21134 12408 21140 12420
rect 21095 12380 21140 12408
rect 21134 12368 21140 12380
rect 21192 12368 21198 12420
rect 21502 12408 21508 12420
rect 21463 12380 21508 12408
rect 21502 12368 21508 12380
rect 21560 12368 21566 12420
rect 21686 12408 21692 12420
rect 21647 12380 21692 12408
rect 21686 12368 21692 12380
rect 21744 12368 21750 12420
rect 25458 12408 25464 12420
rect 25371 12380 25464 12408
rect 25458 12368 25464 12380
rect 25516 12368 25522 12420
rect 27960 12417 27988 12448
rect 28034 12436 28040 12448
rect 28092 12476 28098 12488
rect 28092 12448 28908 12476
rect 28092 12436 28098 12448
rect 27945 12411 28003 12417
rect 27945 12377 27957 12411
rect 27991 12377 28003 12411
rect 27945 12371 28003 12377
rect 28129 12411 28187 12417
rect 28129 12377 28141 12411
rect 28175 12408 28187 12411
rect 28586 12408 28592 12420
rect 28175 12380 28592 12408
rect 28175 12377 28187 12380
rect 28129 12371 28187 12377
rect 28586 12368 28592 12380
rect 28644 12408 28650 12420
rect 28880 12417 28908 12448
rect 28681 12411 28739 12417
rect 28681 12408 28693 12411
rect 28644 12380 28693 12408
rect 28644 12368 28650 12380
rect 28681 12377 28693 12380
rect 28727 12377 28739 12411
rect 28681 12371 28739 12377
rect 28865 12411 28923 12417
rect 28865 12377 28877 12411
rect 28911 12377 28923 12411
rect 28865 12371 28923 12377
rect 16902 12340 16908 12352
rect 16863 12312 16908 12340
rect 16902 12300 16908 12312
rect 16960 12300 16966 12352
rect 21226 12340 21232 12352
rect 21187 12312 21232 12340
rect 21226 12300 21232 12312
rect 21284 12300 21290 12352
rect 22238 12340 22244 12352
rect 22199 12312 22244 12340
rect 22238 12300 22244 12312
rect 22296 12300 22302 12352
rect 22514 12340 22520 12352
rect 22475 12312 22520 12340
rect 22514 12300 22520 12312
rect 22572 12300 22578 12352
rect 24265 12343 24323 12349
rect 24265 12309 24277 12343
rect 24311 12309 24323 12343
rect 25734 12340 25740 12352
rect 25695 12312 25740 12340
rect 24265 12303 24323 12309
rect 15065 12235 15123 12241
rect 15172 12244 16672 12272
rect 13958 12164 13964 12216
rect 14016 12204 14022 12216
rect 15172 12204 15200 12244
rect 16074 12204 16080 12216
rect 14016 12176 15200 12204
rect 16035 12176 16080 12204
rect 14016 12164 14022 12176
rect 16074 12164 16080 12176
rect 16132 12164 16138 12216
rect 18926 12164 18932 12216
rect 18984 12204 18990 12216
rect 19665 12207 19723 12213
rect 19665 12204 19677 12207
rect 18984 12176 19677 12204
rect 18984 12164 18990 12176
rect 19665 12173 19677 12176
rect 19711 12173 19723 12207
rect 19665 12167 19723 12173
rect 22146 12164 22152 12216
rect 22204 12204 22210 12216
rect 24280 12204 24308 12303
rect 25734 12300 25740 12312
rect 25792 12300 25798 12352
rect 22204 12176 24308 12204
rect 22204 12164 22210 12176
rect 11000 12114 30136 12136
rect 11000 12062 14142 12114
rect 14194 12062 14206 12114
rect 14258 12062 14270 12114
rect 14322 12062 14334 12114
rect 14386 12062 24142 12114
rect 24194 12062 24206 12114
rect 24258 12062 24270 12114
rect 24322 12062 24334 12114
rect 24386 12062 30136 12114
rect 11000 12040 30136 12062
rect 11566 11960 11572 12012
rect 11624 12000 11630 12012
rect 11753 12003 11811 12009
rect 11753 12000 11765 12003
rect 11624 11972 11765 12000
rect 11624 11960 11630 11972
rect 11753 11969 11765 11972
rect 11799 11969 11811 12003
rect 12762 12000 12768 12012
rect 12723 11972 12768 12000
rect 11753 11963 11811 11969
rect 12762 11960 12768 11972
rect 12820 11960 12826 12012
rect 14510 11960 14516 12012
rect 14568 12000 14574 12012
rect 20950 12000 20956 12012
rect 14568 11972 20956 12000
rect 14568 11960 14574 11972
rect 20950 11960 20956 11972
rect 21008 11960 21014 12012
rect 21226 11960 21232 12012
rect 21284 12000 21290 12012
rect 21505 12003 21563 12009
rect 21505 12000 21517 12003
rect 21284 11972 21517 12000
rect 21284 11960 21290 11972
rect 21505 11969 21517 11972
rect 21551 11969 21563 12003
rect 21505 11963 21563 11969
rect 26470 11960 26476 12012
rect 26528 12000 26534 12012
rect 26565 12003 26623 12009
rect 26565 12000 26577 12003
rect 26528 11972 26577 12000
rect 26528 11960 26534 11972
rect 26565 11969 26577 11972
rect 26611 11969 26623 12003
rect 28034 12000 28040 12012
rect 27995 11972 28040 12000
rect 26565 11963 26623 11969
rect 28034 11960 28040 11972
rect 28092 11960 28098 12012
rect 16994 11892 17000 11944
rect 17052 11932 17058 11944
rect 21686 11932 21692 11944
rect 17052 11904 18696 11932
rect 17052 11892 17058 11904
rect 13225 11867 13283 11873
rect 13225 11833 13237 11867
rect 13271 11864 13283 11867
rect 13406 11864 13412 11876
rect 13271 11836 13412 11864
rect 13271 11833 13283 11836
rect 13225 11827 13283 11833
rect 13406 11824 13412 11836
rect 13464 11824 13470 11876
rect 14786 11864 14792 11876
rect 13516 11836 14792 11864
rect 10462 11756 10468 11808
rect 10520 11796 10526 11808
rect 11661 11799 11719 11805
rect 11661 11796 11673 11799
rect 10520 11768 11673 11796
rect 10520 11756 10526 11768
rect 11661 11765 11673 11768
rect 11707 11765 11719 11799
rect 11661 11759 11719 11765
rect 13133 11799 13191 11805
rect 13133 11765 13145 11799
rect 13179 11796 13191 11799
rect 13314 11796 13320 11808
rect 13179 11768 13320 11796
rect 13179 11765 13191 11768
rect 13133 11759 13191 11765
rect 13314 11756 13320 11768
rect 13372 11756 13378 11808
rect 13516 11805 13544 11836
rect 14786 11824 14792 11836
rect 14844 11824 14850 11876
rect 14970 11824 14976 11876
rect 15028 11864 15034 11876
rect 16169 11867 16227 11873
rect 16169 11864 16181 11867
rect 15028 11836 16181 11864
rect 15028 11824 15034 11836
rect 16169 11833 16181 11836
rect 16215 11833 16227 11867
rect 16169 11827 16227 11833
rect 16902 11824 16908 11876
rect 16960 11864 16966 11876
rect 18668 11873 18696 11904
rect 21244 11904 21692 11932
rect 17181 11867 17239 11873
rect 17181 11864 17193 11867
rect 16960 11836 17193 11864
rect 16960 11824 16966 11836
rect 17181 11833 17193 11836
rect 17227 11833 17239 11867
rect 17181 11827 17239 11833
rect 18653 11867 18711 11873
rect 18653 11833 18665 11867
rect 18699 11833 18711 11867
rect 18926 11864 18932 11876
rect 18887 11836 18932 11864
rect 18653 11827 18711 11833
rect 18926 11824 18932 11836
rect 18984 11824 18990 11876
rect 20674 11864 20680 11876
rect 20635 11836 20680 11864
rect 20674 11824 20680 11836
rect 20732 11824 20738 11876
rect 21244 11873 21272 11904
rect 21686 11892 21692 11904
rect 21744 11892 21750 11944
rect 22238 11892 22244 11944
rect 22296 11932 22302 11944
rect 22296 11904 23940 11932
rect 22296 11892 22302 11904
rect 21229 11867 21287 11873
rect 21229 11833 21241 11867
rect 21275 11833 21287 11867
rect 21502 11864 21508 11876
rect 21229 11827 21287 11833
rect 21336 11836 21508 11864
rect 13501 11799 13559 11805
rect 13501 11765 13513 11799
rect 13547 11765 13559 11799
rect 13682 11796 13688 11808
rect 13643 11768 13688 11796
rect 13501 11759 13559 11765
rect 13682 11756 13688 11768
rect 13740 11756 13746 11808
rect 14050 11756 14056 11808
rect 14108 11796 14114 11808
rect 14145 11799 14203 11805
rect 14145 11796 14157 11799
rect 14108 11768 14157 11796
rect 14108 11756 14114 11768
rect 14145 11765 14157 11768
rect 14191 11765 14203 11799
rect 16074 11796 16080 11808
rect 15554 11768 16080 11796
rect 14145 11759 14203 11765
rect 16074 11756 16080 11768
rect 16132 11756 16138 11808
rect 17270 11756 17276 11808
rect 17328 11796 17334 11808
rect 17638 11796 17644 11808
rect 17328 11768 17644 11796
rect 17328 11756 17334 11768
rect 17638 11756 17644 11768
rect 17696 11796 17702 11808
rect 17733 11799 17791 11805
rect 17733 11796 17745 11799
rect 17696 11768 17745 11796
rect 17696 11756 17702 11768
rect 17733 11765 17745 11768
rect 17779 11765 17791 11799
rect 17733 11759 17791 11765
rect 18009 11799 18067 11805
rect 18009 11765 18021 11799
rect 18055 11765 18067 11799
rect 18190 11796 18196 11808
rect 18151 11768 18196 11796
rect 18009 11759 18067 11765
rect 14421 11731 14479 11737
rect 14421 11697 14433 11731
rect 14467 11697 14479 11731
rect 18024 11728 18052 11759
rect 18190 11756 18196 11768
rect 18248 11756 18254 11808
rect 21336 11805 21364 11836
rect 21502 11824 21508 11836
rect 21560 11864 21566 11876
rect 23912 11873 23940 11904
rect 22425 11867 22483 11873
rect 22425 11864 22437 11867
rect 21560 11836 22437 11864
rect 21560 11824 21566 11836
rect 22425 11833 22437 11836
rect 22471 11833 22483 11867
rect 22425 11827 22483 11833
rect 23897 11867 23955 11873
rect 23897 11833 23909 11867
rect 23943 11864 23955 11867
rect 25458 11864 25464 11876
rect 23943 11836 25464 11864
rect 23943 11833 23955 11836
rect 23897 11827 23955 11833
rect 25458 11824 25464 11836
rect 25516 11824 25522 11876
rect 25734 11824 25740 11876
rect 25792 11864 25798 11876
rect 25921 11867 25979 11873
rect 25921 11864 25933 11867
rect 25792 11836 25933 11864
rect 25792 11824 25798 11836
rect 25921 11833 25933 11836
rect 25967 11833 25979 11867
rect 25921 11827 25979 11833
rect 21321 11799 21379 11805
rect 21321 11765 21333 11799
rect 21367 11765 21379 11799
rect 22146 11796 22152 11808
rect 21321 11759 21379 11765
rect 21704 11768 22152 11796
rect 19018 11728 19024 11740
rect 18024 11700 19024 11728
rect 14421 11691 14479 11697
rect 14436 11660 14464 11691
rect 19018 11688 19024 11700
rect 19076 11688 19082 11740
rect 19938 11688 19944 11740
rect 19996 11688 20002 11740
rect 20950 11688 20956 11740
rect 21008 11728 21014 11740
rect 21704 11728 21732 11768
rect 22146 11756 22152 11768
rect 22204 11796 22210 11808
rect 22333 11799 22391 11805
rect 22333 11796 22345 11799
rect 22204 11768 22345 11796
rect 22204 11756 22210 11768
rect 22333 11765 22345 11768
rect 22379 11765 22391 11799
rect 26378 11796 26384 11808
rect 26339 11768 26384 11796
rect 22333 11759 22391 11765
rect 26378 11756 26384 11768
rect 26436 11756 26442 11808
rect 27482 11756 27488 11808
rect 27540 11796 27546 11808
rect 27945 11799 28003 11805
rect 27945 11796 27957 11799
rect 27540 11768 27957 11796
rect 27540 11756 27546 11768
rect 27945 11765 27957 11768
rect 27991 11765 28003 11799
rect 27945 11759 28003 11765
rect 24173 11731 24231 11737
rect 24173 11728 24185 11731
rect 21008 11700 21732 11728
rect 23268 11700 24185 11728
rect 21008 11688 21014 11700
rect 16074 11660 16080 11672
rect 14436 11632 16080 11660
rect 16074 11620 16080 11632
rect 16132 11620 16138 11672
rect 18006 11620 18012 11672
rect 18064 11660 18070 11672
rect 23268 11660 23296 11700
rect 24173 11697 24185 11700
rect 24219 11697 24231 11731
rect 25550 11728 25556 11740
rect 25398 11700 25556 11728
rect 24173 11691 24231 11697
rect 25550 11688 25556 11700
rect 25608 11688 25614 11740
rect 18064 11632 23296 11660
rect 18064 11620 18070 11632
rect 23710 11620 23716 11672
rect 23768 11660 23774 11672
rect 24446 11660 24452 11672
rect 23768 11632 24452 11660
rect 23768 11620 23774 11632
rect 24446 11620 24452 11632
rect 24504 11620 24510 11672
rect 11000 11570 30136 11592
rect 11000 11518 19142 11570
rect 19194 11518 19206 11570
rect 19258 11518 19270 11570
rect 19322 11518 19334 11570
rect 19386 11518 29142 11570
rect 29194 11518 29206 11570
rect 29258 11518 29270 11570
rect 29322 11518 29334 11570
rect 29386 11518 30136 11570
rect 11000 11496 30136 11518
rect 16074 11456 16080 11468
rect 16035 11428 16080 11456
rect 16074 11416 16080 11428
rect 16132 11416 16138 11468
rect 17546 11456 17552 11468
rect 17507 11428 17552 11456
rect 17546 11416 17552 11428
rect 17604 11416 17610 11468
rect 18469 11459 18527 11465
rect 18469 11425 18481 11459
rect 18515 11456 18527 11459
rect 18745 11459 18803 11465
rect 18745 11456 18757 11459
rect 18515 11428 18757 11456
rect 18515 11425 18527 11428
rect 18469 11419 18527 11425
rect 18745 11425 18757 11428
rect 18791 11456 18803 11459
rect 19478 11456 19484 11468
rect 18791 11428 19484 11456
rect 18791 11425 18803 11428
rect 18745 11419 18803 11425
rect 19478 11416 19484 11428
rect 19536 11416 19542 11468
rect 19849 11459 19907 11465
rect 19849 11425 19861 11459
rect 19895 11456 19907 11459
rect 19938 11456 19944 11468
rect 19895 11428 19944 11456
rect 19895 11425 19907 11428
rect 19849 11419 19907 11425
rect 19938 11416 19944 11428
rect 19996 11416 20002 11468
rect 25550 11456 25556 11468
rect 25511 11428 25556 11456
rect 25550 11416 25556 11428
rect 25608 11416 25614 11468
rect 15632 11360 16028 11388
rect 15632 11329 15660 11360
rect 15065 11323 15123 11329
rect 15065 11289 15077 11323
rect 15111 11320 15123 11323
rect 15617 11323 15675 11329
rect 15617 11320 15629 11323
rect 15111 11292 15629 11320
rect 15111 11289 15123 11292
rect 15065 11283 15123 11289
rect 15617 11289 15629 11292
rect 15663 11289 15675 11323
rect 15798 11320 15804 11332
rect 15759 11292 15804 11320
rect 15617 11283 15675 11289
rect 15798 11280 15804 11292
rect 15856 11280 15862 11332
rect 14970 11252 14976 11264
rect 14931 11224 14976 11252
rect 14970 11212 14976 11224
rect 15028 11212 15034 11264
rect 16000 11252 16028 11360
rect 17270 11348 17276 11400
rect 17328 11388 17334 11400
rect 20398 11388 20404 11400
rect 17328 11360 20404 11388
rect 17328 11348 17334 11360
rect 20398 11348 20404 11360
rect 20456 11388 20462 11400
rect 21873 11391 21931 11397
rect 20456 11360 21364 11388
rect 20456 11348 20462 11360
rect 17178 11280 17184 11332
rect 17236 11320 17242 11332
rect 17365 11323 17423 11329
rect 17365 11320 17377 11323
rect 17236 11292 17377 11320
rect 17236 11280 17242 11292
rect 17365 11289 17377 11292
rect 17411 11289 17423 11323
rect 17365 11283 17423 11289
rect 17270 11252 17276 11264
rect 16000 11224 17276 11252
rect 17270 11212 17276 11224
rect 17328 11212 17334 11264
rect 17380 11252 17408 11283
rect 18190 11280 18196 11332
rect 18248 11320 18254 11332
rect 20784 11329 20812 11360
rect 18653 11323 18711 11329
rect 18653 11320 18665 11323
rect 18248 11292 18665 11320
rect 18248 11280 18254 11292
rect 18653 11289 18665 11292
rect 18699 11289 18711 11323
rect 18653 11283 18711 11289
rect 19665 11323 19723 11329
rect 19665 11289 19677 11323
rect 19711 11289 19723 11323
rect 19665 11283 19723 11289
rect 20769 11323 20827 11329
rect 20769 11289 20781 11323
rect 20815 11289 20827 11323
rect 20769 11283 20827 11289
rect 20861 11323 20919 11329
rect 20861 11289 20873 11323
rect 20907 11320 20919 11323
rect 20950 11320 20956 11332
rect 20907 11292 20956 11320
rect 20907 11289 20919 11292
rect 20861 11283 20919 11289
rect 19680 11252 19708 11283
rect 20950 11280 20956 11292
rect 21008 11280 21014 11332
rect 21336 11329 21364 11360
rect 21873 11357 21885 11391
rect 21919 11388 21931 11391
rect 22514 11388 22520 11400
rect 21919 11360 22520 11388
rect 21919 11357 21931 11360
rect 21873 11351 21931 11357
rect 22514 11348 22520 11360
rect 22572 11348 22578 11400
rect 21321 11323 21379 11329
rect 21321 11289 21333 11323
rect 21367 11289 21379 11323
rect 21321 11283 21379 11289
rect 21505 11323 21563 11329
rect 21505 11289 21517 11323
rect 21551 11320 21563 11323
rect 21686 11320 21692 11332
rect 21551 11292 21692 11320
rect 21551 11289 21563 11292
rect 21505 11283 21563 11289
rect 21686 11280 21692 11292
rect 21744 11280 21750 11332
rect 23894 11320 23900 11332
rect 23855 11292 23900 11320
rect 23894 11280 23900 11292
rect 23952 11280 23958 11332
rect 25366 11320 25372 11332
rect 25327 11292 25372 11320
rect 25366 11280 25372 11292
rect 25424 11280 25430 11332
rect 17380 11224 19708 11252
rect 15798 11144 15804 11196
rect 15856 11184 15862 11196
rect 18469 11187 18527 11193
rect 18469 11184 18481 11187
rect 15856 11156 18481 11184
rect 15856 11144 15862 11156
rect 18469 11153 18481 11156
rect 18515 11153 18527 11187
rect 18469 11147 18527 11153
rect 21686 11144 21692 11196
rect 21744 11184 21750 11196
rect 23069 11187 23127 11193
rect 23069 11184 23081 11187
rect 21744 11156 23081 11184
rect 21744 11144 21750 11156
rect 23069 11153 23081 11156
rect 23115 11153 23127 11187
rect 23069 11147 23127 11153
rect 11000 11026 30136 11048
rect 11000 10974 14142 11026
rect 14194 10974 14206 11026
rect 14258 10974 14270 11026
rect 14322 10974 14334 11026
rect 14386 10974 24142 11026
rect 24194 10974 24206 11026
rect 24258 10974 24270 11026
rect 24322 10974 24334 11026
rect 24386 10974 30136 11026
rect 11000 10952 30136 10974
<< via1 >>
rect 19142 30014 19194 30066
rect 19206 30014 19258 30066
rect 19270 30014 19322 30066
rect 19334 30014 19386 30066
rect 29142 30014 29194 30066
rect 29206 30014 29258 30066
rect 29270 30014 29322 30066
rect 29334 30014 29386 30066
rect 14976 29819 15028 29828
rect 14976 29785 14985 29819
rect 14985 29785 15019 29819
rect 15019 29785 15028 29819
rect 14976 29776 15028 29785
rect 15068 29776 15120 29828
rect 19760 29776 19812 29828
rect 19852 29819 19904 29828
rect 19852 29785 19861 29819
rect 19861 29785 19895 29819
rect 19895 29785 19904 29819
rect 19852 29776 19904 29785
rect 23348 29776 23400 29828
rect 26384 29819 26436 29828
rect 26384 29785 26393 29819
rect 26393 29785 26427 29819
rect 26427 29785 26436 29819
rect 26384 29776 26436 29785
rect 28684 29776 28736 29828
rect 21140 29751 21192 29760
rect 21140 29717 21149 29751
rect 21149 29717 21183 29751
rect 21183 29717 21192 29751
rect 21140 29708 21192 29717
rect 21968 29640 22020 29692
rect 14700 29572 14752 29624
rect 15988 29572 16040 29624
rect 19024 29615 19076 29624
rect 19024 29581 19033 29615
rect 19033 29581 19067 29615
rect 19067 29581 19076 29615
rect 19024 29572 19076 29581
rect 19668 29615 19720 29624
rect 19668 29581 19677 29615
rect 19677 29581 19711 29615
rect 19711 29581 19720 29615
rect 19668 29572 19720 29581
rect 27488 29572 27540 29624
rect 28868 29572 28920 29624
rect 14142 29470 14194 29522
rect 14206 29470 14258 29522
rect 14270 29470 14322 29522
rect 14334 29470 14386 29522
rect 24142 29470 24194 29522
rect 24206 29470 24258 29522
rect 24270 29470 24322 29522
rect 24334 29470 24386 29522
rect 21324 29368 21376 29420
rect 18380 29300 18432 29352
rect 19760 29300 19812 29352
rect 13504 29232 13556 29284
rect 15160 29207 15212 29216
rect 15160 29173 15169 29207
rect 15169 29173 15203 29207
rect 15203 29173 15212 29207
rect 15160 29164 15212 29173
rect 16356 29232 16408 29284
rect 19668 29232 19720 29284
rect 21140 29232 21192 29284
rect 22060 29232 22112 29284
rect 14056 29096 14108 29148
rect 15436 29096 15488 29148
rect 17644 29164 17696 29216
rect 18564 29096 18616 29148
rect 20036 29164 20088 29216
rect 20680 29207 20732 29216
rect 20680 29173 20689 29207
rect 20689 29173 20723 29207
rect 20723 29173 20732 29207
rect 20680 29164 20732 29173
rect 19852 29096 19904 29148
rect 23532 29232 23584 29284
rect 22704 29207 22756 29216
rect 22704 29173 22713 29207
rect 22713 29173 22747 29207
rect 22747 29173 22756 29207
rect 22704 29164 22756 29173
rect 23348 29207 23400 29216
rect 23348 29173 23357 29207
rect 23357 29173 23391 29207
rect 23391 29173 23400 29207
rect 23348 29164 23400 29173
rect 22152 29096 22204 29148
rect 24452 29164 24504 29216
rect 25464 29207 25516 29216
rect 25464 29173 25473 29207
rect 25473 29173 25507 29207
rect 25507 29173 25516 29207
rect 25464 29164 25516 29173
rect 27396 29164 27448 29216
rect 29512 29164 29564 29216
rect 26384 29139 26436 29148
rect 26384 29105 26393 29139
rect 26393 29105 26427 29139
rect 26427 29105 26436 29139
rect 26384 29096 26436 29105
rect 23716 29028 23768 29080
rect 26292 29028 26344 29080
rect 27120 29071 27172 29080
rect 27120 29037 27129 29071
rect 27129 29037 27163 29071
rect 27163 29037 27172 29071
rect 27120 29028 27172 29037
rect 27212 29071 27264 29080
rect 27212 29037 27221 29071
rect 27221 29037 27255 29071
rect 27255 29037 27264 29071
rect 27212 29028 27264 29037
rect 28776 29028 28828 29080
rect 19142 28926 19194 28978
rect 19206 28926 19258 28978
rect 19270 28926 19322 28978
rect 19334 28926 19386 28978
rect 29142 28926 29194 28978
rect 29206 28926 29258 28978
rect 29270 28926 29322 28978
rect 29334 28926 29386 28978
rect 14516 28824 14568 28876
rect 15068 28756 15120 28808
rect 10652 28688 10704 28740
rect 14056 28731 14108 28740
rect 14056 28697 14065 28731
rect 14065 28697 14099 28731
rect 14099 28697 14108 28731
rect 14056 28688 14108 28697
rect 14976 28731 15028 28740
rect 14976 28697 14985 28731
rect 14985 28697 15019 28731
rect 15019 28697 15028 28731
rect 14976 28688 15028 28697
rect 15436 28731 15488 28740
rect 15436 28697 15445 28731
rect 15445 28697 15479 28731
rect 15479 28697 15488 28731
rect 15436 28688 15488 28697
rect 16724 28731 16776 28740
rect 16724 28697 16733 28731
rect 16733 28697 16767 28731
rect 16767 28697 16776 28731
rect 16724 28688 16776 28697
rect 17644 28620 17696 28672
rect 19024 28756 19076 28808
rect 20680 28824 20732 28876
rect 24452 28867 24504 28876
rect 24452 28833 24461 28867
rect 24461 28833 24495 28867
rect 24495 28833 24504 28867
rect 24452 28824 24504 28833
rect 27764 28824 27816 28876
rect 22704 28756 22756 28808
rect 25464 28756 25516 28808
rect 27488 28799 27540 28808
rect 18196 28688 18248 28740
rect 20312 28688 20364 28740
rect 21140 28688 21192 28740
rect 22152 28731 22204 28740
rect 22152 28697 22161 28731
rect 22161 28697 22195 28731
rect 22195 28697 22204 28731
rect 22152 28688 22204 28697
rect 23624 28731 23676 28740
rect 23624 28697 23633 28731
rect 23633 28697 23667 28731
rect 23667 28697 23676 28731
rect 23624 28688 23676 28697
rect 24728 28688 24780 28740
rect 25280 28688 25332 28740
rect 27488 28765 27497 28799
rect 27497 28765 27531 28799
rect 27531 28765 27540 28799
rect 27488 28756 27540 28765
rect 27396 28731 27448 28740
rect 27396 28697 27405 28731
rect 27405 28697 27439 28731
rect 27439 28697 27448 28731
rect 27396 28688 27448 28697
rect 27856 28688 27908 28740
rect 28960 28688 29012 28740
rect 22612 28620 22664 28672
rect 22796 28663 22848 28672
rect 22796 28629 22805 28663
rect 22805 28629 22839 28663
rect 22839 28629 22848 28663
rect 22796 28620 22848 28629
rect 25464 28663 25516 28672
rect 16632 28552 16684 28604
rect 18380 28595 18432 28604
rect 18380 28561 18389 28595
rect 18389 28561 18423 28595
rect 18423 28561 18432 28595
rect 18380 28552 18432 28561
rect 21968 28595 22020 28604
rect 18288 28484 18340 28536
rect 19668 28484 19720 28536
rect 20220 28484 20272 28536
rect 20772 28484 20824 28536
rect 21968 28561 21977 28595
rect 21977 28561 22011 28595
rect 22011 28561 22020 28595
rect 21968 28552 22020 28561
rect 25464 28629 25473 28663
rect 25473 28629 25507 28663
rect 25507 28629 25516 28663
rect 25464 28620 25516 28629
rect 29604 28620 29656 28672
rect 28592 28484 28644 28536
rect 14142 28382 14194 28434
rect 14206 28382 14258 28434
rect 14270 28382 14322 28434
rect 14334 28382 14386 28434
rect 24142 28382 24194 28434
rect 24206 28382 24258 28434
rect 24270 28382 24322 28434
rect 24334 28382 24386 28434
rect 15160 28280 15212 28332
rect 12492 28212 12544 28264
rect 20680 28280 20732 28332
rect 13964 28144 14016 28196
rect 15068 28144 15120 28196
rect 15436 28187 15488 28196
rect 15436 28153 15445 28187
rect 15445 28153 15479 28187
rect 15479 28153 15488 28187
rect 15436 28144 15488 28153
rect 16632 28144 16684 28196
rect 22520 28212 22572 28264
rect 23348 28212 23400 28264
rect 24728 28212 24780 28264
rect 14700 28119 14752 28128
rect 14700 28085 14709 28119
rect 14709 28085 14743 28119
rect 14743 28085 14752 28119
rect 14700 28076 14752 28085
rect 15988 28119 16040 28128
rect 15988 28085 15997 28119
rect 15997 28085 16031 28119
rect 16031 28085 16040 28119
rect 15988 28076 16040 28085
rect 16724 28076 16776 28128
rect 18012 28076 18064 28128
rect 17828 28051 17880 28060
rect 17828 28017 17837 28051
rect 17837 28017 17871 28051
rect 17871 28017 17880 28051
rect 17828 28008 17880 28017
rect 19760 28144 19812 28196
rect 18564 28119 18616 28128
rect 18564 28085 18573 28119
rect 18573 28085 18607 28119
rect 18607 28085 18616 28119
rect 18564 28076 18616 28085
rect 22704 28144 22756 28196
rect 19944 28076 19996 28128
rect 21784 28076 21836 28128
rect 23716 28076 23768 28128
rect 25372 28119 25424 28128
rect 18380 27940 18432 27992
rect 20036 28008 20088 28060
rect 20588 28051 20640 28060
rect 20588 28017 20597 28051
rect 20597 28017 20631 28051
rect 20631 28017 20640 28051
rect 20588 28008 20640 28017
rect 23808 28008 23860 28060
rect 25372 28085 25381 28119
rect 25381 28085 25415 28119
rect 25415 28085 25424 28119
rect 25372 28076 25424 28085
rect 26292 28008 26344 28060
rect 27396 28008 27448 28060
rect 28224 28008 28276 28060
rect 20496 27940 20548 27992
rect 25372 27940 25424 27992
rect 26384 27940 26436 27992
rect 28316 27940 28368 27992
rect 19142 27838 19194 27890
rect 19206 27838 19258 27890
rect 19270 27838 19322 27890
rect 19334 27838 19386 27890
rect 29142 27838 29194 27890
rect 29206 27838 29258 27890
rect 29270 27838 29322 27890
rect 29334 27838 29386 27890
rect 17644 27736 17696 27788
rect 17828 27736 17880 27788
rect 11940 27600 11992 27652
rect 18840 27668 18892 27720
rect 19484 27668 19536 27720
rect 20312 27711 20364 27720
rect 18288 27643 18340 27652
rect 18288 27609 18297 27643
rect 18297 27609 18331 27643
rect 18331 27609 18340 27643
rect 18288 27600 18340 27609
rect 18012 27575 18064 27584
rect 18012 27541 18021 27575
rect 18021 27541 18055 27575
rect 18055 27541 18064 27575
rect 18012 27532 18064 27541
rect 19024 27600 19076 27652
rect 19760 27643 19812 27652
rect 19760 27609 19769 27643
rect 19769 27609 19803 27643
rect 19803 27609 19812 27643
rect 19760 27600 19812 27609
rect 19392 27532 19444 27584
rect 20312 27677 20321 27711
rect 20321 27677 20355 27711
rect 20355 27677 20364 27711
rect 20312 27668 20364 27677
rect 20496 27736 20548 27788
rect 28224 27736 28276 27788
rect 27396 27711 27448 27720
rect 21784 27643 21836 27652
rect 21784 27609 21793 27643
rect 21793 27609 21827 27643
rect 21827 27609 21836 27643
rect 21784 27600 21836 27609
rect 22612 27643 22664 27652
rect 22612 27609 22621 27643
rect 22621 27609 22655 27643
rect 22655 27609 22664 27643
rect 22612 27600 22664 27609
rect 23072 27600 23124 27652
rect 23532 27600 23584 27652
rect 24912 27600 24964 27652
rect 25280 27600 25332 27652
rect 25832 27643 25884 27652
rect 20680 27532 20732 27584
rect 23256 27532 23308 27584
rect 23348 27575 23400 27584
rect 23348 27541 23357 27575
rect 23357 27541 23391 27575
rect 23391 27541 23400 27575
rect 23348 27532 23400 27541
rect 23900 27532 23952 27584
rect 25832 27609 25841 27643
rect 25841 27609 25875 27643
rect 25875 27609 25884 27643
rect 25832 27600 25884 27609
rect 27396 27677 27405 27711
rect 27405 27677 27439 27711
rect 27439 27677 27448 27711
rect 27396 27668 27448 27677
rect 28408 27600 28460 27652
rect 29512 27600 29564 27652
rect 27764 27532 27816 27584
rect 25096 27464 25148 27516
rect 29144 27507 29196 27516
rect 29144 27473 29153 27507
rect 29153 27473 29187 27507
rect 29187 27473 29196 27507
rect 29144 27464 29196 27473
rect 12308 27396 12360 27448
rect 14792 27396 14844 27448
rect 19576 27396 19628 27448
rect 19668 27396 19720 27448
rect 23348 27396 23400 27448
rect 27028 27396 27080 27448
rect 14142 27294 14194 27346
rect 14206 27294 14258 27346
rect 14270 27294 14322 27346
rect 14334 27294 14386 27346
rect 24142 27294 24194 27346
rect 24206 27294 24258 27346
rect 24270 27294 24322 27346
rect 24334 27294 24386 27346
rect 18012 27192 18064 27244
rect 18748 27192 18800 27244
rect 19668 27192 19720 27244
rect 19392 27124 19444 27176
rect 22152 27192 22204 27244
rect 25740 27192 25792 27244
rect 20036 27124 20088 27176
rect 23992 27124 24044 27176
rect 27396 27124 27448 27176
rect 16908 27056 16960 27108
rect 19024 27056 19076 27108
rect 20588 27056 20640 27108
rect 23808 27099 23860 27108
rect 23808 27065 23817 27099
rect 23817 27065 23851 27099
rect 23851 27065 23860 27099
rect 23808 27056 23860 27065
rect 24452 27056 24504 27108
rect 25832 27056 25884 27108
rect 26384 27056 26436 27108
rect 27212 27099 27264 27108
rect 27212 27065 27221 27099
rect 27221 27065 27255 27099
rect 27255 27065 27264 27099
rect 27212 27056 27264 27065
rect 28408 27099 28460 27108
rect 28408 27065 28417 27099
rect 28417 27065 28451 27099
rect 28451 27065 28460 27099
rect 28408 27056 28460 27065
rect 28868 27056 28920 27108
rect 11296 27031 11348 27040
rect 11296 26997 11305 27031
rect 11305 26997 11339 27031
rect 11339 26997 11348 27031
rect 11296 26988 11348 26997
rect 17736 26988 17788 27040
rect 11572 26963 11624 26972
rect 11572 26929 11581 26963
rect 11581 26929 11615 26963
rect 11615 26929 11624 26963
rect 11572 26920 11624 26929
rect 12308 26920 12360 26972
rect 13228 26920 13280 26972
rect 14056 26963 14108 26972
rect 14056 26929 14065 26963
rect 14065 26929 14099 26963
rect 14099 26929 14108 26963
rect 14056 26920 14108 26929
rect 14792 26920 14844 26972
rect 15804 26963 15856 26972
rect 15804 26929 15813 26963
rect 15813 26929 15847 26963
rect 15847 26929 15856 26963
rect 15804 26920 15856 26929
rect 16724 26963 16776 26972
rect 16724 26929 16733 26963
rect 16733 26929 16767 26963
rect 16767 26929 16776 26963
rect 16724 26920 16776 26929
rect 16908 26895 16960 26904
rect 16908 26861 16917 26895
rect 16917 26861 16951 26895
rect 16951 26861 16960 26895
rect 16908 26852 16960 26861
rect 17828 26852 17880 26904
rect 18748 26988 18800 27040
rect 18932 26963 18984 26972
rect 18932 26929 18941 26963
rect 18941 26929 18975 26963
rect 18975 26929 18984 26963
rect 18932 26920 18984 26929
rect 19024 26920 19076 26972
rect 19576 26988 19628 27040
rect 19944 26988 19996 27040
rect 20220 26988 20272 27040
rect 22060 26988 22112 27040
rect 23716 27031 23768 27040
rect 23716 26997 23725 27031
rect 23725 26997 23759 27031
rect 23759 26997 23768 27031
rect 23716 26988 23768 26997
rect 24912 26988 24964 27040
rect 25556 27031 25608 27040
rect 25556 26997 25565 27031
rect 25565 26997 25599 27031
rect 25599 26997 25608 27031
rect 25556 26988 25608 26997
rect 19484 26852 19536 26904
rect 21600 26920 21652 26972
rect 22520 26963 22572 26972
rect 22520 26929 22529 26963
rect 22529 26929 22563 26963
rect 22563 26929 22572 26963
rect 22520 26920 22572 26929
rect 28500 26920 28552 26972
rect 29144 26920 29196 26972
rect 20312 26895 20364 26904
rect 20312 26861 20321 26895
rect 20321 26861 20355 26895
rect 20355 26861 20364 26895
rect 20312 26852 20364 26861
rect 20404 26895 20456 26904
rect 20404 26861 20413 26895
rect 20413 26861 20447 26895
rect 20447 26861 20456 26895
rect 20404 26852 20456 26861
rect 26476 26852 26528 26904
rect 19142 26750 19194 26802
rect 19206 26750 19258 26802
rect 19270 26750 19322 26802
rect 19334 26750 19386 26802
rect 29142 26750 29194 26802
rect 29206 26750 29258 26802
rect 29270 26750 29322 26802
rect 29334 26750 29386 26802
rect 15804 26648 15856 26700
rect 20312 26691 20364 26700
rect 11572 26580 11624 26632
rect 12584 26512 12636 26564
rect 12676 26555 12728 26564
rect 12676 26521 12685 26555
rect 12685 26521 12719 26555
rect 12719 26521 12728 26555
rect 12860 26555 12912 26564
rect 12676 26512 12728 26521
rect 12860 26521 12869 26555
rect 12869 26521 12903 26555
rect 12903 26521 12912 26555
rect 12860 26512 12912 26521
rect 13228 26555 13280 26564
rect 13228 26521 13237 26555
rect 13237 26521 13271 26555
rect 13271 26521 13280 26555
rect 13228 26512 13280 26521
rect 15252 26555 15304 26564
rect 15252 26521 15261 26555
rect 15261 26521 15295 26555
rect 15295 26521 15304 26555
rect 15252 26512 15304 26521
rect 13136 26444 13188 26496
rect 15344 26444 15396 26496
rect 13228 26376 13280 26428
rect 17552 26512 17604 26564
rect 20312 26657 20321 26691
rect 20321 26657 20355 26691
rect 20355 26657 20364 26691
rect 20312 26648 20364 26657
rect 22520 26648 22572 26700
rect 23624 26648 23676 26700
rect 26384 26691 26436 26700
rect 17828 26623 17880 26632
rect 17828 26589 17837 26623
rect 17837 26589 17871 26623
rect 17871 26589 17880 26623
rect 17828 26580 17880 26589
rect 18012 26580 18064 26632
rect 19944 26580 19996 26632
rect 20404 26623 20456 26632
rect 20404 26589 20413 26623
rect 20413 26589 20447 26623
rect 20447 26589 20456 26623
rect 20404 26580 20456 26589
rect 20680 26580 20732 26632
rect 21600 26580 21652 26632
rect 22060 26623 22112 26632
rect 22060 26589 22069 26623
rect 22069 26589 22103 26623
rect 22103 26589 22112 26623
rect 22060 26580 22112 26589
rect 23716 26623 23768 26632
rect 23716 26589 23725 26623
rect 23725 26589 23759 26623
rect 23759 26589 23768 26623
rect 23716 26580 23768 26589
rect 17736 26555 17788 26564
rect 17736 26521 17745 26555
rect 17745 26521 17779 26555
rect 17779 26521 17788 26555
rect 17736 26512 17788 26521
rect 16724 26444 16776 26496
rect 18932 26512 18984 26564
rect 19484 26512 19536 26564
rect 21692 26555 21744 26564
rect 21692 26521 21701 26555
rect 21701 26521 21735 26555
rect 21735 26521 21744 26555
rect 21692 26512 21744 26521
rect 21876 26512 21928 26564
rect 18472 26444 18524 26496
rect 19944 26444 19996 26496
rect 21784 26444 21836 26496
rect 22888 26512 22940 26564
rect 25832 26512 25884 26564
rect 26384 26657 26393 26691
rect 26393 26657 26427 26691
rect 26427 26657 26436 26691
rect 26384 26648 26436 26657
rect 27120 26580 27172 26632
rect 27764 26580 27816 26632
rect 28500 26623 28552 26632
rect 28500 26589 28509 26623
rect 28509 26589 28543 26623
rect 28543 26589 28552 26623
rect 28500 26580 28552 26589
rect 18288 26376 18340 26428
rect 24912 26444 24964 26496
rect 26476 26512 26528 26564
rect 28960 26512 29012 26564
rect 26384 26376 26436 26428
rect 27580 26376 27632 26428
rect 14976 26308 15028 26360
rect 16724 26308 16776 26360
rect 14142 26206 14194 26258
rect 14206 26206 14258 26258
rect 14270 26206 14322 26258
rect 14334 26206 14386 26258
rect 24142 26206 24194 26258
rect 24206 26206 24258 26258
rect 24270 26206 24322 26258
rect 24334 26206 24386 26258
rect 12584 26147 12636 26156
rect 12584 26113 12593 26147
rect 12593 26113 12627 26147
rect 12627 26113 12636 26147
rect 12584 26104 12636 26113
rect 12860 26036 12912 26088
rect 14056 25968 14108 26020
rect 11664 25943 11716 25952
rect 11664 25909 11673 25943
rect 11673 25909 11707 25943
rect 11707 25909 11716 25943
rect 11664 25900 11716 25909
rect 12768 25943 12820 25952
rect 12768 25909 12777 25943
rect 12777 25909 12811 25943
rect 12811 25909 12820 25943
rect 12768 25900 12820 25909
rect 13504 25900 13556 25952
rect 14516 25900 14568 25952
rect 25556 26104 25608 26156
rect 15252 26011 15304 26020
rect 15252 25977 15261 26011
rect 15261 25977 15295 26011
rect 15295 25977 15304 26011
rect 15252 25968 15304 25977
rect 15344 26011 15396 26020
rect 15344 25977 15353 26011
rect 15353 25977 15387 26011
rect 15387 25977 15396 26011
rect 15344 25968 15396 25977
rect 14884 25900 14936 25952
rect 15712 25832 15764 25884
rect 18012 25968 18064 26020
rect 16908 25943 16960 25952
rect 16724 25875 16776 25884
rect 16724 25841 16733 25875
rect 16733 25841 16767 25875
rect 16767 25841 16776 25875
rect 16724 25832 16776 25841
rect 14884 25764 14936 25816
rect 14976 25764 15028 25816
rect 16908 25909 16917 25943
rect 16917 25909 16951 25943
rect 16951 25909 16960 25943
rect 16908 25900 16960 25909
rect 17184 25900 17236 25952
rect 17736 25900 17788 25952
rect 18564 25968 18616 26020
rect 21784 25968 21836 26020
rect 25372 26011 25424 26020
rect 25372 25977 25381 26011
rect 25381 25977 25415 26011
rect 25415 25977 25424 26011
rect 25372 25968 25424 25977
rect 18196 25900 18248 25952
rect 18932 25900 18984 25952
rect 21416 25943 21468 25952
rect 21416 25909 21425 25943
rect 21425 25909 21459 25943
rect 21459 25909 21468 25943
rect 21416 25900 21468 25909
rect 21692 25900 21744 25952
rect 25280 25943 25332 25952
rect 17276 25832 17328 25884
rect 17552 25832 17604 25884
rect 19024 25832 19076 25884
rect 16908 25764 16960 25816
rect 17000 25807 17052 25816
rect 17000 25773 17009 25807
rect 17009 25773 17043 25807
rect 17043 25773 17052 25807
rect 17000 25764 17052 25773
rect 18104 25764 18156 25816
rect 18380 25764 18432 25816
rect 20588 25832 20640 25884
rect 21232 25875 21284 25884
rect 21232 25841 21241 25875
rect 21241 25841 21275 25875
rect 21275 25841 21284 25875
rect 21232 25832 21284 25841
rect 22520 25832 22572 25884
rect 22888 25832 22940 25884
rect 25280 25909 25289 25943
rect 25289 25909 25323 25943
rect 25323 25909 25332 25943
rect 25280 25900 25332 25909
rect 27120 26036 27172 26088
rect 28684 26036 28736 26088
rect 26476 26011 26528 26020
rect 26476 25977 26485 26011
rect 26485 25977 26519 26011
rect 26519 25977 26528 26011
rect 26476 25968 26528 25977
rect 27028 26011 27080 26020
rect 27028 25977 27037 26011
rect 27037 25977 27071 26011
rect 27071 25977 27080 26011
rect 27028 25968 27080 25977
rect 28776 25968 28828 26020
rect 25740 25943 25792 25952
rect 25740 25909 25749 25943
rect 25749 25909 25783 25943
rect 25783 25909 25792 25943
rect 25740 25900 25792 25909
rect 28040 25900 28092 25952
rect 24176 25832 24228 25884
rect 21692 25764 21744 25816
rect 23440 25764 23492 25816
rect 19142 25662 19194 25714
rect 19206 25662 19258 25714
rect 19270 25662 19322 25714
rect 19334 25662 19386 25714
rect 29142 25662 29194 25714
rect 29206 25662 29258 25714
rect 29270 25662 29322 25714
rect 29334 25662 29386 25714
rect 12676 25560 12728 25612
rect 15712 25603 15764 25612
rect 15712 25569 15721 25603
rect 15721 25569 15755 25603
rect 15755 25569 15764 25603
rect 15712 25560 15764 25569
rect 17184 25560 17236 25612
rect 18840 25603 18892 25612
rect 12768 25535 12820 25544
rect 12768 25501 12777 25535
rect 12777 25501 12811 25535
rect 12811 25501 12820 25535
rect 12768 25492 12820 25501
rect 14608 25492 14660 25544
rect 11940 25467 11992 25476
rect 11940 25433 11949 25467
rect 11949 25433 11983 25467
rect 11983 25433 11992 25467
rect 11940 25424 11992 25433
rect 13504 25424 13556 25476
rect 14792 25467 14844 25476
rect 14792 25433 14801 25467
rect 14801 25433 14835 25467
rect 14835 25433 14844 25467
rect 14792 25424 14844 25433
rect 14884 25424 14936 25476
rect 17000 25492 17052 25544
rect 18840 25569 18849 25603
rect 18849 25569 18883 25603
rect 18883 25569 18892 25603
rect 18840 25560 18892 25569
rect 19760 25560 19812 25612
rect 21508 25560 21560 25612
rect 25280 25560 25332 25612
rect 25464 25560 25516 25612
rect 27948 25560 28000 25612
rect 20220 25492 20272 25544
rect 18380 25467 18432 25476
rect 14516 25399 14568 25408
rect 14516 25365 14525 25399
rect 14525 25365 14559 25399
rect 14559 25365 14568 25399
rect 14516 25356 14568 25365
rect 14976 25399 15028 25408
rect 14976 25365 14985 25399
rect 14985 25365 15019 25399
rect 15019 25365 15028 25399
rect 14976 25356 15028 25365
rect 16264 25356 16316 25408
rect 16724 25356 16776 25408
rect 17552 25356 17604 25408
rect 12124 25263 12176 25272
rect 12124 25229 12133 25263
rect 12133 25229 12167 25263
rect 12167 25229 12176 25263
rect 12124 25220 12176 25229
rect 18380 25433 18386 25467
rect 18386 25433 18432 25467
rect 18380 25424 18432 25433
rect 18472 25424 18524 25476
rect 18564 25399 18616 25408
rect 18564 25365 18573 25399
rect 18573 25365 18607 25399
rect 18607 25365 18616 25399
rect 18564 25356 18616 25365
rect 19484 25356 19536 25408
rect 19852 25424 19904 25476
rect 21600 25492 21652 25544
rect 23164 25492 23216 25544
rect 20404 25399 20456 25408
rect 20404 25365 20413 25399
rect 20413 25365 20447 25399
rect 20447 25365 20456 25399
rect 20404 25356 20456 25365
rect 21048 25356 21100 25408
rect 21876 25399 21928 25408
rect 21876 25365 21885 25399
rect 21885 25365 21919 25399
rect 21919 25365 21928 25399
rect 21876 25356 21928 25365
rect 22428 25356 22480 25408
rect 23900 25424 23952 25476
rect 24820 25424 24872 25476
rect 25740 25492 25792 25544
rect 26936 25492 26988 25544
rect 25464 25424 25516 25476
rect 27580 25467 27632 25476
rect 27580 25433 27589 25467
rect 27589 25433 27623 25467
rect 27623 25433 27632 25467
rect 27580 25424 27632 25433
rect 28684 25492 28736 25544
rect 29512 25492 29564 25544
rect 28040 25424 28092 25476
rect 23532 25356 23584 25408
rect 24176 25399 24228 25408
rect 24176 25365 24185 25399
rect 24185 25365 24219 25399
rect 24219 25365 24228 25399
rect 24176 25356 24228 25365
rect 25004 25356 25056 25408
rect 27028 25399 27080 25408
rect 27028 25365 27037 25399
rect 27037 25365 27071 25399
rect 27071 25365 27080 25399
rect 27028 25356 27080 25365
rect 18840 25288 18892 25340
rect 25924 25288 25976 25340
rect 23808 25220 23860 25272
rect 24636 25220 24688 25272
rect 14142 25118 14194 25170
rect 14206 25118 14258 25170
rect 14270 25118 14322 25170
rect 14334 25118 14386 25170
rect 24142 25118 24194 25170
rect 24206 25118 24258 25170
rect 24270 25118 24322 25170
rect 24334 25118 24386 25170
rect 18564 25016 18616 25068
rect 14516 24948 14568 25000
rect 17552 24948 17604 25000
rect 20404 24948 20456 25000
rect 11296 24855 11348 24864
rect 11296 24821 11305 24855
rect 11305 24821 11339 24855
rect 11339 24821 11348 24855
rect 11296 24812 11348 24821
rect 14884 24880 14936 24932
rect 16724 24880 16776 24932
rect 18288 24880 18340 24932
rect 18932 24923 18984 24932
rect 18932 24889 18941 24923
rect 18941 24889 18975 24923
rect 18975 24889 18984 24923
rect 18932 24880 18984 24889
rect 19484 24880 19536 24932
rect 14516 24855 14568 24864
rect 14516 24821 14525 24855
rect 14525 24821 14559 24855
rect 14559 24821 14568 24855
rect 15804 24855 15856 24864
rect 14516 24812 14568 24821
rect 15804 24821 15813 24855
rect 15813 24821 15847 24855
rect 15847 24821 15856 24855
rect 15804 24812 15856 24821
rect 22336 25016 22388 25068
rect 21048 24948 21100 25000
rect 23440 25016 23492 25068
rect 25464 25016 25516 25068
rect 28040 25059 28092 25068
rect 28040 25025 28049 25059
rect 28049 25025 28083 25059
rect 28083 25025 28092 25059
rect 28040 25016 28092 25025
rect 22428 24812 22480 24864
rect 23164 24880 23216 24932
rect 23532 24948 23584 25000
rect 23440 24812 23492 24864
rect 23808 24812 23860 24864
rect 25004 24880 25056 24932
rect 24544 24812 24596 24864
rect 25556 24948 25608 25000
rect 28316 24948 28368 25000
rect 25924 24923 25976 24932
rect 25924 24889 25933 24923
rect 25933 24889 25967 24923
rect 25967 24889 25976 24923
rect 25924 24880 25976 24889
rect 26752 24880 26804 24932
rect 28960 24880 29012 24932
rect 26016 24855 26068 24864
rect 26016 24821 26025 24855
rect 26025 24821 26059 24855
rect 26059 24821 26068 24855
rect 26016 24812 26068 24821
rect 27948 24855 28000 24864
rect 27948 24821 27957 24855
rect 27957 24821 27991 24855
rect 27991 24821 28000 24855
rect 27948 24812 28000 24821
rect 28592 24855 28644 24864
rect 28592 24821 28601 24855
rect 28601 24821 28635 24855
rect 28635 24821 28644 24855
rect 28592 24812 28644 24821
rect 11572 24787 11624 24796
rect 11572 24753 11581 24787
rect 11581 24753 11615 24787
rect 11615 24753 11624 24787
rect 11572 24744 11624 24753
rect 12124 24744 12176 24796
rect 13412 24744 13464 24796
rect 15620 24787 15672 24796
rect 15620 24753 15629 24787
rect 15629 24753 15663 24787
rect 15663 24753 15672 24787
rect 15620 24744 15672 24753
rect 16816 24744 16868 24796
rect 17184 24744 17236 24796
rect 18104 24744 18156 24796
rect 18840 24744 18892 24796
rect 19760 24787 19812 24796
rect 19760 24753 19769 24787
rect 19769 24753 19803 24787
rect 19803 24753 19812 24787
rect 19760 24744 19812 24753
rect 20588 24787 20640 24796
rect 20588 24753 20597 24787
rect 20597 24753 20631 24787
rect 20631 24753 20640 24787
rect 20588 24744 20640 24753
rect 23348 24744 23400 24796
rect 25372 24744 25424 24796
rect 28132 24744 28184 24796
rect 17000 24676 17052 24728
rect 17368 24719 17420 24728
rect 17368 24685 17377 24719
rect 17377 24685 17411 24719
rect 17411 24685 17420 24719
rect 17368 24676 17420 24685
rect 17552 24676 17604 24728
rect 19668 24719 19720 24728
rect 19668 24685 19677 24719
rect 19677 24685 19711 24719
rect 19711 24685 19720 24719
rect 19668 24676 19720 24685
rect 19852 24676 19904 24728
rect 26568 24676 26620 24728
rect 27028 24719 27080 24728
rect 27028 24685 27037 24719
rect 27037 24685 27071 24719
rect 27071 24685 27080 24719
rect 27028 24676 27080 24685
rect 27212 24676 27264 24728
rect 19142 24574 19194 24626
rect 19206 24574 19258 24626
rect 19270 24574 19322 24626
rect 19334 24574 19386 24626
rect 29142 24574 29194 24626
rect 29206 24574 29258 24626
rect 29270 24574 29322 24626
rect 29334 24574 29386 24626
rect 12124 24336 12176 24388
rect 12400 24336 12452 24388
rect 13412 24336 13464 24388
rect 15988 24472 16040 24524
rect 16724 24472 16776 24524
rect 18012 24472 18064 24524
rect 19668 24472 19720 24524
rect 21508 24515 21560 24524
rect 21508 24481 21517 24515
rect 21517 24481 21551 24515
rect 21551 24481 21560 24515
rect 21508 24472 21560 24481
rect 27212 24472 27264 24524
rect 27764 24515 27816 24524
rect 27764 24481 27773 24515
rect 27773 24481 27807 24515
rect 27807 24481 27816 24515
rect 27764 24472 27816 24481
rect 16816 24336 16868 24388
rect 15988 24311 16040 24320
rect 15988 24277 15994 24311
rect 15994 24277 16040 24311
rect 15988 24268 16040 24277
rect 16172 24311 16224 24320
rect 16172 24277 16181 24311
rect 16181 24277 16215 24311
rect 16215 24277 16224 24311
rect 16172 24268 16224 24277
rect 18196 24404 18248 24456
rect 18380 24404 18432 24456
rect 17276 24379 17328 24388
rect 17276 24345 17285 24379
rect 17285 24345 17319 24379
rect 17319 24345 17328 24379
rect 17276 24336 17328 24345
rect 19760 24336 19812 24388
rect 20128 24336 20180 24388
rect 18564 24243 18616 24252
rect 18564 24209 18573 24243
rect 18573 24209 18607 24243
rect 18607 24209 18616 24243
rect 18564 24200 18616 24209
rect 19668 24268 19720 24320
rect 20956 24336 21008 24388
rect 22060 24336 22112 24388
rect 23164 24379 23216 24388
rect 23164 24345 23173 24379
rect 23173 24345 23207 24379
rect 23207 24345 23216 24379
rect 23164 24336 23216 24345
rect 23808 24404 23860 24456
rect 26752 24404 26804 24456
rect 25556 24336 25608 24388
rect 26016 24336 26068 24388
rect 26476 24379 26528 24388
rect 26476 24345 26485 24379
rect 26485 24345 26519 24379
rect 26519 24345 26528 24379
rect 26476 24336 26528 24345
rect 26844 24379 26896 24388
rect 26844 24345 26853 24379
rect 26853 24345 26887 24379
rect 26887 24345 26896 24379
rect 26844 24336 26896 24345
rect 26936 24379 26988 24388
rect 26936 24345 26945 24379
rect 26945 24345 26979 24379
rect 26979 24345 26988 24379
rect 26936 24336 26988 24345
rect 28132 24379 28184 24388
rect 28132 24345 28141 24379
rect 28141 24345 28175 24379
rect 28175 24345 28184 24379
rect 28132 24336 28184 24345
rect 28500 24379 28552 24388
rect 28500 24345 28509 24379
rect 28509 24345 28543 24379
rect 28543 24345 28552 24379
rect 28500 24336 28552 24345
rect 12032 24132 12084 24184
rect 12952 24132 13004 24184
rect 15988 24132 16040 24184
rect 16172 24132 16224 24184
rect 18196 24132 18248 24184
rect 18472 24132 18524 24184
rect 18656 24132 18708 24184
rect 23164 24200 23216 24252
rect 23624 24200 23676 24252
rect 21232 24132 21284 24184
rect 23440 24175 23492 24184
rect 23440 24141 23449 24175
rect 23449 24141 23483 24175
rect 23483 24141 23492 24175
rect 23440 24132 23492 24141
rect 23808 24175 23860 24184
rect 23808 24141 23817 24175
rect 23817 24141 23851 24175
rect 23851 24141 23860 24175
rect 23808 24132 23860 24141
rect 26108 24175 26160 24184
rect 26108 24141 26117 24175
rect 26117 24141 26151 24175
rect 26151 24141 26160 24175
rect 26108 24132 26160 24141
rect 26844 24200 26896 24252
rect 29328 24404 29380 24456
rect 29512 24472 29564 24524
rect 29512 24336 29564 24388
rect 28500 24132 28552 24184
rect 14142 24030 14194 24082
rect 14206 24030 14258 24082
rect 14270 24030 14322 24082
rect 14334 24030 14386 24082
rect 24142 24030 24194 24082
rect 24206 24030 24258 24082
rect 24270 24030 24322 24082
rect 24334 24030 24386 24082
rect 14884 23928 14936 23980
rect 21048 23928 21100 23980
rect 21508 23928 21560 23980
rect 29328 23928 29380 23980
rect 14792 23860 14844 23912
rect 15988 23860 16040 23912
rect 17184 23860 17236 23912
rect 17552 23860 17604 23912
rect 11572 23835 11624 23844
rect 11572 23801 11581 23835
rect 11581 23801 11615 23835
rect 11615 23801 11624 23835
rect 11572 23792 11624 23801
rect 13412 23792 13464 23844
rect 14700 23835 14752 23844
rect 14700 23801 14709 23835
rect 14709 23801 14743 23835
rect 14743 23801 14752 23835
rect 14700 23792 14752 23801
rect 18748 23860 18800 23912
rect 23624 23860 23676 23912
rect 23716 23860 23768 23912
rect 12032 23767 12084 23776
rect 12032 23733 12041 23767
rect 12041 23733 12075 23767
rect 12075 23733 12084 23767
rect 12032 23724 12084 23733
rect 12216 23767 12268 23776
rect 12216 23733 12225 23767
rect 12225 23733 12259 23767
rect 12259 23733 12268 23767
rect 12216 23724 12268 23733
rect 13044 23767 13096 23776
rect 13044 23733 13053 23767
rect 13053 23733 13087 23767
rect 13087 23733 13096 23767
rect 13044 23724 13096 23733
rect 13504 23767 13556 23776
rect 13504 23733 13513 23767
rect 13513 23733 13547 23767
rect 13547 23733 13556 23767
rect 13504 23724 13556 23733
rect 13964 23724 14016 23776
rect 15068 23724 15120 23776
rect 15252 23792 15304 23844
rect 18288 23792 18340 23844
rect 12584 23656 12636 23708
rect 14976 23656 15028 23708
rect 17368 23724 17420 23776
rect 18656 23724 18708 23776
rect 19024 23792 19076 23844
rect 21048 23792 21100 23844
rect 21876 23792 21928 23844
rect 23348 23792 23400 23844
rect 23900 23835 23952 23844
rect 23900 23801 23909 23835
rect 23909 23801 23943 23835
rect 23943 23801 23952 23835
rect 23900 23792 23952 23801
rect 26016 23860 26068 23912
rect 20128 23767 20180 23776
rect 20128 23733 20137 23767
rect 20137 23733 20171 23767
rect 20171 23733 20180 23767
rect 20128 23724 20180 23733
rect 20956 23724 21008 23776
rect 21324 23724 21376 23776
rect 22060 23724 22112 23776
rect 22980 23724 23032 23776
rect 23532 23767 23584 23776
rect 23532 23733 23541 23767
rect 23541 23733 23575 23767
rect 23575 23733 23584 23767
rect 23532 23724 23584 23733
rect 23716 23724 23768 23776
rect 25924 23792 25976 23844
rect 26108 23767 26160 23776
rect 16172 23656 16224 23708
rect 16816 23656 16868 23708
rect 13596 23631 13648 23640
rect 13596 23597 13605 23631
rect 13605 23597 13639 23631
rect 13639 23597 13648 23631
rect 13596 23588 13648 23597
rect 15620 23588 15672 23640
rect 19484 23656 19536 23708
rect 19576 23588 19628 23640
rect 20864 23656 20916 23708
rect 22428 23588 22480 23640
rect 26108 23733 26117 23767
rect 26117 23733 26151 23767
rect 26151 23733 26160 23767
rect 26108 23724 26160 23733
rect 27764 23792 27816 23844
rect 28500 23835 28552 23844
rect 28500 23801 28509 23835
rect 28509 23801 28543 23835
rect 28543 23801 28552 23835
rect 28500 23792 28552 23801
rect 27396 23724 27448 23776
rect 29144 23767 29196 23776
rect 29144 23733 29153 23767
rect 29153 23733 29187 23767
rect 29187 23733 29196 23767
rect 29144 23724 29196 23733
rect 28408 23699 28460 23708
rect 28408 23665 28417 23699
rect 28417 23665 28451 23699
rect 28451 23665 28460 23699
rect 28408 23656 28460 23665
rect 26200 23631 26252 23640
rect 26200 23597 26209 23631
rect 26209 23597 26243 23631
rect 26243 23597 26252 23631
rect 26200 23588 26252 23597
rect 19142 23486 19194 23538
rect 19206 23486 19258 23538
rect 19270 23486 19322 23538
rect 19334 23486 19386 23538
rect 29142 23486 29194 23538
rect 29206 23486 29258 23538
rect 29270 23486 29322 23538
rect 29334 23486 29386 23538
rect 12124 23316 12176 23368
rect 14792 23384 14844 23436
rect 17092 23384 17144 23436
rect 18196 23427 18248 23436
rect 18196 23393 18205 23427
rect 18205 23393 18239 23427
rect 18239 23393 18248 23427
rect 18196 23384 18248 23393
rect 19668 23427 19720 23436
rect 19668 23393 19677 23427
rect 19677 23393 19711 23427
rect 19711 23393 19720 23427
rect 19668 23384 19720 23393
rect 20864 23427 20916 23436
rect 20864 23393 20873 23427
rect 20873 23393 20907 23427
rect 20907 23393 20916 23427
rect 20864 23384 20916 23393
rect 20956 23384 21008 23436
rect 13596 23316 13648 23368
rect 13228 23291 13280 23300
rect 13228 23257 13237 23291
rect 13237 23257 13271 23291
rect 13271 23257 13280 23291
rect 13228 23248 13280 23257
rect 13412 23291 13464 23300
rect 13412 23257 13421 23291
rect 13421 23257 13455 23291
rect 13455 23257 13464 23291
rect 13412 23248 13464 23257
rect 13872 23248 13924 23300
rect 14516 23291 14568 23300
rect 12952 23223 13004 23232
rect 12952 23189 12961 23223
rect 12961 23189 12995 23223
rect 12995 23189 13004 23223
rect 12952 23180 13004 23189
rect 12400 23112 12452 23164
rect 14516 23257 14525 23291
rect 14525 23257 14559 23291
rect 14559 23257 14568 23291
rect 14516 23248 14568 23257
rect 15988 23316 16040 23368
rect 17000 23316 17052 23368
rect 22244 23316 22296 23368
rect 22520 23316 22572 23368
rect 23440 23316 23492 23368
rect 14884 23291 14936 23300
rect 14884 23257 14893 23291
rect 14893 23257 14927 23291
rect 14927 23257 14936 23291
rect 14884 23248 14936 23257
rect 15436 23291 15488 23300
rect 15436 23257 15445 23291
rect 15445 23257 15479 23291
rect 15479 23257 15488 23291
rect 15436 23248 15488 23257
rect 16172 23291 16224 23300
rect 16172 23257 16181 23291
rect 16181 23257 16215 23291
rect 16215 23257 16224 23291
rect 16172 23248 16224 23257
rect 17092 23248 17144 23300
rect 18012 23291 18064 23300
rect 18012 23257 18021 23291
rect 18021 23257 18055 23291
rect 18055 23257 18064 23291
rect 18012 23248 18064 23257
rect 18380 23291 18432 23300
rect 18380 23257 18389 23291
rect 18389 23257 18423 23291
rect 18423 23257 18432 23291
rect 18380 23248 18432 23257
rect 19576 23291 19628 23300
rect 15068 23223 15120 23232
rect 15068 23189 15077 23223
rect 15077 23189 15111 23223
rect 15111 23189 15120 23223
rect 15068 23180 15120 23189
rect 16264 23180 16316 23232
rect 16540 23180 16592 23232
rect 19576 23257 19585 23291
rect 19585 23257 19619 23291
rect 19619 23257 19628 23291
rect 19576 23248 19628 23257
rect 20036 23248 20088 23300
rect 20864 23248 20916 23300
rect 22060 23248 22112 23300
rect 23716 23316 23768 23368
rect 19760 23180 19812 23232
rect 19944 23180 19996 23232
rect 20404 23223 20456 23232
rect 20404 23189 20410 23223
rect 20410 23189 20456 23223
rect 20404 23180 20456 23189
rect 20496 23180 20548 23232
rect 20680 23180 20732 23232
rect 22888 23223 22940 23232
rect 22888 23189 22897 23223
rect 22897 23189 22931 23223
rect 22931 23189 22940 23223
rect 22888 23180 22940 23189
rect 23624 23248 23676 23300
rect 24544 23316 24596 23368
rect 28408 23316 28460 23368
rect 25096 23248 25148 23300
rect 27396 23291 27448 23300
rect 23440 23180 23492 23232
rect 24544 23180 24596 23232
rect 27396 23257 27405 23291
rect 27405 23257 27439 23291
rect 27439 23257 27448 23291
rect 27396 23248 27448 23257
rect 28224 23248 28276 23300
rect 17552 23044 17604 23096
rect 18196 23044 18248 23096
rect 19300 23044 19352 23096
rect 19760 23044 19812 23096
rect 20864 23044 20916 23096
rect 22428 23044 22480 23096
rect 23808 23112 23860 23164
rect 28316 23112 28368 23164
rect 23532 23044 23584 23096
rect 23900 23044 23952 23096
rect 26660 23044 26712 23096
rect 14142 22942 14194 22994
rect 14206 22942 14258 22994
rect 14270 22942 14322 22994
rect 14334 22942 14386 22994
rect 24142 22942 24194 22994
rect 24206 22942 24258 22994
rect 24270 22942 24322 22994
rect 24334 22942 24386 22994
rect 13228 22840 13280 22892
rect 15068 22840 15120 22892
rect 15252 22840 15304 22892
rect 16632 22840 16684 22892
rect 19668 22840 19720 22892
rect 12216 22747 12268 22756
rect 12216 22713 12225 22747
rect 12225 22713 12259 22747
rect 12259 22713 12268 22747
rect 12216 22704 12268 22713
rect 15436 22704 15488 22756
rect 17000 22704 17052 22756
rect 12124 22679 12176 22688
rect 12124 22645 12133 22679
rect 12133 22645 12167 22679
rect 12167 22645 12176 22679
rect 12124 22636 12176 22645
rect 12400 22679 12452 22688
rect 12400 22645 12409 22679
rect 12409 22645 12443 22679
rect 12443 22645 12452 22679
rect 12400 22636 12452 22645
rect 14792 22636 14844 22688
rect 15252 22679 15304 22688
rect 15252 22645 15261 22679
rect 15261 22645 15295 22679
rect 15295 22645 15304 22679
rect 15252 22636 15304 22645
rect 16632 22636 16684 22688
rect 17092 22679 17144 22688
rect 13688 22568 13740 22620
rect 14700 22568 14752 22620
rect 16172 22568 16224 22620
rect 17092 22645 17101 22679
rect 17101 22645 17135 22679
rect 17135 22645 17144 22679
rect 17092 22636 17144 22645
rect 18380 22704 18432 22756
rect 18748 22704 18800 22756
rect 18012 22636 18064 22688
rect 19300 22679 19352 22688
rect 19300 22645 19309 22679
rect 19309 22645 19343 22679
rect 19343 22645 19352 22679
rect 19300 22636 19352 22645
rect 17276 22568 17328 22620
rect 18104 22568 18156 22620
rect 20128 22772 20180 22824
rect 22796 22840 22848 22892
rect 23348 22840 23400 22892
rect 23532 22840 23584 22892
rect 19484 22704 19536 22756
rect 20404 22704 20456 22756
rect 21048 22772 21100 22824
rect 23440 22772 23492 22824
rect 23716 22772 23768 22824
rect 21508 22704 21560 22756
rect 23164 22704 23216 22756
rect 23900 22747 23952 22756
rect 23900 22713 23909 22747
rect 23909 22713 23943 22747
rect 23943 22713 23952 22747
rect 23900 22704 23952 22713
rect 25096 22840 25148 22892
rect 25004 22704 25056 22756
rect 20220 22636 20272 22688
rect 21048 22679 21100 22688
rect 21048 22645 21057 22679
rect 21057 22645 21091 22679
rect 21091 22645 21100 22679
rect 21048 22636 21100 22645
rect 22520 22636 22572 22688
rect 23256 22636 23308 22688
rect 23808 22636 23860 22688
rect 16448 22500 16500 22552
rect 21232 22568 21284 22620
rect 24544 22636 24596 22688
rect 24912 22636 24964 22688
rect 25372 22679 25424 22688
rect 25372 22645 25381 22679
rect 25381 22645 25415 22679
rect 25415 22645 25424 22679
rect 25372 22636 25424 22645
rect 26200 22704 26252 22756
rect 27028 22704 27080 22756
rect 28592 22636 28644 22688
rect 28960 22636 29012 22688
rect 27396 22568 27448 22620
rect 28224 22568 28276 22620
rect 22336 22500 22388 22552
rect 23256 22500 23308 22552
rect 19142 22398 19194 22450
rect 19206 22398 19258 22450
rect 19270 22398 19322 22450
rect 19334 22398 19386 22450
rect 29142 22398 29194 22450
rect 29206 22398 29258 22450
rect 29270 22398 29322 22450
rect 29334 22398 29386 22450
rect 20680 22296 20732 22348
rect 21968 22296 22020 22348
rect 22612 22296 22664 22348
rect 13964 22271 14016 22280
rect 13964 22237 13973 22271
rect 13973 22237 14007 22271
rect 14007 22237 14016 22271
rect 13964 22228 14016 22237
rect 15068 22228 15120 22280
rect 11940 22160 11992 22212
rect 14792 22203 14844 22212
rect 14792 22169 14801 22203
rect 14801 22169 14835 22203
rect 14835 22169 14844 22203
rect 14792 22160 14844 22169
rect 15252 22160 15304 22212
rect 16264 22160 16316 22212
rect 17000 22228 17052 22280
rect 18104 22203 18156 22212
rect 18104 22169 18113 22203
rect 18113 22169 18147 22203
rect 18147 22169 18156 22203
rect 18104 22160 18156 22169
rect 18380 22203 18432 22212
rect 18380 22169 18389 22203
rect 18389 22169 18423 22203
rect 18423 22169 18432 22203
rect 18380 22160 18432 22169
rect 20220 22228 20272 22280
rect 21416 22228 21468 22280
rect 23900 22228 23952 22280
rect 19760 22160 19812 22212
rect 20496 22203 20548 22212
rect 20496 22169 20505 22203
rect 20505 22169 20539 22203
rect 20539 22169 20548 22203
rect 20496 22160 20548 22169
rect 21692 22160 21744 22212
rect 22980 22203 23032 22212
rect 22980 22169 22986 22203
rect 22986 22169 23032 22203
rect 22980 22160 23032 22169
rect 23256 22160 23308 22212
rect 28592 22228 28644 22280
rect 25096 22160 25148 22212
rect 26200 22160 26252 22212
rect 26384 22160 26436 22212
rect 29880 22160 29932 22212
rect 12032 21999 12084 22008
rect 12032 21965 12041 21999
rect 12041 21965 12075 21999
rect 12075 21965 12084 21999
rect 12032 21956 12084 21965
rect 17184 22092 17236 22144
rect 20404 22092 20456 22144
rect 20588 22092 20640 22144
rect 21876 22092 21928 22144
rect 21968 22135 22020 22144
rect 21968 22101 21977 22135
rect 21977 22101 22011 22135
rect 22011 22101 22020 22135
rect 23164 22135 23216 22144
rect 21968 22092 22020 22101
rect 23164 22101 23173 22135
rect 23173 22101 23207 22135
rect 23207 22101 23216 22135
rect 23164 22092 23216 22101
rect 29328 22135 29380 22144
rect 29328 22101 29337 22135
rect 29337 22101 29371 22135
rect 29371 22101 29380 22135
rect 29328 22092 29380 22101
rect 15804 21956 15856 22008
rect 16816 21956 16868 22008
rect 21232 21956 21284 22008
rect 21968 21956 22020 22008
rect 22336 21956 22388 22008
rect 23624 22024 23676 22076
rect 27396 22067 27448 22076
rect 27396 22033 27405 22067
rect 27405 22033 27439 22067
rect 27439 22033 27448 22067
rect 27396 22024 27448 22033
rect 25280 21999 25332 22008
rect 25280 21965 25289 21999
rect 25289 21965 25323 21999
rect 25323 21965 25332 21999
rect 25280 21956 25332 21965
rect 14142 21854 14194 21906
rect 14206 21854 14258 21906
rect 14270 21854 14322 21906
rect 14334 21854 14386 21906
rect 24142 21854 24194 21906
rect 24206 21854 24258 21906
rect 24270 21854 24322 21906
rect 24334 21854 24386 21906
rect 17000 21795 17052 21804
rect 17000 21761 17009 21795
rect 17009 21761 17043 21795
rect 17043 21761 17052 21795
rect 17000 21752 17052 21761
rect 18012 21795 18064 21804
rect 18012 21761 18021 21795
rect 18021 21761 18055 21795
rect 18055 21761 18064 21795
rect 18012 21752 18064 21761
rect 19576 21752 19628 21804
rect 21692 21795 21744 21804
rect 13044 21616 13096 21668
rect 14516 21684 14568 21736
rect 12216 21548 12268 21600
rect 11848 21523 11900 21532
rect 11848 21489 11857 21523
rect 11857 21489 11891 21523
rect 11891 21489 11900 21523
rect 11848 21480 11900 21489
rect 12676 21591 12728 21600
rect 12676 21557 12685 21591
rect 12685 21557 12719 21591
rect 12719 21557 12728 21591
rect 13136 21591 13188 21600
rect 12676 21548 12728 21557
rect 13136 21557 13145 21591
rect 13145 21557 13179 21591
rect 13179 21557 13188 21591
rect 13136 21548 13188 21557
rect 14516 21591 14568 21600
rect 14516 21557 14525 21591
rect 14525 21557 14559 21591
rect 14559 21557 14568 21591
rect 14516 21548 14568 21557
rect 16816 21684 16868 21736
rect 20036 21684 20088 21736
rect 20588 21684 20640 21736
rect 21692 21761 21701 21795
rect 21701 21761 21735 21795
rect 21735 21761 21744 21795
rect 21692 21752 21744 21761
rect 23808 21752 23860 21804
rect 23164 21684 23216 21736
rect 15068 21616 15120 21668
rect 18748 21616 18800 21668
rect 19024 21616 19076 21668
rect 15528 21591 15580 21600
rect 12768 21480 12820 21532
rect 15528 21557 15537 21591
rect 15537 21557 15571 21591
rect 15571 21557 15580 21591
rect 15528 21548 15580 21557
rect 17828 21548 17880 21600
rect 18104 21548 18156 21600
rect 21508 21616 21560 21668
rect 22704 21616 22756 21668
rect 23440 21616 23492 21668
rect 20404 21591 20456 21600
rect 15436 21480 15488 21532
rect 17736 21523 17788 21532
rect 15252 21412 15304 21464
rect 17736 21489 17745 21523
rect 17745 21489 17779 21523
rect 17779 21489 17788 21523
rect 17736 21480 17788 21489
rect 20404 21557 20413 21591
rect 20413 21557 20447 21591
rect 20447 21557 20456 21591
rect 20404 21548 20456 21557
rect 21140 21548 21192 21600
rect 22612 21591 22664 21600
rect 22612 21557 22621 21591
rect 22621 21557 22655 21591
rect 22655 21557 22664 21591
rect 22612 21548 22664 21557
rect 29696 21616 29748 21668
rect 25556 21591 25608 21600
rect 20220 21480 20272 21532
rect 21416 21480 21468 21532
rect 25556 21557 25565 21591
rect 25565 21557 25599 21591
rect 25599 21557 25608 21591
rect 25556 21548 25608 21557
rect 25648 21548 25700 21600
rect 26384 21548 26436 21600
rect 27948 21591 28000 21600
rect 27948 21557 27957 21591
rect 27957 21557 27991 21591
rect 27991 21557 28000 21591
rect 27948 21548 28000 21557
rect 28776 21548 28828 21600
rect 23348 21523 23400 21532
rect 23348 21489 23357 21523
rect 23357 21489 23391 21523
rect 23391 21489 23400 21523
rect 23348 21480 23400 21489
rect 17276 21412 17328 21464
rect 18564 21412 18616 21464
rect 22704 21412 22756 21464
rect 26568 21480 26620 21532
rect 26752 21480 26804 21532
rect 26844 21480 26896 21532
rect 27396 21480 27448 21532
rect 29604 21480 29656 21532
rect 23900 21412 23952 21464
rect 19142 21310 19194 21362
rect 19206 21310 19258 21362
rect 19270 21310 19322 21362
rect 19334 21310 19386 21362
rect 29142 21310 29194 21362
rect 29206 21310 29258 21362
rect 29270 21310 29322 21362
rect 29334 21310 29386 21362
rect 17092 21208 17144 21260
rect 19852 21208 19904 21260
rect 11848 21140 11900 21192
rect 12032 21140 12084 21192
rect 11296 21115 11348 21124
rect 11296 21081 11305 21115
rect 11305 21081 11339 21115
rect 11339 21081 11348 21115
rect 11296 21072 11348 21081
rect 13136 21072 13188 21124
rect 15252 21140 15304 21192
rect 15528 21140 15580 21192
rect 16264 21115 16316 21124
rect 16264 21081 16273 21115
rect 16273 21081 16307 21115
rect 16307 21081 16316 21115
rect 16264 21072 16316 21081
rect 16448 21115 16500 21124
rect 16448 21081 16457 21115
rect 16457 21081 16491 21115
rect 16491 21081 16500 21115
rect 16448 21072 16500 21081
rect 17828 21140 17880 21192
rect 19576 21140 19628 21192
rect 19668 21140 19720 21192
rect 16908 21115 16960 21124
rect 16908 21081 16917 21115
rect 16917 21081 16951 21115
rect 16951 21081 16960 21115
rect 16908 21072 16960 21081
rect 17184 21115 17236 21124
rect 17184 21081 17204 21115
rect 17204 21081 17236 21115
rect 17184 21072 17236 21081
rect 18564 21072 18616 21124
rect 20220 21115 20272 21124
rect 20220 21081 20229 21115
rect 20229 21081 20263 21115
rect 20263 21081 20272 21115
rect 20220 21072 20272 21081
rect 20404 21072 20456 21124
rect 21508 21072 21560 21124
rect 21876 21115 21928 21124
rect 21876 21081 21885 21115
rect 21885 21081 21919 21115
rect 21919 21081 21928 21115
rect 21876 21072 21928 21081
rect 23992 21140 24044 21192
rect 23348 21072 23400 21124
rect 24912 21208 24964 21260
rect 25464 21140 25516 21192
rect 25556 21140 25608 21192
rect 25188 21072 25240 21124
rect 26752 21140 26804 21192
rect 29512 21140 29564 21192
rect 28592 21072 28644 21124
rect 29604 21072 29656 21124
rect 15252 21004 15304 21056
rect 18104 21004 18156 21056
rect 19024 21004 19076 21056
rect 20128 21047 20180 21056
rect 20128 21013 20137 21047
rect 20137 21013 20171 21047
rect 20171 21013 20180 21047
rect 20128 21004 20180 21013
rect 21140 21004 21192 21056
rect 21692 21047 21744 21056
rect 21692 21013 21701 21047
rect 21701 21013 21735 21047
rect 21735 21013 21744 21047
rect 21692 21004 21744 21013
rect 21968 21004 22020 21056
rect 22152 21047 22204 21056
rect 22152 21013 22161 21047
rect 22161 21013 22195 21047
rect 22195 21013 22204 21047
rect 22152 21004 22204 21013
rect 17184 20936 17236 20988
rect 17552 20936 17604 20988
rect 20404 20936 20456 20988
rect 21784 20936 21836 20988
rect 23532 20936 23584 20988
rect 27212 21047 27264 21056
rect 27212 21013 27221 21047
rect 27221 21013 27255 21047
rect 27255 21013 27264 21047
rect 27212 21004 27264 21013
rect 26844 20936 26896 20988
rect 13872 20868 13924 20920
rect 17736 20868 17788 20920
rect 19944 20868 19996 20920
rect 24636 20868 24688 20920
rect 14142 20766 14194 20818
rect 14206 20766 14258 20818
rect 14270 20766 14322 20818
rect 14334 20766 14386 20818
rect 24142 20766 24194 20818
rect 24206 20766 24258 20818
rect 24270 20766 24322 20818
rect 24334 20766 24386 20818
rect 15436 20707 15488 20716
rect 15436 20673 15445 20707
rect 15445 20673 15479 20707
rect 15479 20673 15488 20707
rect 15436 20664 15488 20673
rect 20128 20664 20180 20716
rect 21876 20664 21928 20716
rect 22704 20664 22756 20716
rect 27212 20664 27264 20716
rect 12216 20571 12268 20580
rect 12216 20537 12225 20571
rect 12225 20537 12259 20571
rect 12259 20537 12268 20571
rect 12216 20528 12268 20537
rect 13136 20571 13188 20580
rect 13136 20537 13145 20571
rect 13145 20537 13179 20571
rect 13179 20537 13188 20571
rect 13136 20528 13188 20537
rect 12952 20460 13004 20512
rect 14516 20596 14568 20648
rect 15712 20596 15764 20648
rect 19668 20596 19720 20648
rect 20404 20596 20456 20648
rect 23440 20596 23492 20648
rect 25556 20596 25608 20648
rect 15068 20528 15120 20580
rect 13688 20503 13740 20512
rect 13688 20469 13697 20503
rect 13697 20469 13731 20503
rect 13731 20469 13740 20503
rect 13688 20460 13740 20469
rect 13872 20503 13924 20512
rect 13872 20469 13881 20503
rect 13881 20469 13915 20503
rect 13915 20469 13924 20503
rect 13872 20460 13924 20469
rect 14608 20460 14660 20512
rect 18012 20528 18064 20580
rect 20588 20528 20640 20580
rect 21600 20528 21652 20580
rect 18104 20503 18156 20512
rect 18104 20469 18113 20503
rect 18113 20469 18147 20503
rect 18147 20469 18156 20503
rect 18104 20460 18156 20469
rect 19944 20503 19996 20512
rect 14424 20392 14476 20444
rect 14884 20435 14936 20444
rect 14884 20401 14893 20435
rect 14893 20401 14927 20435
rect 14927 20401 14936 20435
rect 14884 20392 14936 20401
rect 18932 20435 18984 20444
rect 18932 20401 18941 20435
rect 18941 20401 18975 20435
rect 18975 20401 18984 20435
rect 18932 20392 18984 20401
rect 19944 20469 19953 20503
rect 19953 20469 19987 20503
rect 19987 20469 19996 20503
rect 19944 20460 19996 20469
rect 20220 20460 20272 20512
rect 21508 20460 21560 20512
rect 21784 20460 21836 20512
rect 22336 20503 22388 20512
rect 22336 20469 22345 20503
rect 22345 20469 22379 20503
rect 22379 20469 22388 20503
rect 25648 20528 25700 20580
rect 26844 20571 26896 20580
rect 26844 20537 26853 20571
rect 26853 20537 26887 20571
rect 26887 20537 26896 20571
rect 26844 20528 26896 20537
rect 22336 20460 22388 20469
rect 24636 20503 24688 20512
rect 24636 20469 24645 20503
rect 24645 20469 24679 20503
rect 24679 20469 24688 20503
rect 24636 20460 24688 20469
rect 25188 20460 25240 20512
rect 26476 20503 26528 20512
rect 26476 20469 26485 20503
rect 26485 20469 26519 20503
rect 26519 20469 26528 20503
rect 26476 20460 26528 20469
rect 27948 20503 28000 20512
rect 27948 20469 27957 20503
rect 27957 20469 27991 20503
rect 27991 20469 28000 20503
rect 27948 20460 28000 20469
rect 19668 20392 19720 20444
rect 24544 20392 24596 20444
rect 28776 20392 28828 20444
rect 29604 20392 29656 20444
rect 12676 20324 12728 20376
rect 19760 20324 19812 20376
rect 20220 20324 20272 20376
rect 19142 20222 19194 20274
rect 19206 20222 19258 20274
rect 19270 20222 19322 20274
rect 19334 20222 19386 20274
rect 29142 20222 29194 20274
rect 29206 20222 29258 20274
rect 29270 20222 29322 20274
rect 29334 20222 29386 20274
rect 16448 20120 16500 20172
rect 18196 20120 18248 20172
rect 15804 20095 15856 20104
rect 15804 20061 15813 20095
rect 15813 20061 15847 20095
rect 15847 20061 15856 20095
rect 15804 20052 15856 20061
rect 17000 20095 17052 20104
rect 17000 20061 17009 20095
rect 17009 20061 17043 20095
rect 17043 20061 17052 20095
rect 17552 20095 17604 20104
rect 17000 20052 17052 20061
rect 11664 20027 11716 20036
rect 11664 19993 11673 20027
rect 11673 19993 11707 20027
rect 11707 19993 11716 20027
rect 11664 19984 11716 19993
rect 12676 20027 12728 20036
rect 12676 19993 12685 20027
rect 12685 19993 12719 20027
rect 12719 19993 12728 20027
rect 12952 20027 13004 20036
rect 12676 19984 12728 19993
rect 12952 19993 12961 20027
rect 12961 19993 12995 20027
rect 12995 19993 13004 20027
rect 12952 19984 13004 19993
rect 14424 19984 14476 20036
rect 14608 20027 14660 20036
rect 14608 19993 14617 20027
rect 14617 19993 14651 20027
rect 14651 19993 14660 20027
rect 14608 19984 14660 19993
rect 17184 20027 17236 20036
rect 17184 19993 17193 20027
rect 17193 19993 17227 20027
rect 17227 19993 17236 20027
rect 17184 19984 17236 19993
rect 17552 20061 17561 20095
rect 17561 20061 17595 20095
rect 17595 20061 17604 20095
rect 17552 20052 17604 20061
rect 17828 20052 17880 20104
rect 18932 20095 18984 20104
rect 18932 20061 18941 20095
rect 18941 20061 18975 20095
rect 18975 20061 18984 20095
rect 18932 20052 18984 20061
rect 19208 20052 19260 20104
rect 19852 20120 19904 20172
rect 19760 20095 19812 20104
rect 19760 20061 19769 20095
rect 19769 20061 19803 20095
rect 19803 20061 19812 20095
rect 19760 20052 19812 20061
rect 19944 20095 19996 20104
rect 19944 20061 19953 20095
rect 19953 20061 19987 20095
rect 19987 20061 19996 20095
rect 19944 20052 19996 20061
rect 21508 20052 21560 20104
rect 26476 20052 26528 20104
rect 17736 19984 17788 20036
rect 12768 19959 12820 19968
rect 12768 19925 12777 19959
rect 12777 19925 12811 19959
rect 12811 19925 12820 19959
rect 12768 19916 12820 19925
rect 14700 19916 14752 19968
rect 18012 19916 18064 19968
rect 21048 19984 21100 20036
rect 22152 20027 22204 20036
rect 22152 19993 22161 20027
rect 22161 19993 22195 20027
rect 22195 19993 22204 20027
rect 22152 19984 22204 19993
rect 22244 20027 22296 20036
rect 22244 19993 22253 20027
rect 22253 19993 22287 20027
rect 22287 19993 22296 20027
rect 22244 19984 22296 19993
rect 23532 20027 23584 20036
rect 15712 19848 15764 19900
rect 15896 19848 15948 19900
rect 16264 19848 16316 19900
rect 20220 19916 20272 19968
rect 20404 19916 20456 19968
rect 21692 19959 21744 19968
rect 21692 19925 21701 19959
rect 21701 19925 21735 19959
rect 21735 19925 21744 19959
rect 21692 19916 21744 19925
rect 23532 19993 23541 20027
rect 23541 19993 23575 20027
rect 23575 19993 23584 20027
rect 23532 19984 23584 19993
rect 23992 20027 24044 20036
rect 23992 19993 24001 20027
rect 24001 19993 24035 20027
rect 24035 19993 24044 20027
rect 23992 19984 24044 19993
rect 24636 19984 24688 20036
rect 25556 19984 25608 20036
rect 27948 20120 28000 20172
rect 29512 20052 29564 20104
rect 26016 19916 26068 19968
rect 27304 19984 27356 20036
rect 28592 20027 28644 20036
rect 28592 19993 28601 20027
rect 28601 19993 28635 20027
rect 28635 19993 28644 20027
rect 28592 19984 28644 19993
rect 28868 19916 28920 19968
rect 18932 19848 18984 19900
rect 24912 19848 24964 19900
rect 26200 19848 26252 19900
rect 16080 19823 16132 19832
rect 16080 19789 16089 19823
rect 16089 19789 16123 19823
rect 16123 19789 16132 19823
rect 16080 19780 16132 19789
rect 16724 19780 16776 19832
rect 27764 19823 27816 19832
rect 27764 19789 27773 19823
rect 27773 19789 27807 19823
rect 27807 19789 27816 19823
rect 27764 19780 27816 19789
rect 14142 19678 14194 19730
rect 14206 19678 14258 19730
rect 14270 19678 14322 19730
rect 14334 19678 14386 19730
rect 24142 19678 24194 19730
rect 24206 19678 24258 19730
rect 24270 19678 24322 19730
rect 24334 19678 24386 19730
rect 12768 19440 12820 19492
rect 13872 19440 13924 19492
rect 14608 19440 14660 19492
rect 15252 19440 15304 19492
rect 17184 19508 17236 19560
rect 19944 19508 19996 19560
rect 24268 19551 24320 19560
rect 24268 19517 24277 19551
rect 24277 19517 24311 19551
rect 24311 19517 24320 19551
rect 24268 19508 24320 19517
rect 17828 19483 17880 19492
rect 17828 19449 17837 19483
rect 17837 19449 17871 19483
rect 17871 19449 17880 19483
rect 17828 19440 17880 19449
rect 18932 19483 18984 19492
rect 18932 19449 18941 19483
rect 18941 19449 18975 19483
rect 18975 19449 18984 19483
rect 18932 19440 18984 19449
rect 19668 19483 19720 19492
rect 19668 19449 19677 19483
rect 19677 19449 19711 19483
rect 19711 19449 19720 19483
rect 19668 19440 19720 19449
rect 23992 19440 24044 19492
rect 13688 19372 13740 19424
rect 13964 19372 14016 19424
rect 14516 19304 14568 19356
rect 15068 19236 15120 19288
rect 15344 19236 15396 19288
rect 16080 19372 16132 19424
rect 16724 19415 16776 19424
rect 16724 19381 16733 19415
rect 16733 19381 16767 19415
rect 16767 19381 16776 19415
rect 16724 19372 16776 19381
rect 17184 19372 17236 19424
rect 19208 19415 19260 19424
rect 19208 19381 19217 19415
rect 19217 19381 19251 19415
rect 19251 19381 19260 19415
rect 19208 19372 19260 19381
rect 19484 19372 19536 19424
rect 20220 19372 20272 19424
rect 22980 19415 23032 19424
rect 22980 19381 22989 19415
rect 22989 19381 23023 19415
rect 23023 19381 23032 19415
rect 22980 19372 23032 19381
rect 23072 19372 23124 19424
rect 25280 19508 25332 19560
rect 25464 19508 25516 19560
rect 26476 19576 26528 19628
rect 27304 19576 27356 19628
rect 24636 19440 24688 19492
rect 26660 19508 26712 19560
rect 28592 19508 28644 19560
rect 25464 19415 25516 19424
rect 25464 19381 25473 19415
rect 25473 19381 25507 19415
rect 25507 19381 25516 19415
rect 25464 19372 25516 19381
rect 26200 19415 26252 19424
rect 19760 19304 19812 19356
rect 25556 19304 25608 19356
rect 16816 19279 16868 19288
rect 16816 19245 16825 19279
rect 16825 19245 16859 19279
rect 16859 19245 16868 19279
rect 16816 19236 16868 19245
rect 19024 19236 19076 19288
rect 20312 19236 20364 19288
rect 26200 19381 26209 19415
rect 26209 19381 26243 19415
rect 26243 19381 26252 19415
rect 26200 19372 26252 19381
rect 29880 19440 29932 19492
rect 27028 19347 27080 19356
rect 27028 19313 27037 19347
rect 27037 19313 27071 19347
rect 27071 19313 27080 19347
rect 27028 19304 27080 19313
rect 29512 19372 29564 19424
rect 29972 19304 30024 19356
rect 19142 19134 19194 19186
rect 19206 19134 19258 19186
rect 19270 19134 19322 19186
rect 19334 19134 19386 19186
rect 29142 19134 29194 19186
rect 29206 19134 29258 19186
rect 29270 19134 29322 19186
rect 29334 19134 29386 19186
rect 13872 19032 13924 19084
rect 20312 19075 20364 19084
rect 20312 19041 20321 19075
rect 20321 19041 20355 19075
rect 20355 19041 20364 19075
rect 20312 19032 20364 19041
rect 22152 19032 22204 19084
rect 12860 18964 12912 19016
rect 17460 18964 17512 19016
rect 19760 18964 19812 19016
rect 22796 19032 22848 19084
rect 27028 19032 27080 19084
rect 29696 19032 29748 19084
rect 23072 18964 23124 19016
rect 23992 18964 24044 19016
rect 24268 18964 24320 19016
rect 26016 19007 26068 19016
rect 26016 18973 26025 19007
rect 26025 18973 26059 19007
rect 26059 18973 26068 19007
rect 26016 18964 26068 18973
rect 27764 18964 27816 19016
rect 12952 18939 13004 18948
rect 12952 18905 12961 18939
rect 12961 18905 12995 18939
rect 12995 18905 13004 18939
rect 12952 18896 13004 18905
rect 14700 18939 14752 18948
rect 14700 18905 14709 18939
rect 14709 18905 14743 18939
rect 14743 18905 14752 18939
rect 14700 18896 14752 18905
rect 14884 18939 14936 18948
rect 14884 18905 14893 18939
rect 14893 18905 14927 18939
rect 14927 18905 14936 18939
rect 14884 18896 14936 18905
rect 15068 18939 15120 18948
rect 15068 18905 15077 18939
rect 15077 18905 15111 18939
rect 15111 18905 15120 18939
rect 15068 18896 15120 18905
rect 15252 18896 15304 18948
rect 20956 18896 21008 18948
rect 21968 18939 22020 18948
rect 21968 18905 21977 18939
rect 21977 18905 22011 18939
rect 22011 18905 22020 18939
rect 21968 18896 22020 18905
rect 22980 18896 23032 18948
rect 25556 18939 25608 18948
rect 25556 18905 25565 18939
rect 25565 18905 25599 18939
rect 25599 18905 25608 18939
rect 25556 18896 25608 18905
rect 27948 18939 28000 18948
rect 27948 18905 27957 18939
rect 27957 18905 27991 18939
rect 27991 18905 28000 18939
rect 27948 18896 28000 18905
rect 29604 18896 29656 18948
rect 13320 18828 13372 18880
rect 13044 18760 13096 18812
rect 16448 18828 16500 18880
rect 19484 18828 19536 18880
rect 20220 18828 20272 18880
rect 26568 18871 26620 18880
rect 26568 18837 26577 18871
rect 26577 18837 26611 18871
rect 26611 18837 26620 18871
rect 26568 18828 26620 18837
rect 26936 18803 26988 18812
rect 26936 18769 26945 18803
rect 26945 18769 26979 18803
rect 26979 18769 26988 18803
rect 26936 18760 26988 18769
rect 27856 18760 27908 18812
rect 16908 18692 16960 18744
rect 18564 18692 18616 18744
rect 19024 18692 19076 18744
rect 14142 18590 14194 18642
rect 14206 18590 14258 18642
rect 14270 18590 14322 18642
rect 14334 18590 14386 18642
rect 24142 18590 24194 18642
rect 24206 18590 24258 18642
rect 24270 18590 24322 18642
rect 24334 18590 24386 18642
rect 27948 18531 28000 18540
rect 27948 18497 27957 18531
rect 27957 18497 27991 18531
rect 27991 18497 28000 18531
rect 27948 18488 28000 18497
rect 29696 18488 29748 18540
rect 29972 18488 30024 18540
rect 12584 18420 12636 18472
rect 15068 18420 15120 18472
rect 15896 18463 15948 18472
rect 13320 18395 13372 18404
rect 13320 18361 13329 18395
rect 13329 18361 13363 18395
rect 13363 18361 13372 18395
rect 13320 18352 13372 18361
rect 12860 18327 12912 18336
rect 12860 18293 12869 18327
rect 12869 18293 12903 18327
rect 12903 18293 12912 18327
rect 12860 18284 12912 18293
rect 13872 18284 13924 18336
rect 14608 18284 14660 18336
rect 15896 18429 15905 18463
rect 15905 18429 15939 18463
rect 15939 18429 15948 18463
rect 15896 18420 15948 18429
rect 17460 18463 17512 18472
rect 17460 18429 17469 18463
rect 17469 18429 17503 18463
rect 17503 18429 17512 18463
rect 17460 18420 17512 18429
rect 21968 18420 22020 18472
rect 22244 18420 22296 18472
rect 22796 18463 22848 18472
rect 18564 18352 18616 18404
rect 17000 18284 17052 18336
rect 17920 18284 17972 18336
rect 18656 18327 18708 18336
rect 18656 18293 18665 18327
rect 18665 18293 18699 18327
rect 18699 18293 18708 18327
rect 18656 18284 18708 18293
rect 18840 18284 18892 18336
rect 19484 18284 19536 18336
rect 22796 18429 22805 18463
rect 22805 18429 22839 18463
rect 22839 18429 22848 18463
rect 22796 18420 22848 18429
rect 28868 18463 28920 18472
rect 28868 18429 28877 18463
rect 28877 18429 28911 18463
rect 28911 18429 28920 18463
rect 28868 18420 28920 18429
rect 26936 18352 26988 18404
rect 27028 18352 27080 18404
rect 27764 18352 27816 18404
rect 15436 18259 15488 18268
rect 12492 18148 12544 18200
rect 13964 18148 14016 18200
rect 14516 18148 14568 18200
rect 15436 18225 15445 18259
rect 15445 18225 15479 18259
rect 15479 18225 15488 18259
rect 15436 18216 15488 18225
rect 15344 18148 15396 18200
rect 20128 18259 20180 18268
rect 20128 18225 20137 18259
rect 20137 18225 20171 18259
rect 20171 18225 20180 18259
rect 20128 18216 20180 18225
rect 21140 18216 21192 18268
rect 20772 18148 20824 18200
rect 23072 18216 23124 18268
rect 23992 18284 24044 18336
rect 25004 18327 25056 18336
rect 25004 18293 25013 18327
rect 25013 18293 25047 18327
rect 25047 18293 25056 18327
rect 25004 18284 25056 18293
rect 26568 18284 26620 18336
rect 28776 18327 28828 18336
rect 26384 18216 26436 18268
rect 26660 18259 26712 18268
rect 26660 18225 26669 18259
rect 26669 18225 26703 18259
rect 26703 18225 26712 18259
rect 26660 18216 26712 18225
rect 28776 18293 28785 18327
rect 28785 18293 28819 18327
rect 28819 18293 28828 18327
rect 28776 18284 28828 18293
rect 24820 18191 24872 18200
rect 24820 18157 24829 18191
rect 24829 18157 24863 18191
rect 24863 18157 24872 18191
rect 24820 18148 24872 18157
rect 26200 18148 26252 18200
rect 29880 18216 29932 18268
rect 19142 18046 19194 18098
rect 19206 18046 19258 18098
rect 19270 18046 19322 18098
rect 19334 18046 19386 18098
rect 29142 18046 29194 18098
rect 29206 18046 29258 18098
rect 29270 18046 29322 18098
rect 29334 18046 29386 18098
rect 16540 17944 16592 17996
rect 13964 17919 14016 17928
rect 13964 17885 13973 17919
rect 13973 17885 14007 17919
rect 14007 17885 14016 17919
rect 13964 17876 14016 17885
rect 15436 17876 15488 17928
rect 16816 17944 16868 17996
rect 16908 17987 16960 17996
rect 16908 17953 16917 17987
rect 16917 17953 16951 17987
rect 16951 17953 16960 17987
rect 16908 17944 16960 17953
rect 18840 17944 18892 17996
rect 20496 17944 20548 17996
rect 23348 17944 23400 17996
rect 12584 17851 12636 17860
rect 11664 17783 11716 17792
rect 11664 17749 11673 17783
rect 11673 17749 11707 17783
rect 11707 17749 11716 17783
rect 11664 17740 11716 17749
rect 12584 17817 12593 17851
rect 12593 17817 12627 17851
rect 12627 17817 12636 17851
rect 12584 17808 12636 17817
rect 12860 17851 12912 17860
rect 12860 17817 12869 17851
rect 12869 17817 12903 17851
rect 12903 17817 12912 17851
rect 12860 17808 12912 17817
rect 13044 17851 13096 17860
rect 13044 17817 13053 17851
rect 13053 17817 13087 17851
rect 13087 17817 13096 17851
rect 13044 17808 13096 17817
rect 12952 17740 13004 17792
rect 12768 17672 12820 17724
rect 15344 17808 15396 17860
rect 17920 17876 17972 17928
rect 25004 17876 25056 17928
rect 16816 17851 16868 17860
rect 16816 17817 16825 17851
rect 16825 17817 16859 17851
rect 16859 17817 16868 17851
rect 16816 17808 16868 17817
rect 19944 17851 19996 17860
rect 19944 17817 19953 17851
rect 19953 17817 19987 17851
rect 19987 17817 19996 17851
rect 19944 17808 19996 17817
rect 20772 17808 20824 17860
rect 21140 17851 21192 17860
rect 21140 17817 21149 17851
rect 21149 17817 21183 17851
rect 21183 17817 21192 17851
rect 21140 17808 21192 17817
rect 22336 17808 22388 17860
rect 23440 17851 23492 17860
rect 23440 17817 23449 17851
rect 23449 17817 23483 17851
rect 23483 17817 23492 17851
rect 23440 17808 23492 17817
rect 23992 17808 24044 17860
rect 14976 17672 15028 17724
rect 13320 17604 13372 17656
rect 16724 17740 16776 17792
rect 26568 17876 26620 17928
rect 26660 17808 26712 17860
rect 29604 17876 29656 17928
rect 28500 17851 28552 17860
rect 25740 17783 25792 17792
rect 23716 17672 23768 17724
rect 25740 17749 25749 17783
rect 25749 17749 25783 17783
rect 25783 17749 25792 17783
rect 25740 17740 25792 17749
rect 28500 17817 28509 17851
rect 28509 17817 28543 17851
rect 28543 17817 28552 17851
rect 28500 17808 28552 17817
rect 28592 17808 28644 17860
rect 25556 17672 25608 17724
rect 27764 17715 27816 17724
rect 27764 17681 27773 17715
rect 27773 17681 27807 17715
rect 27807 17681 27816 17715
rect 27764 17672 27816 17681
rect 20680 17604 20732 17656
rect 14142 17502 14194 17554
rect 14206 17502 14258 17554
rect 14270 17502 14322 17554
rect 14334 17502 14386 17554
rect 24142 17502 24194 17554
rect 24206 17502 24258 17554
rect 24270 17502 24322 17554
rect 24334 17502 24386 17554
rect 13320 17400 13372 17452
rect 27120 17400 27172 17452
rect 12952 17264 13004 17316
rect 14608 17307 14660 17316
rect 14608 17273 14617 17307
rect 14617 17273 14651 17307
rect 14651 17273 14660 17307
rect 14608 17264 14660 17273
rect 14976 17307 15028 17316
rect 14976 17273 14985 17307
rect 14985 17273 15019 17307
rect 15019 17273 15028 17307
rect 14976 17264 15028 17273
rect 15068 17264 15120 17316
rect 15436 17307 15488 17316
rect 12492 17239 12544 17248
rect 12492 17205 12501 17239
rect 12501 17205 12535 17239
rect 12535 17205 12544 17239
rect 12492 17196 12544 17205
rect 12768 17239 12820 17248
rect 12768 17205 12777 17239
rect 12777 17205 12811 17239
rect 12811 17205 12820 17239
rect 12768 17196 12820 17205
rect 12860 17196 12912 17248
rect 13320 17196 13372 17248
rect 15436 17273 15445 17307
rect 15445 17273 15479 17307
rect 15479 17273 15488 17307
rect 15436 17264 15488 17273
rect 23900 17332 23952 17384
rect 25556 17375 25608 17384
rect 25556 17341 25565 17375
rect 25565 17341 25599 17375
rect 25599 17341 25608 17375
rect 25556 17332 25608 17341
rect 23532 17264 23584 17316
rect 25372 17264 25424 17316
rect 28500 17307 28552 17316
rect 28500 17273 28509 17307
rect 28509 17273 28543 17307
rect 28543 17273 28552 17307
rect 28500 17264 28552 17273
rect 28960 17264 29012 17316
rect 16724 17239 16776 17248
rect 16724 17205 16733 17239
rect 16733 17205 16767 17239
rect 16767 17205 16776 17239
rect 16724 17196 16776 17205
rect 17000 17239 17052 17248
rect 17000 17205 17009 17239
rect 17009 17205 17043 17239
rect 17043 17205 17052 17239
rect 17000 17196 17052 17205
rect 17920 17239 17972 17248
rect 17920 17205 17929 17239
rect 17929 17205 17963 17239
rect 17963 17205 17972 17239
rect 17920 17196 17972 17205
rect 16816 17128 16868 17180
rect 18104 17103 18156 17112
rect 18104 17069 18113 17103
rect 18113 17069 18147 17103
rect 18147 17069 18156 17103
rect 18104 17060 18156 17069
rect 20680 17196 20732 17248
rect 23348 17239 23400 17248
rect 23348 17205 23357 17239
rect 23357 17205 23391 17239
rect 23391 17205 23400 17239
rect 23348 17196 23400 17205
rect 19576 17171 19628 17180
rect 19576 17137 19585 17171
rect 19585 17137 19619 17171
rect 19619 17137 19628 17171
rect 19576 17128 19628 17137
rect 21324 17171 21376 17180
rect 21324 17137 21333 17171
rect 21333 17137 21367 17171
rect 21367 17137 21376 17171
rect 21324 17128 21376 17137
rect 23716 17196 23768 17248
rect 25004 17239 25056 17248
rect 25004 17205 25013 17239
rect 25013 17205 25047 17239
rect 25047 17205 25056 17239
rect 25004 17196 25056 17205
rect 19484 17060 19536 17112
rect 26476 17128 26528 17180
rect 27212 17196 27264 17248
rect 28316 17196 28368 17248
rect 29880 17196 29932 17248
rect 23440 17060 23492 17112
rect 19142 16958 19194 17010
rect 19206 16958 19258 17010
rect 19270 16958 19322 17010
rect 19334 16958 19386 17010
rect 29142 16958 29194 17010
rect 29206 16958 29258 17010
rect 29270 16958 29322 17010
rect 29334 16958 29386 17010
rect 11664 16788 11716 16840
rect 12124 16788 12176 16840
rect 13320 16831 13372 16840
rect 13320 16797 13329 16831
rect 13329 16797 13363 16831
rect 13363 16797 13372 16831
rect 13320 16788 13372 16797
rect 11296 16763 11348 16772
rect 11296 16729 11305 16763
rect 11305 16729 11339 16763
rect 11339 16729 11348 16763
rect 11296 16720 11348 16729
rect 12952 16720 13004 16772
rect 16448 16856 16500 16908
rect 14516 16788 14568 16840
rect 14700 16788 14752 16840
rect 17644 16856 17696 16908
rect 19484 16856 19536 16908
rect 19576 16856 19628 16908
rect 25740 16856 25792 16908
rect 24820 16788 24872 16840
rect 27764 16788 27816 16840
rect 18104 16720 18156 16772
rect 19576 16720 19628 16772
rect 20772 16720 20824 16772
rect 22520 16720 22572 16772
rect 23440 16720 23492 16772
rect 14976 16652 15028 16704
rect 18012 16652 18064 16704
rect 17184 16516 17236 16568
rect 19484 16652 19536 16704
rect 20864 16695 20916 16704
rect 20864 16661 20873 16695
rect 20873 16661 20907 16695
rect 20907 16661 20916 16695
rect 20864 16652 20916 16661
rect 21140 16695 21192 16704
rect 21140 16661 21149 16695
rect 21149 16661 21183 16695
rect 21183 16661 21192 16695
rect 21140 16652 21192 16661
rect 22244 16584 22296 16636
rect 22336 16584 22388 16636
rect 25832 16720 25884 16772
rect 23992 16695 24044 16704
rect 23992 16661 24001 16695
rect 24001 16661 24035 16695
rect 24035 16661 24044 16695
rect 26476 16720 26528 16772
rect 28500 16720 28552 16772
rect 23992 16652 24044 16661
rect 28776 16652 28828 16704
rect 28868 16652 28920 16704
rect 29604 16584 29656 16636
rect 25372 16559 25424 16568
rect 25372 16525 25381 16559
rect 25381 16525 25415 16559
rect 25415 16525 25424 16559
rect 25372 16516 25424 16525
rect 14142 16414 14194 16466
rect 14206 16414 14258 16466
rect 14270 16414 14322 16466
rect 14334 16414 14386 16466
rect 24142 16414 24194 16466
rect 24206 16414 24258 16466
rect 24270 16414 24322 16466
rect 24334 16414 24386 16466
rect 12124 16355 12176 16364
rect 12124 16321 12133 16355
rect 12133 16321 12167 16355
rect 12167 16321 12176 16355
rect 12124 16312 12176 16321
rect 14700 16312 14752 16364
rect 15436 16312 15488 16364
rect 17000 16312 17052 16364
rect 17920 16312 17972 16364
rect 19576 16355 19628 16364
rect 19576 16321 19585 16355
rect 19585 16321 19619 16355
rect 19619 16321 19628 16355
rect 19576 16312 19628 16321
rect 22520 16355 22572 16364
rect 22520 16321 22529 16355
rect 22529 16321 22563 16355
rect 22563 16321 22572 16355
rect 22520 16312 22572 16321
rect 27120 16355 27172 16364
rect 27120 16321 27129 16355
rect 27129 16321 27163 16355
rect 27163 16321 27172 16355
rect 27120 16312 27172 16321
rect 18012 16287 18064 16296
rect 18012 16253 18021 16287
rect 18021 16253 18055 16287
rect 18055 16253 18064 16287
rect 18012 16244 18064 16253
rect 20864 16244 20916 16296
rect 11940 16151 11992 16160
rect 11940 16117 11949 16151
rect 11949 16117 11983 16151
rect 11983 16117 11992 16151
rect 11940 16108 11992 16117
rect 13780 16108 13832 16160
rect 21140 16176 21192 16228
rect 14976 16108 15028 16160
rect 14884 16040 14936 16092
rect 17184 16151 17236 16160
rect 17184 16117 17193 16151
rect 17193 16117 17227 16151
rect 17227 16117 17236 16151
rect 17644 16151 17696 16160
rect 17184 16108 17236 16117
rect 17644 16117 17653 16151
rect 17653 16117 17687 16151
rect 17687 16117 17696 16151
rect 17644 16108 17696 16117
rect 18288 16108 18340 16160
rect 18932 16108 18984 16160
rect 19024 16040 19076 16092
rect 20772 16108 20824 16160
rect 21416 16151 21468 16160
rect 21416 16117 21425 16151
rect 21425 16117 21459 16151
rect 21459 16117 21468 16151
rect 21416 16108 21468 16117
rect 22336 16151 22388 16160
rect 22336 16117 22345 16151
rect 22345 16117 22379 16151
rect 22379 16117 22388 16151
rect 23164 16176 23216 16228
rect 22336 16108 22388 16117
rect 25372 16108 25424 16160
rect 25832 16108 25884 16160
rect 27028 16151 27080 16160
rect 27028 16117 27037 16151
rect 27037 16117 27071 16151
rect 27071 16117 27080 16151
rect 27028 16108 27080 16117
rect 27856 16108 27908 16160
rect 28960 16108 29012 16160
rect 23900 16083 23952 16092
rect 23900 16049 23909 16083
rect 23909 16049 23943 16083
rect 23943 16049 23952 16083
rect 23900 16040 23952 16049
rect 25280 15972 25332 16024
rect 26292 16015 26344 16024
rect 26292 15981 26301 16015
rect 26301 15981 26335 16015
rect 26335 15981 26344 16015
rect 26292 15972 26344 15981
rect 27948 15972 28000 16024
rect 28592 15972 28644 16024
rect 28684 15972 28736 16024
rect 19142 15870 19194 15922
rect 19206 15870 19258 15922
rect 19270 15870 19322 15922
rect 19334 15870 19386 15922
rect 29142 15870 29194 15922
rect 29206 15870 29258 15922
rect 29270 15870 29322 15922
rect 29334 15870 29386 15922
rect 23900 15768 23952 15820
rect 11756 15675 11808 15684
rect 11756 15641 11765 15675
rect 11765 15641 11799 15675
rect 11799 15641 11808 15675
rect 11756 15632 11808 15641
rect 13044 15675 13096 15684
rect 13044 15641 13053 15675
rect 13053 15641 13087 15675
rect 13087 15641 13096 15675
rect 13044 15632 13096 15641
rect 11664 15607 11716 15616
rect 11664 15573 11673 15607
rect 11673 15573 11707 15607
rect 11707 15573 11716 15607
rect 11664 15564 11716 15573
rect 12676 15564 12728 15616
rect 14792 15675 14844 15684
rect 14792 15641 14801 15675
rect 14801 15641 14835 15675
rect 14835 15641 14844 15675
rect 15252 15675 15304 15684
rect 14792 15632 14844 15641
rect 15252 15641 15261 15675
rect 15261 15641 15295 15675
rect 15295 15641 15304 15675
rect 15252 15632 15304 15641
rect 16080 15632 16132 15684
rect 17184 15675 17236 15684
rect 17184 15641 17193 15675
rect 17193 15641 17227 15675
rect 17227 15641 17236 15675
rect 17184 15632 17236 15641
rect 18196 15632 18248 15684
rect 18288 15632 18340 15684
rect 18564 15675 18616 15684
rect 18564 15641 18573 15675
rect 18573 15641 18607 15675
rect 18607 15641 18616 15675
rect 18564 15632 18616 15641
rect 22244 15675 22296 15684
rect 18932 15607 18984 15616
rect 14700 15496 14752 15548
rect 18932 15573 18941 15607
rect 18941 15573 18975 15607
rect 18975 15573 18984 15607
rect 18932 15564 18984 15573
rect 22244 15641 22253 15675
rect 22253 15641 22287 15675
rect 22287 15641 22296 15675
rect 22244 15632 22296 15641
rect 22520 15632 22572 15684
rect 23164 15564 23216 15616
rect 15252 15496 15304 15548
rect 17644 15496 17696 15548
rect 19852 15539 19904 15548
rect 19852 15505 19861 15539
rect 19861 15505 19895 15539
rect 19895 15505 19904 15539
rect 19852 15496 19904 15505
rect 21324 15496 21376 15548
rect 22428 15496 22480 15548
rect 12032 15428 12084 15480
rect 13228 15428 13280 15480
rect 17184 15428 17236 15480
rect 20312 15471 20364 15480
rect 20312 15437 20321 15471
rect 20321 15437 20355 15471
rect 20355 15437 20364 15471
rect 20312 15428 20364 15437
rect 20404 15428 20456 15480
rect 23808 15675 23860 15684
rect 23808 15641 23817 15675
rect 23817 15641 23851 15675
rect 23851 15641 23860 15675
rect 23808 15632 23860 15641
rect 25924 15632 25976 15684
rect 26016 15675 26068 15684
rect 26016 15641 26025 15675
rect 26025 15641 26059 15675
rect 26059 15641 26068 15675
rect 26016 15632 26068 15641
rect 27948 15700 28000 15752
rect 28684 15700 28736 15752
rect 26016 15496 26068 15548
rect 29144 15564 29196 15616
rect 25556 15428 25608 15480
rect 27396 15428 27448 15480
rect 27764 15428 27816 15480
rect 27856 15428 27908 15480
rect 14142 15326 14194 15378
rect 14206 15326 14258 15378
rect 14270 15326 14322 15378
rect 14334 15326 14386 15378
rect 24142 15326 24194 15378
rect 24206 15326 24258 15378
rect 24270 15326 24322 15378
rect 24334 15326 24386 15378
rect 13964 15224 14016 15276
rect 18656 15224 18708 15276
rect 19024 15224 19076 15276
rect 21416 15224 21468 15276
rect 22520 15224 22572 15276
rect 29144 15267 29196 15276
rect 29144 15233 29153 15267
rect 29153 15233 29187 15267
rect 29187 15233 29196 15267
rect 29144 15224 29196 15233
rect 11940 15131 11992 15140
rect 11940 15097 11949 15131
rect 11949 15097 11983 15131
rect 11983 15097 11992 15131
rect 11940 15088 11992 15097
rect 12952 15131 13004 15140
rect 12952 15097 12961 15131
rect 12961 15097 12995 15131
rect 12995 15097 13004 15131
rect 12952 15088 13004 15097
rect 13228 15131 13280 15140
rect 13228 15097 13237 15131
rect 13237 15097 13271 15131
rect 13271 15097 13280 15131
rect 13228 15088 13280 15097
rect 14792 15088 14844 15140
rect 11664 15063 11716 15072
rect 11664 15029 11673 15063
rect 11673 15029 11707 15063
rect 11707 15029 11716 15063
rect 11664 15020 11716 15029
rect 11756 15020 11808 15072
rect 16080 15088 16132 15140
rect 18564 15088 18616 15140
rect 22980 15156 23032 15208
rect 17184 15020 17236 15072
rect 17368 15020 17420 15072
rect 18196 15063 18248 15072
rect 18196 15029 18205 15063
rect 18205 15029 18239 15063
rect 18239 15029 18248 15063
rect 18196 15020 18248 15029
rect 14240 14952 14292 15004
rect 14608 14952 14660 15004
rect 19852 15020 19904 15072
rect 20312 15020 20364 15072
rect 20588 15063 20640 15072
rect 20588 15029 20597 15063
rect 20597 15029 20631 15063
rect 20631 15029 20640 15063
rect 22336 15088 22388 15140
rect 23808 15088 23860 15140
rect 25556 15131 25608 15140
rect 25556 15097 25565 15131
rect 25565 15097 25599 15131
rect 25599 15097 25608 15131
rect 25556 15088 25608 15097
rect 25924 15088 25976 15140
rect 20588 15020 20640 15029
rect 15344 14884 15396 14936
rect 15528 14927 15580 14936
rect 15528 14893 15537 14927
rect 15537 14893 15571 14927
rect 15571 14893 15580 14927
rect 15528 14884 15580 14893
rect 18288 14927 18340 14936
rect 18288 14893 18297 14927
rect 18297 14893 18331 14927
rect 18331 14893 18340 14927
rect 18288 14884 18340 14893
rect 18932 14952 18984 15004
rect 22244 15020 22296 15072
rect 22428 15063 22480 15072
rect 22428 15029 22437 15063
rect 22437 15029 22471 15063
rect 22471 15029 22480 15063
rect 22428 15020 22480 15029
rect 22612 15020 22664 15072
rect 23992 15063 24044 15072
rect 23992 15029 24001 15063
rect 24001 15029 24035 15063
rect 24035 15029 24044 15063
rect 25280 15063 25332 15072
rect 23992 15020 24044 15029
rect 25280 15029 25289 15063
rect 25289 15029 25323 15063
rect 25323 15029 25332 15063
rect 25280 15020 25332 15029
rect 27948 15063 28000 15072
rect 27948 15029 27957 15063
rect 27957 15029 27991 15063
rect 27991 15029 28000 15063
rect 27948 15020 28000 15029
rect 28592 15063 28644 15072
rect 23808 14952 23860 15004
rect 19024 14884 19076 14936
rect 26292 14952 26344 15004
rect 27764 14952 27816 15004
rect 28592 15029 28601 15063
rect 28601 15029 28635 15063
rect 28635 15029 28644 15063
rect 28592 15020 28644 15029
rect 26568 14884 26620 14936
rect 19142 14782 19194 14834
rect 19206 14782 19258 14834
rect 19270 14782 19322 14834
rect 19334 14782 19386 14834
rect 29142 14782 29194 14834
rect 29206 14782 29258 14834
rect 29270 14782 29322 14834
rect 29334 14782 29386 14834
rect 14240 14680 14292 14732
rect 15344 14680 15396 14732
rect 18564 14680 18616 14732
rect 11940 14587 11992 14596
rect 11940 14553 11949 14587
rect 11949 14553 11983 14587
rect 11983 14553 11992 14587
rect 11940 14544 11992 14553
rect 12032 14519 12084 14528
rect 12032 14485 12041 14519
rect 12041 14485 12075 14519
rect 12075 14485 12084 14519
rect 12032 14476 12084 14485
rect 11572 14408 11624 14460
rect 12952 14587 13004 14596
rect 12952 14553 12969 14587
rect 12969 14553 13003 14587
rect 13003 14553 13004 14587
rect 12952 14544 13004 14553
rect 13780 14544 13832 14596
rect 15528 14544 15580 14596
rect 15896 14587 15948 14596
rect 15896 14553 15905 14587
rect 15905 14553 15939 14587
rect 15939 14553 15948 14587
rect 15896 14544 15948 14553
rect 16080 14587 16132 14596
rect 16080 14553 16089 14587
rect 16089 14553 16123 14587
rect 16123 14553 16132 14587
rect 16080 14544 16132 14553
rect 16448 14544 16500 14596
rect 17184 14587 17236 14596
rect 17184 14553 17193 14587
rect 17193 14553 17227 14587
rect 17227 14553 17236 14587
rect 17184 14544 17236 14553
rect 19852 14612 19904 14664
rect 23992 14680 24044 14732
rect 25924 14680 25976 14732
rect 27948 14680 28000 14732
rect 12400 14519 12452 14528
rect 12400 14485 12409 14519
rect 12409 14485 12443 14519
rect 12443 14485 12452 14519
rect 12400 14476 12452 14485
rect 14608 14476 14660 14528
rect 20312 14544 20364 14596
rect 22612 14544 22664 14596
rect 27028 14612 27080 14664
rect 22980 14587 23032 14596
rect 22980 14553 22989 14587
rect 22989 14553 23023 14587
rect 23023 14553 23032 14587
rect 22980 14544 23032 14553
rect 23164 14544 23216 14596
rect 25280 14587 25332 14596
rect 25280 14553 25289 14587
rect 25289 14553 25323 14587
rect 25323 14553 25332 14587
rect 25280 14544 25332 14553
rect 12952 14408 13004 14460
rect 16264 14451 16316 14460
rect 16264 14417 16273 14451
rect 16273 14417 16307 14451
rect 16307 14417 16316 14451
rect 20036 14476 20088 14528
rect 22520 14519 22572 14528
rect 22520 14485 22529 14519
rect 22529 14485 22563 14519
rect 22563 14485 22572 14519
rect 22520 14476 22572 14485
rect 23900 14476 23952 14528
rect 16264 14408 16316 14417
rect 20588 14408 20640 14460
rect 25924 14408 25976 14460
rect 27764 14612 27816 14664
rect 29512 14612 29564 14664
rect 12768 14340 12820 14392
rect 18932 14340 18984 14392
rect 22060 14383 22112 14392
rect 22060 14349 22069 14383
rect 22069 14349 22103 14383
rect 22103 14349 22112 14383
rect 22060 14340 22112 14349
rect 25464 14383 25516 14392
rect 25464 14349 25473 14383
rect 25473 14349 25507 14383
rect 25507 14349 25516 14383
rect 25464 14340 25516 14349
rect 26568 14476 26620 14528
rect 27396 14519 27448 14528
rect 27396 14485 27405 14519
rect 27405 14485 27439 14519
rect 27439 14485 27448 14519
rect 27396 14476 27448 14485
rect 28224 14476 28276 14528
rect 27856 14340 27908 14392
rect 14142 14238 14194 14290
rect 14206 14238 14258 14290
rect 14270 14238 14322 14290
rect 14334 14238 14386 14290
rect 24142 14238 24194 14290
rect 24206 14238 24258 14290
rect 24270 14238 24322 14290
rect 24334 14238 24386 14290
rect 13044 14179 13096 14188
rect 13044 14145 13053 14179
rect 13053 14145 13087 14179
rect 13087 14145 13096 14179
rect 13044 14136 13096 14145
rect 13872 14136 13924 14188
rect 16816 14136 16868 14188
rect 17920 14136 17972 14188
rect 22428 14136 22480 14188
rect 28224 14179 28276 14188
rect 28224 14145 28233 14179
rect 28233 14145 28267 14179
rect 28267 14145 28276 14179
rect 28224 14136 28276 14145
rect 28868 14136 28920 14188
rect 11572 13975 11624 13984
rect 11572 13941 11581 13975
rect 11581 13941 11615 13975
rect 11615 13941 11624 13975
rect 11572 13932 11624 13941
rect 12400 14000 12452 14052
rect 25464 14068 25516 14120
rect 12768 13932 12820 13984
rect 27948 14000 28000 14052
rect 13688 13975 13740 13984
rect 13688 13941 13697 13975
rect 13697 13941 13731 13975
rect 13731 13941 13740 13975
rect 13688 13932 13740 13941
rect 13872 13932 13924 13984
rect 14240 13864 14292 13916
rect 13964 13796 14016 13848
rect 14792 13975 14844 13984
rect 14792 13941 14801 13975
rect 14801 13941 14835 13975
rect 14835 13941 14844 13975
rect 14792 13932 14844 13941
rect 16816 13975 16868 13984
rect 16816 13941 16825 13975
rect 16825 13941 16859 13975
rect 16859 13941 16868 13975
rect 16816 13932 16868 13941
rect 16908 13932 16960 13984
rect 17552 13975 17604 13984
rect 17552 13941 17561 13975
rect 17561 13941 17595 13975
rect 17595 13941 17604 13975
rect 17552 13932 17604 13941
rect 19116 13932 19168 13984
rect 20036 13975 20088 13984
rect 20036 13941 20045 13975
rect 20045 13941 20079 13975
rect 20079 13941 20088 13975
rect 20036 13932 20088 13941
rect 20312 13932 20364 13984
rect 20772 13975 20824 13984
rect 20772 13941 20781 13975
rect 20781 13941 20815 13975
rect 20815 13941 20824 13975
rect 20772 13932 20824 13941
rect 22336 13975 22388 13984
rect 22336 13941 22345 13975
rect 22345 13941 22379 13975
rect 22379 13941 22388 13975
rect 22336 13932 22388 13941
rect 22612 13932 22664 13984
rect 23808 13932 23860 13984
rect 25096 13975 25148 13984
rect 17276 13864 17328 13916
rect 17736 13864 17788 13916
rect 20404 13907 20456 13916
rect 14976 13796 15028 13848
rect 20404 13873 20413 13907
rect 20413 13873 20447 13907
rect 20447 13873 20456 13907
rect 20404 13864 20456 13873
rect 18748 13796 18800 13848
rect 24268 13796 24320 13848
rect 25096 13941 25105 13975
rect 25105 13941 25139 13975
rect 25139 13941 25148 13975
rect 25096 13932 25148 13941
rect 24912 13864 24964 13916
rect 25464 13932 25516 13984
rect 28500 13932 28552 13984
rect 27856 13864 27908 13916
rect 25188 13796 25240 13848
rect 19142 13694 19194 13746
rect 19206 13694 19258 13746
rect 19270 13694 19322 13746
rect 19334 13694 19386 13746
rect 29142 13694 29194 13746
rect 29206 13694 29258 13746
rect 29270 13694 29322 13746
rect 29334 13694 29386 13746
rect 12768 13524 12820 13576
rect 13872 13524 13924 13576
rect 14884 13524 14936 13576
rect 15896 13524 15948 13576
rect 17736 13567 17788 13576
rect 12032 13456 12084 13508
rect 13136 13456 13188 13508
rect 13964 13499 14016 13508
rect 13964 13465 13973 13499
rect 13973 13465 14007 13499
rect 14007 13465 14016 13499
rect 13964 13456 14016 13465
rect 17736 13533 17745 13567
rect 17745 13533 17779 13567
rect 17779 13533 17788 13567
rect 17736 13524 17788 13533
rect 19576 13592 19628 13644
rect 22612 13592 22664 13644
rect 23900 13592 23952 13644
rect 29512 13592 29564 13644
rect 14976 13388 15028 13440
rect 16264 13431 16316 13440
rect 16264 13397 16273 13431
rect 16273 13397 16307 13431
rect 16307 13397 16316 13431
rect 16264 13388 16316 13397
rect 14240 13363 14292 13372
rect 14240 13329 14249 13363
rect 14249 13329 14283 13363
rect 14283 13329 14292 13363
rect 14240 13320 14292 13329
rect 18380 13499 18432 13508
rect 18380 13465 18389 13499
rect 18389 13465 18423 13499
rect 18423 13465 18432 13499
rect 18380 13456 18432 13465
rect 18748 13499 18800 13508
rect 18748 13465 18757 13499
rect 18757 13465 18791 13499
rect 18791 13465 18800 13499
rect 18748 13456 18800 13465
rect 18932 13499 18984 13508
rect 18932 13465 18941 13499
rect 18941 13465 18975 13499
rect 18975 13465 18984 13499
rect 18932 13456 18984 13465
rect 20036 13456 20088 13508
rect 20312 13456 20364 13508
rect 21140 13456 21192 13508
rect 16448 13431 16500 13440
rect 16448 13397 16457 13431
rect 16457 13397 16491 13431
rect 16491 13397 16500 13431
rect 18288 13431 18340 13440
rect 16448 13388 16500 13397
rect 18288 13397 18297 13431
rect 18297 13397 18331 13431
rect 18331 13397 18340 13431
rect 18288 13388 18340 13397
rect 21232 13431 21284 13440
rect 21232 13397 21241 13431
rect 21241 13397 21275 13431
rect 21275 13397 21284 13431
rect 22060 13456 22112 13508
rect 28132 13524 28184 13576
rect 23808 13456 23860 13508
rect 24268 13499 24320 13508
rect 24268 13465 24277 13499
rect 24277 13465 24311 13499
rect 24311 13465 24320 13499
rect 24268 13456 24320 13465
rect 25464 13499 25516 13508
rect 25464 13465 25473 13499
rect 25473 13465 25507 13499
rect 25507 13465 25516 13499
rect 26568 13499 26620 13508
rect 25464 13456 25516 13465
rect 26568 13465 26577 13499
rect 26577 13465 26611 13499
rect 26611 13465 26620 13499
rect 26568 13456 26620 13465
rect 28960 13456 29012 13508
rect 21232 13388 21284 13397
rect 25280 13388 25332 13440
rect 27488 13388 27540 13440
rect 28592 13431 28644 13440
rect 28592 13397 28601 13431
rect 28601 13397 28635 13431
rect 28635 13397 28644 13431
rect 28592 13388 28644 13397
rect 17184 13320 17236 13372
rect 17276 13320 17328 13372
rect 12952 13252 13004 13304
rect 13688 13252 13740 13304
rect 24912 13252 24964 13304
rect 14142 13150 14194 13202
rect 14206 13150 14258 13202
rect 14270 13150 14322 13202
rect 14334 13150 14386 13202
rect 24142 13150 24194 13202
rect 24206 13150 24258 13202
rect 24270 13150 24322 13202
rect 24334 13150 24386 13202
rect 18380 13048 18432 13100
rect 12952 12955 13004 12964
rect 12952 12921 12961 12955
rect 12961 12921 12995 12955
rect 12995 12921 13004 12955
rect 12952 12912 13004 12921
rect 12032 12844 12084 12896
rect 12584 12844 12636 12896
rect 13412 12955 13464 12964
rect 13412 12921 13421 12955
rect 13421 12921 13455 12955
rect 13455 12921 13464 12955
rect 13412 12912 13464 12921
rect 13320 12708 13372 12760
rect 14148 12887 14200 12896
rect 14148 12853 14157 12887
rect 14157 12853 14191 12887
rect 14191 12853 14200 12887
rect 14148 12844 14200 12853
rect 14332 12844 14384 12896
rect 18840 12912 18892 12964
rect 20588 13048 20640 13100
rect 25280 13048 25332 13100
rect 28132 13091 28184 13100
rect 28132 13057 28141 13091
rect 28141 13057 28175 13091
rect 28175 13057 28184 13091
rect 28132 13048 28184 13057
rect 19024 12980 19076 13032
rect 14976 12844 15028 12896
rect 19300 12912 19352 12964
rect 21232 12980 21284 13032
rect 20036 12912 20088 12964
rect 20680 12912 20732 12964
rect 19392 12887 19444 12896
rect 19392 12853 19401 12887
rect 19401 12853 19435 12887
rect 19435 12853 19444 12887
rect 19392 12844 19444 12853
rect 21232 12887 21284 12896
rect 21232 12853 21241 12887
rect 21241 12853 21275 12887
rect 21275 12853 21284 12887
rect 21232 12844 21284 12853
rect 22152 12844 22204 12896
rect 25188 12912 25240 12964
rect 27396 12912 27448 12964
rect 28776 12955 28828 12964
rect 28776 12921 28785 12955
rect 28785 12921 28819 12955
rect 28819 12921 28828 12955
rect 28776 12912 28828 12921
rect 24728 12844 24780 12896
rect 24912 12887 24964 12896
rect 24912 12853 24921 12887
rect 24921 12853 24955 12887
rect 24955 12853 24964 12887
rect 24912 12844 24964 12853
rect 25096 12887 25148 12896
rect 25096 12853 25105 12887
rect 25105 12853 25139 12887
rect 25139 12853 25148 12887
rect 25924 12887 25976 12896
rect 25096 12844 25148 12853
rect 25924 12853 25933 12887
rect 25933 12853 25967 12887
rect 25967 12853 25976 12887
rect 25924 12844 25976 12853
rect 26016 12887 26068 12896
rect 26016 12853 26025 12887
rect 26025 12853 26059 12887
rect 26059 12853 26068 12887
rect 26016 12844 26068 12853
rect 19576 12776 19628 12828
rect 27764 12776 27816 12828
rect 29604 12844 29656 12896
rect 14148 12708 14200 12760
rect 14792 12708 14844 12760
rect 15988 12708 16040 12760
rect 19944 12708 19996 12760
rect 21692 12708 21744 12760
rect 23900 12751 23952 12760
rect 23900 12717 23909 12751
rect 23909 12717 23943 12751
rect 23943 12717 23952 12751
rect 23900 12708 23952 12717
rect 25372 12708 25424 12760
rect 26384 12708 26436 12760
rect 28960 12776 29012 12828
rect 19142 12606 19194 12658
rect 19206 12606 19258 12658
rect 19270 12606 19322 12658
rect 19334 12606 19386 12658
rect 29142 12606 29194 12658
rect 29206 12606 29258 12658
rect 29270 12606 29322 12658
rect 29334 12606 29386 12658
rect 12308 12504 12360 12556
rect 13136 12479 13188 12488
rect 13136 12445 13145 12479
rect 13145 12445 13179 12479
rect 13179 12445 13188 12479
rect 13136 12436 13188 12445
rect 12032 12411 12084 12420
rect 12032 12377 12041 12411
rect 12041 12377 12075 12411
rect 12075 12377 12084 12411
rect 12032 12368 12084 12377
rect 12584 12411 12636 12420
rect 12584 12377 12593 12411
rect 12593 12377 12627 12411
rect 12627 12377 12636 12411
rect 12584 12368 12636 12377
rect 12768 12368 12820 12420
rect 14148 12504 14200 12556
rect 13688 12368 13740 12420
rect 14792 12368 14844 12420
rect 15804 12368 15856 12420
rect 16540 12368 16592 12420
rect 16908 12436 16960 12488
rect 17552 12436 17604 12488
rect 18196 12436 18248 12488
rect 18748 12436 18800 12488
rect 19852 12504 19904 12556
rect 23532 12504 23584 12556
rect 25372 12436 25424 12488
rect 26568 12504 26620 12556
rect 27856 12504 27908 12556
rect 26476 12436 26528 12488
rect 27488 12479 27540 12488
rect 27488 12445 27497 12479
rect 27497 12445 27531 12479
rect 27531 12445 27540 12479
rect 27488 12436 27540 12445
rect 19576 12411 19628 12420
rect 14332 12300 14384 12352
rect 13412 12232 13464 12284
rect 19576 12377 19585 12411
rect 19585 12377 19619 12411
rect 19619 12377 19628 12411
rect 19576 12368 19628 12377
rect 21140 12411 21192 12420
rect 21140 12377 21149 12411
rect 21149 12377 21183 12411
rect 21183 12377 21192 12411
rect 21140 12368 21192 12377
rect 21508 12411 21560 12420
rect 21508 12377 21517 12411
rect 21517 12377 21551 12411
rect 21551 12377 21560 12411
rect 21508 12368 21560 12377
rect 21692 12411 21744 12420
rect 21692 12377 21701 12411
rect 21701 12377 21735 12411
rect 21735 12377 21744 12411
rect 21692 12368 21744 12377
rect 25464 12411 25516 12420
rect 25464 12377 25473 12411
rect 25473 12377 25507 12411
rect 25507 12377 25516 12411
rect 25464 12368 25516 12377
rect 28040 12436 28092 12488
rect 28592 12368 28644 12420
rect 16908 12343 16960 12352
rect 16908 12309 16917 12343
rect 16917 12309 16951 12343
rect 16951 12309 16960 12343
rect 16908 12300 16960 12309
rect 21232 12343 21284 12352
rect 21232 12309 21241 12343
rect 21241 12309 21275 12343
rect 21275 12309 21284 12343
rect 21232 12300 21284 12309
rect 22244 12343 22296 12352
rect 22244 12309 22253 12343
rect 22253 12309 22287 12343
rect 22287 12309 22296 12343
rect 22244 12300 22296 12309
rect 22520 12343 22572 12352
rect 22520 12309 22529 12343
rect 22529 12309 22563 12343
rect 22563 12309 22572 12343
rect 22520 12300 22572 12309
rect 25740 12343 25792 12352
rect 13964 12164 14016 12216
rect 16080 12207 16132 12216
rect 16080 12173 16089 12207
rect 16089 12173 16123 12207
rect 16123 12173 16132 12207
rect 16080 12164 16132 12173
rect 18932 12164 18984 12216
rect 22152 12164 22204 12216
rect 25740 12309 25749 12343
rect 25749 12309 25783 12343
rect 25783 12309 25792 12343
rect 25740 12300 25792 12309
rect 14142 12062 14194 12114
rect 14206 12062 14258 12114
rect 14270 12062 14322 12114
rect 14334 12062 14386 12114
rect 24142 12062 24194 12114
rect 24206 12062 24258 12114
rect 24270 12062 24322 12114
rect 24334 12062 24386 12114
rect 11572 11960 11624 12012
rect 12768 12003 12820 12012
rect 12768 11969 12777 12003
rect 12777 11969 12811 12003
rect 12811 11969 12820 12003
rect 12768 11960 12820 11969
rect 14516 11960 14568 12012
rect 20956 11960 21008 12012
rect 21232 11960 21284 12012
rect 26476 11960 26528 12012
rect 28040 12003 28092 12012
rect 28040 11969 28049 12003
rect 28049 11969 28083 12003
rect 28083 11969 28092 12003
rect 28040 11960 28092 11969
rect 17000 11892 17052 11944
rect 13412 11824 13464 11876
rect 10468 11756 10520 11808
rect 13320 11756 13372 11808
rect 14792 11824 14844 11876
rect 14976 11824 15028 11876
rect 16908 11824 16960 11876
rect 18932 11867 18984 11876
rect 18932 11833 18941 11867
rect 18941 11833 18975 11867
rect 18975 11833 18984 11867
rect 18932 11824 18984 11833
rect 20680 11867 20732 11876
rect 20680 11833 20689 11867
rect 20689 11833 20723 11867
rect 20723 11833 20732 11867
rect 20680 11824 20732 11833
rect 21692 11892 21744 11944
rect 22244 11892 22296 11944
rect 13688 11799 13740 11808
rect 13688 11765 13697 11799
rect 13697 11765 13731 11799
rect 13731 11765 13740 11799
rect 13688 11756 13740 11765
rect 14056 11756 14108 11808
rect 16080 11756 16132 11808
rect 17276 11756 17328 11808
rect 17644 11756 17696 11808
rect 18196 11799 18248 11808
rect 18196 11765 18205 11799
rect 18205 11765 18239 11799
rect 18239 11765 18248 11799
rect 18196 11756 18248 11765
rect 21508 11824 21560 11876
rect 25464 11824 25516 11876
rect 25740 11824 25792 11876
rect 19024 11688 19076 11740
rect 19944 11688 19996 11740
rect 20956 11688 21008 11740
rect 22152 11756 22204 11808
rect 26384 11799 26436 11808
rect 26384 11765 26393 11799
rect 26393 11765 26427 11799
rect 26427 11765 26436 11799
rect 26384 11756 26436 11765
rect 27488 11756 27540 11808
rect 16080 11620 16132 11672
rect 18012 11620 18064 11672
rect 25556 11688 25608 11740
rect 23716 11620 23768 11672
rect 24452 11620 24504 11672
rect 19142 11518 19194 11570
rect 19206 11518 19258 11570
rect 19270 11518 19322 11570
rect 19334 11518 19386 11570
rect 29142 11518 29194 11570
rect 29206 11518 29258 11570
rect 29270 11518 29322 11570
rect 29334 11518 29386 11570
rect 16080 11459 16132 11468
rect 16080 11425 16089 11459
rect 16089 11425 16123 11459
rect 16123 11425 16132 11459
rect 16080 11416 16132 11425
rect 17552 11459 17604 11468
rect 17552 11425 17561 11459
rect 17561 11425 17595 11459
rect 17595 11425 17604 11459
rect 17552 11416 17604 11425
rect 19484 11416 19536 11468
rect 19944 11416 19996 11468
rect 25556 11459 25608 11468
rect 25556 11425 25565 11459
rect 25565 11425 25599 11459
rect 25599 11425 25608 11459
rect 25556 11416 25608 11425
rect 15804 11323 15856 11332
rect 15804 11289 15813 11323
rect 15813 11289 15847 11323
rect 15847 11289 15856 11323
rect 15804 11280 15856 11289
rect 14976 11255 15028 11264
rect 14976 11221 14985 11255
rect 14985 11221 15019 11255
rect 15019 11221 15028 11255
rect 14976 11212 15028 11221
rect 17276 11348 17328 11400
rect 20404 11348 20456 11400
rect 17184 11280 17236 11332
rect 17276 11212 17328 11264
rect 18196 11280 18248 11332
rect 20956 11280 21008 11332
rect 22520 11348 22572 11400
rect 21692 11280 21744 11332
rect 23900 11323 23952 11332
rect 23900 11289 23909 11323
rect 23909 11289 23943 11323
rect 23943 11289 23952 11323
rect 23900 11280 23952 11289
rect 25372 11323 25424 11332
rect 25372 11289 25381 11323
rect 25381 11289 25415 11323
rect 25415 11289 25424 11323
rect 25372 11280 25424 11289
rect 15804 11144 15856 11196
rect 21692 11144 21744 11196
rect 14142 10974 14194 11026
rect 14206 10974 14258 11026
rect 14270 10974 14322 11026
rect 14334 10974 14386 11026
rect 24142 10974 24194 11026
rect 24206 10974 24258 11026
rect 24270 10974 24322 11026
rect 24334 10974 24386 11026
<< metal2 >>
rect 10650 31576 10706 32376
rect 12490 31576 12546 32376
rect 14514 31576 14570 32376
rect 16354 31576 16410 32376
rect 18194 31576 18250 32376
rect 20218 31576 20274 32376
rect 22058 31576 22114 32376
rect 23898 31576 23954 32376
rect 25922 31576 25978 32376
rect 27762 31576 27818 32376
rect 29602 31576 29658 32376
rect 10664 28746 10692 31576
rect 10652 28740 10704 28746
rect 10652 28682 10704 28688
rect 12504 28270 12532 31576
rect 14116 29524 14412 29544
rect 14172 29522 14196 29524
rect 14252 29522 14276 29524
rect 14332 29522 14356 29524
rect 14194 29470 14196 29522
rect 14258 29470 14270 29522
rect 14332 29470 14334 29522
rect 14172 29468 14196 29470
rect 14252 29468 14276 29470
rect 14332 29468 14356 29470
rect 14116 29448 14412 29468
rect 13502 29320 13558 29329
rect 13502 29255 13504 29264
rect 13556 29255 13558 29264
rect 13504 29226 13556 29232
rect 14056 29148 14108 29154
rect 14056 29090 14108 29096
rect 14068 28746 14096 29090
rect 14528 28882 14556 31576
rect 14976 29828 15028 29834
rect 14976 29770 15028 29776
rect 15068 29828 15120 29834
rect 15068 29770 15120 29776
rect 14700 29624 14752 29630
rect 14700 29566 14752 29572
rect 14516 28876 14568 28882
rect 14516 28818 14568 28824
rect 14056 28740 14108 28746
rect 14056 28682 14108 28688
rect 14068 28626 14096 28682
rect 13976 28598 14096 28626
rect 12492 28264 12544 28270
rect 12492 28206 12544 28212
rect 13976 28202 14004 28598
rect 14116 28436 14412 28456
rect 14172 28434 14196 28436
rect 14252 28434 14276 28436
rect 14332 28434 14356 28436
rect 14194 28382 14196 28434
rect 14258 28382 14270 28434
rect 14332 28382 14334 28434
rect 14172 28380 14196 28382
rect 14252 28380 14276 28382
rect 14332 28380 14356 28382
rect 14116 28360 14412 28380
rect 13964 28196 14016 28202
rect 13964 28138 14016 28144
rect 14712 28134 14740 29566
rect 14988 28746 15016 29770
rect 15080 28814 15108 29770
rect 15988 29624 16040 29630
rect 15988 29566 16040 29572
rect 15160 29216 15212 29222
rect 15160 29158 15212 29164
rect 15068 28808 15120 28814
rect 15068 28750 15120 28756
rect 14976 28740 15028 28746
rect 14976 28682 15028 28688
rect 15080 28202 15108 28750
rect 15172 28338 15200 29158
rect 15436 29148 15488 29154
rect 15436 29090 15488 29096
rect 15448 28746 15476 29090
rect 15436 28740 15488 28746
rect 15436 28682 15488 28688
rect 15160 28332 15212 28338
rect 15160 28274 15212 28280
rect 15448 28202 15476 28682
rect 15068 28196 15120 28202
rect 15068 28138 15120 28144
rect 15436 28196 15488 28202
rect 15436 28138 15488 28144
rect 16000 28134 16028 29566
rect 16368 29290 16396 31576
rect 16356 29284 16408 29290
rect 16356 29226 16408 29232
rect 17644 29216 17696 29222
rect 17644 29158 17696 29164
rect 16724 28740 16776 28746
rect 16724 28682 16776 28688
rect 16632 28604 16684 28610
rect 16632 28546 16684 28552
rect 16644 28202 16672 28546
rect 16632 28196 16684 28202
rect 16632 28138 16684 28144
rect 16736 28134 16764 28682
rect 17656 28678 17684 29158
rect 18208 28746 18236 31576
rect 19116 30068 19412 30088
rect 19172 30066 19196 30068
rect 19252 30066 19276 30068
rect 19332 30066 19356 30068
rect 19194 30014 19196 30066
rect 19258 30014 19270 30066
rect 19332 30014 19334 30066
rect 19172 30012 19196 30014
rect 19252 30012 19276 30014
rect 19332 30012 19356 30014
rect 19116 29992 19412 30012
rect 19760 29828 19812 29834
rect 19760 29770 19812 29776
rect 19852 29828 19904 29834
rect 19852 29770 19904 29776
rect 19024 29624 19076 29630
rect 19024 29566 19076 29572
rect 19668 29624 19720 29630
rect 19668 29566 19720 29572
rect 18380 29352 18432 29358
rect 18380 29294 18432 29300
rect 18196 28740 18248 28746
rect 18196 28682 18248 28688
rect 17644 28672 17696 28678
rect 17644 28614 17696 28620
rect 14700 28128 14752 28134
rect 14700 28070 14752 28076
rect 15988 28128 16040 28134
rect 15988 28070 16040 28076
rect 16724 28128 16776 28134
rect 16724 28070 16776 28076
rect 17656 27794 17684 28614
rect 18392 28610 18420 29294
rect 18564 29148 18616 29154
rect 18564 29090 18616 29096
rect 18380 28604 18432 28610
rect 18380 28546 18432 28552
rect 18288 28536 18340 28542
rect 18288 28478 18340 28484
rect 18012 28128 18064 28134
rect 18012 28070 18064 28076
rect 17828 28060 17880 28066
rect 17828 28002 17880 28008
rect 17840 27794 17868 28002
rect 17644 27788 17696 27794
rect 17644 27730 17696 27736
rect 17828 27788 17880 27794
rect 17828 27730 17880 27736
rect 11940 27652 11992 27658
rect 11940 27594 11992 27600
rect 11296 27040 11348 27046
rect 11296 26982 11348 26988
rect 11308 24870 11336 26982
rect 11572 26972 11624 26978
rect 11572 26914 11624 26920
rect 11584 26638 11612 26914
rect 11572 26632 11624 26638
rect 11572 26574 11624 26580
rect 11662 26328 11718 26337
rect 11662 26263 11718 26272
rect 11676 25958 11704 26263
rect 11664 25952 11716 25958
rect 11664 25894 11716 25900
rect 11952 25482 11980 27594
rect 18024 27590 18052 28070
rect 18300 27658 18328 28478
rect 18392 27998 18420 28546
rect 18576 28134 18604 29090
rect 19036 28814 19064 29566
rect 19680 29290 19708 29566
rect 19772 29358 19800 29770
rect 19760 29352 19812 29358
rect 19760 29294 19812 29300
rect 19668 29284 19720 29290
rect 19668 29226 19720 29232
rect 19116 28980 19412 29000
rect 19172 28978 19196 28980
rect 19252 28978 19276 28980
rect 19332 28978 19356 28980
rect 19194 28926 19196 28978
rect 19258 28926 19270 28978
rect 19332 28926 19334 28978
rect 19172 28924 19196 28926
rect 19252 28924 19276 28926
rect 19332 28924 19356 28926
rect 19116 28904 19412 28924
rect 19024 28808 19076 28814
rect 19024 28750 19076 28756
rect 19668 28536 19720 28542
rect 19668 28478 19720 28484
rect 18564 28128 18616 28134
rect 18564 28070 18616 28076
rect 18380 27992 18432 27998
rect 18380 27934 18432 27940
rect 19116 27892 19412 27912
rect 19172 27890 19196 27892
rect 19252 27890 19276 27892
rect 19332 27890 19356 27892
rect 19194 27838 19196 27890
rect 19258 27838 19270 27890
rect 19332 27838 19334 27890
rect 19172 27836 19196 27838
rect 19252 27836 19276 27838
rect 19332 27836 19356 27838
rect 19116 27816 19412 27836
rect 18840 27720 18892 27726
rect 18840 27662 18892 27668
rect 19484 27720 19536 27726
rect 19484 27662 19536 27668
rect 18288 27652 18340 27658
rect 18288 27594 18340 27600
rect 18012 27584 18064 27590
rect 18012 27526 18064 27532
rect 12308 27448 12360 27454
rect 12308 27390 12360 27396
rect 14792 27448 14844 27454
rect 14792 27390 14844 27396
rect 12320 26978 12348 27390
rect 14116 27348 14412 27368
rect 14172 27346 14196 27348
rect 14252 27346 14276 27348
rect 14332 27346 14356 27348
rect 14194 27294 14196 27346
rect 14258 27294 14270 27346
rect 14332 27294 14334 27346
rect 14172 27292 14196 27294
rect 14252 27292 14276 27294
rect 14332 27292 14356 27294
rect 14116 27272 14412 27292
rect 14804 26978 14832 27390
rect 18024 27250 18052 27526
rect 18012 27244 18064 27250
rect 18012 27186 18064 27192
rect 18748 27244 18800 27250
rect 18748 27186 18800 27192
rect 16908 27108 16960 27114
rect 16908 27050 16960 27056
rect 12308 26972 12360 26978
rect 12308 26914 12360 26920
rect 13228 26972 13280 26978
rect 13228 26914 13280 26920
rect 14056 26972 14108 26978
rect 14056 26914 14108 26920
rect 14792 26972 14844 26978
rect 14792 26914 14844 26920
rect 15804 26972 15856 26978
rect 15804 26914 15856 26920
rect 16724 26972 16776 26978
rect 16724 26914 16776 26920
rect 13240 26570 13268 26914
rect 12584 26564 12636 26570
rect 12584 26506 12636 26512
rect 12676 26564 12728 26570
rect 12676 26506 12728 26512
rect 12860 26564 12912 26570
rect 12860 26506 12912 26512
rect 13228 26564 13280 26570
rect 13228 26506 13280 26512
rect 12596 26162 12624 26506
rect 12584 26156 12636 26162
rect 12584 26098 12636 26104
rect 12688 25618 12716 26506
rect 12872 26094 12900 26506
rect 13136 26496 13188 26502
rect 13136 26438 13188 26444
rect 12860 26088 12912 26094
rect 12860 26030 12912 26036
rect 12768 25952 12820 25958
rect 12768 25894 12820 25900
rect 12676 25612 12728 25618
rect 12676 25554 12728 25560
rect 12780 25550 12808 25894
rect 12768 25544 12820 25550
rect 12768 25486 12820 25492
rect 11940 25476 11992 25482
rect 11940 25418 11992 25424
rect 11296 24864 11348 24870
rect 11296 24806 11348 24812
rect 11308 21130 11336 24806
rect 11572 24796 11624 24802
rect 11572 24738 11624 24744
rect 11584 23850 11612 24738
rect 11572 23844 11624 23850
rect 11572 23786 11624 23792
rect 11952 22218 11980 25418
rect 12124 25272 12176 25278
rect 12124 25214 12176 25220
rect 12136 24802 12164 25214
rect 12124 24796 12176 24802
rect 12124 24738 12176 24744
rect 12124 24388 12176 24394
rect 12124 24330 12176 24336
rect 12400 24388 12452 24394
rect 12400 24330 12452 24336
rect 12032 24184 12084 24190
rect 12032 24126 12084 24132
rect 12044 23782 12072 24126
rect 12032 23776 12084 23782
rect 12032 23718 12084 23724
rect 12136 23374 12164 24330
rect 12216 23776 12268 23782
rect 12216 23718 12268 23724
rect 12124 23368 12176 23374
rect 12124 23310 12176 23316
rect 12136 22694 12164 23310
rect 12228 22762 12256 23718
rect 12412 23170 12440 24330
rect 12584 23708 12636 23714
rect 12872 23696 12900 26030
rect 12952 24184 13004 24190
rect 12952 24126 13004 24132
rect 12636 23668 12900 23696
rect 12584 23650 12636 23656
rect 12400 23164 12452 23170
rect 12400 23106 12452 23112
rect 12216 22756 12268 22762
rect 12216 22698 12268 22704
rect 12412 22694 12440 23106
rect 12124 22688 12176 22694
rect 12124 22630 12176 22636
rect 12400 22688 12452 22694
rect 12400 22630 12452 22636
rect 11940 22212 11992 22218
rect 11940 22154 11992 22160
rect 11848 21532 11900 21538
rect 11848 21474 11900 21480
rect 11860 21198 11888 21474
rect 11848 21192 11900 21198
rect 11848 21134 11900 21140
rect 11296 21124 11348 21130
rect 11296 21066 11348 21072
rect 11308 16778 11336 21066
rect 11662 20888 11718 20897
rect 11662 20823 11718 20832
rect 11676 20042 11704 20823
rect 11664 20036 11716 20042
rect 11664 19978 11716 19984
rect 11664 17792 11716 17798
rect 11664 17734 11716 17740
rect 11676 16846 11704 17734
rect 11664 16840 11716 16846
rect 11664 16782 11716 16788
rect 11296 16772 11348 16778
rect 11296 16714 11348 16720
rect 11952 16166 11980 22154
rect 12032 22008 12084 22014
rect 12032 21950 12084 21956
rect 12044 21198 12072 21950
rect 12216 21600 12268 21606
rect 12216 21542 12268 21548
rect 12596 21588 12624 23650
rect 12964 23238 12992 24126
rect 13044 23776 13096 23782
rect 13148 23764 13176 26438
rect 13240 26434 13268 26506
rect 14068 26450 14096 26914
rect 15816 26706 15844 26914
rect 15804 26700 15856 26706
rect 15804 26642 15856 26648
rect 15252 26564 15304 26570
rect 15252 26506 15304 26512
rect 13228 26428 13280 26434
rect 13228 26370 13280 26376
rect 13976 26422 14096 26450
rect 13976 26144 14004 26422
rect 14976 26360 15028 26366
rect 14976 26302 15028 26308
rect 14116 26260 14412 26280
rect 14172 26258 14196 26260
rect 14252 26258 14276 26260
rect 14332 26258 14356 26260
rect 14194 26206 14196 26258
rect 14258 26206 14270 26258
rect 14332 26206 14334 26258
rect 14172 26204 14196 26206
rect 14252 26204 14276 26206
rect 14332 26204 14356 26206
rect 14116 26184 14412 26204
rect 13976 26116 14096 26144
rect 14068 26026 14096 26116
rect 14056 26020 14108 26026
rect 14056 25962 14108 25968
rect 13504 25952 13556 25958
rect 13504 25894 13556 25900
rect 14516 25952 14568 25958
rect 14516 25894 14568 25900
rect 14884 25952 14936 25958
rect 14884 25894 14936 25900
rect 13516 25482 13544 25894
rect 13504 25476 13556 25482
rect 13504 25418 13556 25424
rect 13412 24796 13464 24802
rect 13412 24738 13464 24744
rect 13424 24394 13452 24738
rect 13412 24388 13464 24394
rect 13412 24330 13464 24336
rect 13424 23850 13452 24330
rect 13412 23844 13464 23850
rect 13412 23786 13464 23792
rect 13096 23736 13176 23764
rect 13044 23718 13096 23724
rect 12952 23232 13004 23238
rect 12952 23174 13004 23180
rect 13056 21674 13084 23718
rect 13424 23306 13452 23786
rect 13516 23782 13544 25418
rect 14528 25414 14556 25894
rect 14896 25822 14924 25894
rect 14988 25822 15016 26302
rect 15264 26026 15292 26506
rect 16736 26502 16764 26914
rect 16920 26910 16948 27050
rect 18760 27046 18788 27186
rect 17736 27040 17788 27046
rect 17736 26982 17788 26988
rect 18748 27040 18800 27046
rect 18748 26982 18800 26988
rect 16908 26904 16960 26910
rect 16908 26846 16960 26852
rect 15344 26496 15396 26502
rect 15344 26438 15396 26444
rect 16724 26496 16776 26502
rect 16724 26438 16776 26444
rect 15356 26026 15384 26438
rect 16736 26366 16764 26438
rect 16724 26360 16776 26366
rect 16724 26302 16776 26308
rect 15252 26020 15304 26026
rect 15252 25962 15304 25968
rect 15344 26020 15396 26026
rect 15344 25962 15396 25968
rect 16736 25890 16764 26302
rect 16920 25958 16948 26846
rect 17748 26570 17776 26982
rect 17828 26904 17880 26910
rect 17828 26846 17880 26852
rect 17840 26638 17868 26846
rect 17828 26632 17880 26638
rect 17828 26574 17880 26580
rect 18012 26632 18064 26638
rect 18012 26574 18064 26580
rect 17552 26564 17604 26570
rect 17552 26506 17604 26512
rect 17736 26564 17788 26570
rect 17736 26506 17788 26512
rect 16908 25952 16960 25958
rect 16908 25894 16960 25900
rect 17184 25952 17236 25958
rect 17184 25894 17236 25900
rect 15712 25884 15764 25890
rect 15712 25826 15764 25832
rect 16724 25884 16776 25890
rect 16724 25826 16776 25832
rect 14884 25816 14936 25822
rect 14884 25758 14936 25764
rect 14976 25816 15028 25822
rect 14976 25758 15028 25764
rect 14608 25544 14660 25550
rect 14608 25486 14660 25492
rect 14516 25408 14568 25414
rect 14516 25350 14568 25356
rect 14116 25172 14412 25192
rect 14172 25170 14196 25172
rect 14252 25170 14276 25172
rect 14332 25170 14356 25172
rect 14194 25118 14196 25170
rect 14258 25118 14270 25170
rect 14332 25118 14334 25170
rect 14172 25116 14196 25118
rect 14252 25116 14276 25118
rect 14332 25116 14356 25118
rect 14116 25096 14412 25116
rect 14528 25006 14556 25350
rect 14516 25000 14568 25006
rect 14516 24942 14568 24948
rect 14516 24864 14568 24870
rect 14620 24852 14648 25486
rect 14792 25476 14844 25482
rect 14792 25418 14844 25424
rect 14884 25476 14936 25482
rect 14884 25418 14936 25424
rect 14568 24824 14648 24852
rect 14516 24806 14568 24812
rect 14116 24084 14412 24104
rect 14172 24082 14196 24084
rect 14252 24082 14276 24084
rect 14332 24082 14356 24084
rect 14194 24030 14196 24082
rect 14258 24030 14270 24082
rect 14332 24030 14334 24082
rect 14172 24028 14196 24030
rect 14252 24028 14276 24030
rect 14332 24028 14356 24030
rect 14116 24008 14412 24028
rect 13504 23776 13556 23782
rect 13504 23718 13556 23724
rect 13964 23776 14016 23782
rect 13964 23718 14016 23724
rect 13596 23640 13648 23646
rect 13596 23582 13648 23588
rect 13870 23608 13926 23617
rect 13608 23374 13636 23582
rect 13870 23543 13926 23552
rect 13596 23368 13648 23374
rect 13596 23310 13648 23316
rect 13884 23306 13912 23543
rect 13228 23300 13280 23306
rect 13228 23242 13280 23248
rect 13412 23300 13464 23306
rect 13412 23242 13464 23248
rect 13872 23300 13924 23306
rect 13872 23242 13924 23248
rect 13240 22898 13268 23242
rect 13228 22892 13280 22898
rect 13228 22834 13280 22840
rect 13688 22620 13740 22626
rect 13688 22562 13740 22568
rect 13044 21668 13096 21674
rect 13044 21610 13096 21616
rect 12676 21600 12728 21606
rect 12596 21560 12676 21588
rect 12032 21192 12084 21198
rect 12032 21134 12084 21140
rect 12228 20586 12256 21542
rect 12216 20580 12268 20586
rect 12216 20522 12268 20528
rect 12596 18478 12624 21560
rect 12676 21542 12728 21548
rect 12768 21532 12820 21538
rect 12768 21474 12820 21480
rect 12676 20376 12728 20382
rect 12676 20318 12728 20324
rect 12688 20042 12716 20318
rect 12676 20036 12728 20042
rect 12676 19978 12728 19984
rect 12780 19974 12808 21474
rect 12952 20512 13004 20518
rect 12952 20454 13004 20460
rect 12964 20042 12992 20454
rect 12952 20036 13004 20042
rect 12872 19996 12952 20024
rect 12768 19968 12820 19974
rect 12768 19910 12820 19916
rect 12780 19498 12808 19910
rect 12768 19492 12820 19498
rect 12768 19434 12820 19440
rect 12872 19022 12900 19996
rect 12952 19978 13004 19984
rect 12860 19016 12912 19022
rect 12860 18958 12912 18964
rect 12952 18948 13004 18954
rect 12952 18890 13004 18896
rect 12584 18472 12636 18478
rect 12584 18414 12636 18420
rect 12492 18200 12544 18206
rect 12492 18142 12544 18148
rect 12504 17254 12532 18142
rect 12596 17866 12624 18414
rect 12860 18336 12912 18342
rect 12860 18278 12912 18284
rect 12674 17896 12730 17905
rect 12584 17860 12636 17866
rect 12872 17866 12900 18278
rect 12674 17831 12730 17840
rect 12860 17860 12912 17866
rect 12584 17802 12636 17808
rect 12492 17248 12544 17254
rect 12492 17190 12544 17196
rect 12124 16840 12176 16846
rect 12124 16782 12176 16788
rect 12136 16370 12164 16782
rect 12124 16364 12176 16370
rect 12124 16306 12176 16312
rect 11940 16160 11992 16166
rect 11940 16102 11992 16108
rect 11756 15684 11808 15690
rect 11756 15626 11808 15632
rect 11664 15616 11716 15622
rect 11664 15558 11716 15564
rect 11676 15078 11704 15558
rect 11768 15078 11796 15626
rect 12688 15622 12716 17831
rect 12860 17802 12912 17808
rect 12768 17724 12820 17730
rect 12768 17666 12820 17672
rect 12780 17254 12808 17666
rect 12872 17254 12900 17802
rect 12964 17798 12992 18890
rect 13056 18818 13084 21610
rect 13136 21600 13188 21606
rect 13136 21542 13188 21548
rect 13148 21130 13176 21542
rect 13136 21124 13188 21130
rect 13136 21066 13188 21072
rect 13148 20586 13176 21066
rect 13136 20580 13188 20586
rect 13136 20522 13188 20528
rect 13700 20518 13728 22562
rect 13976 22286 14004 23718
rect 14528 23306 14556 24806
rect 14804 23918 14832 25418
rect 14896 24938 14924 25418
rect 14988 25414 15016 25758
rect 15724 25618 15752 25826
rect 15712 25612 15764 25618
rect 15712 25554 15764 25560
rect 16736 25414 16764 25826
rect 16908 25816 16960 25822
rect 16908 25758 16960 25764
rect 17000 25816 17052 25822
rect 17000 25758 17052 25764
rect 14976 25408 15028 25414
rect 14976 25350 15028 25356
rect 16264 25408 16316 25414
rect 16264 25350 16316 25356
rect 16724 25408 16776 25414
rect 16724 25350 16776 25356
rect 14884 24932 14936 24938
rect 14884 24874 14936 24880
rect 14896 23986 14924 24874
rect 14884 23980 14936 23986
rect 14884 23922 14936 23928
rect 14792 23912 14844 23918
rect 14792 23854 14844 23860
rect 14700 23844 14752 23850
rect 14700 23786 14752 23792
rect 14516 23300 14568 23306
rect 14516 23242 14568 23248
rect 14116 22996 14412 23016
rect 14172 22994 14196 22996
rect 14252 22994 14276 22996
rect 14332 22994 14356 22996
rect 14194 22942 14196 22994
rect 14258 22942 14270 22994
rect 14332 22942 14334 22994
rect 14172 22940 14196 22942
rect 14252 22940 14276 22942
rect 14332 22940 14356 22942
rect 14116 22920 14412 22940
rect 13964 22280 14016 22286
rect 13964 22222 14016 22228
rect 14116 21908 14412 21928
rect 14172 21906 14196 21908
rect 14252 21906 14276 21908
rect 14332 21906 14356 21908
rect 14194 21854 14196 21906
rect 14258 21854 14270 21906
rect 14332 21854 14334 21906
rect 14172 21852 14196 21854
rect 14252 21852 14276 21854
rect 14332 21852 14356 21854
rect 14116 21832 14412 21852
rect 14528 21742 14556 23242
rect 14712 22626 14740 23786
rect 14804 23442 14832 23854
rect 14792 23436 14844 23442
rect 14792 23378 14844 23384
rect 14804 22694 14832 23378
rect 14896 23306 14924 23922
rect 14988 23714 15016 25350
rect 15804 24864 15856 24870
rect 15802 24832 15804 24841
rect 15856 24832 15858 24841
rect 15620 24796 15672 24802
rect 15802 24767 15858 24776
rect 15620 24738 15672 24744
rect 15252 23844 15304 23850
rect 15252 23786 15304 23792
rect 15068 23776 15120 23782
rect 15068 23718 15120 23724
rect 14976 23708 15028 23714
rect 14976 23650 15028 23656
rect 14884 23300 14936 23306
rect 14884 23242 14936 23248
rect 15080 23238 15108 23718
rect 15068 23232 15120 23238
rect 15068 23174 15120 23180
rect 15080 22898 15108 23174
rect 15264 22898 15292 23786
rect 15632 23646 15660 24738
rect 15988 24524 16040 24530
rect 15988 24466 16040 24472
rect 16000 24326 16028 24466
rect 15988 24320 16040 24326
rect 15988 24262 16040 24268
rect 16172 24320 16224 24326
rect 16276 24274 16304 25350
rect 16724 24932 16776 24938
rect 16920 24920 16948 25758
rect 17012 25550 17040 25758
rect 17196 25618 17224 25894
rect 17564 25890 17592 26506
rect 17748 25958 17776 26506
rect 18024 26026 18052 26574
rect 18472 26496 18524 26502
rect 18472 26438 18524 26444
rect 18288 26428 18340 26434
rect 18288 26370 18340 26376
rect 18300 26042 18328 26370
rect 18012 26020 18064 26026
rect 18012 25962 18064 25968
rect 18116 26014 18328 26042
rect 17736 25952 17788 25958
rect 17736 25894 17788 25900
rect 17276 25884 17328 25890
rect 17276 25826 17328 25832
rect 17552 25884 17604 25890
rect 17552 25826 17604 25832
rect 17184 25612 17236 25618
rect 17184 25554 17236 25560
rect 17000 25544 17052 25550
rect 17000 25486 17052 25492
rect 16776 24892 16948 24920
rect 16724 24874 16776 24880
rect 16736 24530 16764 24874
rect 17012 24818 17040 25486
rect 16816 24796 16868 24802
rect 17012 24790 17132 24818
rect 17196 24802 17224 25554
rect 16816 24738 16868 24744
rect 16724 24524 16776 24530
rect 16724 24466 16776 24472
rect 16828 24394 16856 24738
rect 17000 24728 17052 24734
rect 17000 24670 17052 24676
rect 16816 24388 16868 24394
rect 16816 24330 16868 24336
rect 16224 24268 16304 24274
rect 16172 24262 16304 24268
rect 16184 24246 16304 24262
rect 15988 24184 16040 24190
rect 15988 24126 16040 24132
rect 16172 24184 16224 24190
rect 16172 24126 16224 24132
rect 16000 23918 16028 24126
rect 15988 23912 16040 23918
rect 15988 23854 16040 23860
rect 15620 23640 15672 23646
rect 15620 23582 15672 23588
rect 16000 23374 16028 23854
rect 16184 23714 16212 24126
rect 16172 23708 16224 23714
rect 16172 23650 16224 23656
rect 15988 23368 16040 23374
rect 15988 23310 16040 23316
rect 16184 23306 16212 23650
rect 15436 23300 15488 23306
rect 15436 23242 15488 23248
rect 16172 23300 16224 23306
rect 16172 23242 16224 23248
rect 15068 22892 15120 22898
rect 15068 22834 15120 22840
rect 15252 22892 15304 22898
rect 15252 22834 15304 22840
rect 14792 22688 14844 22694
rect 14792 22630 14844 22636
rect 14700 22620 14752 22626
rect 14700 22562 14752 22568
rect 14804 22218 14832 22630
rect 15080 22286 15108 22834
rect 15264 22694 15292 22834
rect 15448 22762 15476 23242
rect 15436 22756 15488 22762
rect 15436 22698 15488 22704
rect 15252 22688 15304 22694
rect 15252 22630 15304 22636
rect 15068 22280 15120 22286
rect 15068 22222 15120 22228
rect 14792 22212 14844 22218
rect 14792 22154 14844 22160
rect 14516 21736 14568 21742
rect 14516 21678 14568 21684
rect 15080 21674 15108 22222
rect 15264 22218 15292 22630
rect 16184 22626 16212 23242
rect 16276 23238 16304 24246
rect 16828 23714 16856 24330
rect 16816 23708 16868 23714
rect 16816 23650 16868 23656
rect 16264 23232 16316 23238
rect 16264 23174 16316 23180
rect 16540 23232 16592 23238
rect 16540 23174 16592 23180
rect 16172 22620 16224 22626
rect 16172 22562 16224 22568
rect 16276 22218 16304 23174
rect 16448 22552 16500 22558
rect 16448 22494 16500 22500
rect 15252 22212 15304 22218
rect 15252 22154 15304 22160
rect 16264 22212 16316 22218
rect 16264 22154 16316 22160
rect 15804 22008 15856 22014
rect 15804 21950 15856 21956
rect 15068 21668 15120 21674
rect 15068 21610 15120 21616
rect 14516 21600 14568 21606
rect 14516 21542 14568 21548
rect 13872 20920 13924 20926
rect 13872 20862 13924 20868
rect 13884 20518 13912 20862
rect 14116 20820 14412 20840
rect 14172 20818 14196 20820
rect 14252 20818 14276 20820
rect 14332 20818 14356 20820
rect 14194 20766 14196 20818
rect 14258 20766 14270 20818
rect 14332 20766 14334 20818
rect 14172 20764 14196 20766
rect 14252 20764 14276 20766
rect 14332 20764 14356 20766
rect 14116 20744 14412 20764
rect 14528 20654 14556 21542
rect 14516 20648 14568 20654
rect 14516 20590 14568 20596
rect 15080 20586 15108 21610
rect 15528 21600 15580 21606
rect 15528 21542 15580 21548
rect 15436 21532 15488 21538
rect 15436 21474 15488 21480
rect 15252 21464 15304 21470
rect 15252 21406 15304 21412
rect 15264 21198 15292 21406
rect 15252 21192 15304 21198
rect 15252 21134 15304 21140
rect 15252 21056 15304 21062
rect 15252 20998 15304 21004
rect 15068 20580 15120 20586
rect 15068 20522 15120 20528
rect 13688 20512 13740 20518
rect 13688 20454 13740 20460
rect 13872 20512 13924 20518
rect 13872 20454 13924 20460
rect 14608 20512 14660 20518
rect 14608 20454 14660 20460
rect 13700 19430 13728 20454
rect 13884 19498 13912 20454
rect 14424 20444 14476 20450
rect 14424 20386 14476 20392
rect 14436 20042 14464 20386
rect 14620 20042 14648 20454
rect 14884 20444 14936 20450
rect 14884 20386 14936 20392
rect 14424 20036 14476 20042
rect 14608 20036 14660 20042
rect 14476 19996 14556 20024
rect 14424 19978 14476 19984
rect 14116 19732 14412 19752
rect 14172 19730 14196 19732
rect 14252 19730 14276 19732
rect 14332 19730 14356 19732
rect 14194 19678 14196 19730
rect 14258 19678 14270 19730
rect 14332 19678 14334 19730
rect 14172 19676 14196 19678
rect 14252 19676 14276 19678
rect 14332 19676 14356 19678
rect 14116 19656 14412 19676
rect 13872 19492 13924 19498
rect 13872 19434 13924 19440
rect 13688 19424 13740 19430
rect 13964 19424 14016 19430
rect 13688 19366 13740 19372
rect 13884 19372 13964 19378
rect 13884 19366 14016 19372
rect 13884 19350 14004 19366
rect 14528 19362 14556 19996
rect 14608 19978 14660 19984
rect 14620 19498 14648 19978
rect 14700 19968 14752 19974
rect 14700 19910 14752 19916
rect 14608 19492 14660 19498
rect 14608 19434 14660 19440
rect 14516 19356 14568 19362
rect 13884 19090 13912 19350
rect 14516 19298 14568 19304
rect 13872 19084 13924 19090
rect 13872 19026 13924 19032
rect 13320 18880 13372 18886
rect 13320 18822 13372 18828
rect 13044 18812 13096 18818
rect 13044 18754 13096 18760
rect 13056 17866 13084 18754
rect 13332 18410 13360 18822
rect 13320 18404 13372 18410
rect 13320 18346 13372 18352
rect 13044 17860 13096 17866
rect 13044 17802 13096 17808
rect 12952 17792 13004 17798
rect 12952 17734 13004 17740
rect 12964 17322 12992 17734
rect 13332 17662 13360 18346
rect 13884 18342 13912 19026
rect 14712 18954 14740 19910
rect 14896 18954 14924 20386
rect 15080 19294 15108 20522
rect 15264 19498 15292 20998
rect 15448 20722 15476 21474
rect 15540 21198 15568 21542
rect 15528 21192 15580 21198
rect 15528 21134 15580 21140
rect 15436 20716 15488 20722
rect 15436 20658 15488 20664
rect 15712 20648 15764 20654
rect 15712 20590 15764 20596
rect 15724 19906 15752 20590
rect 15816 20110 15844 21950
rect 16276 21130 16304 22154
rect 16460 21130 16488 22494
rect 16264 21124 16316 21130
rect 16264 21066 16316 21072
rect 16448 21124 16500 21130
rect 16448 21066 16500 21072
rect 15804 20104 15856 20110
rect 15804 20046 15856 20052
rect 16276 19906 16304 21066
rect 16460 20178 16488 21066
rect 16448 20172 16500 20178
rect 16448 20114 16500 20120
rect 15712 19900 15764 19906
rect 15712 19842 15764 19848
rect 15896 19900 15948 19906
rect 15896 19842 15948 19848
rect 16264 19900 16316 19906
rect 16264 19842 16316 19848
rect 15252 19492 15304 19498
rect 15252 19434 15304 19440
rect 15068 19288 15120 19294
rect 15068 19230 15120 19236
rect 15264 18954 15292 19434
rect 15344 19288 15396 19294
rect 15344 19230 15396 19236
rect 14700 18948 14752 18954
rect 14700 18890 14752 18896
rect 14884 18948 14936 18954
rect 14884 18890 14936 18896
rect 15068 18948 15120 18954
rect 15068 18890 15120 18896
rect 15252 18948 15304 18954
rect 15252 18890 15304 18896
rect 14116 18644 14412 18664
rect 14172 18642 14196 18644
rect 14252 18642 14276 18644
rect 14332 18642 14356 18644
rect 14194 18590 14196 18642
rect 14258 18590 14270 18642
rect 14332 18590 14334 18642
rect 14172 18588 14196 18590
rect 14252 18588 14276 18590
rect 14332 18588 14356 18590
rect 14116 18568 14412 18588
rect 15080 18478 15108 18890
rect 15068 18472 15120 18478
rect 15068 18414 15120 18420
rect 13872 18336 13924 18342
rect 13872 18278 13924 18284
rect 14608 18336 14660 18342
rect 14608 18278 14660 18284
rect 13320 17656 13372 17662
rect 13320 17598 13372 17604
rect 13332 17458 13360 17598
rect 13320 17452 13372 17458
rect 13320 17394 13372 17400
rect 12952 17316 13004 17322
rect 12952 17258 13004 17264
rect 12768 17248 12820 17254
rect 12768 17190 12820 17196
rect 12860 17248 12912 17254
rect 12860 17190 12912 17196
rect 13320 17248 13372 17254
rect 13320 17190 13372 17196
rect 13332 16846 13360 17190
rect 13320 16840 13372 16846
rect 13320 16782 13372 16788
rect 12952 16772 13004 16778
rect 12952 16714 13004 16720
rect 12676 15616 12728 15622
rect 12676 15558 12728 15564
rect 12032 15480 12084 15486
rect 12032 15422 12084 15428
rect 11940 15140 11992 15146
rect 11940 15082 11992 15088
rect 11664 15072 11716 15078
rect 11664 15014 11716 15020
rect 11756 15072 11808 15078
rect 11756 15014 11808 15020
rect 11952 14602 11980 15082
rect 11940 14596 11992 14602
rect 11940 14538 11992 14544
rect 12044 14534 12072 15422
rect 12964 15146 12992 16714
rect 13780 16160 13832 16166
rect 13780 16102 13832 16108
rect 13044 15684 13096 15690
rect 13044 15626 13096 15632
rect 12952 15140 13004 15146
rect 12952 15082 13004 15088
rect 12952 14596 13004 14602
rect 12952 14538 13004 14544
rect 12032 14528 12084 14534
rect 12032 14470 12084 14476
rect 12400 14528 12452 14534
rect 12400 14470 12452 14476
rect 11572 14460 11624 14466
rect 11572 14402 11624 14408
rect 11584 13990 11612 14402
rect 11572 13984 11624 13990
rect 11572 13926 11624 13932
rect 11584 12018 11612 13926
rect 12044 13514 12072 14470
rect 12412 14058 12440 14470
rect 12964 14466 12992 14538
rect 12952 14460 13004 14466
rect 12952 14402 13004 14408
rect 12768 14392 12820 14398
rect 12768 14334 12820 14340
rect 12400 14052 12452 14058
rect 12400 13994 12452 14000
rect 12780 13990 12808 14334
rect 13056 14194 13084 15626
rect 13228 15480 13280 15486
rect 13228 15422 13280 15428
rect 13240 15146 13268 15422
rect 13228 15140 13280 15146
rect 13228 15082 13280 15088
rect 13792 14602 13820 16102
rect 13780 14596 13832 14602
rect 13780 14538 13832 14544
rect 13884 14194 13912 18278
rect 13964 18200 14016 18206
rect 13964 18142 14016 18148
rect 14516 18200 14568 18206
rect 14516 18142 14568 18148
rect 13976 17934 14004 18142
rect 13964 17928 14016 17934
rect 13964 17870 14016 17876
rect 14116 17556 14412 17576
rect 14172 17554 14196 17556
rect 14252 17554 14276 17556
rect 14332 17554 14356 17556
rect 14194 17502 14196 17554
rect 14258 17502 14270 17554
rect 14332 17502 14334 17554
rect 14172 17500 14196 17502
rect 14252 17500 14276 17502
rect 14332 17500 14356 17502
rect 14116 17480 14412 17500
rect 14528 16846 14556 18142
rect 14620 17322 14648 18278
rect 14976 17724 15028 17730
rect 14976 17666 15028 17672
rect 14988 17322 15016 17666
rect 15080 17322 15108 18414
rect 15356 18206 15384 19230
rect 15908 18478 15936 19842
rect 16080 19832 16132 19838
rect 16080 19774 16132 19780
rect 16092 19430 16120 19774
rect 16080 19424 16132 19430
rect 16080 19366 16132 19372
rect 16448 18880 16500 18886
rect 16448 18822 16500 18828
rect 15896 18472 15948 18478
rect 15896 18414 15948 18420
rect 15436 18268 15488 18274
rect 15436 18210 15488 18216
rect 15344 18200 15396 18206
rect 15344 18142 15396 18148
rect 15356 17866 15384 18142
rect 15448 17934 15476 18210
rect 15436 17928 15488 17934
rect 15436 17870 15488 17876
rect 15344 17860 15396 17866
rect 15344 17802 15396 17808
rect 15448 17322 15476 17870
rect 14608 17316 14660 17322
rect 14608 17258 14660 17264
rect 14976 17316 15028 17322
rect 14976 17258 15028 17264
rect 15068 17316 15120 17322
rect 15068 17258 15120 17264
rect 15436 17316 15488 17322
rect 15436 17258 15488 17264
rect 14516 16840 14568 16846
rect 14516 16782 14568 16788
rect 14700 16840 14752 16846
rect 14700 16782 14752 16788
rect 14116 16468 14412 16488
rect 14172 16466 14196 16468
rect 14252 16466 14276 16468
rect 14332 16466 14356 16468
rect 14194 16414 14196 16466
rect 14258 16414 14270 16466
rect 14332 16414 14334 16466
rect 14172 16412 14196 16414
rect 14252 16412 14276 16414
rect 14332 16412 14356 16414
rect 14116 16392 14412 16412
rect 14712 16370 14740 16782
rect 14988 16710 15016 17258
rect 14976 16704 15028 16710
rect 14976 16646 15028 16652
rect 14700 16364 14752 16370
rect 14700 16306 14752 16312
rect 14988 16166 15016 16646
rect 15448 16370 15476 17258
rect 16460 16914 16488 18822
rect 16552 18002 16580 23174
rect 16632 22892 16684 22898
rect 16632 22834 16684 22840
rect 16644 22694 16672 22834
rect 16632 22688 16684 22694
rect 16632 22630 16684 22636
rect 16828 22014 16856 23650
rect 17012 23374 17040 24670
rect 17104 23442 17132 24790
rect 17184 24796 17236 24802
rect 17184 24738 17236 24744
rect 17196 23918 17224 24738
rect 17288 24394 17316 25826
rect 17564 25414 17592 25826
rect 18116 25822 18144 26014
rect 18196 25952 18248 25958
rect 18196 25894 18248 25900
rect 18104 25816 18156 25822
rect 18104 25758 18156 25764
rect 17552 25408 17604 25414
rect 17552 25350 17604 25356
rect 17564 25006 17592 25350
rect 17552 25000 17604 25006
rect 17552 24942 17604 24948
rect 17564 24734 17592 24942
rect 18104 24796 18156 24802
rect 18104 24738 18156 24744
rect 17368 24728 17420 24734
rect 17368 24670 17420 24676
rect 17552 24728 17604 24734
rect 17552 24670 17604 24676
rect 17276 24388 17328 24394
rect 17276 24330 17328 24336
rect 17184 23912 17236 23918
rect 17184 23854 17236 23860
rect 17380 23782 17408 24670
rect 17564 23918 17592 24670
rect 18012 24524 18064 24530
rect 18012 24466 18064 24472
rect 17552 23912 17604 23918
rect 17552 23854 17604 23860
rect 17368 23776 17420 23782
rect 17368 23718 17420 23724
rect 17092 23436 17144 23442
rect 17092 23378 17144 23384
rect 17000 23368 17052 23374
rect 17000 23310 17052 23316
rect 17092 23300 17144 23306
rect 17092 23242 17144 23248
rect 17000 22756 17052 22762
rect 16920 22716 17000 22744
rect 16816 22008 16868 22014
rect 16816 21950 16868 21956
rect 16828 21742 16856 21950
rect 16816 21736 16868 21742
rect 16816 21678 16868 21684
rect 16920 21130 16948 22716
rect 17000 22698 17052 22704
rect 17104 22694 17132 23242
rect 17564 23102 17592 23854
rect 18024 23306 18052 24466
rect 18012 23300 18064 23306
rect 18012 23242 18064 23248
rect 17552 23096 17604 23102
rect 17552 23038 17604 23044
rect 17092 22688 17144 22694
rect 17092 22630 17144 22636
rect 18012 22688 18064 22694
rect 18012 22630 18064 22636
rect 17000 22280 17052 22286
rect 17000 22222 17052 22228
rect 17012 21810 17040 22222
rect 17000 21804 17052 21810
rect 17000 21746 17052 21752
rect 17104 21266 17132 22630
rect 17276 22620 17328 22626
rect 17276 22562 17328 22568
rect 17184 22144 17236 22150
rect 17184 22086 17236 22092
rect 17092 21260 17144 21266
rect 17092 21202 17144 21208
rect 17196 21130 17224 22086
rect 17288 21470 17316 22562
rect 18024 21810 18052 22630
rect 18116 22626 18144 24738
rect 18208 24462 18236 25894
rect 18300 24938 18328 26014
rect 18380 25816 18432 25822
rect 18380 25758 18432 25764
rect 18484 25770 18512 26438
rect 18564 26020 18616 26026
rect 18616 25980 18696 26008
rect 18564 25962 18616 25968
rect 18392 25482 18420 25758
rect 18484 25742 18604 25770
rect 18380 25476 18432 25482
rect 18380 25418 18432 25424
rect 18472 25476 18524 25482
rect 18472 25418 18524 25424
rect 18288 24932 18340 24938
rect 18288 24874 18340 24880
rect 18196 24456 18248 24462
rect 18196 24398 18248 24404
rect 18196 24184 18248 24190
rect 18196 24126 18248 24132
rect 18208 23442 18236 24126
rect 18300 23850 18328 24874
rect 18392 24462 18420 25418
rect 18380 24456 18432 24462
rect 18380 24398 18432 24404
rect 18484 24190 18512 25418
rect 18576 25414 18604 25742
rect 18564 25408 18616 25414
rect 18564 25350 18616 25356
rect 18564 25068 18616 25074
rect 18564 25010 18616 25016
rect 18576 24258 18604 25010
rect 18564 24252 18616 24258
rect 18564 24194 18616 24200
rect 18668 24190 18696 25980
rect 18852 25618 18880 27662
rect 19024 27652 19076 27658
rect 19024 27594 19076 27600
rect 19036 27114 19064 27594
rect 19392 27584 19444 27590
rect 19392 27526 19444 27532
rect 19404 27182 19432 27526
rect 19392 27176 19444 27182
rect 19392 27118 19444 27124
rect 19024 27108 19076 27114
rect 19024 27050 19076 27056
rect 19036 26978 19064 27050
rect 18932 26972 18984 26978
rect 18932 26914 18984 26920
rect 19024 26972 19076 26978
rect 19024 26914 19076 26920
rect 18944 26570 18972 26914
rect 19496 26910 19524 27662
rect 19680 27454 19708 28478
rect 19772 28202 19800 29294
rect 19864 29154 19892 29770
rect 20036 29216 20088 29222
rect 20036 29158 20088 29164
rect 19852 29148 19904 29154
rect 19852 29090 19904 29096
rect 19864 28218 19892 29090
rect 19760 28196 19812 28202
rect 19864 28190 19984 28218
rect 19760 28138 19812 28144
rect 19956 28134 19984 28190
rect 19944 28128 19996 28134
rect 19944 28070 19996 28076
rect 20048 28066 20076 29158
rect 20232 28542 20260 31576
rect 21140 29760 21192 29766
rect 21140 29702 21192 29708
rect 21152 29290 21180 29702
rect 21968 29692 22020 29698
rect 21968 29634 22020 29640
rect 21324 29420 21376 29426
rect 21324 29362 21376 29368
rect 21140 29284 21192 29290
rect 21140 29226 21192 29232
rect 20680 29216 20732 29222
rect 20680 29158 20732 29164
rect 20692 28882 20720 29158
rect 20680 28876 20732 28882
rect 20680 28818 20732 28824
rect 20312 28740 20364 28746
rect 20312 28682 20364 28688
rect 20220 28536 20272 28542
rect 20220 28478 20272 28484
rect 20036 28060 20088 28066
rect 20036 28002 20088 28008
rect 19760 27652 19812 27658
rect 19760 27594 19812 27600
rect 19576 27448 19628 27454
rect 19576 27390 19628 27396
rect 19668 27448 19720 27454
rect 19668 27390 19720 27396
rect 19588 27046 19616 27390
rect 19680 27250 19708 27390
rect 19668 27244 19720 27250
rect 19668 27186 19720 27192
rect 19576 27040 19628 27046
rect 19576 26982 19628 26988
rect 19484 26904 19536 26910
rect 19484 26846 19536 26852
rect 19116 26804 19412 26824
rect 19172 26802 19196 26804
rect 19252 26802 19276 26804
rect 19332 26802 19356 26804
rect 19194 26750 19196 26802
rect 19258 26750 19270 26802
rect 19332 26750 19334 26802
rect 19172 26748 19196 26750
rect 19252 26748 19276 26750
rect 19332 26748 19356 26750
rect 19116 26728 19412 26748
rect 19496 26570 19524 26846
rect 18932 26564 18984 26570
rect 18932 26506 18984 26512
rect 19484 26564 19536 26570
rect 19484 26506 19536 26512
rect 18932 25952 18984 25958
rect 18932 25894 18984 25900
rect 18840 25612 18892 25618
rect 18840 25554 18892 25560
rect 18840 25340 18892 25346
rect 18840 25282 18892 25288
rect 18852 24802 18880 25282
rect 18944 24938 18972 25894
rect 19024 25884 19076 25890
rect 19024 25826 19076 25832
rect 18932 24932 18984 24938
rect 18932 24874 18984 24880
rect 19036 24841 19064 25826
rect 19116 25716 19412 25736
rect 19172 25714 19196 25716
rect 19252 25714 19276 25716
rect 19332 25714 19356 25716
rect 19194 25662 19196 25714
rect 19258 25662 19270 25714
rect 19332 25662 19334 25714
rect 19172 25660 19196 25662
rect 19252 25660 19276 25662
rect 19332 25660 19356 25662
rect 19116 25640 19412 25660
rect 19496 25414 19524 26506
rect 19772 25618 19800 27594
rect 20048 27182 20076 28002
rect 20324 27726 20352 28682
rect 20692 28338 20720 28818
rect 21152 28746 21180 29226
rect 21140 28740 21192 28746
rect 21140 28682 21192 28688
rect 20772 28536 20824 28542
rect 20772 28478 20824 28484
rect 20680 28332 20732 28338
rect 20680 28274 20732 28280
rect 20588 28060 20640 28066
rect 20588 28002 20640 28008
rect 20496 27992 20548 27998
rect 20496 27934 20548 27940
rect 20508 27794 20536 27934
rect 20496 27788 20548 27794
rect 20496 27730 20548 27736
rect 20312 27720 20364 27726
rect 20312 27662 20364 27668
rect 20036 27176 20088 27182
rect 20036 27118 20088 27124
rect 20600 27114 20628 28002
rect 20680 27584 20732 27590
rect 20680 27526 20732 27532
rect 20588 27108 20640 27114
rect 20588 27050 20640 27056
rect 19944 27040 19996 27046
rect 19944 26982 19996 26988
rect 20220 27040 20272 27046
rect 20220 26982 20272 26988
rect 19956 26638 19984 26982
rect 19944 26632 19996 26638
rect 19944 26574 19996 26580
rect 19944 26496 19996 26502
rect 19944 26438 19996 26444
rect 19760 25612 19812 25618
rect 19760 25554 19812 25560
rect 19852 25476 19904 25482
rect 19852 25418 19904 25424
rect 19484 25408 19536 25414
rect 19484 25350 19536 25356
rect 19496 24938 19524 25350
rect 19484 24932 19536 24938
rect 19484 24874 19536 24880
rect 19022 24832 19078 24841
rect 18840 24796 18892 24802
rect 19022 24767 19078 24776
rect 19760 24796 19812 24802
rect 18840 24738 18892 24744
rect 18472 24184 18524 24190
rect 18472 24126 18524 24132
rect 18656 24184 18708 24190
rect 18656 24126 18708 24132
rect 18288 23844 18340 23850
rect 18288 23786 18340 23792
rect 18668 23782 18696 24126
rect 18748 23912 18800 23918
rect 18748 23854 18800 23860
rect 18656 23776 18708 23782
rect 18656 23718 18708 23724
rect 18196 23436 18248 23442
rect 18196 23378 18248 23384
rect 18380 23300 18432 23306
rect 18380 23242 18432 23248
rect 18196 23096 18248 23102
rect 18196 23038 18248 23044
rect 18104 22620 18156 22626
rect 18104 22562 18156 22568
rect 18116 22218 18144 22562
rect 18104 22212 18156 22218
rect 18104 22154 18156 22160
rect 18012 21804 18064 21810
rect 18012 21746 18064 21752
rect 18116 21606 18144 22154
rect 17828 21600 17880 21606
rect 17828 21542 17880 21548
rect 18104 21600 18156 21606
rect 18104 21542 18156 21548
rect 17736 21532 17788 21538
rect 17736 21474 17788 21480
rect 17276 21464 17328 21470
rect 17276 21406 17328 21412
rect 16908 21124 16960 21130
rect 16908 21066 16960 21072
rect 17184 21124 17236 21130
rect 17184 21066 17236 21072
rect 17196 20994 17224 21066
rect 17184 20988 17236 20994
rect 17184 20930 17236 20936
rect 17552 20988 17604 20994
rect 17552 20930 17604 20936
rect 17564 20110 17592 20930
rect 17748 20926 17776 21474
rect 17840 21198 17868 21542
rect 17828 21192 17880 21198
rect 18116 21146 18144 21542
rect 17828 21134 17880 21140
rect 17736 20920 17788 20926
rect 17736 20862 17788 20868
rect 17000 20104 17052 20110
rect 17000 20046 17052 20052
rect 17552 20104 17604 20110
rect 17552 20046 17604 20052
rect 16724 19832 16776 19838
rect 16724 19774 16776 19780
rect 16736 19430 16764 19774
rect 16724 19424 16776 19430
rect 16724 19366 16776 19372
rect 16816 19288 16868 19294
rect 16816 19230 16868 19236
rect 16828 18002 16856 19230
rect 16908 18744 16960 18750
rect 16908 18686 16960 18692
rect 16920 18002 16948 18686
rect 17012 18342 17040 20046
rect 17748 20042 17776 20862
rect 17840 20110 17868 21134
rect 18024 21118 18144 21146
rect 18024 20586 18052 21118
rect 18104 21056 18156 21062
rect 18104 20998 18156 21004
rect 18012 20580 18064 20586
rect 18012 20522 18064 20528
rect 17828 20104 17880 20110
rect 17828 20046 17880 20052
rect 17184 20036 17236 20042
rect 17184 19978 17236 19984
rect 17736 20036 17788 20042
rect 17736 19978 17788 19984
rect 17196 19566 17224 19978
rect 17184 19560 17236 19566
rect 17184 19502 17236 19508
rect 17196 19430 17224 19502
rect 17840 19498 17868 20046
rect 18024 19974 18052 20522
rect 18116 20518 18144 20998
rect 18104 20512 18156 20518
rect 18104 20454 18156 20460
rect 18208 20178 18236 23038
rect 18392 22762 18420 23242
rect 18760 22762 18788 23854
rect 19036 23850 19064 24767
rect 19760 24738 19812 24744
rect 19668 24728 19720 24734
rect 19668 24670 19720 24676
rect 19116 24628 19412 24648
rect 19172 24626 19196 24628
rect 19252 24626 19276 24628
rect 19332 24626 19356 24628
rect 19194 24574 19196 24626
rect 19258 24574 19270 24626
rect 19332 24574 19334 24626
rect 19172 24572 19196 24574
rect 19252 24572 19276 24574
rect 19332 24572 19356 24574
rect 19116 24552 19412 24572
rect 19680 24530 19708 24670
rect 19668 24524 19720 24530
rect 19668 24466 19720 24472
rect 19772 24394 19800 24738
rect 19864 24734 19892 25418
rect 19852 24728 19904 24734
rect 19852 24670 19904 24676
rect 19760 24388 19812 24394
rect 19760 24330 19812 24336
rect 19668 24320 19720 24326
rect 19668 24262 19720 24268
rect 19024 23844 19076 23850
rect 19024 23786 19076 23792
rect 19484 23708 19536 23714
rect 19484 23650 19536 23656
rect 19116 23540 19412 23560
rect 19172 23538 19196 23540
rect 19252 23538 19276 23540
rect 19332 23538 19356 23540
rect 19194 23486 19196 23538
rect 19258 23486 19270 23538
rect 19332 23486 19334 23538
rect 19172 23484 19196 23486
rect 19252 23484 19276 23486
rect 19332 23484 19356 23486
rect 19116 23464 19412 23484
rect 19300 23096 19352 23102
rect 19300 23038 19352 23044
rect 18380 22756 18432 22762
rect 18380 22698 18432 22704
rect 18748 22756 18800 22762
rect 18748 22698 18800 22704
rect 18392 22218 18420 22698
rect 18380 22212 18432 22218
rect 18380 22154 18432 22160
rect 18760 21674 18788 22698
rect 19312 22694 19340 23038
rect 19496 22762 19524 23650
rect 19576 23640 19628 23646
rect 19576 23582 19628 23588
rect 19588 23306 19616 23582
rect 19680 23442 19708 24262
rect 19668 23436 19720 23442
rect 19668 23378 19720 23384
rect 19576 23300 19628 23306
rect 19576 23242 19628 23248
rect 19680 22898 19708 23378
rect 19760 23232 19812 23238
rect 19760 23174 19812 23180
rect 19772 23102 19800 23174
rect 19760 23096 19812 23102
rect 19760 23038 19812 23044
rect 19668 22892 19720 22898
rect 19668 22834 19720 22840
rect 19484 22756 19536 22762
rect 19484 22698 19536 22704
rect 19300 22688 19352 22694
rect 19300 22630 19352 22636
rect 19116 22452 19412 22472
rect 19172 22450 19196 22452
rect 19252 22450 19276 22452
rect 19332 22450 19356 22452
rect 19194 22398 19196 22450
rect 19258 22398 19270 22450
rect 19332 22398 19334 22450
rect 19172 22396 19196 22398
rect 19252 22396 19276 22398
rect 19332 22396 19356 22398
rect 19116 22376 19412 22396
rect 19772 22218 19800 23038
rect 19760 22212 19812 22218
rect 19760 22154 19812 22160
rect 19576 21804 19628 21810
rect 19576 21746 19628 21752
rect 18748 21668 18800 21674
rect 18748 21610 18800 21616
rect 19024 21668 19076 21674
rect 19024 21610 19076 21616
rect 18564 21464 18616 21470
rect 18564 21406 18616 21412
rect 18576 21130 18604 21406
rect 18564 21124 18616 21130
rect 18564 21066 18616 21072
rect 18196 20172 18248 20178
rect 18196 20114 18248 20120
rect 18208 20081 18236 20114
rect 18194 20072 18250 20081
rect 18194 20007 18250 20016
rect 18012 19968 18064 19974
rect 18012 19910 18064 19916
rect 17828 19492 17880 19498
rect 17828 19434 17880 19440
rect 17184 19424 17236 19430
rect 17184 19366 17236 19372
rect 17460 19016 17512 19022
rect 17460 18958 17512 18964
rect 17472 18478 17500 18958
rect 18576 18750 18604 21066
rect 19036 21062 19064 21610
rect 19116 21364 19412 21384
rect 19172 21362 19196 21364
rect 19252 21362 19276 21364
rect 19332 21362 19356 21364
rect 19194 21310 19196 21362
rect 19258 21310 19270 21362
rect 19332 21310 19334 21362
rect 19172 21308 19196 21310
rect 19252 21308 19276 21310
rect 19332 21308 19356 21310
rect 19116 21288 19412 21308
rect 19588 21198 19616 21746
rect 19864 21266 19892 24670
rect 19956 23238 19984 26438
rect 20232 25550 20260 26982
rect 20312 26904 20364 26910
rect 20312 26846 20364 26852
rect 20404 26904 20456 26910
rect 20404 26846 20456 26852
rect 20324 26706 20352 26846
rect 20312 26700 20364 26706
rect 20312 26642 20364 26648
rect 20416 26638 20444 26846
rect 20692 26638 20720 27526
rect 20404 26632 20456 26638
rect 20404 26574 20456 26580
rect 20680 26632 20732 26638
rect 20680 26574 20732 26580
rect 20588 25884 20640 25890
rect 20588 25826 20640 25832
rect 20220 25544 20272 25550
rect 20220 25486 20272 25492
rect 20232 24546 20260 25486
rect 20404 25408 20456 25414
rect 20404 25350 20456 25356
rect 20416 25006 20444 25350
rect 20404 25000 20456 25006
rect 20404 24942 20456 24948
rect 20600 24802 20628 25826
rect 20588 24796 20640 24802
rect 20588 24738 20640 24744
rect 20048 24518 20260 24546
rect 20048 23306 20076 24518
rect 20128 24388 20180 24394
rect 20128 24330 20180 24336
rect 20140 23782 20168 24330
rect 20128 23776 20180 23782
rect 20128 23718 20180 23724
rect 20036 23300 20088 23306
rect 20036 23242 20088 23248
rect 19944 23232 19996 23238
rect 19944 23174 19996 23180
rect 20048 21742 20076 23242
rect 20140 22830 20168 23718
rect 20692 23238 20720 26574
rect 20404 23232 20456 23238
rect 20404 23174 20456 23180
rect 20496 23232 20548 23238
rect 20496 23174 20548 23180
rect 20680 23232 20732 23238
rect 20680 23174 20732 23180
rect 20128 22824 20180 22830
rect 20128 22766 20180 22772
rect 20416 22762 20444 23174
rect 20404 22756 20456 22762
rect 20404 22698 20456 22704
rect 20220 22688 20272 22694
rect 20220 22630 20272 22636
rect 20232 22286 20260 22630
rect 20220 22280 20272 22286
rect 20220 22222 20272 22228
rect 20416 22150 20444 22698
rect 20508 22218 20536 23174
rect 20692 22354 20720 23174
rect 20680 22348 20732 22354
rect 20680 22290 20732 22296
rect 20496 22212 20548 22218
rect 20496 22154 20548 22160
rect 20404 22144 20456 22150
rect 20404 22086 20456 22092
rect 20036 21736 20088 21742
rect 20036 21678 20088 21684
rect 20404 21600 20456 21606
rect 20404 21542 20456 21548
rect 20220 21532 20272 21538
rect 20220 21474 20272 21480
rect 19852 21260 19904 21266
rect 19852 21202 19904 21208
rect 19576 21192 19628 21198
rect 19576 21134 19628 21140
rect 19668 21192 19720 21198
rect 19668 21134 19720 21140
rect 19024 21056 19076 21062
rect 19024 20998 19076 21004
rect 19680 20654 19708 21134
rect 19668 20648 19720 20654
rect 19668 20590 19720 20596
rect 18932 20444 18984 20450
rect 18932 20386 18984 20392
rect 19668 20444 19720 20450
rect 19668 20386 19720 20392
rect 18944 20110 18972 20386
rect 19116 20276 19412 20296
rect 19172 20274 19196 20276
rect 19252 20274 19276 20276
rect 19332 20274 19356 20276
rect 19194 20222 19196 20274
rect 19258 20222 19270 20274
rect 19332 20222 19334 20274
rect 19172 20220 19196 20222
rect 19252 20220 19276 20222
rect 19332 20220 19356 20222
rect 19116 20200 19412 20220
rect 18932 20104 18984 20110
rect 18932 20046 18984 20052
rect 19208 20104 19260 20110
rect 19208 20046 19260 20052
rect 18932 19900 18984 19906
rect 18932 19842 18984 19848
rect 18944 19498 18972 19842
rect 18932 19492 18984 19498
rect 18932 19434 18984 19440
rect 19220 19430 19248 20046
rect 19680 19498 19708 20386
rect 19760 20376 19812 20382
rect 19760 20318 19812 20324
rect 19772 20110 19800 20318
rect 19864 20178 19892 21202
rect 20232 21130 20260 21474
rect 20416 21130 20444 21542
rect 20220 21124 20272 21130
rect 20220 21066 20272 21072
rect 20404 21124 20456 21130
rect 20404 21066 20456 21072
rect 20128 21056 20180 21062
rect 20128 20998 20180 21004
rect 19944 20920 19996 20926
rect 19944 20862 19996 20868
rect 19956 20518 19984 20862
rect 20140 20722 20168 20998
rect 20416 20994 20444 21066
rect 20404 20988 20456 20994
rect 20404 20930 20456 20936
rect 20128 20716 20180 20722
rect 20128 20658 20180 20664
rect 20404 20648 20456 20654
rect 20404 20590 20456 20596
rect 19944 20512 19996 20518
rect 19944 20454 19996 20460
rect 20220 20512 20272 20518
rect 20220 20454 20272 20460
rect 20232 20382 20260 20454
rect 20220 20376 20272 20382
rect 20220 20318 20272 20324
rect 19852 20172 19904 20178
rect 19852 20114 19904 20120
rect 19760 20104 19812 20110
rect 19944 20104 19996 20110
rect 19760 20046 19812 20052
rect 19942 20072 19944 20081
rect 19996 20072 19998 20081
rect 19668 19492 19720 19498
rect 19668 19434 19720 19440
rect 19208 19424 19260 19430
rect 19208 19366 19260 19372
rect 19484 19424 19536 19430
rect 19484 19366 19536 19372
rect 19024 19288 19076 19294
rect 19024 19230 19076 19236
rect 19036 18750 19064 19230
rect 19116 19188 19412 19208
rect 19172 19186 19196 19188
rect 19252 19186 19276 19188
rect 19332 19186 19356 19188
rect 19194 19134 19196 19186
rect 19258 19134 19270 19186
rect 19332 19134 19334 19186
rect 19172 19132 19196 19134
rect 19252 19132 19276 19134
rect 19332 19132 19356 19134
rect 19116 19112 19412 19132
rect 19496 18886 19524 19366
rect 19772 19362 19800 20046
rect 19942 20007 19998 20016
rect 19956 19566 19984 20007
rect 20416 19974 20444 20590
rect 20220 19968 20272 19974
rect 20220 19910 20272 19916
rect 20404 19968 20456 19974
rect 20404 19910 20456 19916
rect 19944 19560 19996 19566
rect 19944 19502 19996 19508
rect 20232 19430 20260 19910
rect 20220 19424 20272 19430
rect 20220 19366 20272 19372
rect 19760 19356 19812 19362
rect 19760 19298 19812 19304
rect 19772 19022 19800 19298
rect 19760 19016 19812 19022
rect 19760 18958 19812 18964
rect 20232 18886 20260 19366
rect 20312 19288 20364 19294
rect 20312 19230 20364 19236
rect 20324 19090 20352 19230
rect 20312 19084 20364 19090
rect 20312 19026 20364 19032
rect 19484 18880 19536 18886
rect 19484 18822 19536 18828
rect 20220 18880 20272 18886
rect 20220 18822 20272 18828
rect 18564 18744 18616 18750
rect 18564 18686 18616 18692
rect 19024 18744 19076 18750
rect 19024 18686 19076 18692
rect 17460 18472 17512 18478
rect 17460 18414 17512 18420
rect 18576 18410 18604 18686
rect 18564 18404 18616 18410
rect 18564 18346 18616 18352
rect 19496 18342 19524 18822
rect 17000 18336 17052 18342
rect 17000 18278 17052 18284
rect 17920 18336 17972 18342
rect 17920 18278 17972 18284
rect 18656 18336 18708 18342
rect 18656 18278 18708 18284
rect 18840 18336 18892 18342
rect 18840 18278 18892 18284
rect 19484 18336 19536 18342
rect 19484 18278 19536 18284
rect 16540 17996 16592 18002
rect 16540 17938 16592 17944
rect 16816 17996 16868 18002
rect 16816 17938 16868 17944
rect 16908 17996 16960 18002
rect 16908 17938 16960 17944
rect 17932 17934 17960 18278
rect 17920 17928 17972 17934
rect 17920 17870 17972 17876
rect 16816 17860 16868 17866
rect 16816 17802 16868 17808
rect 16724 17792 16776 17798
rect 16724 17734 16776 17740
rect 16736 17254 16764 17734
rect 16724 17248 16776 17254
rect 16724 17190 16776 17196
rect 16828 17186 16856 17802
rect 17932 17254 17960 17870
rect 17000 17248 17052 17254
rect 17000 17190 17052 17196
rect 17920 17248 17972 17254
rect 17920 17190 17972 17196
rect 16816 17180 16868 17186
rect 16816 17122 16868 17128
rect 16448 16908 16500 16914
rect 16448 16850 16500 16856
rect 17012 16370 17040 17190
rect 17644 16908 17696 16914
rect 17644 16850 17696 16856
rect 17184 16568 17236 16574
rect 17184 16510 17236 16516
rect 15436 16364 15488 16370
rect 15436 16306 15488 16312
rect 17000 16364 17052 16370
rect 17000 16306 17052 16312
rect 17196 16166 17224 16510
rect 17656 16250 17684 16850
rect 17932 16370 17960 17190
rect 18104 17112 18156 17118
rect 18104 17054 18156 17060
rect 18116 16778 18144 17054
rect 18104 16772 18156 16778
rect 18104 16714 18156 16720
rect 18012 16704 18064 16710
rect 18012 16646 18064 16652
rect 17920 16364 17972 16370
rect 17920 16306 17972 16312
rect 17564 16222 17684 16250
rect 14976 16160 15028 16166
rect 14976 16102 15028 16108
rect 17184 16160 17236 16166
rect 17184 16102 17236 16108
rect 14884 16092 14936 16098
rect 14884 16034 14936 16040
rect 14792 15684 14844 15690
rect 14792 15626 14844 15632
rect 14700 15548 14752 15554
rect 14700 15490 14752 15496
rect 14116 15380 14412 15400
rect 14172 15378 14196 15380
rect 14252 15378 14276 15380
rect 14332 15378 14356 15380
rect 14194 15326 14196 15378
rect 14258 15326 14270 15378
rect 14332 15326 14334 15378
rect 14172 15324 14196 15326
rect 14252 15324 14276 15326
rect 14332 15324 14356 15326
rect 14116 15304 14412 15324
rect 13964 15276 14016 15282
rect 13964 15218 14016 15224
rect 13976 15185 14004 15218
rect 13962 15176 14018 15185
rect 13962 15111 14018 15120
rect 14240 15004 14292 15010
rect 14240 14946 14292 14952
rect 14608 15004 14660 15010
rect 14608 14946 14660 14952
rect 14252 14738 14280 14946
rect 14240 14732 14292 14738
rect 14240 14674 14292 14680
rect 14620 14534 14648 14946
rect 14608 14528 14660 14534
rect 14608 14470 14660 14476
rect 14116 14292 14412 14312
rect 14172 14290 14196 14292
rect 14252 14290 14276 14292
rect 14332 14290 14356 14292
rect 14194 14238 14196 14290
rect 14258 14238 14270 14290
rect 14332 14238 14334 14290
rect 14172 14236 14196 14238
rect 14252 14236 14276 14238
rect 14332 14236 14356 14238
rect 14116 14216 14412 14236
rect 13044 14188 13096 14194
rect 13044 14130 13096 14136
rect 13872 14188 13924 14194
rect 13872 14130 13924 14136
rect 12768 13984 12820 13990
rect 12768 13926 12820 13932
rect 13688 13984 13740 13990
rect 13688 13926 13740 13932
rect 13872 13984 13924 13990
rect 14712 13972 14740 15490
rect 14804 15146 14832 15626
rect 14792 15140 14844 15146
rect 14792 15082 14844 15088
rect 14792 13984 14844 13990
rect 14712 13944 14792 13972
rect 13872 13926 13924 13932
rect 14792 13926 14844 13932
rect 12780 13582 12808 13926
rect 12768 13576 12820 13582
rect 12768 13518 12820 13524
rect 12032 13508 12084 13514
rect 12032 13450 12084 13456
rect 13136 13508 13188 13514
rect 13136 13450 13188 13456
rect 12952 13304 13004 13310
rect 12952 13246 13004 13252
rect 12964 12970 12992 13246
rect 12952 12964 13004 12970
rect 12952 12906 13004 12912
rect 12032 12896 12084 12902
rect 12032 12838 12084 12844
rect 12584 12896 12636 12902
rect 12584 12838 12636 12844
rect 12044 12465 12072 12838
rect 12308 12556 12360 12562
rect 12308 12498 12360 12504
rect 12030 12456 12086 12465
rect 12030 12391 12032 12400
rect 12084 12391 12086 12400
rect 12032 12362 12084 12368
rect 11572 12012 11624 12018
rect 11572 11954 11624 11960
rect 10468 11808 10520 11814
rect 10468 11750 10520 11756
rect 10480 9624 10508 11750
rect 12320 9624 12348 12498
rect 12596 12426 12624 12838
rect 13148 12494 13176 13450
rect 13700 13310 13728 13926
rect 13884 13582 13912 13926
rect 14240 13916 14292 13922
rect 14240 13858 14292 13864
rect 13964 13848 14016 13854
rect 13964 13790 14016 13796
rect 13872 13576 13924 13582
rect 13872 13518 13924 13524
rect 13976 13514 14004 13790
rect 13964 13508 14016 13514
rect 13964 13450 14016 13456
rect 14252 13378 14280 13858
rect 14896 13582 14924 16034
rect 17196 15690 17224 16102
rect 15252 15684 15304 15690
rect 15252 15626 15304 15632
rect 16080 15684 16132 15690
rect 16080 15626 16132 15632
rect 17184 15684 17236 15690
rect 17236 15644 17408 15672
rect 17184 15626 17236 15632
rect 15264 15554 15292 15626
rect 15252 15548 15304 15554
rect 15252 15490 15304 15496
rect 16092 15146 16120 15626
rect 17184 15480 17236 15486
rect 17184 15422 17236 15428
rect 16080 15140 16132 15146
rect 16080 15082 16132 15088
rect 15344 14936 15396 14942
rect 15344 14878 15396 14884
rect 15528 14936 15580 14942
rect 15528 14878 15580 14884
rect 15356 14738 15384 14878
rect 15344 14732 15396 14738
rect 15344 14674 15396 14680
rect 15540 14602 15568 14878
rect 16092 14602 16120 15082
rect 17196 15078 17224 15422
rect 17380 15078 17408 15644
rect 17184 15072 17236 15078
rect 17184 15014 17236 15020
rect 17368 15072 17420 15078
rect 17368 15014 17420 15020
rect 17196 14602 17224 15014
rect 15528 14596 15580 14602
rect 15528 14538 15580 14544
rect 15896 14596 15948 14602
rect 15896 14538 15948 14544
rect 16080 14596 16132 14602
rect 16080 14538 16132 14544
rect 16448 14596 16500 14602
rect 16448 14538 16500 14544
rect 17184 14596 17236 14602
rect 17184 14538 17236 14544
rect 14976 13848 15028 13854
rect 14976 13790 15028 13796
rect 14884 13576 14936 13582
rect 14884 13518 14936 13524
rect 14988 13446 15016 13790
rect 15908 13582 15936 14538
rect 16264 14460 16316 14466
rect 16264 14402 16316 14408
rect 15896 13576 15948 13582
rect 15896 13518 15948 13524
rect 16276 13446 16304 14402
rect 16460 13446 16488 14538
rect 16816 14188 16868 14194
rect 16816 14130 16868 14136
rect 16828 13990 16856 14130
rect 16816 13984 16868 13990
rect 16816 13926 16868 13932
rect 16908 13984 16960 13990
rect 16908 13926 16960 13932
rect 14976 13440 15028 13446
rect 14976 13382 15028 13388
rect 16264 13440 16316 13446
rect 16264 13382 16316 13388
rect 16448 13440 16500 13446
rect 16448 13382 16500 13388
rect 14240 13372 14292 13378
rect 14240 13314 14292 13320
rect 13688 13304 13740 13310
rect 13688 13246 13740 13252
rect 14116 13204 14412 13224
rect 14172 13202 14196 13204
rect 14252 13202 14276 13204
rect 14332 13202 14356 13204
rect 14194 13150 14196 13202
rect 14258 13150 14270 13202
rect 14332 13150 14334 13202
rect 14172 13148 14196 13150
rect 14252 13148 14276 13150
rect 14332 13148 14356 13150
rect 14116 13128 14412 13148
rect 13412 12964 13464 12970
rect 13412 12906 13464 12912
rect 13320 12760 13372 12766
rect 13320 12702 13372 12708
rect 13136 12488 13188 12494
rect 13136 12430 13188 12436
rect 12584 12420 12636 12426
rect 12584 12362 12636 12368
rect 12768 12420 12820 12426
rect 12768 12362 12820 12368
rect 12780 12018 12808 12362
rect 12768 12012 12820 12018
rect 12768 11954 12820 11960
rect 13332 11814 13360 12702
rect 13424 12290 13452 12906
rect 14148 12896 14200 12902
rect 14148 12838 14200 12844
rect 14332 12896 14384 12902
rect 14332 12838 14384 12844
rect 14976 12896 15028 12902
rect 14976 12838 15028 12844
rect 14160 12766 14188 12838
rect 14148 12760 14200 12766
rect 14148 12702 14200 12708
rect 14160 12562 14188 12702
rect 14148 12556 14200 12562
rect 14148 12498 14200 12504
rect 13688 12420 13740 12426
rect 13688 12362 13740 12368
rect 13412 12284 13464 12290
rect 13412 12226 13464 12232
rect 13424 11882 13452 12226
rect 13412 11876 13464 11882
rect 13412 11818 13464 11824
rect 13700 11814 13728 12362
rect 14344 12358 14372 12838
rect 14792 12760 14844 12766
rect 14792 12702 14844 12708
rect 14804 12426 14832 12702
rect 14792 12420 14844 12426
rect 14792 12362 14844 12368
rect 14332 12352 14384 12358
rect 14332 12294 14384 12300
rect 13964 12216 14016 12222
rect 13964 12158 14016 12164
rect 13976 11898 14004 12158
rect 14116 12116 14412 12136
rect 14172 12114 14196 12116
rect 14252 12114 14276 12116
rect 14332 12114 14356 12116
rect 14194 12062 14196 12114
rect 14258 12062 14270 12114
rect 14332 12062 14334 12114
rect 14172 12060 14196 12062
rect 14252 12060 14276 12062
rect 14332 12060 14356 12062
rect 14116 12040 14412 12060
rect 14516 12012 14568 12018
rect 14516 11954 14568 11960
rect 13976 11870 14096 11898
rect 14068 11814 14096 11870
rect 13320 11808 13372 11814
rect 13320 11750 13372 11756
rect 13688 11808 13740 11814
rect 13688 11750 13740 11756
rect 14056 11808 14108 11814
rect 14056 11750 14108 11756
rect 14116 11028 14412 11048
rect 14172 11026 14196 11028
rect 14252 11026 14276 11028
rect 14332 11026 14356 11028
rect 14194 10974 14196 11026
rect 14258 10974 14270 11026
rect 14332 10974 14334 11026
rect 14172 10972 14196 10974
rect 14252 10972 14276 10974
rect 14332 10972 14356 10974
rect 14116 10952 14412 10972
rect 14528 10810 14556 11954
rect 14804 11882 14832 12362
rect 14988 11882 15016 12838
rect 15988 12760 16040 12766
rect 15988 12702 16040 12708
rect 15804 12420 15856 12426
rect 15804 12362 15856 12368
rect 14792 11876 14844 11882
rect 14792 11818 14844 11824
rect 14976 11876 15028 11882
rect 14976 11818 15028 11824
rect 14988 11270 15016 11818
rect 15816 11338 15844 12362
rect 15804 11332 15856 11338
rect 15804 11274 15856 11280
rect 14976 11264 15028 11270
rect 14976 11206 15028 11212
rect 15816 11202 15844 11274
rect 15804 11196 15856 11202
rect 15804 11138 15856 11144
rect 14160 10782 14556 10810
rect 14160 9624 14188 10782
rect 16000 9624 16028 12702
rect 16828 12442 16856 13926
rect 16920 12494 16948 13926
rect 17196 13378 17224 14538
rect 17564 13990 17592 16222
rect 17644 16160 17696 16166
rect 17644 16102 17696 16108
rect 17656 15554 17684 16102
rect 17644 15548 17696 15554
rect 17644 15490 17696 15496
rect 17552 13984 17604 13990
rect 17552 13926 17604 13932
rect 17276 13916 17328 13922
rect 17276 13858 17328 13864
rect 17288 13378 17316 13858
rect 17184 13372 17236 13378
rect 17184 13314 17236 13320
rect 17276 13372 17328 13378
rect 17276 13314 17328 13320
rect 16552 12426 16856 12442
rect 16908 12488 16960 12494
rect 17552 12488 17604 12494
rect 16960 12436 17040 12442
rect 16908 12430 17040 12436
rect 17552 12430 17604 12436
rect 16540 12420 16856 12426
rect 16592 12414 16856 12420
rect 16920 12414 17040 12430
rect 16540 12362 16592 12368
rect 16080 12216 16132 12222
rect 16080 12158 16132 12164
rect 16092 11814 16120 12158
rect 16080 11808 16132 11814
rect 16080 11750 16132 11756
rect 16828 11762 16856 12414
rect 16908 12352 16960 12358
rect 16908 12294 16960 12300
rect 16920 11882 16948 12294
rect 17012 11950 17040 12414
rect 17000 11944 17052 11950
rect 17000 11886 17052 11892
rect 16908 11876 16960 11882
rect 16908 11818 16960 11824
rect 17276 11808 17328 11814
rect 16828 11734 17224 11762
rect 17276 11750 17328 11756
rect 16080 11672 16132 11678
rect 16080 11614 16132 11620
rect 16092 11474 16120 11614
rect 16080 11468 16132 11474
rect 16080 11410 16132 11416
rect 17196 11338 17224 11734
rect 17288 11406 17316 11750
rect 17564 11474 17592 12430
rect 17656 11814 17684 15490
rect 17932 14194 17960 16306
rect 18024 16302 18052 16646
rect 18012 16296 18064 16302
rect 18012 16238 18064 16244
rect 18288 16160 18340 16166
rect 18288 16102 18340 16108
rect 18300 15690 18328 16102
rect 18196 15684 18248 15690
rect 18196 15626 18248 15632
rect 18288 15684 18340 15690
rect 18288 15626 18340 15632
rect 18564 15684 18616 15690
rect 18564 15626 18616 15632
rect 18208 15078 18236 15626
rect 18196 15072 18248 15078
rect 18196 15014 18248 15020
rect 18300 14942 18328 15626
rect 18576 15146 18604 15626
rect 18668 15282 18696 18278
rect 18852 18002 18880 18278
rect 20128 18268 20180 18274
rect 20128 18210 20180 18216
rect 19116 18100 19412 18120
rect 19172 18098 19196 18100
rect 19252 18098 19276 18100
rect 19332 18098 19356 18100
rect 19194 18046 19196 18098
rect 19258 18046 19270 18098
rect 19332 18046 19334 18098
rect 19172 18044 19196 18046
rect 19252 18044 19276 18046
rect 19332 18044 19356 18046
rect 19116 18024 19412 18044
rect 18840 17996 18892 18002
rect 18840 17938 18892 17944
rect 18656 15276 18708 15282
rect 18656 15218 18708 15224
rect 18564 15140 18616 15146
rect 18564 15082 18616 15088
rect 18288 14936 18340 14942
rect 18288 14878 18340 14884
rect 17920 14188 17972 14194
rect 17920 14130 17972 14136
rect 17736 13916 17788 13922
rect 17736 13858 17788 13864
rect 17748 13582 17776 13858
rect 17736 13576 17788 13582
rect 17736 13518 17788 13524
rect 18300 13446 18328 14878
rect 18576 14738 18604 15082
rect 18564 14732 18616 14738
rect 18564 14674 18616 14680
rect 18748 13848 18800 13854
rect 18748 13790 18800 13796
rect 18760 13514 18788 13790
rect 18380 13508 18432 13514
rect 18380 13450 18432 13456
rect 18748 13508 18800 13514
rect 18748 13450 18800 13456
rect 18288 13440 18340 13446
rect 18288 13382 18340 13388
rect 18392 13106 18420 13450
rect 18380 13100 18432 13106
rect 18380 13042 18432 13048
rect 18760 12494 18788 13450
rect 18852 12970 18880 17938
rect 19944 17860 19996 17866
rect 20140 17848 20168 18210
rect 20508 18002 20536 22154
rect 20588 22144 20640 22150
rect 20588 22086 20640 22092
rect 20600 21742 20628 22086
rect 20588 21736 20640 21742
rect 20588 21678 20640 21684
rect 20600 20586 20628 21678
rect 20588 20580 20640 20586
rect 20588 20522 20640 20528
rect 20784 18206 20812 28478
rect 21232 25884 21284 25890
rect 21232 25826 21284 25832
rect 21048 25408 21100 25414
rect 21048 25350 21100 25356
rect 21060 25006 21088 25350
rect 21048 25000 21100 25006
rect 21048 24942 21100 24948
rect 20956 24388 21008 24394
rect 20956 24330 21008 24336
rect 20968 23782 20996 24330
rect 21060 23986 21088 24942
rect 21244 24190 21272 25826
rect 21232 24184 21284 24190
rect 21232 24126 21284 24132
rect 21048 23980 21100 23986
rect 21048 23922 21100 23928
rect 21048 23844 21100 23850
rect 21048 23786 21100 23792
rect 20956 23776 21008 23782
rect 20956 23718 21008 23724
rect 20864 23708 20916 23714
rect 20864 23650 20916 23656
rect 20876 23442 20904 23650
rect 20968 23442 20996 23718
rect 20864 23436 20916 23442
rect 20864 23378 20916 23384
rect 20956 23436 21008 23442
rect 20956 23378 21008 23384
rect 20864 23300 20916 23306
rect 20864 23242 20916 23248
rect 20876 23102 20904 23242
rect 20864 23096 20916 23102
rect 20864 23038 20916 23044
rect 21060 22830 21088 23786
rect 21048 22824 21100 22830
rect 21048 22766 21100 22772
rect 21048 22688 21100 22694
rect 21048 22630 21100 22636
rect 21060 20042 21088 22630
rect 21244 22626 21272 24126
rect 21336 23782 21364 29362
rect 21980 28610 22008 29634
rect 22072 29290 22100 31576
rect 23348 29828 23400 29834
rect 23348 29770 23400 29776
rect 22060 29284 22112 29290
rect 22060 29226 22112 29232
rect 23360 29222 23388 29770
rect 23532 29284 23584 29290
rect 23532 29226 23584 29232
rect 22704 29216 22756 29222
rect 22704 29158 22756 29164
rect 23348 29216 23400 29222
rect 23348 29158 23400 29164
rect 22152 29148 22204 29154
rect 22152 29090 22204 29096
rect 22164 28746 22192 29090
rect 22716 28814 22744 29158
rect 22704 28808 22756 28814
rect 22704 28750 22756 28756
rect 22152 28740 22204 28746
rect 22152 28682 22204 28688
rect 22612 28672 22664 28678
rect 22612 28614 22664 28620
rect 21968 28604 22020 28610
rect 21968 28546 22020 28552
rect 22520 28264 22572 28270
rect 22520 28206 22572 28212
rect 21784 28128 21836 28134
rect 21784 28070 21836 28076
rect 21796 27658 21824 28070
rect 21784 27652 21836 27658
rect 21784 27594 21836 27600
rect 21600 26972 21652 26978
rect 21600 26914 21652 26920
rect 21612 26638 21640 26914
rect 21600 26632 21652 26638
rect 21600 26574 21652 26580
rect 21416 25952 21468 25958
rect 21416 25894 21468 25900
rect 21324 23776 21376 23782
rect 21324 23718 21376 23724
rect 21232 22620 21284 22626
rect 21232 22562 21284 22568
rect 21244 22014 21272 22562
rect 21428 22286 21456 25894
rect 21508 25612 21560 25618
rect 21508 25554 21560 25560
rect 21520 24530 21548 25554
rect 21612 25550 21640 26574
rect 21692 26564 21744 26570
rect 21692 26506 21744 26512
rect 21704 25958 21732 26506
rect 21796 26502 21824 27594
rect 22152 27244 22204 27250
rect 22152 27186 22204 27192
rect 22060 27040 22112 27046
rect 22060 26982 22112 26988
rect 22072 26638 22100 26982
rect 22060 26632 22112 26638
rect 22060 26574 22112 26580
rect 21876 26564 21928 26570
rect 21876 26506 21928 26512
rect 21784 26496 21836 26502
rect 21784 26438 21836 26444
rect 21796 26026 21824 26438
rect 21784 26020 21836 26026
rect 21784 25962 21836 25968
rect 21692 25952 21744 25958
rect 21692 25894 21744 25900
rect 21692 25816 21744 25822
rect 21692 25758 21744 25764
rect 21600 25544 21652 25550
rect 21600 25486 21652 25492
rect 21508 24524 21560 24530
rect 21508 24466 21560 24472
rect 21520 23986 21548 24466
rect 21508 23980 21560 23986
rect 21508 23922 21560 23928
rect 21704 23764 21732 25758
rect 21888 25414 21916 26506
rect 21876 25408 21928 25414
rect 21876 25350 21928 25356
rect 21888 23850 21916 25350
rect 22072 24394 22100 26574
rect 22060 24388 22112 24394
rect 22060 24330 22112 24336
rect 21876 23844 21928 23850
rect 21876 23786 21928 23792
rect 21612 23736 21732 23764
rect 21508 22756 21560 22762
rect 21508 22698 21560 22704
rect 21416 22280 21468 22286
rect 21416 22222 21468 22228
rect 21232 22008 21284 22014
rect 21232 21950 21284 21956
rect 21140 21600 21192 21606
rect 21140 21542 21192 21548
rect 21152 21062 21180 21542
rect 21428 21538 21456 22222
rect 21520 21674 21548 22698
rect 21508 21668 21560 21674
rect 21508 21610 21560 21616
rect 21416 21532 21468 21538
rect 21416 21474 21468 21480
rect 21520 21130 21548 21610
rect 21508 21124 21560 21130
rect 21508 21066 21560 21072
rect 21140 21056 21192 21062
rect 21140 20998 21192 21004
rect 21520 20518 21548 21066
rect 21612 20586 21640 23736
rect 21692 22212 21744 22218
rect 21692 22154 21744 22160
rect 21704 21810 21732 22154
rect 21888 22150 21916 23786
rect 22072 23782 22100 24330
rect 22060 23776 22112 23782
rect 22060 23718 22112 23724
rect 22072 23306 22100 23718
rect 22060 23300 22112 23306
rect 22060 23242 22112 23248
rect 21968 22348 22020 22354
rect 21968 22290 22020 22296
rect 21980 22150 22008 22290
rect 21876 22144 21928 22150
rect 21876 22086 21928 22092
rect 21968 22144 22020 22150
rect 21968 22086 22020 22092
rect 21968 22008 22020 22014
rect 21968 21950 22020 21956
rect 21692 21804 21744 21810
rect 21692 21746 21744 21752
rect 21876 21124 21928 21130
rect 21876 21066 21928 21072
rect 21692 21056 21744 21062
rect 21692 20998 21744 21004
rect 21600 20580 21652 20586
rect 21600 20522 21652 20528
rect 21508 20512 21560 20518
rect 21508 20454 21560 20460
rect 21520 20110 21548 20454
rect 21508 20104 21560 20110
rect 21508 20046 21560 20052
rect 21048 20036 21100 20042
rect 21048 19978 21100 19984
rect 21704 19974 21732 20998
rect 21784 20988 21836 20994
rect 21784 20930 21836 20936
rect 21796 20518 21824 20930
rect 21888 20722 21916 21066
rect 21980 21062 22008 21950
rect 22164 21062 22192 27186
rect 22532 26978 22560 28206
rect 22624 27658 22652 28614
rect 22716 28202 22744 28750
rect 22796 28672 22848 28678
rect 22796 28614 22848 28620
rect 22704 28196 22756 28202
rect 22704 28138 22756 28144
rect 22612 27652 22664 27658
rect 22612 27594 22664 27600
rect 22520 26972 22572 26978
rect 22520 26914 22572 26920
rect 22532 26706 22560 26914
rect 22520 26700 22572 26706
rect 22520 26642 22572 26648
rect 22520 25884 22572 25890
rect 22520 25826 22572 25832
rect 22428 25408 22480 25414
rect 22428 25350 22480 25356
rect 22440 25090 22468 25350
rect 22348 25074 22468 25090
rect 22336 25068 22468 25074
rect 22388 25062 22468 25068
rect 22336 25010 22388 25016
rect 22532 24954 22560 25826
rect 22440 24926 22560 24954
rect 22440 24870 22468 24926
rect 22428 24864 22480 24870
rect 22428 24806 22480 24812
rect 22808 24002 22836 28614
rect 23360 28270 23388 29158
rect 23544 28728 23572 29226
rect 23716 29080 23768 29086
rect 23716 29022 23768 29028
rect 23624 28740 23676 28746
rect 23544 28700 23624 28728
rect 23348 28264 23400 28270
rect 23348 28206 23400 28212
rect 23544 27674 23572 28700
rect 23624 28682 23676 28688
rect 23728 28134 23756 29022
rect 23716 28128 23768 28134
rect 23716 28070 23768 28076
rect 23808 28060 23860 28066
rect 23808 28002 23860 28008
rect 23268 27658 23572 27674
rect 23072 27652 23124 27658
rect 23072 27594 23124 27600
rect 23268 27652 23584 27658
rect 23268 27646 23532 27652
rect 22888 26564 22940 26570
rect 22888 26506 22940 26512
rect 22900 25890 22928 26506
rect 22888 25884 22940 25890
rect 22888 25826 22940 25832
rect 22624 23974 22836 24002
rect 22428 23640 22480 23646
rect 22428 23582 22480 23588
rect 22244 23368 22296 23374
rect 22296 23316 22376 23322
rect 22244 23310 22376 23316
rect 22256 23294 22376 23310
rect 22348 22558 22376 23294
rect 22440 23102 22468 23582
rect 22520 23368 22572 23374
rect 22520 23310 22572 23316
rect 22428 23096 22480 23102
rect 22428 23038 22480 23044
rect 22532 22694 22560 23310
rect 22520 22688 22572 22694
rect 22520 22630 22572 22636
rect 22336 22552 22388 22558
rect 22336 22494 22388 22500
rect 22624 22354 22652 23974
rect 22900 23238 22928 25826
rect 22980 23776 23032 23782
rect 22980 23718 23032 23724
rect 22888 23232 22940 23238
rect 22888 23174 22940 23180
rect 22900 22914 22928 23174
rect 22808 22898 22928 22914
rect 22796 22892 22928 22898
rect 22848 22886 22928 22892
rect 22796 22834 22848 22840
rect 22612 22348 22664 22354
rect 22612 22290 22664 22296
rect 22336 22008 22388 22014
rect 22336 21950 22388 21956
rect 21968 21056 22020 21062
rect 21968 20998 22020 21004
rect 22152 21056 22204 21062
rect 22204 21016 22284 21044
rect 22152 20998 22204 21004
rect 21876 20716 21928 20722
rect 21876 20658 21928 20664
rect 21784 20512 21836 20518
rect 21784 20454 21836 20460
rect 22256 20042 22284 21016
rect 22348 20518 22376 21950
rect 22624 21606 22652 22290
rect 22992 22218 23020 23718
rect 22980 22212 23032 22218
rect 22980 22154 23032 22160
rect 23084 22098 23112 27594
rect 23268 27590 23296 27646
rect 23532 27594 23584 27600
rect 23256 27584 23308 27590
rect 23256 27526 23308 27532
rect 23348 27584 23400 27590
rect 23348 27526 23400 27532
rect 23360 27454 23388 27526
rect 23348 27448 23400 27454
rect 23348 27390 23400 27396
rect 23164 25544 23216 25550
rect 23164 25486 23216 25492
rect 23176 24938 23204 25486
rect 23164 24932 23216 24938
rect 23164 24874 23216 24880
rect 23360 24802 23388 27390
rect 23820 27114 23848 28002
rect 23912 27590 23940 31576
rect 24116 29524 24412 29544
rect 24172 29522 24196 29524
rect 24252 29522 24276 29524
rect 24332 29522 24356 29524
rect 24194 29470 24196 29522
rect 24258 29470 24270 29522
rect 24332 29470 24334 29522
rect 24172 29468 24196 29470
rect 24252 29468 24276 29470
rect 24332 29468 24356 29470
rect 24116 29448 24412 29468
rect 24452 29216 24504 29222
rect 24452 29158 24504 29164
rect 25464 29216 25516 29222
rect 25464 29158 25516 29164
rect 24464 28882 24492 29158
rect 24452 28876 24504 28882
rect 24452 28818 24504 28824
rect 25476 28814 25504 29158
rect 25464 28808 25516 28814
rect 25464 28750 25516 28756
rect 24728 28740 24780 28746
rect 24728 28682 24780 28688
rect 25280 28740 25332 28746
rect 25280 28682 25332 28688
rect 24116 28436 24412 28456
rect 24172 28434 24196 28436
rect 24252 28434 24276 28436
rect 24332 28434 24356 28436
rect 24194 28382 24196 28434
rect 24258 28382 24270 28434
rect 24332 28382 24334 28434
rect 24172 28380 24196 28382
rect 24252 28380 24276 28382
rect 24332 28380 24356 28382
rect 24116 28360 24412 28380
rect 24740 28270 24768 28682
rect 24728 28264 24780 28270
rect 24728 28206 24780 28212
rect 23900 27584 23952 27590
rect 23900 27526 23952 27532
rect 24116 27348 24412 27368
rect 24172 27346 24196 27348
rect 24252 27346 24276 27348
rect 24332 27346 24356 27348
rect 24194 27294 24196 27346
rect 24258 27294 24270 27346
rect 24332 27294 24334 27346
rect 24172 27292 24196 27294
rect 24252 27292 24276 27294
rect 24332 27292 24356 27294
rect 24116 27272 24412 27292
rect 23992 27176 24044 27182
rect 23992 27118 24044 27124
rect 23808 27108 23860 27114
rect 23808 27050 23860 27056
rect 23716 27040 23768 27046
rect 23716 26982 23768 26988
rect 23624 26700 23676 26706
rect 23624 26642 23676 26648
rect 23440 25816 23492 25822
rect 23440 25758 23492 25764
rect 23452 25074 23480 25758
rect 23532 25408 23584 25414
rect 23532 25350 23584 25356
rect 23440 25068 23492 25074
rect 23440 25010 23492 25016
rect 23544 25006 23572 25350
rect 23532 25000 23584 25006
rect 23532 24942 23584 24948
rect 23440 24864 23492 24870
rect 23440 24806 23492 24812
rect 23348 24796 23400 24802
rect 23348 24738 23400 24744
rect 23164 24388 23216 24394
rect 23360 24376 23388 24738
rect 23216 24348 23388 24376
rect 23164 24330 23216 24336
rect 23452 24308 23480 24806
rect 23360 24280 23480 24308
rect 23164 24252 23216 24258
rect 23164 24194 23216 24200
rect 23176 22762 23204 24194
rect 23360 23850 23388 24280
rect 23440 24184 23492 24190
rect 23440 24126 23492 24132
rect 23348 23844 23400 23850
rect 23348 23786 23400 23792
rect 23452 23374 23480 24126
rect 23544 23782 23572 24942
rect 23636 24258 23664 26642
rect 23728 26638 23756 26982
rect 23716 26632 23768 26638
rect 23716 26574 23768 26580
rect 23900 25476 23952 25482
rect 23900 25418 23952 25424
rect 23808 25272 23860 25278
rect 23808 25214 23860 25220
rect 23820 24870 23848 25214
rect 23808 24864 23860 24870
rect 23808 24806 23860 24812
rect 23820 24462 23848 24806
rect 23808 24456 23860 24462
rect 23808 24398 23860 24404
rect 23624 24252 23676 24258
rect 23624 24194 23676 24200
rect 23636 24002 23664 24194
rect 23808 24184 23860 24190
rect 23808 24126 23860 24132
rect 23636 23974 23756 24002
rect 23728 23918 23756 23974
rect 23624 23912 23676 23918
rect 23624 23854 23676 23860
rect 23716 23912 23768 23918
rect 23716 23854 23768 23860
rect 23532 23776 23584 23782
rect 23532 23718 23584 23724
rect 23440 23368 23492 23374
rect 23440 23310 23492 23316
rect 23636 23306 23664 23854
rect 23716 23776 23768 23782
rect 23716 23718 23768 23724
rect 23728 23374 23756 23718
rect 23716 23368 23768 23374
rect 23716 23310 23768 23316
rect 23624 23300 23676 23306
rect 23624 23242 23676 23248
rect 23440 23232 23492 23238
rect 23440 23174 23492 23180
rect 23348 22892 23400 22898
rect 23348 22834 23400 22840
rect 23164 22756 23216 22762
rect 23164 22698 23216 22704
rect 23256 22688 23308 22694
rect 23256 22630 23308 22636
rect 23268 22558 23296 22630
rect 23256 22552 23308 22558
rect 23256 22494 23308 22500
rect 23268 22218 23296 22494
rect 23360 22234 23388 22834
rect 23452 22830 23480 23174
rect 23532 23096 23584 23102
rect 23532 23038 23584 23044
rect 23544 22898 23572 23038
rect 23532 22892 23584 22898
rect 23532 22834 23584 22840
rect 23440 22824 23492 22830
rect 23440 22766 23492 22772
rect 23256 22212 23308 22218
rect 23360 22206 23480 22234
rect 23256 22154 23308 22160
rect 22992 22070 23112 22098
rect 23164 22144 23216 22150
rect 23164 22086 23216 22092
rect 22704 21668 22756 21674
rect 22704 21610 22756 21616
rect 22612 21600 22664 21606
rect 22612 21542 22664 21548
rect 22716 21470 22744 21610
rect 22704 21464 22756 21470
rect 22704 21406 22756 21412
rect 22716 20722 22744 21406
rect 22704 20716 22756 20722
rect 22704 20658 22756 20664
rect 22336 20512 22388 20518
rect 22336 20454 22388 20460
rect 22152 20036 22204 20042
rect 22152 19978 22204 19984
rect 22244 20036 22296 20042
rect 22244 19978 22296 19984
rect 21692 19968 21744 19974
rect 21692 19910 21744 19916
rect 22164 19090 22192 19978
rect 22152 19084 22204 19090
rect 22152 19026 22204 19032
rect 20956 18948 21008 18954
rect 20956 18890 21008 18896
rect 21968 18948 22020 18954
rect 21968 18890 22020 18896
rect 20772 18200 20824 18206
rect 20772 18142 20824 18148
rect 20496 17996 20548 18002
rect 20496 17938 20548 17944
rect 20784 17866 20812 18142
rect 19996 17820 20168 17848
rect 20772 17860 20824 17866
rect 19944 17802 19996 17808
rect 20772 17802 20824 17808
rect 19576 17180 19628 17186
rect 19576 17122 19628 17128
rect 19484 17112 19536 17118
rect 19484 17054 19536 17060
rect 19116 17012 19412 17032
rect 19172 17010 19196 17012
rect 19252 17010 19276 17012
rect 19332 17010 19356 17012
rect 19194 16958 19196 17010
rect 19258 16958 19270 17010
rect 19332 16958 19334 17010
rect 19172 16956 19196 16958
rect 19252 16956 19276 16958
rect 19332 16956 19356 16958
rect 19116 16936 19412 16956
rect 19496 16914 19524 17054
rect 19588 16914 19616 17122
rect 19484 16908 19536 16914
rect 19484 16850 19536 16856
rect 19576 16908 19628 16914
rect 19576 16850 19628 16856
rect 19496 16710 19524 16850
rect 19576 16772 19628 16778
rect 19576 16714 19628 16720
rect 19484 16704 19536 16710
rect 19484 16646 19536 16652
rect 19588 16370 19616 16714
rect 19576 16364 19628 16370
rect 19576 16306 19628 16312
rect 18932 16160 18984 16166
rect 18932 16102 18984 16108
rect 18944 15622 18972 16102
rect 19024 16092 19076 16098
rect 19024 16034 19076 16040
rect 18932 15616 18984 15622
rect 18932 15558 18984 15564
rect 18944 15010 18972 15558
rect 19036 15282 19064 16034
rect 19116 15924 19412 15944
rect 19172 15922 19196 15924
rect 19252 15922 19276 15924
rect 19332 15922 19356 15924
rect 19194 15870 19196 15922
rect 19258 15870 19270 15922
rect 19332 15870 19334 15922
rect 19172 15868 19196 15870
rect 19252 15868 19276 15870
rect 19332 15868 19356 15870
rect 19116 15848 19412 15868
rect 19852 15548 19904 15554
rect 19852 15490 19904 15496
rect 19024 15276 19076 15282
rect 19024 15218 19076 15224
rect 19864 15078 19892 15490
rect 19852 15072 19904 15078
rect 19852 15014 19904 15020
rect 18932 15004 18984 15010
rect 18932 14946 18984 14952
rect 19024 14936 19076 14942
rect 19024 14878 19076 14884
rect 18932 14392 18984 14398
rect 18932 14334 18984 14340
rect 18944 13514 18972 14334
rect 19036 13972 19064 14878
rect 19116 14836 19412 14856
rect 19172 14834 19196 14836
rect 19252 14834 19276 14836
rect 19332 14834 19356 14836
rect 19194 14782 19196 14834
rect 19258 14782 19270 14834
rect 19332 14782 19334 14834
rect 19172 14780 19196 14782
rect 19252 14780 19276 14782
rect 19332 14780 19356 14782
rect 19116 14760 19412 14780
rect 19864 14670 19892 15014
rect 19852 14664 19904 14670
rect 19852 14606 19904 14612
rect 19116 13984 19168 13990
rect 19036 13944 19116 13972
rect 19116 13926 19168 13932
rect 19116 13748 19412 13768
rect 19172 13746 19196 13748
rect 19252 13746 19276 13748
rect 19332 13746 19356 13748
rect 19194 13694 19196 13746
rect 19258 13694 19270 13746
rect 19332 13694 19334 13746
rect 19172 13692 19196 13694
rect 19252 13692 19276 13694
rect 19332 13692 19356 13694
rect 19116 13672 19412 13692
rect 19576 13644 19628 13650
rect 19576 13586 19628 13592
rect 18932 13508 18984 13514
rect 18932 13450 18984 13456
rect 18944 13122 18972 13450
rect 18944 13094 19064 13122
rect 19036 13038 19064 13094
rect 19024 13032 19076 13038
rect 19588 12986 19616 13586
rect 19024 12974 19076 12980
rect 18840 12964 18892 12970
rect 18840 12906 18892 12912
rect 18196 12488 18248 12494
rect 18196 12430 18248 12436
rect 18748 12488 18800 12494
rect 18748 12430 18800 12436
rect 18208 11814 18236 12430
rect 18932 12216 18984 12222
rect 18932 12158 18984 12164
rect 18944 11882 18972 12158
rect 18932 11876 18984 11882
rect 18932 11818 18984 11824
rect 17644 11808 17696 11814
rect 17644 11750 17696 11756
rect 18196 11808 18248 11814
rect 18196 11750 18248 11756
rect 18012 11672 18064 11678
rect 18012 11614 18064 11620
rect 17552 11468 17604 11474
rect 17552 11410 17604 11416
rect 17276 11400 17328 11406
rect 17276 11342 17328 11348
rect 17184 11332 17236 11338
rect 17184 11274 17236 11280
rect 17288 11270 17316 11342
rect 17276 11264 17328 11270
rect 17276 11206 17328 11212
rect 18024 9624 18052 11614
rect 18208 11338 18236 11750
rect 19036 11746 19064 12974
rect 19312 12970 19616 12986
rect 19300 12964 19616 12970
rect 19352 12958 19616 12964
rect 19300 12906 19352 12912
rect 19392 12896 19444 12902
rect 19444 12856 19524 12884
rect 19392 12838 19444 12844
rect 19116 12660 19412 12680
rect 19172 12658 19196 12660
rect 19252 12658 19276 12660
rect 19332 12658 19356 12660
rect 19194 12606 19196 12658
rect 19258 12606 19270 12658
rect 19332 12606 19334 12658
rect 19172 12604 19196 12606
rect 19252 12604 19276 12606
rect 19332 12604 19356 12606
rect 19116 12584 19412 12604
rect 19024 11740 19076 11746
rect 19024 11682 19076 11688
rect 19116 11572 19412 11592
rect 19172 11570 19196 11572
rect 19252 11570 19276 11572
rect 19332 11570 19356 11572
rect 19194 11518 19196 11570
rect 19258 11518 19270 11570
rect 19332 11518 19334 11570
rect 19172 11516 19196 11518
rect 19252 11516 19276 11518
rect 19332 11516 19356 11518
rect 19116 11496 19412 11516
rect 19496 11474 19524 12856
rect 19576 12828 19628 12834
rect 19576 12770 19628 12776
rect 19588 12426 19616 12770
rect 19956 12766 19984 17802
rect 20680 17656 20732 17662
rect 20680 17598 20732 17604
rect 20692 17254 20720 17598
rect 20680 17248 20732 17254
rect 20680 17190 20732 17196
rect 20772 16772 20824 16778
rect 20772 16714 20824 16720
rect 20784 16166 20812 16714
rect 20864 16704 20916 16710
rect 20864 16646 20916 16652
rect 20876 16302 20904 16646
rect 20864 16296 20916 16302
rect 20864 16238 20916 16244
rect 20772 16160 20824 16166
rect 20772 16102 20824 16108
rect 20312 15480 20364 15486
rect 20312 15422 20364 15428
rect 20404 15480 20456 15486
rect 20404 15422 20456 15428
rect 20324 15078 20352 15422
rect 20312 15072 20364 15078
rect 20312 15014 20364 15020
rect 20324 14602 20352 15014
rect 20312 14596 20364 14602
rect 20312 14538 20364 14544
rect 20036 14528 20088 14534
rect 20036 14470 20088 14476
rect 20048 13990 20076 14470
rect 20324 13990 20352 14538
rect 20036 13984 20088 13990
rect 20036 13926 20088 13932
rect 20312 13984 20364 13990
rect 20312 13926 20364 13932
rect 20048 13514 20076 13926
rect 20324 13514 20352 13926
rect 20416 13922 20444 15422
rect 20588 15072 20640 15078
rect 20588 15014 20640 15020
rect 20600 14466 20628 15014
rect 20588 14460 20640 14466
rect 20588 14402 20640 14408
rect 20404 13916 20456 13922
rect 20404 13858 20456 13864
rect 20036 13508 20088 13514
rect 20036 13450 20088 13456
rect 20312 13508 20364 13514
rect 20312 13450 20364 13456
rect 20048 12970 20076 13450
rect 20036 12964 20088 12970
rect 20036 12906 20088 12912
rect 19944 12760 19996 12766
rect 19944 12702 19996 12708
rect 19852 12556 19904 12562
rect 19852 12498 19904 12504
rect 19576 12420 19628 12426
rect 19576 12362 19628 12368
rect 19484 11468 19536 11474
rect 19484 11410 19536 11416
rect 18196 11332 18248 11338
rect 18196 11274 18248 11280
rect 19864 9624 19892 12498
rect 19944 11740 19996 11746
rect 19944 11682 19996 11688
rect 19956 11474 19984 11682
rect 19944 11468 19996 11474
rect 19944 11410 19996 11416
rect 20416 11406 20444 13858
rect 20600 13106 20628 14402
rect 20784 13990 20812 16102
rect 20772 13984 20824 13990
rect 20772 13926 20824 13932
rect 20588 13100 20640 13106
rect 20588 13042 20640 13048
rect 20680 12964 20732 12970
rect 20680 12906 20732 12912
rect 20692 11882 20720 12906
rect 20968 12018 20996 18890
rect 21980 18478 22008 18890
rect 22256 18478 22284 19978
rect 22992 19430 23020 22070
rect 23176 21742 23204 22086
rect 23164 21736 23216 21742
rect 23164 21678 23216 21684
rect 23452 21674 23480 22206
rect 23636 22082 23664 23242
rect 23820 23170 23848 24126
rect 23912 23850 23940 25418
rect 23900 23844 23952 23850
rect 23900 23786 23952 23792
rect 23808 23164 23860 23170
rect 23808 23106 23860 23112
rect 23900 23096 23952 23102
rect 23900 23038 23952 23044
rect 23716 22824 23768 22830
rect 23716 22766 23768 22772
rect 23624 22076 23676 22082
rect 23624 22018 23676 22024
rect 23440 21668 23492 21674
rect 23440 21610 23492 21616
rect 23348 21532 23400 21538
rect 23348 21474 23400 21480
rect 23360 21130 23388 21474
rect 23348 21124 23400 21130
rect 23348 21066 23400 21072
rect 23452 20654 23480 21610
rect 23532 20988 23584 20994
rect 23532 20930 23584 20936
rect 23440 20648 23492 20654
rect 23440 20590 23492 20596
rect 23544 20042 23572 20930
rect 23532 20036 23584 20042
rect 23532 19978 23584 19984
rect 22980 19424 23032 19430
rect 22980 19366 23032 19372
rect 23072 19424 23124 19430
rect 23072 19366 23124 19372
rect 22796 19084 22848 19090
rect 22796 19026 22848 19032
rect 22808 18478 22836 19026
rect 22992 18954 23020 19366
rect 23084 19022 23112 19366
rect 23072 19016 23124 19022
rect 23072 18958 23124 18964
rect 22980 18948 23032 18954
rect 22980 18890 23032 18896
rect 21968 18472 22020 18478
rect 21968 18414 22020 18420
rect 22244 18472 22296 18478
rect 22244 18414 22296 18420
rect 22796 18472 22848 18478
rect 22796 18414 22848 18420
rect 23084 18274 23112 18958
rect 21140 18268 21192 18274
rect 21140 18210 21192 18216
rect 23072 18268 23124 18274
rect 23072 18210 23124 18216
rect 21152 17866 21180 18210
rect 23348 17996 23400 18002
rect 23348 17938 23400 17944
rect 21140 17860 21192 17866
rect 21140 17802 21192 17808
rect 22336 17860 22388 17866
rect 22336 17802 22388 17808
rect 21324 17180 21376 17186
rect 21324 17122 21376 17128
rect 21140 16704 21192 16710
rect 21140 16646 21192 16652
rect 21152 16234 21180 16646
rect 21140 16228 21192 16234
rect 21140 16170 21192 16176
rect 21336 15554 21364 17122
rect 22348 16642 22376 17802
rect 23360 17254 23388 17938
rect 23440 17860 23492 17866
rect 23440 17802 23492 17808
rect 23348 17248 23400 17254
rect 23348 17190 23400 17196
rect 23452 17118 23480 17802
rect 23728 17730 23756 22766
rect 23912 22762 23940 23038
rect 23900 22756 23952 22762
rect 23900 22698 23952 22704
rect 23808 22688 23860 22694
rect 23808 22630 23860 22636
rect 23820 21810 23848 22630
rect 23912 22286 23940 22698
rect 23900 22280 23952 22286
rect 23900 22222 23952 22228
rect 23808 21804 23860 21810
rect 23808 21746 23860 21752
rect 23900 21464 23952 21470
rect 23900 21406 23952 21412
rect 23716 17724 23768 17730
rect 23716 17666 23768 17672
rect 23532 17316 23584 17322
rect 23532 17258 23584 17264
rect 23440 17112 23492 17118
rect 23440 17054 23492 17060
rect 23452 16778 23480 17054
rect 22520 16772 22572 16778
rect 22520 16714 22572 16720
rect 23440 16772 23492 16778
rect 23440 16714 23492 16720
rect 22244 16636 22296 16642
rect 22244 16578 22296 16584
rect 22336 16636 22388 16642
rect 22336 16578 22388 16584
rect 21416 16160 21468 16166
rect 21416 16102 21468 16108
rect 21324 15548 21376 15554
rect 21324 15490 21376 15496
rect 21428 15282 21456 16102
rect 22256 15690 22284 16578
rect 22348 16166 22376 16578
rect 22532 16370 22560 16714
rect 22520 16364 22572 16370
rect 22520 16306 22572 16312
rect 23164 16228 23216 16234
rect 23164 16170 23216 16176
rect 22336 16160 22388 16166
rect 22336 16102 22388 16108
rect 22244 15684 22296 15690
rect 22244 15626 22296 15632
rect 22520 15684 22572 15690
rect 22520 15626 22572 15632
rect 21416 15276 21468 15282
rect 21416 15218 21468 15224
rect 22256 15078 22284 15626
rect 22428 15548 22480 15554
rect 22428 15490 22480 15496
rect 22440 15434 22468 15490
rect 22348 15406 22468 15434
rect 22348 15146 22376 15406
rect 22532 15282 22560 15626
rect 23176 15622 23204 16170
rect 23164 15616 23216 15622
rect 23164 15558 23216 15564
rect 22520 15276 22572 15282
rect 22520 15218 22572 15224
rect 22336 15140 22388 15146
rect 22336 15082 22388 15088
rect 22244 15072 22296 15078
rect 22244 15014 22296 15020
rect 22060 14392 22112 14398
rect 22060 14334 22112 14340
rect 22072 13514 22100 14334
rect 22348 13990 22376 15082
rect 22428 15072 22480 15078
rect 22428 15014 22480 15020
rect 22440 14194 22468 15014
rect 22532 14534 22560 15218
rect 22980 15208 23032 15214
rect 22980 15150 23032 15156
rect 22612 15072 22664 15078
rect 22612 15014 22664 15020
rect 22624 14602 22652 15014
rect 22992 14602 23020 15150
rect 23176 14602 23204 15558
rect 22612 14596 22664 14602
rect 22612 14538 22664 14544
rect 22980 14596 23032 14602
rect 22980 14538 23032 14544
rect 23164 14596 23216 14602
rect 23164 14538 23216 14544
rect 22520 14528 22572 14534
rect 22520 14470 22572 14476
rect 22428 14188 22480 14194
rect 22428 14130 22480 14136
rect 22624 13990 22652 14538
rect 22336 13984 22388 13990
rect 22336 13926 22388 13932
rect 22612 13984 22664 13990
rect 22612 13926 22664 13932
rect 22624 13650 22652 13926
rect 22612 13644 22664 13650
rect 22612 13586 22664 13592
rect 21140 13508 21192 13514
rect 21140 13450 21192 13456
rect 22060 13508 22112 13514
rect 22060 13450 22112 13456
rect 21152 12426 21180 13450
rect 21232 13440 21284 13446
rect 21232 13382 21284 13388
rect 21244 13038 21272 13382
rect 21232 13032 21284 13038
rect 21232 12974 21284 12980
rect 21232 12896 21284 12902
rect 21232 12838 21284 12844
rect 22152 12896 22204 12902
rect 22152 12838 22204 12844
rect 21140 12420 21192 12426
rect 21140 12362 21192 12368
rect 21244 12358 21272 12838
rect 21692 12760 21744 12766
rect 21692 12702 21744 12708
rect 21704 12426 21732 12702
rect 21508 12420 21560 12426
rect 21508 12362 21560 12368
rect 21692 12420 21744 12426
rect 21692 12362 21744 12368
rect 21232 12352 21284 12358
rect 21232 12294 21284 12300
rect 21244 12018 21272 12294
rect 20956 12012 21008 12018
rect 20956 11954 21008 11960
rect 21232 12012 21284 12018
rect 21232 11954 21284 11960
rect 21520 11882 21548 12362
rect 21704 11950 21732 12362
rect 22164 12222 22192 12838
rect 23544 12562 23572 17258
rect 23728 17254 23756 17666
rect 23912 17390 23940 21406
rect 24004 21198 24032 27118
rect 24452 27108 24504 27114
rect 24452 27050 24504 27056
rect 24116 26260 24412 26280
rect 24172 26258 24196 26260
rect 24252 26258 24276 26260
rect 24332 26258 24356 26260
rect 24194 26206 24196 26258
rect 24258 26206 24270 26258
rect 24332 26206 24334 26258
rect 24172 26204 24196 26206
rect 24252 26204 24276 26206
rect 24332 26204 24356 26206
rect 24116 26184 24412 26204
rect 24176 25884 24228 25890
rect 24176 25826 24228 25832
rect 24188 25414 24216 25826
rect 24176 25408 24228 25414
rect 24176 25350 24228 25356
rect 24116 25172 24412 25192
rect 24172 25170 24196 25172
rect 24252 25170 24276 25172
rect 24332 25170 24356 25172
rect 24194 25118 24196 25170
rect 24258 25118 24270 25170
rect 24332 25118 24334 25170
rect 24172 25116 24196 25118
rect 24252 25116 24276 25118
rect 24332 25116 24356 25118
rect 24116 25096 24412 25116
rect 24116 24084 24412 24104
rect 24172 24082 24196 24084
rect 24252 24082 24276 24084
rect 24332 24082 24356 24084
rect 24194 24030 24196 24082
rect 24258 24030 24270 24082
rect 24332 24030 24334 24082
rect 24172 24028 24196 24030
rect 24252 24028 24276 24030
rect 24332 24028 24356 24030
rect 24116 24008 24412 24028
rect 24116 22996 24412 23016
rect 24172 22994 24196 22996
rect 24252 22994 24276 22996
rect 24332 22994 24356 22996
rect 24194 22942 24196 22994
rect 24258 22942 24270 22994
rect 24332 22942 24334 22994
rect 24172 22940 24196 22942
rect 24252 22940 24276 22942
rect 24332 22940 24356 22942
rect 24116 22920 24412 22940
rect 24116 21908 24412 21928
rect 24172 21906 24196 21908
rect 24252 21906 24276 21908
rect 24332 21906 24356 21908
rect 24194 21854 24196 21906
rect 24258 21854 24270 21906
rect 24332 21854 24334 21906
rect 24172 21852 24196 21854
rect 24252 21852 24276 21854
rect 24332 21852 24356 21854
rect 24116 21832 24412 21852
rect 23992 21192 24044 21198
rect 23992 21134 24044 21140
rect 24116 20820 24412 20840
rect 24172 20818 24196 20820
rect 24252 20818 24276 20820
rect 24332 20818 24356 20820
rect 24194 20766 24196 20818
rect 24258 20766 24270 20818
rect 24332 20766 24334 20818
rect 24172 20764 24196 20766
rect 24252 20764 24276 20766
rect 24332 20764 24356 20766
rect 24116 20744 24412 20764
rect 23992 20036 24044 20042
rect 23992 19978 24044 19984
rect 24004 19498 24032 19978
rect 24116 19732 24412 19752
rect 24172 19730 24196 19732
rect 24252 19730 24276 19732
rect 24332 19730 24356 19732
rect 24194 19678 24196 19730
rect 24258 19678 24270 19730
rect 24332 19678 24334 19730
rect 24172 19676 24196 19678
rect 24252 19676 24276 19678
rect 24332 19676 24356 19678
rect 24116 19656 24412 19676
rect 24268 19560 24320 19566
rect 24268 19502 24320 19508
rect 23992 19492 24044 19498
rect 23992 19434 24044 19440
rect 24280 19022 24308 19502
rect 23992 19016 24044 19022
rect 23992 18958 24044 18964
rect 24268 19016 24320 19022
rect 24268 18958 24320 18964
rect 24004 18342 24032 18958
rect 24116 18644 24412 18664
rect 24172 18642 24196 18644
rect 24252 18642 24276 18644
rect 24332 18642 24356 18644
rect 24194 18590 24196 18642
rect 24258 18590 24270 18642
rect 24332 18590 24334 18642
rect 24172 18588 24196 18590
rect 24252 18588 24276 18590
rect 24332 18588 24356 18590
rect 24116 18568 24412 18588
rect 23992 18336 24044 18342
rect 23992 18278 24044 18284
rect 23992 17860 24044 17866
rect 23992 17802 24044 17808
rect 23900 17384 23952 17390
rect 23900 17326 23952 17332
rect 23716 17248 23768 17254
rect 23716 17190 23768 17196
rect 24004 16710 24032 17802
rect 24116 17556 24412 17576
rect 24172 17554 24196 17556
rect 24252 17554 24276 17556
rect 24332 17554 24356 17556
rect 24194 17502 24196 17554
rect 24258 17502 24270 17554
rect 24332 17502 24334 17554
rect 24172 17500 24196 17502
rect 24252 17500 24276 17502
rect 24332 17500 24356 17502
rect 24116 17480 24412 17500
rect 23992 16704 24044 16710
rect 23992 16646 24044 16652
rect 24116 16468 24412 16488
rect 24172 16466 24196 16468
rect 24252 16466 24276 16468
rect 24332 16466 24356 16468
rect 24194 16414 24196 16466
rect 24258 16414 24270 16466
rect 24332 16414 24334 16466
rect 24172 16412 24196 16414
rect 24252 16412 24276 16414
rect 24332 16412 24356 16414
rect 24116 16392 24412 16412
rect 23900 16092 23952 16098
rect 23900 16034 23952 16040
rect 23912 15826 23940 16034
rect 23900 15820 23952 15826
rect 23900 15762 23952 15768
rect 23808 15684 23860 15690
rect 23808 15626 23860 15632
rect 23820 15146 23848 15626
rect 24116 15380 24412 15400
rect 24172 15378 24196 15380
rect 24252 15378 24276 15380
rect 24332 15378 24356 15380
rect 24194 15326 24196 15378
rect 24258 15326 24270 15378
rect 24332 15326 24334 15378
rect 24172 15324 24196 15326
rect 24252 15324 24276 15326
rect 24332 15324 24356 15326
rect 24116 15304 24412 15324
rect 23808 15140 23860 15146
rect 23808 15082 23860 15088
rect 23992 15072 24044 15078
rect 23992 15014 24044 15020
rect 23808 15004 23860 15010
rect 23808 14946 23860 14952
rect 23820 13990 23848 14946
rect 24004 14738 24032 15014
rect 23992 14732 24044 14738
rect 23992 14674 24044 14680
rect 23900 14528 23952 14534
rect 23900 14470 23952 14476
rect 23808 13984 23860 13990
rect 23808 13926 23860 13932
rect 23820 13514 23848 13926
rect 23912 13650 23940 14470
rect 24116 14292 24412 14312
rect 24172 14290 24196 14292
rect 24252 14290 24276 14292
rect 24332 14290 24356 14292
rect 24194 14238 24196 14290
rect 24258 14238 24270 14290
rect 24332 14238 24334 14290
rect 24172 14236 24196 14238
rect 24252 14236 24276 14238
rect 24332 14236 24356 14238
rect 24116 14216 24412 14236
rect 24268 13848 24320 13854
rect 24268 13790 24320 13796
rect 23900 13644 23952 13650
rect 23900 13586 23952 13592
rect 24280 13514 24308 13790
rect 23808 13508 23860 13514
rect 23808 13450 23860 13456
rect 24268 13508 24320 13514
rect 24268 13450 24320 13456
rect 24116 13204 24412 13224
rect 24172 13202 24196 13204
rect 24252 13202 24276 13204
rect 24332 13202 24356 13204
rect 24194 13150 24196 13202
rect 24258 13150 24270 13202
rect 24332 13150 24334 13202
rect 24172 13148 24196 13150
rect 24252 13148 24276 13150
rect 24332 13148 24356 13150
rect 24116 13128 24412 13148
rect 23900 12760 23952 12766
rect 23900 12702 23952 12708
rect 23532 12556 23584 12562
rect 23532 12498 23584 12504
rect 22244 12352 22296 12358
rect 22244 12294 22296 12300
rect 22520 12352 22572 12358
rect 22520 12294 22572 12300
rect 22152 12216 22204 12222
rect 22152 12158 22204 12164
rect 21692 11944 21744 11950
rect 21692 11886 21744 11892
rect 20680 11876 20732 11882
rect 20680 11818 20732 11824
rect 21508 11876 21560 11882
rect 21508 11818 21560 11824
rect 20956 11740 21008 11746
rect 20956 11682 21008 11688
rect 20404 11400 20456 11406
rect 20404 11342 20456 11348
rect 20968 11338 20996 11682
rect 21704 11338 21732 11886
rect 22164 11814 22192 12158
rect 22256 11950 22284 12294
rect 22244 11944 22296 11950
rect 22244 11886 22296 11892
rect 22152 11808 22204 11814
rect 22152 11750 22204 11756
rect 22532 11406 22560 12294
rect 23716 11672 23768 11678
rect 23716 11614 23768 11620
rect 22520 11400 22572 11406
rect 22520 11342 22572 11348
rect 20956 11332 21008 11338
rect 20956 11274 21008 11280
rect 21692 11332 21744 11338
rect 21692 11274 21744 11280
rect 21692 11196 21744 11202
rect 21692 11138 21744 11144
rect 21704 9624 21732 11138
rect 23728 9624 23756 11614
rect 23912 11338 23940 12702
rect 24116 12116 24412 12136
rect 24172 12114 24196 12116
rect 24252 12114 24276 12116
rect 24332 12114 24356 12116
rect 24194 12062 24196 12114
rect 24258 12062 24270 12114
rect 24332 12062 24334 12114
rect 24172 12060 24196 12062
rect 24252 12060 24276 12062
rect 24332 12060 24356 12062
rect 24116 12040 24412 12060
rect 24464 11678 24492 27050
rect 24636 25272 24688 25278
rect 24636 25214 24688 25220
rect 24544 24864 24596 24870
rect 24544 24806 24596 24812
rect 24556 23374 24584 24806
rect 24544 23368 24596 23374
rect 24544 23310 24596 23316
rect 24544 23232 24596 23238
rect 24544 23174 24596 23180
rect 24556 22694 24584 23174
rect 24544 22688 24596 22694
rect 24544 22630 24596 22636
rect 24648 21010 24676 25214
rect 24556 20982 24676 21010
rect 24556 20450 24584 20982
rect 24636 20920 24688 20926
rect 24636 20862 24688 20868
rect 24648 20518 24676 20862
rect 24636 20512 24688 20518
rect 24636 20454 24688 20460
rect 24544 20444 24596 20450
rect 24544 20386 24596 20392
rect 24636 20036 24688 20042
rect 24636 19978 24688 19984
rect 24648 19498 24676 19978
rect 24636 19492 24688 19498
rect 24636 19434 24688 19440
rect 24740 12902 24768 28206
rect 25292 27658 25320 28682
rect 25464 28672 25516 28678
rect 25464 28614 25516 28620
rect 25372 28128 25424 28134
rect 25372 28070 25424 28076
rect 25384 27998 25412 28070
rect 25372 27992 25424 27998
rect 25372 27934 25424 27940
rect 24912 27652 24964 27658
rect 24912 27594 24964 27600
rect 25280 27652 25332 27658
rect 25280 27594 25332 27600
rect 24924 27046 24952 27594
rect 25096 27516 25148 27522
rect 25148 27476 25228 27504
rect 25096 27458 25148 27464
rect 24912 27040 24964 27046
rect 24912 26982 24964 26988
rect 24924 26502 24952 26982
rect 24912 26496 24964 26502
rect 24912 26438 24964 26444
rect 24818 25512 24874 25521
rect 24818 25447 24820 25456
rect 24872 25447 24874 25456
rect 24820 25418 24872 25424
rect 24924 22694 24952 26438
rect 25004 25408 25056 25414
rect 25004 25350 25056 25356
rect 25016 24938 25044 25350
rect 25004 24932 25056 24938
rect 25004 24874 25056 24880
rect 25016 22762 25044 24874
rect 25096 23300 25148 23306
rect 25096 23242 25148 23248
rect 25108 22898 25136 23242
rect 25096 22892 25148 22898
rect 25096 22834 25148 22840
rect 25004 22756 25056 22762
rect 25004 22698 25056 22704
rect 24912 22688 24964 22694
rect 24912 22630 24964 22636
rect 24924 21266 24952 22630
rect 25108 22218 25136 22834
rect 25096 22212 25148 22218
rect 25096 22154 25148 22160
rect 24912 21260 24964 21266
rect 24912 21202 24964 21208
rect 24924 19906 24952 21202
rect 25200 21130 25228 27476
rect 25372 26020 25424 26026
rect 25372 25962 25424 25968
rect 25280 25952 25332 25958
rect 25280 25894 25332 25900
rect 25292 25618 25320 25894
rect 25280 25612 25332 25618
rect 25280 25554 25332 25560
rect 25384 24802 25412 25962
rect 25476 25618 25504 28614
rect 25832 27652 25884 27658
rect 25832 27594 25884 27600
rect 25740 27244 25792 27250
rect 25740 27186 25792 27192
rect 25556 27040 25608 27046
rect 25556 26982 25608 26988
rect 25568 26162 25596 26982
rect 25556 26156 25608 26162
rect 25556 26098 25608 26104
rect 25752 25958 25780 27186
rect 25844 27114 25872 27594
rect 25832 27108 25884 27114
rect 25832 27050 25884 27056
rect 25832 26564 25884 26570
rect 25936 26552 25964 31576
rect 26384 29828 26436 29834
rect 26384 29770 26436 29776
rect 26396 29154 26424 29770
rect 27488 29624 27540 29630
rect 27488 29566 27540 29572
rect 27396 29216 27448 29222
rect 27396 29158 27448 29164
rect 26384 29148 26436 29154
rect 26384 29090 26436 29096
rect 26292 29080 26344 29086
rect 26292 29022 26344 29028
rect 26304 28066 26332 29022
rect 26292 28060 26344 28066
rect 26292 28002 26344 28008
rect 26396 27998 26424 29090
rect 27120 29080 27172 29086
rect 27120 29022 27172 29028
rect 27212 29080 27264 29086
rect 27212 29022 27264 29028
rect 26384 27992 26436 27998
rect 26384 27934 26436 27940
rect 27028 27448 27080 27454
rect 27028 27390 27080 27396
rect 26384 27108 26436 27114
rect 26384 27050 26436 27056
rect 26396 26706 26424 27050
rect 26476 26904 26528 26910
rect 26476 26846 26528 26852
rect 26384 26700 26436 26706
rect 26384 26642 26436 26648
rect 26488 26570 26516 26846
rect 25884 26524 25964 26552
rect 26476 26564 26528 26570
rect 25832 26506 25884 26512
rect 26476 26506 26528 26512
rect 26384 26428 26436 26434
rect 26384 26370 26436 26376
rect 25740 25952 25792 25958
rect 25740 25894 25792 25900
rect 25464 25612 25516 25618
rect 25464 25554 25516 25560
rect 25752 25550 25780 25894
rect 25740 25544 25792 25550
rect 25740 25486 25792 25492
rect 25464 25476 25516 25482
rect 25464 25418 25516 25424
rect 25476 25074 25504 25418
rect 25924 25340 25976 25346
rect 25924 25282 25976 25288
rect 25464 25068 25516 25074
rect 25464 25010 25516 25016
rect 25556 25000 25608 25006
rect 25556 24942 25608 24948
rect 25372 24796 25424 24802
rect 25372 24738 25424 24744
rect 25384 22694 25412 24738
rect 25568 24394 25596 24942
rect 25936 24938 25964 25282
rect 26396 24954 26424 26370
rect 26488 26026 26516 26506
rect 27040 26026 27068 27390
rect 27132 26638 27160 29022
rect 27224 27114 27252 29022
rect 27408 28746 27436 29158
rect 27500 28814 27528 29566
rect 27776 28882 27804 31576
rect 29116 30068 29412 30088
rect 29172 30066 29196 30068
rect 29252 30066 29276 30068
rect 29332 30066 29356 30068
rect 29194 30014 29196 30066
rect 29258 30014 29270 30066
rect 29332 30014 29334 30066
rect 29172 30012 29196 30014
rect 29252 30012 29276 30014
rect 29332 30012 29356 30014
rect 29116 29992 29412 30012
rect 28958 29864 29014 29873
rect 28684 29828 28736 29834
rect 28958 29799 29014 29808
rect 28684 29770 28736 29776
rect 27764 28876 27816 28882
rect 27764 28818 27816 28824
rect 27488 28808 27540 28814
rect 27488 28750 27540 28756
rect 27396 28740 27448 28746
rect 27396 28682 27448 28688
rect 27856 28740 27908 28746
rect 27856 28682 27908 28688
rect 27396 28060 27448 28066
rect 27396 28002 27448 28008
rect 27408 27726 27436 28002
rect 27396 27720 27448 27726
rect 27396 27662 27448 27668
rect 27408 27182 27436 27662
rect 27764 27584 27816 27590
rect 27764 27526 27816 27532
rect 27396 27176 27448 27182
rect 27396 27118 27448 27124
rect 27212 27108 27264 27114
rect 27212 27050 27264 27056
rect 27776 26638 27804 27526
rect 27120 26632 27172 26638
rect 27120 26574 27172 26580
rect 27764 26632 27816 26638
rect 27764 26574 27816 26580
rect 27132 26094 27160 26574
rect 27580 26428 27632 26434
rect 27580 26370 27632 26376
rect 27120 26088 27172 26094
rect 27120 26030 27172 26036
rect 26476 26020 26528 26026
rect 26476 25962 26528 25968
rect 27028 26020 27080 26026
rect 27028 25962 27080 25968
rect 26936 25544 26988 25550
rect 26936 25486 26988 25492
rect 27026 25512 27082 25521
rect 25924 24932 25976 24938
rect 26396 24926 26516 24954
rect 25924 24874 25976 24880
rect 25556 24388 25608 24394
rect 25556 24330 25608 24336
rect 25936 23850 25964 24874
rect 26016 24864 26068 24870
rect 26016 24806 26068 24812
rect 26028 24394 26056 24806
rect 26488 24394 26516 24926
rect 26752 24932 26804 24938
rect 26752 24874 26804 24880
rect 26568 24728 26620 24734
rect 26568 24670 26620 24676
rect 26016 24388 26068 24394
rect 26016 24330 26068 24336
rect 26476 24388 26528 24394
rect 26476 24330 26528 24336
rect 26028 23918 26056 24330
rect 26108 24184 26160 24190
rect 26108 24126 26160 24132
rect 26016 23912 26068 23918
rect 26016 23854 26068 23860
rect 25924 23844 25976 23850
rect 25924 23786 25976 23792
rect 26120 23782 26148 24126
rect 26108 23776 26160 23782
rect 26108 23718 26160 23724
rect 26200 23640 26252 23646
rect 26200 23582 26252 23588
rect 26212 22762 26240 23582
rect 26200 22756 26252 22762
rect 26200 22698 26252 22704
rect 25372 22688 25424 22694
rect 25372 22630 25424 22636
rect 25280 22008 25332 22014
rect 25280 21950 25332 21956
rect 25188 21124 25240 21130
rect 25188 21066 25240 21072
rect 25200 20518 25228 21066
rect 25188 20512 25240 20518
rect 25188 20454 25240 20460
rect 24912 19900 24964 19906
rect 24912 19842 24964 19848
rect 25292 19566 25320 21950
rect 25280 19560 25332 19566
rect 25280 19502 25332 19508
rect 25004 18336 25056 18342
rect 25004 18278 25056 18284
rect 24820 18200 24872 18206
rect 24820 18142 24872 18148
rect 24832 16846 24860 18142
rect 25016 17934 25044 18278
rect 25004 17928 25056 17934
rect 25004 17870 25056 17876
rect 25016 17254 25044 17870
rect 25384 17322 25412 22630
rect 26212 22218 26240 22698
rect 26200 22212 26252 22218
rect 26200 22154 26252 22160
rect 26384 22212 26436 22218
rect 26384 22154 26436 22160
rect 26396 21606 26424 22154
rect 25556 21600 25608 21606
rect 25556 21542 25608 21548
rect 25648 21600 25700 21606
rect 25648 21542 25700 21548
rect 26384 21600 26436 21606
rect 26384 21542 26436 21548
rect 25568 21198 25596 21542
rect 25464 21192 25516 21198
rect 25464 21134 25516 21140
rect 25556 21192 25608 21198
rect 25556 21134 25608 21140
rect 25476 20194 25504 21134
rect 25568 20654 25596 21134
rect 25556 20648 25608 20654
rect 25556 20590 25608 20596
rect 25660 20586 25688 21542
rect 26580 21538 26608 24670
rect 26764 24462 26792 24874
rect 26752 24456 26804 24462
rect 26752 24398 26804 24404
rect 26948 24394 26976 25486
rect 27592 25482 27620 26370
rect 27026 25447 27082 25456
rect 27580 25476 27632 25482
rect 27040 25414 27068 25447
rect 27580 25418 27632 25424
rect 27028 25408 27080 25414
rect 27028 25350 27080 25356
rect 27028 24728 27080 24734
rect 27028 24670 27080 24676
rect 27212 24728 27264 24734
rect 27212 24670 27264 24676
rect 26844 24388 26896 24394
rect 26844 24330 26896 24336
rect 26936 24388 26988 24394
rect 26936 24330 26988 24336
rect 26856 24258 26884 24330
rect 26844 24252 26896 24258
rect 26844 24194 26896 24200
rect 26660 23096 26712 23102
rect 26660 23038 26712 23044
rect 26568 21532 26620 21538
rect 26568 21474 26620 21480
rect 25648 20580 25700 20586
rect 25648 20522 25700 20528
rect 26476 20512 26528 20518
rect 26476 20454 26528 20460
rect 25476 20166 25688 20194
rect 25556 20036 25608 20042
rect 25556 19978 25608 19984
rect 25464 19560 25516 19566
rect 25464 19502 25516 19508
rect 25476 19430 25504 19502
rect 25464 19424 25516 19430
rect 25464 19366 25516 19372
rect 25568 19362 25596 19978
rect 25556 19356 25608 19362
rect 25556 19298 25608 19304
rect 25568 18954 25596 19298
rect 25556 18948 25608 18954
rect 25556 18890 25608 18896
rect 25556 17724 25608 17730
rect 25556 17666 25608 17672
rect 25568 17390 25596 17666
rect 25556 17384 25608 17390
rect 25556 17326 25608 17332
rect 25372 17316 25424 17322
rect 25372 17258 25424 17264
rect 25004 17248 25056 17254
rect 25004 17190 25056 17196
rect 24820 16840 24872 16846
rect 24820 16782 24872 16788
rect 25372 16568 25424 16574
rect 25372 16510 25424 16516
rect 25384 16166 25412 16510
rect 25372 16160 25424 16166
rect 25372 16102 25424 16108
rect 25280 16024 25332 16030
rect 25280 15966 25332 15972
rect 25292 15078 25320 15966
rect 25556 15480 25608 15486
rect 25556 15422 25608 15428
rect 25568 15146 25596 15422
rect 25556 15140 25608 15146
rect 25556 15082 25608 15088
rect 25280 15072 25332 15078
rect 25280 15014 25332 15020
rect 25280 14596 25332 14602
rect 25280 14538 25332 14544
rect 25096 13984 25148 13990
rect 25096 13926 25148 13932
rect 24912 13916 24964 13922
rect 24912 13858 24964 13864
rect 24924 13310 24952 13858
rect 24912 13304 24964 13310
rect 24912 13246 24964 13252
rect 24924 12902 24952 13246
rect 25108 12902 25136 13926
rect 25188 13848 25240 13854
rect 25188 13790 25240 13796
rect 25200 12970 25228 13790
rect 25292 13446 25320 14538
rect 25464 14392 25516 14398
rect 25464 14334 25516 14340
rect 25476 14126 25504 14334
rect 25464 14120 25516 14126
rect 25464 14062 25516 14068
rect 25464 13984 25516 13990
rect 25464 13926 25516 13932
rect 25476 13514 25504 13926
rect 25464 13508 25516 13514
rect 25464 13450 25516 13456
rect 25280 13440 25332 13446
rect 25280 13382 25332 13388
rect 25292 13106 25320 13382
rect 25280 13100 25332 13106
rect 25280 13042 25332 13048
rect 25188 12964 25240 12970
rect 25188 12906 25240 12912
rect 24728 12896 24780 12902
rect 24728 12838 24780 12844
rect 24912 12896 24964 12902
rect 24912 12838 24964 12844
rect 25096 12896 25148 12902
rect 25096 12838 25148 12844
rect 25372 12760 25424 12766
rect 25372 12702 25424 12708
rect 25384 12494 25412 12702
rect 25372 12488 25424 12494
rect 25372 12430 25424 12436
rect 24452 11672 24504 11678
rect 24452 11614 24504 11620
rect 25384 11338 25412 12430
rect 25464 12420 25516 12426
rect 25464 12362 25516 12368
rect 25476 11882 25504 12362
rect 25464 11876 25516 11882
rect 25464 11818 25516 11824
rect 25660 11762 25688 20166
rect 26488 20110 26516 20454
rect 26476 20104 26528 20110
rect 26476 20046 26528 20052
rect 26016 19968 26068 19974
rect 26016 19910 26068 19916
rect 26028 19022 26056 19910
rect 26200 19900 26252 19906
rect 26200 19842 26252 19848
rect 26212 19430 26240 19842
rect 26488 19634 26516 20046
rect 26476 19628 26528 19634
rect 26476 19570 26528 19576
rect 26672 19566 26700 23038
rect 27040 22762 27068 24670
rect 27224 24530 27252 24670
rect 27212 24524 27264 24530
rect 27212 24466 27264 24472
rect 27764 24524 27816 24530
rect 27764 24466 27816 24472
rect 27776 23850 27804 24466
rect 27764 23844 27816 23850
rect 27764 23786 27816 23792
rect 27396 23776 27448 23782
rect 27396 23718 27448 23724
rect 27408 23306 27436 23718
rect 27396 23300 27448 23306
rect 27396 23242 27448 23248
rect 27028 22756 27080 22762
rect 27028 22698 27080 22704
rect 27396 22620 27448 22626
rect 27396 22562 27448 22568
rect 27408 22082 27436 22562
rect 27396 22076 27448 22082
rect 27396 22018 27448 22024
rect 27408 21538 27436 22018
rect 26752 21532 26804 21538
rect 26752 21474 26804 21480
rect 26844 21532 26896 21538
rect 26844 21474 26896 21480
rect 27396 21532 27448 21538
rect 27396 21474 27448 21480
rect 26764 21198 26792 21474
rect 26752 21192 26804 21198
rect 26752 21134 26804 21140
rect 26856 20994 26884 21474
rect 27212 21056 27264 21062
rect 27212 20998 27264 21004
rect 26844 20988 26896 20994
rect 26844 20930 26896 20936
rect 26856 20586 26884 20930
rect 27224 20722 27252 20998
rect 27212 20716 27264 20722
rect 27212 20658 27264 20664
rect 26844 20580 26896 20586
rect 26844 20522 26896 20528
rect 27304 20036 27356 20042
rect 27304 19978 27356 19984
rect 27316 19634 27344 19978
rect 27764 19832 27816 19838
rect 27764 19774 27816 19780
rect 27304 19628 27356 19634
rect 27304 19570 27356 19576
rect 26660 19560 26712 19566
rect 26660 19502 26712 19508
rect 26200 19424 26252 19430
rect 26200 19366 26252 19372
rect 26016 19016 26068 19022
rect 26016 18958 26068 18964
rect 26212 18206 26240 19366
rect 27028 19356 27080 19362
rect 27028 19298 27080 19304
rect 27040 19090 27068 19298
rect 27028 19084 27080 19090
rect 27028 19026 27080 19032
rect 26568 18880 26620 18886
rect 26568 18822 26620 18828
rect 26580 18342 26608 18822
rect 26936 18812 26988 18818
rect 26936 18754 26988 18760
rect 26948 18410 26976 18754
rect 27040 18410 27068 19026
rect 27776 19022 27804 19774
rect 27764 19016 27816 19022
rect 27764 18958 27816 18964
rect 27868 18818 27896 28682
rect 28592 28536 28644 28542
rect 28592 28478 28644 28484
rect 28224 28060 28276 28066
rect 28224 28002 28276 28008
rect 28236 27794 28264 28002
rect 28316 27992 28368 27998
rect 28316 27934 28368 27940
rect 28224 27788 28276 27794
rect 28224 27730 28276 27736
rect 28040 25952 28092 25958
rect 28040 25894 28092 25900
rect 27948 25612 28000 25618
rect 27948 25554 28000 25560
rect 27960 24870 27988 25554
rect 28052 25482 28080 25894
rect 28040 25476 28092 25482
rect 28040 25418 28092 25424
rect 28052 25074 28080 25418
rect 28040 25068 28092 25074
rect 28040 25010 28092 25016
rect 28328 25006 28356 27934
rect 28408 27652 28460 27658
rect 28408 27594 28460 27600
rect 28420 27114 28448 27594
rect 28408 27108 28460 27114
rect 28408 27050 28460 27056
rect 28500 26972 28552 26978
rect 28500 26914 28552 26920
rect 28512 26638 28540 26914
rect 28500 26632 28552 26638
rect 28500 26574 28552 26580
rect 28604 26450 28632 28478
rect 28512 26422 28632 26450
rect 28316 25000 28368 25006
rect 28316 24942 28368 24948
rect 27948 24864 28000 24870
rect 27948 24806 28000 24812
rect 28132 24796 28184 24802
rect 28132 24738 28184 24744
rect 28144 24394 28172 24738
rect 28132 24388 28184 24394
rect 28132 24330 28184 24336
rect 28328 24274 28356 24942
rect 28512 24394 28540 26422
rect 28696 26094 28724 29770
rect 28868 29624 28920 29630
rect 28868 29566 28920 29572
rect 28776 29080 28828 29086
rect 28776 29022 28828 29028
rect 28684 26088 28736 26094
rect 28684 26030 28736 26036
rect 28696 25550 28724 26030
rect 28788 26026 28816 29022
rect 28880 27114 28908 29566
rect 28972 28746 29000 29799
rect 29512 29216 29564 29222
rect 29512 29158 29564 29164
rect 29116 28980 29412 29000
rect 29172 28978 29196 28980
rect 29252 28978 29276 28980
rect 29332 28978 29356 28980
rect 29194 28926 29196 28978
rect 29258 28926 29270 28978
rect 29332 28926 29334 28978
rect 29172 28924 29196 28926
rect 29252 28924 29276 28926
rect 29332 28924 29356 28926
rect 29116 28904 29412 28924
rect 28960 28740 29012 28746
rect 28960 28682 29012 28688
rect 29116 27892 29412 27912
rect 29172 27890 29196 27892
rect 29252 27890 29276 27892
rect 29332 27890 29356 27892
rect 29194 27838 29196 27890
rect 29258 27838 29270 27890
rect 29332 27838 29334 27890
rect 29172 27836 29196 27838
rect 29252 27836 29276 27838
rect 29332 27836 29356 27838
rect 29116 27816 29412 27836
rect 29524 27658 29552 29158
rect 29616 28678 29644 31576
rect 29604 28672 29656 28678
rect 29604 28614 29656 28620
rect 29512 27652 29564 27658
rect 29512 27594 29564 27600
rect 29144 27516 29196 27522
rect 29144 27458 29196 27464
rect 28958 27416 29014 27425
rect 28958 27351 29014 27360
rect 28868 27108 28920 27114
rect 28868 27050 28920 27056
rect 28972 26570 29000 27351
rect 29156 26978 29184 27458
rect 29144 26972 29196 26978
rect 29144 26914 29196 26920
rect 29116 26804 29412 26824
rect 29172 26802 29196 26804
rect 29252 26802 29276 26804
rect 29332 26802 29356 26804
rect 29194 26750 29196 26802
rect 29258 26750 29270 26802
rect 29332 26750 29334 26802
rect 29172 26748 29196 26750
rect 29252 26748 29276 26750
rect 29332 26748 29356 26750
rect 29116 26728 29412 26748
rect 28960 26564 29012 26570
rect 28960 26506 29012 26512
rect 28776 26020 28828 26026
rect 28776 25962 28828 25968
rect 29116 25716 29412 25736
rect 29172 25714 29196 25716
rect 29252 25714 29276 25716
rect 29332 25714 29356 25716
rect 29194 25662 29196 25714
rect 29258 25662 29270 25714
rect 29332 25662 29334 25714
rect 29172 25660 29196 25662
rect 29252 25660 29276 25662
rect 29332 25660 29356 25662
rect 29116 25640 29412 25660
rect 29524 25550 29552 27594
rect 28684 25544 28736 25550
rect 28684 25486 28736 25492
rect 29512 25544 29564 25550
rect 29512 25486 29564 25492
rect 28960 24932 29012 24938
rect 28960 24874 29012 24880
rect 28592 24864 28644 24870
rect 28592 24806 28644 24812
rect 28500 24388 28552 24394
rect 28500 24330 28552 24336
rect 28236 24246 28356 24274
rect 28236 23306 28264 24246
rect 28500 24184 28552 24190
rect 28500 24126 28552 24132
rect 28512 23850 28540 24126
rect 28500 23844 28552 23850
rect 28500 23786 28552 23792
rect 28408 23708 28460 23714
rect 28408 23650 28460 23656
rect 28420 23374 28448 23650
rect 28408 23368 28460 23374
rect 28408 23310 28460 23316
rect 28224 23300 28276 23306
rect 28224 23242 28276 23248
rect 28236 22626 28264 23242
rect 28316 23164 28368 23170
rect 28316 23106 28368 23112
rect 28224 22620 28276 22626
rect 28224 22562 28276 22568
rect 27948 21600 28000 21606
rect 27948 21542 28000 21548
rect 27960 20518 27988 21542
rect 27948 20512 28000 20518
rect 27948 20454 28000 20460
rect 27960 20178 27988 20454
rect 27948 20172 28000 20178
rect 27948 20114 28000 20120
rect 27948 18948 28000 18954
rect 27948 18890 28000 18896
rect 27856 18812 27908 18818
rect 27856 18754 27908 18760
rect 26936 18404 26988 18410
rect 26936 18346 26988 18352
rect 27028 18404 27080 18410
rect 27028 18346 27080 18352
rect 27764 18404 27816 18410
rect 27764 18346 27816 18352
rect 26568 18336 26620 18342
rect 26568 18278 26620 18284
rect 26384 18268 26436 18274
rect 26384 18210 26436 18216
rect 26200 18200 26252 18206
rect 26200 18142 26252 18148
rect 26396 18154 26424 18210
rect 26396 18126 26516 18154
rect 25740 17792 25792 17798
rect 25740 17734 25792 17740
rect 25752 16914 25780 17734
rect 26488 17186 26516 18126
rect 26580 17934 26608 18278
rect 26660 18268 26712 18274
rect 26660 18210 26712 18216
rect 26568 17928 26620 17934
rect 26568 17870 26620 17876
rect 26672 17866 26700 18210
rect 26660 17860 26712 17866
rect 26660 17802 26712 17808
rect 27776 17730 27804 18346
rect 27764 17724 27816 17730
rect 27764 17666 27816 17672
rect 27120 17452 27172 17458
rect 27120 17394 27172 17400
rect 26476 17180 26528 17186
rect 26476 17122 26528 17128
rect 25740 16908 25792 16914
rect 25740 16850 25792 16856
rect 26488 16778 26516 17122
rect 25832 16772 25884 16778
rect 25832 16714 25884 16720
rect 26476 16772 26528 16778
rect 26476 16714 26528 16720
rect 25844 16166 25872 16714
rect 27132 16370 27160 17394
rect 27212 17248 27264 17254
rect 27212 17190 27264 17196
rect 27120 16364 27172 16370
rect 27120 16306 27172 16312
rect 25832 16160 25884 16166
rect 25832 16102 25884 16108
rect 27028 16160 27080 16166
rect 27028 16102 27080 16108
rect 26292 16024 26344 16030
rect 26292 15966 26344 15972
rect 25924 15684 25976 15690
rect 25924 15626 25976 15632
rect 26016 15684 26068 15690
rect 26016 15626 26068 15632
rect 25936 15146 25964 15626
rect 26028 15554 26056 15626
rect 26016 15548 26068 15554
rect 26016 15490 26068 15496
rect 25924 15140 25976 15146
rect 25924 15082 25976 15088
rect 25936 14738 25964 15082
rect 25924 14732 25976 14738
rect 25924 14674 25976 14680
rect 25924 14460 25976 14466
rect 25924 14402 25976 14408
rect 25936 12902 25964 14402
rect 26028 12902 26056 15490
rect 26304 15010 26332 15966
rect 26292 15004 26344 15010
rect 26292 14946 26344 14952
rect 26568 14936 26620 14942
rect 26568 14878 26620 14884
rect 26580 14534 26608 14878
rect 27040 14670 27068 16102
rect 27028 14664 27080 14670
rect 27028 14606 27080 14612
rect 26568 14528 26620 14534
rect 26568 14470 26620 14476
rect 26580 13514 26608 14470
rect 26568 13508 26620 13514
rect 26568 13450 26620 13456
rect 25924 12896 25976 12902
rect 25924 12838 25976 12844
rect 26016 12896 26068 12902
rect 26016 12838 26068 12844
rect 26384 12760 26436 12766
rect 26384 12702 26436 12708
rect 25740 12352 25792 12358
rect 25740 12294 25792 12300
rect 25752 11882 25780 12294
rect 25740 11876 25792 11882
rect 25740 11818 25792 11824
rect 26396 11814 26424 12702
rect 26580 12562 26608 13450
rect 27224 13281 27252 17190
rect 27776 16846 27804 17666
rect 27764 16840 27816 16846
rect 27764 16782 27816 16788
rect 27868 16250 27896 18754
rect 27960 18546 27988 18890
rect 27948 18540 28000 18546
rect 27948 18482 28000 18488
rect 28328 17254 28356 23106
rect 28604 22694 28632 24806
rect 28972 22694 29000 24874
rect 29116 24628 29412 24648
rect 29172 24626 29196 24628
rect 29252 24626 29276 24628
rect 29332 24626 29356 24628
rect 29194 24574 29196 24626
rect 29258 24574 29270 24626
rect 29332 24574 29334 24626
rect 29172 24572 29196 24574
rect 29252 24572 29276 24574
rect 29332 24572 29356 24574
rect 29116 24552 29412 24572
rect 29524 24530 29552 25486
rect 29512 24524 29564 24530
rect 29512 24466 29564 24472
rect 29328 24456 29380 24462
rect 29142 24424 29198 24433
rect 29328 24398 29380 24404
rect 29142 24359 29198 24368
rect 29156 23782 29184 24359
rect 29340 23986 29368 24398
rect 29512 24388 29564 24394
rect 29512 24330 29564 24336
rect 29328 23980 29380 23986
rect 29328 23922 29380 23928
rect 29144 23776 29196 23782
rect 29144 23718 29196 23724
rect 29116 23540 29412 23560
rect 29172 23538 29196 23540
rect 29252 23538 29276 23540
rect 29332 23538 29356 23540
rect 29194 23486 29196 23538
rect 29258 23486 29270 23538
rect 29332 23486 29334 23538
rect 29172 23484 29196 23486
rect 29252 23484 29276 23486
rect 29332 23484 29356 23486
rect 29116 23464 29412 23484
rect 28592 22688 28644 22694
rect 28592 22630 28644 22636
rect 28960 22688 29012 22694
rect 28960 22630 29012 22636
rect 28604 22286 28632 22630
rect 29116 22452 29412 22472
rect 29172 22450 29196 22452
rect 29252 22450 29276 22452
rect 29332 22450 29356 22452
rect 29194 22398 29196 22450
rect 29258 22398 29270 22450
rect 29332 22398 29334 22450
rect 29172 22396 29196 22398
rect 29252 22396 29276 22398
rect 29332 22396 29356 22398
rect 29116 22376 29412 22396
rect 28592 22280 28644 22286
rect 28592 22222 28644 22228
rect 29328 22144 29380 22150
rect 29328 22086 29380 22092
rect 29340 21713 29368 22086
rect 29326 21704 29382 21713
rect 29326 21639 29382 21648
rect 28776 21600 28828 21606
rect 28776 21542 28828 21548
rect 28592 21124 28644 21130
rect 28592 21066 28644 21072
rect 28604 20042 28632 21066
rect 28788 20450 28816 21542
rect 29116 21364 29412 21384
rect 29172 21362 29196 21364
rect 29252 21362 29276 21364
rect 29332 21362 29356 21364
rect 29194 21310 29196 21362
rect 29258 21310 29270 21362
rect 29332 21310 29334 21362
rect 29172 21308 29196 21310
rect 29252 21308 29276 21310
rect 29332 21308 29356 21310
rect 29116 21288 29412 21308
rect 29524 21198 29552 24330
rect 29880 22212 29932 22218
rect 29880 22154 29932 22160
rect 29696 21668 29748 21674
rect 29696 21610 29748 21616
rect 29604 21532 29656 21538
rect 29604 21474 29656 21480
rect 29512 21192 29564 21198
rect 29512 21134 29564 21140
rect 28776 20444 28828 20450
rect 28776 20386 28828 20392
rect 28592 20036 28644 20042
rect 28592 19978 28644 19984
rect 28604 19566 28632 19978
rect 28592 19560 28644 19566
rect 28592 19502 28644 19508
rect 28788 18342 28816 20386
rect 29116 20276 29412 20296
rect 29172 20274 29196 20276
rect 29252 20274 29276 20276
rect 29332 20274 29356 20276
rect 29194 20222 29196 20274
rect 29258 20222 29270 20274
rect 29332 20222 29334 20274
rect 29172 20220 29196 20222
rect 29252 20220 29276 20222
rect 29332 20220 29356 20222
rect 29116 20200 29412 20220
rect 29524 20110 29552 21134
rect 29616 21130 29644 21474
rect 29604 21124 29656 21130
rect 29604 21066 29656 21072
rect 29616 20450 29644 21066
rect 29604 20444 29656 20450
rect 29604 20386 29656 20392
rect 29512 20104 29564 20110
rect 29512 20046 29564 20052
rect 28868 19968 28920 19974
rect 28868 19910 28920 19916
rect 28880 18478 28908 19910
rect 29512 19424 29564 19430
rect 29512 19366 29564 19372
rect 29116 19188 29412 19208
rect 29172 19186 29196 19188
rect 29252 19186 29276 19188
rect 29332 19186 29356 19188
rect 29194 19134 29196 19186
rect 29258 19134 29270 19186
rect 29332 19134 29334 19186
rect 29172 19132 29196 19134
rect 29252 19132 29276 19134
rect 29332 19132 29356 19134
rect 29116 19112 29412 19132
rect 29524 18993 29552 19366
rect 29510 18984 29566 18993
rect 29616 18954 29644 20386
rect 29708 19090 29736 21610
rect 29892 19498 29920 22154
rect 29880 19492 29932 19498
rect 29880 19434 29932 19440
rect 29696 19084 29748 19090
rect 29696 19026 29748 19032
rect 29510 18919 29566 18928
rect 29604 18948 29656 18954
rect 29604 18890 29656 18896
rect 29696 18540 29748 18546
rect 29696 18482 29748 18488
rect 28868 18472 28920 18478
rect 28868 18414 28920 18420
rect 28776 18336 28828 18342
rect 28776 18278 28828 18284
rect 29116 18100 29412 18120
rect 29172 18098 29196 18100
rect 29252 18098 29276 18100
rect 29332 18098 29356 18100
rect 29194 18046 29196 18098
rect 29258 18046 29270 18098
rect 29332 18046 29334 18098
rect 29172 18044 29196 18046
rect 29252 18044 29276 18046
rect 29332 18044 29356 18046
rect 29116 18024 29412 18044
rect 29604 17928 29656 17934
rect 29604 17870 29656 17876
rect 28500 17860 28552 17866
rect 28500 17802 28552 17808
rect 28592 17860 28644 17866
rect 28592 17802 28644 17808
rect 28512 17322 28540 17802
rect 28500 17316 28552 17322
rect 28500 17258 28552 17264
rect 28316 17248 28368 17254
rect 28316 17190 28368 17196
rect 28512 16778 28540 17258
rect 28500 16772 28552 16778
rect 28500 16714 28552 16720
rect 28604 16658 28632 17802
rect 28960 17316 29012 17322
rect 28960 17258 29012 17264
rect 27776 16222 27896 16250
rect 28512 16630 28632 16658
rect 28776 16704 28828 16710
rect 28776 16646 28828 16652
rect 28868 16704 28920 16710
rect 28868 16646 28920 16652
rect 27776 15486 27804 16222
rect 27856 16160 27908 16166
rect 27856 16102 27908 16108
rect 27868 15486 27896 16102
rect 27948 16024 28000 16030
rect 27948 15966 28000 15972
rect 27960 15758 27988 15966
rect 27948 15752 28000 15758
rect 27948 15694 28000 15700
rect 27396 15480 27448 15486
rect 27396 15422 27448 15428
rect 27764 15480 27816 15486
rect 27764 15422 27816 15428
rect 27856 15480 27908 15486
rect 27856 15422 27908 15428
rect 27408 14534 27436 15422
rect 27764 15004 27816 15010
rect 27764 14946 27816 14952
rect 27776 14670 27804 14946
rect 27764 14664 27816 14670
rect 27764 14606 27816 14612
rect 27396 14528 27448 14534
rect 27396 14470 27448 14476
rect 27776 14210 27804 14606
rect 27868 14398 27896 15422
rect 27948 15072 28000 15078
rect 27948 15014 28000 15020
rect 27960 14738 27988 15014
rect 27948 14732 28000 14738
rect 27948 14674 28000 14680
rect 27856 14392 27908 14398
rect 27856 14334 27908 14340
rect 27776 14182 27896 14210
rect 27868 13922 27896 14182
rect 27960 14058 27988 14674
rect 28224 14528 28276 14534
rect 28224 14470 28276 14476
rect 28236 14194 28264 14470
rect 28224 14188 28276 14194
rect 28224 14130 28276 14136
rect 27948 14052 28000 14058
rect 27948 13994 28000 14000
rect 28512 13990 28540 16630
rect 28592 16024 28644 16030
rect 28592 15966 28644 15972
rect 28684 16024 28736 16030
rect 28684 15966 28736 15972
rect 28604 15078 28632 15966
rect 28696 15758 28724 15966
rect 28684 15752 28736 15758
rect 28684 15694 28736 15700
rect 28592 15072 28644 15078
rect 28592 15014 28644 15020
rect 28500 13984 28552 13990
rect 28500 13926 28552 13932
rect 27856 13916 27908 13922
rect 27856 13858 27908 13864
rect 27488 13440 27540 13446
rect 27488 13382 27540 13388
rect 27210 13272 27266 13281
rect 27210 13207 27266 13216
rect 27396 12964 27448 12970
rect 27396 12906 27448 12912
rect 26568 12556 26620 12562
rect 26568 12498 26620 12504
rect 26476 12488 26528 12494
rect 26476 12430 26528 12436
rect 26488 12018 26516 12430
rect 26476 12012 26528 12018
rect 26476 11954 26528 11960
rect 26384 11808 26436 11814
rect 25556 11740 25608 11746
rect 25660 11734 25780 11762
rect 26384 11750 26436 11756
rect 25556 11682 25608 11688
rect 25568 11474 25596 11682
rect 25556 11468 25608 11474
rect 25556 11410 25608 11416
rect 23900 11332 23952 11338
rect 23900 11274 23952 11280
rect 25372 11332 25424 11338
rect 25372 11274 25424 11280
rect 24116 11028 24412 11048
rect 24172 11026 24196 11028
rect 24252 11026 24276 11028
rect 24332 11026 24356 11028
rect 24194 10974 24196 11026
rect 24258 10974 24270 11026
rect 24332 10974 24334 11026
rect 24172 10972 24196 10974
rect 24252 10972 24276 10974
rect 24332 10972 24356 10974
rect 24116 10952 24412 10972
rect 25752 10130 25780 11734
rect 25568 10102 25780 10130
rect 25568 9624 25596 10102
rect 27408 9624 27436 12906
rect 27500 12494 27528 13382
rect 27764 12828 27816 12834
rect 27764 12770 27816 12776
rect 27488 12488 27540 12494
rect 27488 12430 27540 12436
rect 27500 11814 27528 12430
rect 27488 11808 27540 11814
rect 27488 11750 27540 11756
rect 27776 10561 27804 12770
rect 27868 12562 27896 13858
rect 28132 13576 28184 13582
rect 28132 13518 28184 13524
rect 28144 13106 28172 13518
rect 28592 13440 28644 13446
rect 28592 13382 28644 13388
rect 28132 13100 28184 13106
rect 28132 13042 28184 13048
rect 27856 12556 27908 12562
rect 27856 12498 27908 12504
rect 28040 12488 28092 12494
rect 28040 12430 28092 12436
rect 28052 12018 28080 12430
rect 28604 12426 28632 13382
rect 28788 12970 28816 16646
rect 28880 14194 28908 16646
rect 28972 16273 29000 17258
rect 29116 17012 29412 17032
rect 29172 17010 29196 17012
rect 29252 17010 29276 17012
rect 29332 17010 29356 17012
rect 29194 16958 29196 17010
rect 29258 16958 29270 17010
rect 29332 16958 29334 17010
rect 29172 16956 29196 16958
rect 29252 16956 29276 16958
rect 29332 16956 29356 16958
rect 29116 16936 29412 16956
rect 29616 16642 29644 17870
rect 29604 16636 29656 16642
rect 29604 16578 29656 16584
rect 28958 16264 29014 16273
rect 28958 16199 29014 16208
rect 28960 16160 29012 16166
rect 28960 16102 29012 16108
rect 28868 14188 28920 14194
rect 28868 14130 28920 14136
rect 28972 13514 29000 16102
rect 29116 15924 29412 15944
rect 29172 15922 29196 15924
rect 29252 15922 29276 15924
rect 29332 15922 29356 15924
rect 29194 15870 29196 15922
rect 29258 15870 29270 15922
rect 29332 15870 29334 15922
rect 29172 15868 29196 15870
rect 29252 15868 29276 15870
rect 29332 15868 29356 15870
rect 29116 15848 29412 15868
rect 29144 15616 29196 15622
rect 29144 15558 29196 15564
rect 29156 15282 29184 15558
rect 29144 15276 29196 15282
rect 29144 15218 29196 15224
rect 29116 14836 29412 14856
rect 29172 14834 29196 14836
rect 29252 14834 29276 14836
rect 29332 14834 29356 14836
rect 29194 14782 29196 14834
rect 29258 14782 29270 14834
rect 29332 14782 29334 14834
rect 29172 14780 29196 14782
rect 29252 14780 29276 14782
rect 29332 14780 29356 14782
rect 29116 14760 29412 14780
rect 29512 14664 29564 14670
rect 29512 14606 29564 14612
rect 29116 13748 29412 13768
rect 29172 13746 29196 13748
rect 29252 13746 29276 13748
rect 29332 13746 29356 13748
rect 29194 13694 29196 13746
rect 29258 13694 29270 13746
rect 29332 13694 29334 13746
rect 29172 13692 29196 13694
rect 29252 13692 29276 13694
rect 29332 13692 29356 13694
rect 29116 13672 29412 13692
rect 29524 13650 29552 14606
rect 29512 13644 29564 13650
rect 29512 13586 29564 13592
rect 28960 13508 29012 13514
rect 28960 13450 29012 13456
rect 28776 12964 28828 12970
rect 28776 12906 28828 12912
rect 28972 12834 29000 13450
rect 29616 12902 29644 16578
rect 29604 12896 29656 12902
rect 29604 12838 29656 12844
rect 28960 12828 29012 12834
rect 28960 12770 29012 12776
rect 29708 12714 29736 18482
rect 29892 18274 29920 19434
rect 29972 19356 30024 19362
rect 29972 19298 30024 19304
rect 29984 18546 30012 19298
rect 29972 18540 30024 18546
rect 29972 18482 30024 18488
rect 29880 18268 29932 18274
rect 29880 18210 29932 18216
rect 29892 17254 29920 18210
rect 29880 17248 29932 17254
rect 29880 17190 29932 17196
rect 29524 12686 29736 12714
rect 29116 12660 29412 12680
rect 29172 12658 29196 12660
rect 29252 12658 29276 12660
rect 29332 12658 29356 12660
rect 29194 12606 29196 12658
rect 29258 12606 29270 12658
rect 29332 12606 29334 12658
rect 29172 12604 29196 12606
rect 29252 12604 29276 12606
rect 29332 12604 29356 12606
rect 29116 12584 29412 12604
rect 28592 12420 28644 12426
rect 28592 12362 28644 12368
rect 28040 12012 28092 12018
rect 28040 11954 28092 11960
rect 29116 11572 29412 11592
rect 29172 11570 29196 11572
rect 29252 11570 29276 11572
rect 29332 11570 29356 11572
rect 29194 11518 29196 11570
rect 29258 11518 29270 11570
rect 29332 11518 29334 11570
rect 29172 11516 29196 11518
rect 29252 11516 29276 11518
rect 29332 11516 29356 11518
rect 29116 11496 29412 11516
rect 27762 10552 27818 10561
rect 27762 10487 27818 10496
rect 29524 9722 29552 12686
rect 29432 9694 29552 9722
rect 29432 9624 29460 9694
rect 10466 8824 10522 9624
rect 12306 8824 12362 9624
rect 14146 8824 14202 9624
rect 15986 8824 16042 9624
rect 18010 8824 18066 9624
rect 19850 8824 19906 9624
rect 21690 8824 21746 9624
rect 23714 8824 23770 9624
rect 25554 8824 25610 9624
rect 27394 8824 27450 9624
rect 29418 8824 29474 9624
<< via2 >>
rect 14116 29522 14172 29524
rect 14196 29522 14252 29524
rect 14276 29522 14332 29524
rect 14356 29522 14412 29524
rect 14116 29470 14142 29522
rect 14142 29470 14172 29522
rect 14196 29470 14206 29522
rect 14206 29470 14252 29522
rect 14276 29470 14322 29522
rect 14322 29470 14332 29522
rect 14356 29470 14386 29522
rect 14386 29470 14412 29522
rect 14116 29468 14172 29470
rect 14196 29468 14252 29470
rect 14276 29468 14332 29470
rect 14356 29468 14412 29470
rect 13502 29284 13558 29320
rect 13502 29264 13504 29284
rect 13504 29264 13556 29284
rect 13556 29264 13558 29284
rect 14116 28434 14172 28436
rect 14196 28434 14252 28436
rect 14276 28434 14332 28436
rect 14356 28434 14412 28436
rect 14116 28382 14142 28434
rect 14142 28382 14172 28434
rect 14196 28382 14206 28434
rect 14206 28382 14252 28434
rect 14276 28382 14322 28434
rect 14322 28382 14332 28434
rect 14356 28382 14386 28434
rect 14386 28382 14412 28434
rect 14116 28380 14172 28382
rect 14196 28380 14252 28382
rect 14276 28380 14332 28382
rect 14356 28380 14412 28382
rect 19116 30066 19172 30068
rect 19196 30066 19252 30068
rect 19276 30066 19332 30068
rect 19356 30066 19412 30068
rect 19116 30014 19142 30066
rect 19142 30014 19172 30066
rect 19196 30014 19206 30066
rect 19206 30014 19252 30066
rect 19276 30014 19322 30066
rect 19322 30014 19332 30066
rect 19356 30014 19386 30066
rect 19386 30014 19412 30066
rect 19116 30012 19172 30014
rect 19196 30012 19252 30014
rect 19276 30012 19332 30014
rect 19356 30012 19412 30014
rect 11662 26272 11718 26328
rect 19116 28978 19172 28980
rect 19196 28978 19252 28980
rect 19276 28978 19332 28980
rect 19356 28978 19412 28980
rect 19116 28926 19142 28978
rect 19142 28926 19172 28978
rect 19196 28926 19206 28978
rect 19206 28926 19252 28978
rect 19276 28926 19322 28978
rect 19322 28926 19332 28978
rect 19356 28926 19386 28978
rect 19386 28926 19412 28978
rect 19116 28924 19172 28926
rect 19196 28924 19252 28926
rect 19276 28924 19332 28926
rect 19356 28924 19412 28926
rect 19116 27890 19172 27892
rect 19196 27890 19252 27892
rect 19276 27890 19332 27892
rect 19356 27890 19412 27892
rect 19116 27838 19142 27890
rect 19142 27838 19172 27890
rect 19196 27838 19206 27890
rect 19206 27838 19252 27890
rect 19276 27838 19322 27890
rect 19322 27838 19332 27890
rect 19356 27838 19386 27890
rect 19386 27838 19412 27890
rect 19116 27836 19172 27838
rect 19196 27836 19252 27838
rect 19276 27836 19332 27838
rect 19356 27836 19412 27838
rect 14116 27346 14172 27348
rect 14196 27346 14252 27348
rect 14276 27346 14332 27348
rect 14356 27346 14412 27348
rect 14116 27294 14142 27346
rect 14142 27294 14172 27346
rect 14196 27294 14206 27346
rect 14206 27294 14252 27346
rect 14276 27294 14322 27346
rect 14322 27294 14332 27346
rect 14356 27294 14386 27346
rect 14386 27294 14412 27346
rect 14116 27292 14172 27294
rect 14196 27292 14252 27294
rect 14276 27292 14332 27294
rect 14356 27292 14412 27294
rect 11662 20832 11718 20888
rect 14116 26258 14172 26260
rect 14196 26258 14252 26260
rect 14276 26258 14332 26260
rect 14356 26258 14412 26260
rect 14116 26206 14142 26258
rect 14142 26206 14172 26258
rect 14196 26206 14206 26258
rect 14206 26206 14252 26258
rect 14276 26206 14322 26258
rect 14322 26206 14332 26258
rect 14356 26206 14386 26258
rect 14386 26206 14412 26258
rect 14116 26204 14172 26206
rect 14196 26204 14252 26206
rect 14276 26204 14332 26206
rect 14356 26204 14412 26206
rect 14116 25170 14172 25172
rect 14196 25170 14252 25172
rect 14276 25170 14332 25172
rect 14356 25170 14412 25172
rect 14116 25118 14142 25170
rect 14142 25118 14172 25170
rect 14196 25118 14206 25170
rect 14206 25118 14252 25170
rect 14276 25118 14322 25170
rect 14322 25118 14332 25170
rect 14356 25118 14386 25170
rect 14386 25118 14412 25170
rect 14116 25116 14172 25118
rect 14196 25116 14252 25118
rect 14276 25116 14332 25118
rect 14356 25116 14412 25118
rect 14116 24082 14172 24084
rect 14196 24082 14252 24084
rect 14276 24082 14332 24084
rect 14356 24082 14412 24084
rect 14116 24030 14142 24082
rect 14142 24030 14172 24082
rect 14196 24030 14206 24082
rect 14206 24030 14252 24082
rect 14276 24030 14322 24082
rect 14322 24030 14332 24082
rect 14356 24030 14386 24082
rect 14386 24030 14412 24082
rect 14116 24028 14172 24030
rect 14196 24028 14252 24030
rect 14276 24028 14332 24030
rect 14356 24028 14412 24030
rect 13870 23552 13926 23608
rect 12674 17840 12730 17896
rect 14116 22994 14172 22996
rect 14196 22994 14252 22996
rect 14276 22994 14332 22996
rect 14356 22994 14412 22996
rect 14116 22942 14142 22994
rect 14142 22942 14172 22994
rect 14196 22942 14206 22994
rect 14206 22942 14252 22994
rect 14276 22942 14322 22994
rect 14322 22942 14332 22994
rect 14356 22942 14386 22994
rect 14386 22942 14412 22994
rect 14116 22940 14172 22942
rect 14196 22940 14252 22942
rect 14276 22940 14332 22942
rect 14356 22940 14412 22942
rect 14116 21906 14172 21908
rect 14196 21906 14252 21908
rect 14276 21906 14332 21908
rect 14356 21906 14412 21908
rect 14116 21854 14142 21906
rect 14142 21854 14172 21906
rect 14196 21854 14206 21906
rect 14206 21854 14252 21906
rect 14276 21854 14322 21906
rect 14322 21854 14332 21906
rect 14356 21854 14386 21906
rect 14386 21854 14412 21906
rect 14116 21852 14172 21854
rect 14196 21852 14252 21854
rect 14276 21852 14332 21854
rect 14356 21852 14412 21854
rect 15802 24812 15804 24832
rect 15804 24812 15856 24832
rect 15856 24812 15858 24832
rect 15802 24776 15858 24812
rect 14116 20818 14172 20820
rect 14196 20818 14252 20820
rect 14276 20818 14332 20820
rect 14356 20818 14412 20820
rect 14116 20766 14142 20818
rect 14142 20766 14172 20818
rect 14196 20766 14206 20818
rect 14206 20766 14252 20818
rect 14276 20766 14322 20818
rect 14322 20766 14332 20818
rect 14356 20766 14386 20818
rect 14386 20766 14412 20818
rect 14116 20764 14172 20766
rect 14196 20764 14252 20766
rect 14276 20764 14332 20766
rect 14356 20764 14412 20766
rect 14116 19730 14172 19732
rect 14196 19730 14252 19732
rect 14276 19730 14332 19732
rect 14356 19730 14412 19732
rect 14116 19678 14142 19730
rect 14142 19678 14172 19730
rect 14196 19678 14206 19730
rect 14206 19678 14252 19730
rect 14276 19678 14322 19730
rect 14322 19678 14332 19730
rect 14356 19678 14386 19730
rect 14386 19678 14412 19730
rect 14116 19676 14172 19678
rect 14196 19676 14252 19678
rect 14276 19676 14332 19678
rect 14356 19676 14412 19678
rect 14116 18642 14172 18644
rect 14196 18642 14252 18644
rect 14276 18642 14332 18644
rect 14356 18642 14412 18644
rect 14116 18590 14142 18642
rect 14142 18590 14172 18642
rect 14196 18590 14206 18642
rect 14206 18590 14252 18642
rect 14276 18590 14322 18642
rect 14322 18590 14332 18642
rect 14356 18590 14386 18642
rect 14386 18590 14412 18642
rect 14116 18588 14172 18590
rect 14196 18588 14252 18590
rect 14276 18588 14332 18590
rect 14356 18588 14412 18590
rect 14116 17554 14172 17556
rect 14196 17554 14252 17556
rect 14276 17554 14332 17556
rect 14356 17554 14412 17556
rect 14116 17502 14142 17554
rect 14142 17502 14172 17554
rect 14196 17502 14206 17554
rect 14206 17502 14252 17554
rect 14276 17502 14322 17554
rect 14322 17502 14332 17554
rect 14356 17502 14386 17554
rect 14386 17502 14412 17554
rect 14116 17500 14172 17502
rect 14196 17500 14252 17502
rect 14276 17500 14332 17502
rect 14356 17500 14412 17502
rect 14116 16466 14172 16468
rect 14196 16466 14252 16468
rect 14276 16466 14332 16468
rect 14356 16466 14412 16468
rect 14116 16414 14142 16466
rect 14142 16414 14172 16466
rect 14196 16414 14206 16466
rect 14206 16414 14252 16466
rect 14276 16414 14322 16466
rect 14322 16414 14332 16466
rect 14356 16414 14386 16466
rect 14386 16414 14412 16466
rect 14116 16412 14172 16414
rect 14196 16412 14252 16414
rect 14276 16412 14332 16414
rect 14356 16412 14412 16414
rect 19116 26802 19172 26804
rect 19196 26802 19252 26804
rect 19276 26802 19332 26804
rect 19356 26802 19412 26804
rect 19116 26750 19142 26802
rect 19142 26750 19172 26802
rect 19196 26750 19206 26802
rect 19206 26750 19252 26802
rect 19276 26750 19322 26802
rect 19322 26750 19332 26802
rect 19356 26750 19386 26802
rect 19386 26750 19412 26802
rect 19116 26748 19172 26750
rect 19196 26748 19252 26750
rect 19276 26748 19332 26750
rect 19356 26748 19412 26750
rect 19116 25714 19172 25716
rect 19196 25714 19252 25716
rect 19276 25714 19332 25716
rect 19356 25714 19412 25716
rect 19116 25662 19142 25714
rect 19142 25662 19172 25714
rect 19196 25662 19206 25714
rect 19206 25662 19252 25714
rect 19276 25662 19322 25714
rect 19322 25662 19332 25714
rect 19356 25662 19386 25714
rect 19386 25662 19412 25714
rect 19116 25660 19172 25662
rect 19196 25660 19252 25662
rect 19276 25660 19332 25662
rect 19356 25660 19412 25662
rect 19022 24776 19078 24832
rect 19116 24626 19172 24628
rect 19196 24626 19252 24628
rect 19276 24626 19332 24628
rect 19356 24626 19412 24628
rect 19116 24574 19142 24626
rect 19142 24574 19172 24626
rect 19196 24574 19206 24626
rect 19206 24574 19252 24626
rect 19276 24574 19322 24626
rect 19322 24574 19332 24626
rect 19356 24574 19386 24626
rect 19386 24574 19412 24626
rect 19116 24572 19172 24574
rect 19196 24572 19252 24574
rect 19276 24572 19332 24574
rect 19356 24572 19412 24574
rect 19116 23538 19172 23540
rect 19196 23538 19252 23540
rect 19276 23538 19332 23540
rect 19356 23538 19412 23540
rect 19116 23486 19142 23538
rect 19142 23486 19172 23538
rect 19196 23486 19206 23538
rect 19206 23486 19252 23538
rect 19276 23486 19322 23538
rect 19322 23486 19332 23538
rect 19356 23486 19386 23538
rect 19386 23486 19412 23538
rect 19116 23484 19172 23486
rect 19196 23484 19252 23486
rect 19276 23484 19332 23486
rect 19356 23484 19412 23486
rect 19116 22450 19172 22452
rect 19196 22450 19252 22452
rect 19276 22450 19332 22452
rect 19356 22450 19412 22452
rect 19116 22398 19142 22450
rect 19142 22398 19172 22450
rect 19196 22398 19206 22450
rect 19206 22398 19252 22450
rect 19276 22398 19322 22450
rect 19322 22398 19332 22450
rect 19356 22398 19386 22450
rect 19386 22398 19412 22450
rect 19116 22396 19172 22398
rect 19196 22396 19252 22398
rect 19276 22396 19332 22398
rect 19356 22396 19412 22398
rect 18194 20016 18250 20072
rect 19116 21362 19172 21364
rect 19196 21362 19252 21364
rect 19276 21362 19332 21364
rect 19356 21362 19412 21364
rect 19116 21310 19142 21362
rect 19142 21310 19172 21362
rect 19196 21310 19206 21362
rect 19206 21310 19252 21362
rect 19276 21310 19322 21362
rect 19322 21310 19332 21362
rect 19356 21310 19386 21362
rect 19386 21310 19412 21362
rect 19116 21308 19172 21310
rect 19196 21308 19252 21310
rect 19276 21308 19332 21310
rect 19356 21308 19412 21310
rect 19116 20274 19172 20276
rect 19196 20274 19252 20276
rect 19276 20274 19332 20276
rect 19356 20274 19412 20276
rect 19116 20222 19142 20274
rect 19142 20222 19172 20274
rect 19196 20222 19206 20274
rect 19206 20222 19252 20274
rect 19276 20222 19322 20274
rect 19322 20222 19332 20274
rect 19356 20222 19386 20274
rect 19386 20222 19412 20274
rect 19116 20220 19172 20222
rect 19196 20220 19252 20222
rect 19276 20220 19332 20222
rect 19356 20220 19412 20222
rect 19942 20052 19944 20072
rect 19944 20052 19996 20072
rect 19996 20052 19998 20072
rect 19116 19186 19172 19188
rect 19196 19186 19252 19188
rect 19276 19186 19332 19188
rect 19356 19186 19412 19188
rect 19116 19134 19142 19186
rect 19142 19134 19172 19186
rect 19196 19134 19206 19186
rect 19206 19134 19252 19186
rect 19276 19134 19322 19186
rect 19322 19134 19332 19186
rect 19356 19134 19386 19186
rect 19386 19134 19412 19186
rect 19116 19132 19172 19134
rect 19196 19132 19252 19134
rect 19276 19132 19332 19134
rect 19356 19132 19412 19134
rect 19942 20016 19998 20052
rect 14116 15378 14172 15380
rect 14196 15378 14252 15380
rect 14276 15378 14332 15380
rect 14356 15378 14412 15380
rect 14116 15326 14142 15378
rect 14142 15326 14172 15378
rect 14196 15326 14206 15378
rect 14206 15326 14252 15378
rect 14276 15326 14322 15378
rect 14322 15326 14332 15378
rect 14356 15326 14386 15378
rect 14386 15326 14412 15378
rect 14116 15324 14172 15326
rect 14196 15324 14252 15326
rect 14276 15324 14332 15326
rect 14356 15324 14412 15326
rect 13962 15120 14018 15176
rect 14116 14290 14172 14292
rect 14196 14290 14252 14292
rect 14276 14290 14332 14292
rect 14356 14290 14412 14292
rect 14116 14238 14142 14290
rect 14142 14238 14172 14290
rect 14196 14238 14206 14290
rect 14206 14238 14252 14290
rect 14276 14238 14322 14290
rect 14322 14238 14332 14290
rect 14356 14238 14386 14290
rect 14386 14238 14412 14290
rect 14116 14236 14172 14238
rect 14196 14236 14252 14238
rect 14276 14236 14332 14238
rect 14356 14236 14412 14238
rect 12030 12420 12086 12456
rect 12030 12400 12032 12420
rect 12032 12400 12084 12420
rect 12084 12400 12086 12420
rect 14116 13202 14172 13204
rect 14196 13202 14252 13204
rect 14276 13202 14332 13204
rect 14356 13202 14412 13204
rect 14116 13150 14142 13202
rect 14142 13150 14172 13202
rect 14196 13150 14206 13202
rect 14206 13150 14252 13202
rect 14276 13150 14322 13202
rect 14322 13150 14332 13202
rect 14356 13150 14386 13202
rect 14386 13150 14412 13202
rect 14116 13148 14172 13150
rect 14196 13148 14252 13150
rect 14276 13148 14332 13150
rect 14356 13148 14412 13150
rect 14116 12114 14172 12116
rect 14196 12114 14252 12116
rect 14276 12114 14332 12116
rect 14356 12114 14412 12116
rect 14116 12062 14142 12114
rect 14142 12062 14172 12114
rect 14196 12062 14206 12114
rect 14206 12062 14252 12114
rect 14276 12062 14322 12114
rect 14322 12062 14332 12114
rect 14356 12062 14386 12114
rect 14386 12062 14412 12114
rect 14116 12060 14172 12062
rect 14196 12060 14252 12062
rect 14276 12060 14332 12062
rect 14356 12060 14412 12062
rect 14116 11026 14172 11028
rect 14196 11026 14252 11028
rect 14276 11026 14332 11028
rect 14356 11026 14412 11028
rect 14116 10974 14142 11026
rect 14142 10974 14172 11026
rect 14196 10974 14206 11026
rect 14206 10974 14252 11026
rect 14276 10974 14322 11026
rect 14322 10974 14332 11026
rect 14356 10974 14386 11026
rect 14386 10974 14412 11026
rect 14116 10972 14172 10974
rect 14196 10972 14252 10974
rect 14276 10972 14332 10974
rect 14356 10972 14412 10974
rect 19116 18098 19172 18100
rect 19196 18098 19252 18100
rect 19276 18098 19332 18100
rect 19356 18098 19412 18100
rect 19116 18046 19142 18098
rect 19142 18046 19172 18098
rect 19196 18046 19206 18098
rect 19206 18046 19252 18098
rect 19276 18046 19322 18098
rect 19322 18046 19332 18098
rect 19356 18046 19386 18098
rect 19386 18046 19412 18098
rect 19116 18044 19172 18046
rect 19196 18044 19252 18046
rect 19276 18044 19332 18046
rect 19356 18044 19412 18046
rect 24116 29522 24172 29524
rect 24196 29522 24252 29524
rect 24276 29522 24332 29524
rect 24356 29522 24412 29524
rect 24116 29470 24142 29522
rect 24142 29470 24172 29522
rect 24196 29470 24206 29522
rect 24206 29470 24252 29522
rect 24276 29470 24322 29522
rect 24322 29470 24332 29522
rect 24356 29470 24386 29522
rect 24386 29470 24412 29522
rect 24116 29468 24172 29470
rect 24196 29468 24252 29470
rect 24276 29468 24332 29470
rect 24356 29468 24412 29470
rect 24116 28434 24172 28436
rect 24196 28434 24252 28436
rect 24276 28434 24332 28436
rect 24356 28434 24412 28436
rect 24116 28382 24142 28434
rect 24142 28382 24172 28434
rect 24196 28382 24206 28434
rect 24206 28382 24252 28434
rect 24276 28382 24322 28434
rect 24322 28382 24332 28434
rect 24356 28382 24386 28434
rect 24386 28382 24412 28434
rect 24116 28380 24172 28382
rect 24196 28380 24252 28382
rect 24276 28380 24332 28382
rect 24356 28380 24412 28382
rect 24116 27346 24172 27348
rect 24196 27346 24252 27348
rect 24276 27346 24332 27348
rect 24356 27346 24412 27348
rect 24116 27294 24142 27346
rect 24142 27294 24172 27346
rect 24196 27294 24206 27346
rect 24206 27294 24252 27346
rect 24276 27294 24322 27346
rect 24322 27294 24332 27346
rect 24356 27294 24386 27346
rect 24386 27294 24412 27346
rect 24116 27292 24172 27294
rect 24196 27292 24252 27294
rect 24276 27292 24332 27294
rect 24356 27292 24412 27294
rect 19116 17010 19172 17012
rect 19196 17010 19252 17012
rect 19276 17010 19332 17012
rect 19356 17010 19412 17012
rect 19116 16958 19142 17010
rect 19142 16958 19172 17010
rect 19196 16958 19206 17010
rect 19206 16958 19252 17010
rect 19276 16958 19322 17010
rect 19322 16958 19332 17010
rect 19356 16958 19386 17010
rect 19386 16958 19412 17010
rect 19116 16956 19172 16958
rect 19196 16956 19252 16958
rect 19276 16956 19332 16958
rect 19356 16956 19412 16958
rect 19116 15922 19172 15924
rect 19196 15922 19252 15924
rect 19276 15922 19332 15924
rect 19356 15922 19412 15924
rect 19116 15870 19142 15922
rect 19142 15870 19172 15922
rect 19196 15870 19206 15922
rect 19206 15870 19252 15922
rect 19276 15870 19322 15922
rect 19322 15870 19332 15922
rect 19356 15870 19386 15922
rect 19386 15870 19412 15922
rect 19116 15868 19172 15870
rect 19196 15868 19252 15870
rect 19276 15868 19332 15870
rect 19356 15868 19412 15870
rect 19116 14834 19172 14836
rect 19196 14834 19252 14836
rect 19276 14834 19332 14836
rect 19356 14834 19412 14836
rect 19116 14782 19142 14834
rect 19142 14782 19172 14834
rect 19196 14782 19206 14834
rect 19206 14782 19252 14834
rect 19276 14782 19322 14834
rect 19322 14782 19332 14834
rect 19356 14782 19386 14834
rect 19386 14782 19412 14834
rect 19116 14780 19172 14782
rect 19196 14780 19252 14782
rect 19276 14780 19332 14782
rect 19356 14780 19412 14782
rect 19116 13746 19172 13748
rect 19196 13746 19252 13748
rect 19276 13746 19332 13748
rect 19356 13746 19412 13748
rect 19116 13694 19142 13746
rect 19142 13694 19172 13746
rect 19196 13694 19206 13746
rect 19206 13694 19252 13746
rect 19276 13694 19322 13746
rect 19322 13694 19332 13746
rect 19356 13694 19386 13746
rect 19386 13694 19412 13746
rect 19116 13692 19172 13694
rect 19196 13692 19252 13694
rect 19276 13692 19332 13694
rect 19356 13692 19412 13694
rect 19116 12658 19172 12660
rect 19196 12658 19252 12660
rect 19276 12658 19332 12660
rect 19356 12658 19412 12660
rect 19116 12606 19142 12658
rect 19142 12606 19172 12658
rect 19196 12606 19206 12658
rect 19206 12606 19252 12658
rect 19276 12606 19322 12658
rect 19322 12606 19332 12658
rect 19356 12606 19386 12658
rect 19386 12606 19412 12658
rect 19116 12604 19172 12606
rect 19196 12604 19252 12606
rect 19276 12604 19332 12606
rect 19356 12604 19412 12606
rect 19116 11570 19172 11572
rect 19196 11570 19252 11572
rect 19276 11570 19332 11572
rect 19356 11570 19412 11572
rect 19116 11518 19142 11570
rect 19142 11518 19172 11570
rect 19196 11518 19206 11570
rect 19206 11518 19252 11570
rect 19276 11518 19322 11570
rect 19322 11518 19332 11570
rect 19356 11518 19386 11570
rect 19386 11518 19412 11570
rect 19116 11516 19172 11518
rect 19196 11516 19252 11518
rect 19276 11516 19332 11518
rect 19356 11516 19412 11518
rect 24116 26258 24172 26260
rect 24196 26258 24252 26260
rect 24276 26258 24332 26260
rect 24356 26258 24412 26260
rect 24116 26206 24142 26258
rect 24142 26206 24172 26258
rect 24196 26206 24206 26258
rect 24206 26206 24252 26258
rect 24276 26206 24322 26258
rect 24322 26206 24332 26258
rect 24356 26206 24386 26258
rect 24386 26206 24412 26258
rect 24116 26204 24172 26206
rect 24196 26204 24252 26206
rect 24276 26204 24332 26206
rect 24356 26204 24412 26206
rect 24116 25170 24172 25172
rect 24196 25170 24252 25172
rect 24276 25170 24332 25172
rect 24356 25170 24412 25172
rect 24116 25118 24142 25170
rect 24142 25118 24172 25170
rect 24196 25118 24206 25170
rect 24206 25118 24252 25170
rect 24276 25118 24322 25170
rect 24322 25118 24332 25170
rect 24356 25118 24386 25170
rect 24386 25118 24412 25170
rect 24116 25116 24172 25118
rect 24196 25116 24252 25118
rect 24276 25116 24332 25118
rect 24356 25116 24412 25118
rect 24116 24082 24172 24084
rect 24196 24082 24252 24084
rect 24276 24082 24332 24084
rect 24356 24082 24412 24084
rect 24116 24030 24142 24082
rect 24142 24030 24172 24082
rect 24196 24030 24206 24082
rect 24206 24030 24252 24082
rect 24276 24030 24322 24082
rect 24322 24030 24332 24082
rect 24356 24030 24386 24082
rect 24386 24030 24412 24082
rect 24116 24028 24172 24030
rect 24196 24028 24252 24030
rect 24276 24028 24332 24030
rect 24356 24028 24412 24030
rect 24116 22994 24172 22996
rect 24196 22994 24252 22996
rect 24276 22994 24332 22996
rect 24356 22994 24412 22996
rect 24116 22942 24142 22994
rect 24142 22942 24172 22994
rect 24196 22942 24206 22994
rect 24206 22942 24252 22994
rect 24276 22942 24322 22994
rect 24322 22942 24332 22994
rect 24356 22942 24386 22994
rect 24386 22942 24412 22994
rect 24116 22940 24172 22942
rect 24196 22940 24252 22942
rect 24276 22940 24332 22942
rect 24356 22940 24412 22942
rect 24116 21906 24172 21908
rect 24196 21906 24252 21908
rect 24276 21906 24332 21908
rect 24356 21906 24412 21908
rect 24116 21854 24142 21906
rect 24142 21854 24172 21906
rect 24196 21854 24206 21906
rect 24206 21854 24252 21906
rect 24276 21854 24322 21906
rect 24322 21854 24332 21906
rect 24356 21854 24386 21906
rect 24386 21854 24412 21906
rect 24116 21852 24172 21854
rect 24196 21852 24252 21854
rect 24276 21852 24332 21854
rect 24356 21852 24412 21854
rect 24116 20818 24172 20820
rect 24196 20818 24252 20820
rect 24276 20818 24332 20820
rect 24356 20818 24412 20820
rect 24116 20766 24142 20818
rect 24142 20766 24172 20818
rect 24196 20766 24206 20818
rect 24206 20766 24252 20818
rect 24276 20766 24322 20818
rect 24322 20766 24332 20818
rect 24356 20766 24386 20818
rect 24386 20766 24412 20818
rect 24116 20764 24172 20766
rect 24196 20764 24252 20766
rect 24276 20764 24332 20766
rect 24356 20764 24412 20766
rect 24116 19730 24172 19732
rect 24196 19730 24252 19732
rect 24276 19730 24332 19732
rect 24356 19730 24412 19732
rect 24116 19678 24142 19730
rect 24142 19678 24172 19730
rect 24196 19678 24206 19730
rect 24206 19678 24252 19730
rect 24276 19678 24322 19730
rect 24322 19678 24332 19730
rect 24356 19678 24386 19730
rect 24386 19678 24412 19730
rect 24116 19676 24172 19678
rect 24196 19676 24252 19678
rect 24276 19676 24332 19678
rect 24356 19676 24412 19678
rect 24116 18642 24172 18644
rect 24196 18642 24252 18644
rect 24276 18642 24332 18644
rect 24356 18642 24412 18644
rect 24116 18590 24142 18642
rect 24142 18590 24172 18642
rect 24196 18590 24206 18642
rect 24206 18590 24252 18642
rect 24276 18590 24322 18642
rect 24322 18590 24332 18642
rect 24356 18590 24386 18642
rect 24386 18590 24412 18642
rect 24116 18588 24172 18590
rect 24196 18588 24252 18590
rect 24276 18588 24332 18590
rect 24356 18588 24412 18590
rect 24116 17554 24172 17556
rect 24196 17554 24252 17556
rect 24276 17554 24332 17556
rect 24356 17554 24412 17556
rect 24116 17502 24142 17554
rect 24142 17502 24172 17554
rect 24196 17502 24206 17554
rect 24206 17502 24252 17554
rect 24276 17502 24322 17554
rect 24322 17502 24332 17554
rect 24356 17502 24386 17554
rect 24386 17502 24412 17554
rect 24116 17500 24172 17502
rect 24196 17500 24252 17502
rect 24276 17500 24332 17502
rect 24356 17500 24412 17502
rect 24116 16466 24172 16468
rect 24196 16466 24252 16468
rect 24276 16466 24332 16468
rect 24356 16466 24412 16468
rect 24116 16414 24142 16466
rect 24142 16414 24172 16466
rect 24196 16414 24206 16466
rect 24206 16414 24252 16466
rect 24276 16414 24322 16466
rect 24322 16414 24332 16466
rect 24356 16414 24386 16466
rect 24386 16414 24412 16466
rect 24116 16412 24172 16414
rect 24196 16412 24252 16414
rect 24276 16412 24332 16414
rect 24356 16412 24412 16414
rect 24116 15378 24172 15380
rect 24196 15378 24252 15380
rect 24276 15378 24332 15380
rect 24356 15378 24412 15380
rect 24116 15326 24142 15378
rect 24142 15326 24172 15378
rect 24196 15326 24206 15378
rect 24206 15326 24252 15378
rect 24276 15326 24322 15378
rect 24322 15326 24332 15378
rect 24356 15326 24386 15378
rect 24386 15326 24412 15378
rect 24116 15324 24172 15326
rect 24196 15324 24252 15326
rect 24276 15324 24332 15326
rect 24356 15324 24412 15326
rect 24116 14290 24172 14292
rect 24196 14290 24252 14292
rect 24276 14290 24332 14292
rect 24356 14290 24412 14292
rect 24116 14238 24142 14290
rect 24142 14238 24172 14290
rect 24196 14238 24206 14290
rect 24206 14238 24252 14290
rect 24276 14238 24322 14290
rect 24322 14238 24332 14290
rect 24356 14238 24386 14290
rect 24386 14238 24412 14290
rect 24116 14236 24172 14238
rect 24196 14236 24252 14238
rect 24276 14236 24332 14238
rect 24356 14236 24412 14238
rect 24116 13202 24172 13204
rect 24196 13202 24252 13204
rect 24276 13202 24332 13204
rect 24356 13202 24412 13204
rect 24116 13150 24142 13202
rect 24142 13150 24172 13202
rect 24196 13150 24206 13202
rect 24206 13150 24252 13202
rect 24276 13150 24322 13202
rect 24322 13150 24332 13202
rect 24356 13150 24386 13202
rect 24386 13150 24412 13202
rect 24116 13148 24172 13150
rect 24196 13148 24252 13150
rect 24276 13148 24332 13150
rect 24356 13148 24412 13150
rect 24116 12114 24172 12116
rect 24196 12114 24252 12116
rect 24276 12114 24332 12116
rect 24356 12114 24412 12116
rect 24116 12062 24142 12114
rect 24142 12062 24172 12114
rect 24196 12062 24206 12114
rect 24206 12062 24252 12114
rect 24276 12062 24322 12114
rect 24322 12062 24332 12114
rect 24356 12062 24386 12114
rect 24386 12062 24412 12114
rect 24116 12060 24172 12062
rect 24196 12060 24252 12062
rect 24276 12060 24332 12062
rect 24356 12060 24412 12062
rect 24818 25476 24874 25512
rect 24818 25456 24820 25476
rect 24820 25456 24872 25476
rect 24872 25456 24874 25476
rect 29116 30066 29172 30068
rect 29196 30066 29252 30068
rect 29276 30066 29332 30068
rect 29356 30066 29412 30068
rect 29116 30014 29142 30066
rect 29142 30014 29172 30066
rect 29196 30014 29206 30066
rect 29206 30014 29252 30066
rect 29276 30014 29322 30066
rect 29322 30014 29332 30066
rect 29356 30014 29386 30066
rect 29386 30014 29412 30066
rect 29116 30012 29172 30014
rect 29196 30012 29252 30014
rect 29276 30012 29332 30014
rect 29356 30012 29412 30014
rect 28958 29808 29014 29864
rect 27026 25456 27082 25512
rect 29116 28978 29172 28980
rect 29196 28978 29252 28980
rect 29276 28978 29332 28980
rect 29356 28978 29412 28980
rect 29116 28926 29142 28978
rect 29142 28926 29172 28978
rect 29196 28926 29206 28978
rect 29206 28926 29252 28978
rect 29276 28926 29322 28978
rect 29322 28926 29332 28978
rect 29356 28926 29386 28978
rect 29386 28926 29412 28978
rect 29116 28924 29172 28926
rect 29196 28924 29252 28926
rect 29276 28924 29332 28926
rect 29356 28924 29412 28926
rect 29116 27890 29172 27892
rect 29196 27890 29252 27892
rect 29276 27890 29332 27892
rect 29356 27890 29412 27892
rect 29116 27838 29142 27890
rect 29142 27838 29172 27890
rect 29196 27838 29206 27890
rect 29206 27838 29252 27890
rect 29276 27838 29322 27890
rect 29322 27838 29332 27890
rect 29356 27838 29386 27890
rect 29386 27838 29412 27890
rect 29116 27836 29172 27838
rect 29196 27836 29252 27838
rect 29276 27836 29332 27838
rect 29356 27836 29412 27838
rect 28958 27360 29014 27416
rect 29116 26802 29172 26804
rect 29196 26802 29252 26804
rect 29276 26802 29332 26804
rect 29356 26802 29412 26804
rect 29116 26750 29142 26802
rect 29142 26750 29172 26802
rect 29196 26750 29206 26802
rect 29206 26750 29252 26802
rect 29276 26750 29322 26802
rect 29322 26750 29332 26802
rect 29356 26750 29386 26802
rect 29386 26750 29412 26802
rect 29116 26748 29172 26750
rect 29196 26748 29252 26750
rect 29276 26748 29332 26750
rect 29356 26748 29412 26750
rect 29116 25714 29172 25716
rect 29196 25714 29252 25716
rect 29276 25714 29332 25716
rect 29356 25714 29412 25716
rect 29116 25662 29142 25714
rect 29142 25662 29172 25714
rect 29196 25662 29206 25714
rect 29206 25662 29252 25714
rect 29276 25662 29322 25714
rect 29322 25662 29332 25714
rect 29356 25662 29386 25714
rect 29386 25662 29412 25714
rect 29116 25660 29172 25662
rect 29196 25660 29252 25662
rect 29276 25660 29332 25662
rect 29356 25660 29412 25662
rect 29116 24626 29172 24628
rect 29196 24626 29252 24628
rect 29276 24626 29332 24628
rect 29356 24626 29412 24628
rect 29116 24574 29142 24626
rect 29142 24574 29172 24626
rect 29196 24574 29206 24626
rect 29206 24574 29252 24626
rect 29276 24574 29322 24626
rect 29322 24574 29332 24626
rect 29356 24574 29386 24626
rect 29386 24574 29412 24626
rect 29116 24572 29172 24574
rect 29196 24572 29252 24574
rect 29276 24572 29332 24574
rect 29356 24572 29412 24574
rect 29142 24368 29198 24424
rect 29116 23538 29172 23540
rect 29196 23538 29252 23540
rect 29276 23538 29332 23540
rect 29356 23538 29412 23540
rect 29116 23486 29142 23538
rect 29142 23486 29172 23538
rect 29196 23486 29206 23538
rect 29206 23486 29252 23538
rect 29276 23486 29322 23538
rect 29322 23486 29332 23538
rect 29356 23486 29386 23538
rect 29386 23486 29412 23538
rect 29116 23484 29172 23486
rect 29196 23484 29252 23486
rect 29276 23484 29332 23486
rect 29356 23484 29412 23486
rect 29116 22450 29172 22452
rect 29196 22450 29252 22452
rect 29276 22450 29332 22452
rect 29356 22450 29412 22452
rect 29116 22398 29142 22450
rect 29142 22398 29172 22450
rect 29196 22398 29206 22450
rect 29206 22398 29252 22450
rect 29276 22398 29322 22450
rect 29322 22398 29332 22450
rect 29356 22398 29386 22450
rect 29386 22398 29412 22450
rect 29116 22396 29172 22398
rect 29196 22396 29252 22398
rect 29276 22396 29332 22398
rect 29356 22396 29412 22398
rect 29326 21648 29382 21704
rect 29116 21362 29172 21364
rect 29196 21362 29252 21364
rect 29276 21362 29332 21364
rect 29356 21362 29412 21364
rect 29116 21310 29142 21362
rect 29142 21310 29172 21362
rect 29196 21310 29206 21362
rect 29206 21310 29252 21362
rect 29276 21310 29322 21362
rect 29322 21310 29332 21362
rect 29356 21310 29386 21362
rect 29386 21310 29412 21362
rect 29116 21308 29172 21310
rect 29196 21308 29252 21310
rect 29276 21308 29332 21310
rect 29356 21308 29412 21310
rect 29116 20274 29172 20276
rect 29196 20274 29252 20276
rect 29276 20274 29332 20276
rect 29356 20274 29412 20276
rect 29116 20222 29142 20274
rect 29142 20222 29172 20274
rect 29196 20222 29206 20274
rect 29206 20222 29252 20274
rect 29276 20222 29322 20274
rect 29322 20222 29332 20274
rect 29356 20222 29386 20274
rect 29386 20222 29412 20274
rect 29116 20220 29172 20222
rect 29196 20220 29252 20222
rect 29276 20220 29332 20222
rect 29356 20220 29412 20222
rect 29116 19186 29172 19188
rect 29196 19186 29252 19188
rect 29276 19186 29332 19188
rect 29356 19186 29412 19188
rect 29116 19134 29142 19186
rect 29142 19134 29172 19186
rect 29196 19134 29206 19186
rect 29206 19134 29252 19186
rect 29276 19134 29322 19186
rect 29322 19134 29332 19186
rect 29356 19134 29386 19186
rect 29386 19134 29412 19186
rect 29116 19132 29172 19134
rect 29196 19132 29252 19134
rect 29276 19132 29332 19134
rect 29356 19132 29412 19134
rect 29510 18928 29566 18984
rect 29116 18098 29172 18100
rect 29196 18098 29252 18100
rect 29276 18098 29332 18100
rect 29356 18098 29412 18100
rect 29116 18046 29142 18098
rect 29142 18046 29172 18098
rect 29196 18046 29206 18098
rect 29206 18046 29252 18098
rect 29276 18046 29322 18098
rect 29322 18046 29332 18098
rect 29356 18046 29386 18098
rect 29386 18046 29412 18098
rect 29116 18044 29172 18046
rect 29196 18044 29252 18046
rect 29276 18044 29332 18046
rect 29356 18044 29412 18046
rect 27210 13216 27266 13272
rect 24116 11026 24172 11028
rect 24196 11026 24252 11028
rect 24276 11026 24332 11028
rect 24356 11026 24412 11028
rect 24116 10974 24142 11026
rect 24142 10974 24172 11026
rect 24196 10974 24206 11026
rect 24206 10974 24252 11026
rect 24276 10974 24322 11026
rect 24322 10974 24332 11026
rect 24356 10974 24386 11026
rect 24386 10974 24412 11026
rect 24116 10972 24172 10974
rect 24196 10972 24252 10974
rect 24276 10972 24332 10974
rect 24356 10972 24412 10974
rect 29116 17010 29172 17012
rect 29196 17010 29252 17012
rect 29276 17010 29332 17012
rect 29356 17010 29412 17012
rect 29116 16958 29142 17010
rect 29142 16958 29172 17010
rect 29196 16958 29206 17010
rect 29206 16958 29252 17010
rect 29276 16958 29322 17010
rect 29322 16958 29332 17010
rect 29356 16958 29386 17010
rect 29386 16958 29412 17010
rect 29116 16956 29172 16958
rect 29196 16956 29252 16958
rect 29276 16956 29332 16958
rect 29356 16956 29412 16958
rect 28958 16208 29014 16264
rect 29116 15922 29172 15924
rect 29196 15922 29252 15924
rect 29276 15922 29332 15924
rect 29356 15922 29412 15924
rect 29116 15870 29142 15922
rect 29142 15870 29172 15922
rect 29196 15870 29206 15922
rect 29206 15870 29252 15922
rect 29276 15870 29322 15922
rect 29322 15870 29332 15922
rect 29356 15870 29386 15922
rect 29386 15870 29412 15922
rect 29116 15868 29172 15870
rect 29196 15868 29252 15870
rect 29276 15868 29332 15870
rect 29356 15868 29412 15870
rect 29116 14834 29172 14836
rect 29196 14834 29252 14836
rect 29276 14834 29332 14836
rect 29356 14834 29412 14836
rect 29116 14782 29142 14834
rect 29142 14782 29172 14834
rect 29196 14782 29206 14834
rect 29206 14782 29252 14834
rect 29276 14782 29322 14834
rect 29322 14782 29332 14834
rect 29356 14782 29386 14834
rect 29386 14782 29412 14834
rect 29116 14780 29172 14782
rect 29196 14780 29252 14782
rect 29276 14780 29332 14782
rect 29356 14780 29412 14782
rect 29116 13746 29172 13748
rect 29196 13746 29252 13748
rect 29276 13746 29332 13748
rect 29356 13746 29412 13748
rect 29116 13694 29142 13746
rect 29142 13694 29172 13746
rect 29196 13694 29206 13746
rect 29206 13694 29252 13746
rect 29276 13694 29322 13746
rect 29322 13694 29332 13746
rect 29356 13694 29386 13746
rect 29386 13694 29412 13746
rect 29116 13692 29172 13694
rect 29196 13692 29252 13694
rect 29276 13692 29332 13694
rect 29356 13692 29412 13694
rect 29116 12658 29172 12660
rect 29196 12658 29252 12660
rect 29276 12658 29332 12660
rect 29356 12658 29412 12660
rect 29116 12606 29142 12658
rect 29142 12606 29172 12658
rect 29196 12606 29206 12658
rect 29206 12606 29252 12658
rect 29276 12606 29322 12658
rect 29322 12606 29332 12658
rect 29356 12606 29386 12658
rect 29386 12606 29412 12658
rect 29116 12604 29172 12606
rect 29196 12604 29252 12606
rect 29276 12604 29332 12606
rect 29356 12604 29412 12606
rect 29116 11570 29172 11572
rect 29196 11570 29252 11572
rect 29276 11570 29332 11572
rect 29356 11570 29412 11572
rect 29116 11518 29142 11570
rect 29142 11518 29172 11570
rect 29196 11518 29206 11570
rect 29206 11518 29252 11570
rect 29276 11518 29322 11570
rect 29322 11518 29332 11570
rect 29356 11518 29386 11570
rect 29386 11518 29412 11570
rect 29116 11516 29172 11518
rect 29196 11516 29252 11518
rect 29276 11516 29332 11518
rect 29356 11516 29412 11518
rect 27762 10496 27818 10552
<< metal3 >>
rect 0 41032 41136 41040
rect 0 37048 8 41032
rect 3992 37048 19112 41032
rect 19416 37048 29112 41032
rect 29416 37048 37144 41032
rect 41128 37048 41136 41032
rect 0 37040 41136 37048
rect 5000 36032 36136 36040
rect 5000 32048 5008 36032
rect 8992 32048 14112 36032
rect 14416 32048 24112 36032
rect 24416 32048 32144 36032
rect 36128 32048 36136 36032
rect 5000 32040 36136 32048
rect 30504 30138 31304 30168
rect 29646 30078 31304 30138
rect 19104 30072 19424 30073
rect 19104 30008 19112 30072
rect 19176 30008 19192 30072
rect 19256 30008 19272 30072
rect 19336 30008 19352 30072
rect 19416 30008 19424 30072
rect 19104 30007 19424 30008
rect 29104 30072 29424 30073
rect 29104 30008 29112 30072
rect 29176 30008 29192 30072
rect 29256 30008 29272 30072
rect 29336 30008 29352 30072
rect 29416 30008 29424 30072
rect 29104 30007 29424 30008
rect 28953 29866 29019 29869
rect 29646 29866 29706 30078
rect 30504 30048 31304 30078
rect 28953 29864 29706 29866
rect 28953 29808 28958 29864
rect 29014 29808 29706 29864
rect 28953 29806 29706 29808
rect 28953 29803 29019 29806
rect 14104 29528 14424 29529
rect 14104 29464 14112 29528
rect 14176 29464 14192 29528
rect 14256 29464 14272 29528
rect 14336 29464 14352 29528
rect 14416 29464 14424 29528
rect 14104 29463 14424 29464
rect 24104 29528 24424 29529
rect 24104 29464 24112 29528
rect 24176 29464 24192 29528
rect 24256 29464 24272 29528
rect 24336 29464 24352 29528
rect 24416 29464 24424 29528
rect 24104 29463 24424 29464
rect 9896 29322 10696 29352
rect 13497 29322 13563 29325
rect 9896 29320 13563 29322
rect 9896 29264 13502 29320
rect 13558 29264 13563 29320
rect 9896 29262 13563 29264
rect 9896 29232 10696 29262
rect 13497 29259 13563 29262
rect 19104 28984 19424 28985
rect 19104 28920 19112 28984
rect 19176 28920 19192 28984
rect 19256 28920 19272 28984
rect 19336 28920 19352 28984
rect 19416 28920 19424 28984
rect 19104 28919 19424 28920
rect 29104 28984 29424 28985
rect 29104 28920 29112 28984
rect 29176 28920 29192 28984
rect 29256 28920 29272 28984
rect 29336 28920 29352 28984
rect 29416 28920 29424 28984
rect 29104 28919 29424 28920
rect 14104 28440 14424 28441
rect 14104 28376 14112 28440
rect 14176 28376 14192 28440
rect 14256 28376 14272 28440
rect 14336 28376 14352 28440
rect 14416 28376 14424 28440
rect 14104 28375 14424 28376
rect 24104 28440 24424 28441
rect 24104 28376 24112 28440
rect 24176 28376 24192 28440
rect 24256 28376 24272 28440
rect 24336 28376 24352 28440
rect 24416 28376 24424 28440
rect 24104 28375 24424 28376
rect 19104 27896 19424 27897
rect 19104 27832 19112 27896
rect 19176 27832 19192 27896
rect 19256 27832 19272 27896
rect 19336 27832 19352 27896
rect 19416 27832 19424 27896
rect 19104 27831 19424 27832
rect 29104 27896 29424 27897
rect 29104 27832 29112 27896
rect 29176 27832 29192 27896
rect 29256 27832 29272 27896
rect 29336 27832 29352 27896
rect 29416 27832 29424 27896
rect 29104 27831 29424 27832
rect 28953 27418 29019 27421
rect 30504 27418 31304 27448
rect 28953 27416 31304 27418
rect 28953 27360 28958 27416
rect 29014 27360 31304 27416
rect 28953 27358 31304 27360
rect 28953 27355 29019 27358
rect 14104 27352 14424 27353
rect 14104 27288 14112 27352
rect 14176 27288 14192 27352
rect 14256 27288 14272 27352
rect 14336 27288 14352 27352
rect 14416 27288 14424 27352
rect 14104 27287 14424 27288
rect 24104 27352 24424 27353
rect 24104 27288 24112 27352
rect 24176 27288 24192 27352
rect 24256 27288 24272 27352
rect 24336 27288 24352 27352
rect 24416 27288 24424 27352
rect 30504 27328 31304 27358
rect 24104 27287 24424 27288
rect 19104 26808 19424 26809
rect 19104 26744 19112 26808
rect 19176 26744 19192 26808
rect 19256 26744 19272 26808
rect 19336 26744 19352 26808
rect 19416 26744 19424 26808
rect 19104 26743 19424 26744
rect 29104 26808 29424 26809
rect 29104 26744 29112 26808
rect 29176 26744 29192 26808
rect 29256 26744 29272 26808
rect 29336 26744 29352 26808
rect 29416 26744 29424 26808
rect 29104 26743 29424 26744
rect 9896 26330 10696 26360
rect 11657 26330 11723 26333
rect 9896 26328 11723 26330
rect 9896 26272 11662 26328
rect 11718 26272 11723 26328
rect 9896 26270 11723 26272
rect 9896 26240 10696 26270
rect 11657 26267 11723 26270
rect 14104 26264 14424 26265
rect 14104 26200 14112 26264
rect 14176 26200 14192 26264
rect 14256 26200 14272 26264
rect 14336 26200 14352 26264
rect 14416 26200 14424 26264
rect 14104 26199 14424 26200
rect 24104 26264 24424 26265
rect 24104 26200 24112 26264
rect 24176 26200 24192 26264
rect 24256 26200 24272 26264
rect 24336 26200 24352 26264
rect 24416 26200 24424 26264
rect 24104 26199 24424 26200
rect 19104 25720 19424 25721
rect 19104 25656 19112 25720
rect 19176 25656 19192 25720
rect 19256 25656 19272 25720
rect 19336 25656 19352 25720
rect 19416 25656 19424 25720
rect 19104 25655 19424 25656
rect 29104 25720 29424 25721
rect 29104 25656 29112 25720
rect 29176 25656 29192 25720
rect 29256 25656 29272 25720
rect 29336 25656 29352 25720
rect 29416 25656 29424 25720
rect 29104 25655 29424 25656
rect 24813 25514 24879 25517
rect 27021 25514 27087 25517
rect 24813 25512 27087 25514
rect 24813 25456 24818 25512
rect 24874 25456 27026 25512
rect 27082 25456 27087 25512
rect 24813 25454 27087 25456
rect 24813 25451 24879 25454
rect 27021 25451 27087 25454
rect 14104 25176 14424 25177
rect 14104 25112 14112 25176
rect 14176 25112 14192 25176
rect 14256 25112 14272 25176
rect 14336 25112 14352 25176
rect 14416 25112 14424 25176
rect 14104 25111 14424 25112
rect 24104 25176 24424 25177
rect 24104 25112 24112 25176
rect 24176 25112 24192 25176
rect 24256 25112 24272 25176
rect 24336 25112 24352 25176
rect 24416 25112 24424 25176
rect 24104 25111 24424 25112
rect 15797 24834 15863 24837
rect 19017 24834 19083 24837
rect 15797 24832 19083 24834
rect 15797 24776 15802 24832
rect 15858 24776 19022 24832
rect 19078 24776 19083 24832
rect 15797 24774 19083 24776
rect 15797 24771 15863 24774
rect 19017 24771 19083 24774
rect 30504 24698 31304 24728
rect 29646 24638 31304 24698
rect 19104 24632 19424 24633
rect 19104 24568 19112 24632
rect 19176 24568 19192 24632
rect 19256 24568 19272 24632
rect 19336 24568 19352 24632
rect 19416 24568 19424 24632
rect 19104 24567 19424 24568
rect 29104 24632 29424 24633
rect 29104 24568 29112 24632
rect 29176 24568 29192 24632
rect 29256 24568 29272 24632
rect 29336 24568 29352 24632
rect 29416 24568 29424 24632
rect 29104 24567 29424 24568
rect 29137 24426 29203 24429
rect 29646 24426 29706 24638
rect 30504 24608 31304 24638
rect 29137 24424 29706 24426
rect 29137 24368 29142 24424
rect 29198 24368 29706 24424
rect 29137 24366 29706 24368
rect 29137 24363 29203 24366
rect 14104 24088 14424 24089
rect 14104 24024 14112 24088
rect 14176 24024 14192 24088
rect 14256 24024 14272 24088
rect 14336 24024 14352 24088
rect 14416 24024 14424 24088
rect 14104 24023 14424 24024
rect 24104 24088 24424 24089
rect 24104 24024 24112 24088
rect 24176 24024 24192 24088
rect 24256 24024 24272 24088
rect 24336 24024 24352 24088
rect 24416 24024 24424 24088
rect 24104 24023 24424 24024
rect 9896 23610 10696 23640
rect 13865 23610 13931 23613
rect 9896 23608 13931 23610
rect 9896 23552 13870 23608
rect 13926 23552 13931 23608
rect 9896 23550 13931 23552
rect 9896 23520 10696 23550
rect 13865 23547 13931 23550
rect 19104 23544 19424 23545
rect 19104 23480 19112 23544
rect 19176 23480 19192 23544
rect 19256 23480 19272 23544
rect 19336 23480 19352 23544
rect 19416 23480 19424 23544
rect 19104 23479 19424 23480
rect 29104 23544 29424 23545
rect 29104 23480 29112 23544
rect 29176 23480 29192 23544
rect 29256 23480 29272 23544
rect 29336 23480 29352 23544
rect 29416 23480 29424 23544
rect 29104 23479 29424 23480
rect 14104 23000 14424 23001
rect 14104 22936 14112 23000
rect 14176 22936 14192 23000
rect 14256 22936 14272 23000
rect 14336 22936 14352 23000
rect 14416 22936 14424 23000
rect 14104 22935 14424 22936
rect 24104 23000 24424 23001
rect 24104 22936 24112 23000
rect 24176 22936 24192 23000
rect 24256 22936 24272 23000
rect 24336 22936 24352 23000
rect 24416 22936 24424 23000
rect 24104 22935 24424 22936
rect 19104 22456 19424 22457
rect 19104 22392 19112 22456
rect 19176 22392 19192 22456
rect 19256 22392 19272 22456
rect 19336 22392 19352 22456
rect 19416 22392 19424 22456
rect 19104 22391 19424 22392
rect 29104 22456 29424 22457
rect 29104 22392 29112 22456
rect 29176 22392 29192 22456
rect 29256 22392 29272 22456
rect 29336 22392 29352 22456
rect 29416 22392 29424 22456
rect 29104 22391 29424 22392
rect 14104 21912 14424 21913
rect 14104 21848 14112 21912
rect 14176 21848 14192 21912
rect 14256 21848 14272 21912
rect 14336 21848 14352 21912
rect 14416 21848 14424 21912
rect 14104 21847 14424 21848
rect 24104 21912 24424 21913
rect 24104 21848 24112 21912
rect 24176 21848 24192 21912
rect 24256 21848 24272 21912
rect 24336 21848 24352 21912
rect 24416 21848 24424 21912
rect 24104 21847 24424 21848
rect 29321 21706 29387 21709
rect 30504 21706 31304 21736
rect 29321 21704 31304 21706
rect 29321 21648 29326 21704
rect 29382 21648 31304 21704
rect 29321 21646 31304 21648
rect 29321 21643 29387 21646
rect 30504 21616 31304 21646
rect 19104 21368 19424 21369
rect 19104 21304 19112 21368
rect 19176 21304 19192 21368
rect 19256 21304 19272 21368
rect 19336 21304 19352 21368
rect 19416 21304 19424 21368
rect 19104 21303 19424 21304
rect 29104 21368 29424 21369
rect 29104 21304 29112 21368
rect 29176 21304 29192 21368
rect 29256 21304 29272 21368
rect 29336 21304 29352 21368
rect 29416 21304 29424 21368
rect 29104 21303 29424 21304
rect 9896 20890 10696 20920
rect 11657 20890 11723 20893
rect 9896 20888 11723 20890
rect 9896 20832 11662 20888
rect 11718 20832 11723 20888
rect 9896 20830 11723 20832
rect 9896 20800 10696 20830
rect 11657 20827 11723 20830
rect 14104 20824 14424 20825
rect 14104 20760 14112 20824
rect 14176 20760 14192 20824
rect 14256 20760 14272 20824
rect 14336 20760 14352 20824
rect 14416 20760 14424 20824
rect 14104 20759 14424 20760
rect 24104 20824 24424 20825
rect 24104 20760 24112 20824
rect 24176 20760 24192 20824
rect 24256 20760 24272 20824
rect 24336 20760 24352 20824
rect 24416 20760 24424 20824
rect 24104 20759 24424 20760
rect 19104 20280 19424 20281
rect 19104 20216 19112 20280
rect 19176 20216 19192 20280
rect 19256 20216 19272 20280
rect 19336 20216 19352 20280
rect 19416 20216 19424 20280
rect 19104 20215 19424 20216
rect 29104 20280 29424 20281
rect 29104 20216 29112 20280
rect 29176 20216 29192 20280
rect 29256 20216 29272 20280
rect 29336 20216 29352 20280
rect 29416 20216 29424 20280
rect 29104 20215 29424 20216
rect 18189 20074 18255 20077
rect 19937 20074 20003 20077
rect 18189 20072 20003 20074
rect 18189 20016 18194 20072
rect 18250 20016 19942 20072
rect 19998 20016 20003 20072
rect 18189 20014 20003 20016
rect 18189 20011 18255 20014
rect 19937 20011 20003 20014
rect 14104 19736 14424 19737
rect 14104 19672 14112 19736
rect 14176 19672 14192 19736
rect 14256 19672 14272 19736
rect 14336 19672 14352 19736
rect 14416 19672 14424 19736
rect 14104 19671 14424 19672
rect 24104 19736 24424 19737
rect 24104 19672 24112 19736
rect 24176 19672 24192 19736
rect 24256 19672 24272 19736
rect 24336 19672 24352 19736
rect 24416 19672 24424 19736
rect 24104 19671 24424 19672
rect 19104 19192 19424 19193
rect 19104 19128 19112 19192
rect 19176 19128 19192 19192
rect 19256 19128 19272 19192
rect 19336 19128 19352 19192
rect 19416 19128 19424 19192
rect 19104 19127 19424 19128
rect 29104 19192 29424 19193
rect 29104 19128 29112 19192
rect 29176 19128 29192 19192
rect 29256 19128 29272 19192
rect 29336 19128 29352 19192
rect 29416 19128 29424 19192
rect 29104 19127 29424 19128
rect 29505 18986 29571 18989
rect 30504 18986 31304 19016
rect 29505 18984 31304 18986
rect 29505 18928 29510 18984
rect 29566 18928 31304 18984
rect 29505 18926 31304 18928
rect 29505 18923 29571 18926
rect 30504 18896 31304 18926
rect 14104 18648 14424 18649
rect 14104 18584 14112 18648
rect 14176 18584 14192 18648
rect 14256 18584 14272 18648
rect 14336 18584 14352 18648
rect 14416 18584 14424 18648
rect 14104 18583 14424 18584
rect 24104 18648 24424 18649
rect 24104 18584 24112 18648
rect 24176 18584 24192 18648
rect 24256 18584 24272 18648
rect 24336 18584 24352 18648
rect 24416 18584 24424 18648
rect 24104 18583 24424 18584
rect 19104 18104 19424 18105
rect 19104 18040 19112 18104
rect 19176 18040 19192 18104
rect 19256 18040 19272 18104
rect 19336 18040 19352 18104
rect 19416 18040 19424 18104
rect 19104 18039 19424 18040
rect 29104 18104 29424 18105
rect 29104 18040 29112 18104
rect 29176 18040 29192 18104
rect 29256 18040 29272 18104
rect 29336 18040 29352 18104
rect 29416 18040 29424 18104
rect 29104 18039 29424 18040
rect 9896 17898 10696 17928
rect 12669 17898 12735 17901
rect 9896 17896 12735 17898
rect 9896 17840 12674 17896
rect 12730 17840 12735 17896
rect 9896 17838 12735 17840
rect 9896 17808 10696 17838
rect 12669 17835 12735 17838
rect 14104 17560 14424 17561
rect 14104 17496 14112 17560
rect 14176 17496 14192 17560
rect 14256 17496 14272 17560
rect 14336 17496 14352 17560
rect 14416 17496 14424 17560
rect 14104 17495 14424 17496
rect 24104 17560 24424 17561
rect 24104 17496 24112 17560
rect 24176 17496 24192 17560
rect 24256 17496 24272 17560
rect 24336 17496 24352 17560
rect 24416 17496 24424 17560
rect 24104 17495 24424 17496
rect 19104 17016 19424 17017
rect 19104 16952 19112 17016
rect 19176 16952 19192 17016
rect 19256 16952 19272 17016
rect 19336 16952 19352 17016
rect 19416 16952 19424 17016
rect 19104 16951 19424 16952
rect 29104 17016 29424 17017
rect 29104 16952 29112 17016
rect 29176 16952 29192 17016
rect 29256 16952 29272 17016
rect 29336 16952 29352 17016
rect 29416 16952 29424 17016
rect 29104 16951 29424 16952
rect 14104 16472 14424 16473
rect 14104 16408 14112 16472
rect 14176 16408 14192 16472
rect 14256 16408 14272 16472
rect 14336 16408 14352 16472
rect 14416 16408 14424 16472
rect 14104 16407 14424 16408
rect 24104 16472 24424 16473
rect 24104 16408 24112 16472
rect 24176 16408 24192 16472
rect 24256 16408 24272 16472
rect 24336 16408 24352 16472
rect 24416 16408 24424 16472
rect 24104 16407 24424 16408
rect 28953 16266 29019 16269
rect 30504 16266 31304 16296
rect 28953 16264 31304 16266
rect 28953 16208 28958 16264
rect 29014 16208 31304 16264
rect 28953 16206 31304 16208
rect 28953 16203 29019 16206
rect 30504 16176 31304 16206
rect 19104 15928 19424 15929
rect 19104 15864 19112 15928
rect 19176 15864 19192 15928
rect 19256 15864 19272 15928
rect 19336 15864 19352 15928
rect 19416 15864 19424 15928
rect 19104 15863 19424 15864
rect 29104 15928 29424 15929
rect 29104 15864 29112 15928
rect 29176 15864 29192 15928
rect 29256 15864 29272 15928
rect 29336 15864 29352 15928
rect 29416 15864 29424 15928
rect 29104 15863 29424 15864
rect 14104 15384 14424 15385
rect 14104 15320 14112 15384
rect 14176 15320 14192 15384
rect 14256 15320 14272 15384
rect 14336 15320 14352 15384
rect 14416 15320 14424 15384
rect 14104 15319 14424 15320
rect 24104 15384 24424 15385
rect 24104 15320 24112 15384
rect 24176 15320 24192 15384
rect 24256 15320 24272 15384
rect 24336 15320 24352 15384
rect 24416 15320 24424 15384
rect 24104 15319 24424 15320
rect 9896 15178 10696 15208
rect 13957 15178 14023 15181
rect 9896 15176 14023 15178
rect 9896 15120 13962 15176
rect 14018 15120 14023 15176
rect 9896 15118 14023 15120
rect 9896 15088 10696 15118
rect 13957 15115 14023 15118
rect 19104 14840 19424 14841
rect 19104 14776 19112 14840
rect 19176 14776 19192 14840
rect 19256 14776 19272 14840
rect 19336 14776 19352 14840
rect 19416 14776 19424 14840
rect 19104 14775 19424 14776
rect 29104 14840 29424 14841
rect 29104 14776 29112 14840
rect 29176 14776 29192 14840
rect 29256 14776 29272 14840
rect 29336 14776 29352 14840
rect 29416 14776 29424 14840
rect 29104 14775 29424 14776
rect 14104 14296 14424 14297
rect 14104 14232 14112 14296
rect 14176 14232 14192 14296
rect 14256 14232 14272 14296
rect 14336 14232 14352 14296
rect 14416 14232 14424 14296
rect 14104 14231 14424 14232
rect 24104 14296 24424 14297
rect 24104 14232 24112 14296
rect 24176 14232 24192 14296
rect 24256 14232 24272 14296
rect 24336 14232 24352 14296
rect 24416 14232 24424 14296
rect 24104 14231 24424 14232
rect 19104 13752 19424 13753
rect 19104 13688 19112 13752
rect 19176 13688 19192 13752
rect 19256 13688 19272 13752
rect 19336 13688 19352 13752
rect 19416 13688 19424 13752
rect 19104 13687 19424 13688
rect 29104 13752 29424 13753
rect 29104 13688 29112 13752
rect 29176 13688 29192 13752
rect 29256 13688 29272 13752
rect 29336 13688 29352 13752
rect 29416 13688 29424 13752
rect 29104 13687 29424 13688
rect 27205 13274 27271 13277
rect 30504 13274 31304 13304
rect 27205 13272 31304 13274
rect 27205 13216 27210 13272
rect 27266 13216 31304 13272
rect 27205 13214 31304 13216
rect 27205 13211 27271 13214
rect 14104 13208 14424 13209
rect 14104 13144 14112 13208
rect 14176 13144 14192 13208
rect 14256 13144 14272 13208
rect 14336 13144 14352 13208
rect 14416 13144 14424 13208
rect 14104 13143 14424 13144
rect 24104 13208 24424 13209
rect 24104 13144 24112 13208
rect 24176 13144 24192 13208
rect 24256 13144 24272 13208
rect 24336 13144 24352 13208
rect 24416 13144 24424 13208
rect 30504 13184 31304 13214
rect 24104 13143 24424 13144
rect 19104 12664 19424 12665
rect 19104 12600 19112 12664
rect 19176 12600 19192 12664
rect 19256 12600 19272 12664
rect 19336 12600 19352 12664
rect 19416 12600 19424 12664
rect 19104 12599 19424 12600
rect 29104 12664 29424 12665
rect 29104 12600 29112 12664
rect 29176 12600 29192 12664
rect 29256 12600 29272 12664
rect 29336 12600 29352 12664
rect 29416 12600 29424 12664
rect 29104 12599 29424 12600
rect 9896 12458 10696 12488
rect 12025 12458 12091 12461
rect 9896 12456 12091 12458
rect 9896 12400 12030 12456
rect 12086 12400 12091 12456
rect 9896 12398 12091 12400
rect 9896 12368 10696 12398
rect 12025 12395 12091 12398
rect 14104 12120 14424 12121
rect 14104 12056 14112 12120
rect 14176 12056 14192 12120
rect 14256 12056 14272 12120
rect 14336 12056 14352 12120
rect 14416 12056 14424 12120
rect 14104 12055 14424 12056
rect 24104 12120 24424 12121
rect 24104 12056 24112 12120
rect 24176 12056 24192 12120
rect 24256 12056 24272 12120
rect 24336 12056 24352 12120
rect 24416 12056 24424 12120
rect 24104 12055 24424 12056
rect 19104 11576 19424 11577
rect 19104 11512 19112 11576
rect 19176 11512 19192 11576
rect 19256 11512 19272 11576
rect 19336 11512 19352 11576
rect 19416 11512 19424 11576
rect 19104 11511 19424 11512
rect 29104 11576 29424 11577
rect 29104 11512 29112 11576
rect 29176 11512 29192 11576
rect 29256 11512 29272 11576
rect 29336 11512 29352 11576
rect 29416 11512 29424 11576
rect 29104 11511 29424 11512
rect 14104 11032 14424 11033
rect 14104 10968 14112 11032
rect 14176 10968 14192 11032
rect 14256 10968 14272 11032
rect 14336 10968 14352 11032
rect 14416 10968 14424 11032
rect 14104 10967 14424 10968
rect 24104 11032 24424 11033
rect 24104 10968 24112 11032
rect 24176 10968 24192 11032
rect 24256 10968 24272 11032
rect 24336 10968 24352 11032
rect 24416 10968 24424 11032
rect 24104 10967 24424 10968
rect 27757 10554 27823 10557
rect 30504 10554 31304 10584
rect 27757 10552 31304 10554
rect 27757 10496 27762 10552
rect 27818 10496 31304 10552
rect 27757 10494 31304 10496
rect 27757 10491 27823 10494
rect 30504 10464 31304 10494
rect 5000 8992 36136 9000
rect 5000 5008 5008 8992
rect 8992 5008 14112 8992
rect 14416 5008 24112 8992
rect 24416 5008 32144 8992
rect 36128 5008 36136 8992
rect 5000 5000 36136 5008
rect 0 3992 41136 4000
rect 0 8 8 3992
rect 3992 8 19112 3992
rect 19416 8 29112 3992
rect 29416 8 37144 3992
rect 41128 8 41136 3992
rect 0 0 41136 8
<< via3 >>
rect 8 37048 3992 41032
rect 19112 37048 19416 41032
rect 29112 37048 29416 41032
rect 37144 37048 41128 41032
rect 5008 32048 8992 36032
rect 14112 32048 14416 36032
rect 24112 32048 24416 36032
rect 32144 32048 36128 36032
rect 19112 30068 19176 30072
rect 19112 30012 19116 30068
rect 19116 30012 19172 30068
rect 19172 30012 19176 30068
rect 19112 30008 19176 30012
rect 19192 30068 19256 30072
rect 19192 30012 19196 30068
rect 19196 30012 19252 30068
rect 19252 30012 19256 30068
rect 19192 30008 19256 30012
rect 19272 30068 19336 30072
rect 19272 30012 19276 30068
rect 19276 30012 19332 30068
rect 19332 30012 19336 30068
rect 19272 30008 19336 30012
rect 19352 30068 19416 30072
rect 19352 30012 19356 30068
rect 19356 30012 19412 30068
rect 19412 30012 19416 30068
rect 19352 30008 19416 30012
rect 29112 30068 29176 30072
rect 29112 30012 29116 30068
rect 29116 30012 29172 30068
rect 29172 30012 29176 30068
rect 29112 30008 29176 30012
rect 29192 30068 29256 30072
rect 29192 30012 29196 30068
rect 29196 30012 29252 30068
rect 29252 30012 29256 30068
rect 29192 30008 29256 30012
rect 29272 30068 29336 30072
rect 29272 30012 29276 30068
rect 29276 30012 29332 30068
rect 29332 30012 29336 30068
rect 29272 30008 29336 30012
rect 29352 30068 29416 30072
rect 29352 30012 29356 30068
rect 29356 30012 29412 30068
rect 29412 30012 29416 30068
rect 29352 30008 29416 30012
rect 14112 29524 14176 29528
rect 14112 29468 14116 29524
rect 14116 29468 14172 29524
rect 14172 29468 14176 29524
rect 14112 29464 14176 29468
rect 14192 29524 14256 29528
rect 14192 29468 14196 29524
rect 14196 29468 14252 29524
rect 14252 29468 14256 29524
rect 14192 29464 14256 29468
rect 14272 29524 14336 29528
rect 14272 29468 14276 29524
rect 14276 29468 14332 29524
rect 14332 29468 14336 29524
rect 14272 29464 14336 29468
rect 14352 29524 14416 29528
rect 14352 29468 14356 29524
rect 14356 29468 14412 29524
rect 14412 29468 14416 29524
rect 14352 29464 14416 29468
rect 24112 29524 24176 29528
rect 24112 29468 24116 29524
rect 24116 29468 24172 29524
rect 24172 29468 24176 29524
rect 24112 29464 24176 29468
rect 24192 29524 24256 29528
rect 24192 29468 24196 29524
rect 24196 29468 24252 29524
rect 24252 29468 24256 29524
rect 24192 29464 24256 29468
rect 24272 29524 24336 29528
rect 24272 29468 24276 29524
rect 24276 29468 24332 29524
rect 24332 29468 24336 29524
rect 24272 29464 24336 29468
rect 24352 29524 24416 29528
rect 24352 29468 24356 29524
rect 24356 29468 24412 29524
rect 24412 29468 24416 29524
rect 24352 29464 24416 29468
rect 19112 28980 19176 28984
rect 19112 28924 19116 28980
rect 19116 28924 19172 28980
rect 19172 28924 19176 28980
rect 19112 28920 19176 28924
rect 19192 28980 19256 28984
rect 19192 28924 19196 28980
rect 19196 28924 19252 28980
rect 19252 28924 19256 28980
rect 19192 28920 19256 28924
rect 19272 28980 19336 28984
rect 19272 28924 19276 28980
rect 19276 28924 19332 28980
rect 19332 28924 19336 28980
rect 19272 28920 19336 28924
rect 19352 28980 19416 28984
rect 19352 28924 19356 28980
rect 19356 28924 19412 28980
rect 19412 28924 19416 28980
rect 19352 28920 19416 28924
rect 29112 28980 29176 28984
rect 29112 28924 29116 28980
rect 29116 28924 29172 28980
rect 29172 28924 29176 28980
rect 29112 28920 29176 28924
rect 29192 28980 29256 28984
rect 29192 28924 29196 28980
rect 29196 28924 29252 28980
rect 29252 28924 29256 28980
rect 29192 28920 29256 28924
rect 29272 28980 29336 28984
rect 29272 28924 29276 28980
rect 29276 28924 29332 28980
rect 29332 28924 29336 28980
rect 29272 28920 29336 28924
rect 29352 28980 29416 28984
rect 29352 28924 29356 28980
rect 29356 28924 29412 28980
rect 29412 28924 29416 28980
rect 29352 28920 29416 28924
rect 14112 28436 14176 28440
rect 14112 28380 14116 28436
rect 14116 28380 14172 28436
rect 14172 28380 14176 28436
rect 14112 28376 14176 28380
rect 14192 28436 14256 28440
rect 14192 28380 14196 28436
rect 14196 28380 14252 28436
rect 14252 28380 14256 28436
rect 14192 28376 14256 28380
rect 14272 28436 14336 28440
rect 14272 28380 14276 28436
rect 14276 28380 14332 28436
rect 14332 28380 14336 28436
rect 14272 28376 14336 28380
rect 14352 28436 14416 28440
rect 14352 28380 14356 28436
rect 14356 28380 14412 28436
rect 14412 28380 14416 28436
rect 14352 28376 14416 28380
rect 24112 28436 24176 28440
rect 24112 28380 24116 28436
rect 24116 28380 24172 28436
rect 24172 28380 24176 28436
rect 24112 28376 24176 28380
rect 24192 28436 24256 28440
rect 24192 28380 24196 28436
rect 24196 28380 24252 28436
rect 24252 28380 24256 28436
rect 24192 28376 24256 28380
rect 24272 28436 24336 28440
rect 24272 28380 24276 28436
rect 24276 28380 24332 28436
rect 24332 28380 24336 28436
rect 24272 28376 24336 28380
rect 24352 28436 24416 28440
rect 24352 28380 24356 28436
rect 24356 28380 24412 28436
rect 24412 28380 24416 28436
rect 24352 28376 24416 28380
rect 19112 27892 19176 27896
rect 19112 27836 19116 27892
rect 19116 27836 19172 27892
rect 19172 27836 19176 27892
rect 19112 27832 19176 27836
rect 19192 27892 19256 27896
rect 19192 27836 19196 27892
rect 19196 27836 19252 27892
rect 19252 27836 19256 27892
rect 19192 27832 19256 27836
rect 19272 27892 19336 27896
rect 19272 27836 19276 27892
rect 19276 27836 19332 27892
rect 19332 27836 19336 27892
rect 19272 27832 19336 27836
rect 19352 27892 19416 27896
rect 19352 27836 19356 27892
rect 19356 27836 19412 27892
rect 19412 27836 19416 27892
rect 19352 27832 19416 27836
rect 29112 27892 29176 27896
rect 29112 27836 29116 27892
rect 29116 27836 29172 27892
rect 29172 27836 29176 27892
rect 29112 27832 29176 27836
rect 29192 27892 29256 27896
rect 29192 27836 29196 27892
rect 29196 27836 29252 27892
rect 29252 27836 29256 27892
rect 29192 27832 29256 27836
rect 29272 27892 29336 27896
rect 29272 27836 29276 27892
rect 29276 27836 29332 27892
rect 29332 27836 29336 27892
rect 29272 27832 29336 27836
rect 29352 27892 29416 27896
rect 29352 27836 29356 27892
rect 29356 27836 29412 27892
rect 29412 27836 29416 27892
rect 29352 27832 29416 27836
rect 14112 27348 14176 27352
rect 14112 27292 14116 27348
rect 14116 27292 14172 27348
rect 14172 27292 14176 27348
rect 14112 27288 14176 27292
rect 14192 27348 14256 27352
rect 14192 27292 14196 27348
rect 14196 27292 14252 27348
rect 14252 27292 14256 27348
rect 14192 27288 14256 27292
rect 14272 27348 14336 27352
rect 14272 27292 14276 27348
rect 14276 27292 14332 27348
rect 14332 27292 14336 27348
rect 14272 27288 14336 27292
rect 14352 27348 14416 27352
rect 14352 27292 14356 27348
rect 14356 27292 14412 27348
rect 14412 27292 14416 27348
rect 14352 27288 14416 27292
rect 24112 27348 24176 27352
rect 24112 27292 24116 27348
rect 24116 27292 24172 27348
rect 24172 27292 24176 27348
rect 24112 27288 24176 27292
rect 24192 27348 24256 27352
rect 24192 27292 24196 27348
rect 24196 27292 24252 27348
rect 24252 27292 24256 27348
rect 24192 27288 24256 27292
rect 24272 27348 24336 27352
rect 24272 27292 24276 27348
rect 24276 27292 24332 27348
rect 24332 27292 24336 27348
rect 24272 27288 24336 27292
rect 24352 27348 24416 27352
rect 24352 27292 24356 27348
rect 24356 27292 24412 27348
rect 24412 27292 24416 27348
rect 24352 27288 24416 27292
rect 19112 26804 19176 26808
rect 19112 26748 19116 26804
rect 19116 26748 19172 26804
rect 19172 26748 19176 26804
rect 19112 26744 19176 26748
rect 19192 26804 19256 26808
rect 19192 26748 19196 26804
rect 19196 26748 19252 26804
rect 19252 26748 19256 26804
rect 19192 26744 19256 26748
rect 19272 26804 19336 26808
rect 19272 26748 19276 26804
rect 19276 26748 19332 26804
rect 19332 26748 19336 26804
rect 19272 26744 19336 26748
rect 19352 26804 19416 26808
rect 19352 26748 19356 26804
rect 19356 26748 19412 26804
rect 19412 26748 19416 26804
rect 19352 26744 19416 26748
rect 29112 26804 29176 26808
rect 29112 26748 29116 26804
rect 29116 26748 29172 26804
rect 29172 26748 29176 26804
rect 29112 26744 29176 26748
rect 29192 26804 29256 26808
rect 29192 26748 29196 26804
rect 29196 26748 29252 26804
rect 29252 26748 29256 26804
rect 29192 26744 29256 26748
rect 29272 26804 29336 26808
rect 29272 26748 29276 26804
rect 29276 26748 29332 26804
rect 29332 26748 29336 26804
rect 29272 26744 29336 26748
rect 29352 26804 29416 26808
rect 29352 26748 29356 26804
rect 29356 26748 29412 26804
rect 29412 26748 29416 26804
rect 29352 26744 29416 26748
rect 14112 26260 14176 26264
rect 14112 26204 14116 26260
rect 14116 26204 14172 26260
rect 14172 26204 14176 26260
rect 14112 26200 14176 26204
rect 14192 26260 14256 26264
rect 14192 26204 14196 26260
rect 14196 26204 14252 26260
rect 14252 26204 14256 26260
rect 14192 26200 14256 26204
rect 14272 26260 14336 26264
rect 14272 26204 14276 26260
rect 14276 26204 14332 26260
rect 14332 26204 14336 26260
rect 14272 26200 14336 26204
rect 14352 26260 14416 26264
rect 14352 26204 14356 26260
rect 14356 26204 14412 26260
rect 14412 26204 14416 26260
rect 14352 26200 14416 26204
rect 24112 26260 24176 26264
rect 24112 26204 24116 26260
rect 24116 26204 24172 26260
rect 24172 26204 24176 26260
rect 24112 26200 24176 26204
rect 24192 26260 24256 26264
rect 24192 26204 24196 26260
rect 24196 26204 24252 26260
rect 24252 26204 24256 26260
rect 24192 26200 24256 26204
rect 24272 26260 24336 26264
rect 24272 26204 24276 26260
rect 24276 26204 24332 26260
rect 24332 26204 24336 26260
rect 24272 26200 24336 26204
rect 24352 26260 24416 26264
rect 24352 26204 24356 26260
rect 24356 26204 24412 26260
rect 24412 26204 24416 26260
rect 24352 26200 24416 26204
rect 19112 25716 19176 25720
rect 19112 25660 19116 25716
rect 19116 25660 19172 25716
rect 19172 25660 19176 25716
rect 19112 25656 19176 25660
rect 19192 25716 19256 25720
rect 19192 25660 19196 25716
rect 19196 25660 19252 25716
rect 19252 25660 19256 25716
rect 19192 25656 19256 25660
rect 19272 25716 19336 25720
rect 19272 25660 19276 25716
rect 19276 25660 19332 25716
rect 19332 25660 19336 25716
rect 19272 25656 19336 25660
rect 19352 25716 19416 25720
rect 19352 25660 19356 25716
rect 19356 25660 19412 25716
rect 19412 25660 19416 25716
rect 19352 25656 19416 25660
rect 29112 25716 29176 25720
rect 29112 25660 29116 25716
rect 29116 25660 29172 25716
rect 29172 25660 29176 25716
rect 29112 25656 29176 25660
rect 29192 25716 29256 25720
rect 29192 25660 29196 25716
rect 29196 25660 29252 25716
rect 29252 25660 29256 25716
rect 29192 25656 29256 25660
rect 29272 25716 29336 25720
rect 29272 25660 29276 25716
rect 29276 25660 29332 25716
rect 29332 25660 29336 25716
rect 29272 25656 29336 25660
rect 29352 25716 29416 25720
rect 29352 25660 29356 25716
rect 29356 25660 29412 25716
rect 29412 25660 29416 25716
rect 29352 25656 29416 25660
rect 14112 25172 14176 25176
rect 14112 25116 14116 25172
rect 14116 25116 14172 25172
rect 14172 25116 14176 25172
rect 14112 25112 14176 25116
rect 14192 25172 14256 25176
rect 14192 25116 14196 25172
rect 14196 25116 14252 25172
rect 14252 25116 14256 25172
rect 14192 25112 14256 25116
rect 14272 25172 14336 25176
rect 14272 25116 14276 25172
rect 14276 25116 14332 25172
rect 14332 25116 14336 25172
rect 14272 25112 14336 25116
rect 14352 25172 14416 25176
rect 14352 25116 14356 25172
rect 14356 25116 14412 25172
rect 14412 25116 14416 25172
rect 14352 25112 14416 25116
rect 24112 25172 24176 25176
rect 24112 25116 24116 25172
rect 24116 25116 24172 25172
rect 24172 25116 24176 25172
rect 24112 25112 24176 25116
rect 24192 25172 24256 25176
rect 24192 25116 24196 25172
rect 24196 25116 24252 25172
rect 24252 25116 24256 25172
rect 24192 25112 24256 25116
rect 24272 25172 24336 25176
rect 24272 25116 24276 25172
rect 24276 25116 24332 25172
rect 24332 25116 24336 25172
rect 24272 25112 24336 25116
rect 24352 25172 24416 25176
rect 24352 25116 24356 25172
rect 24356 25116 24412 25172
rect 24412 25116 24416 25172
rect 24352 25112 24416 25116
rect 19112 24628 19176 24632
rect 19112 24572 19116 24628
rect 19116 24572 19172 24628
rect 19172 24572 19176 24628
rect 19112 24568 19176 24572
rect 19192 24628 19256 24632
rect 19192 24572 19196 24628
rect 19196 24572 19252 24628
rect 19252 24572 19256 24628
rect 19192 24568 19256 24572
rect 19272 24628 19336 24632
rect 19272 24572 19276 24628
rect 19276 24572 19332 24628
rect 19332 24572 19336 24628
rect 19272 24568 19336 24572
rect 19352 24628 19416 24632
rect 19352 24572 19356 24628
rect 19356 24572 19412 24628
rect 19412 24572 19416 24628
rect 19352 24568 19416 24572
rect 29112 24628 29176 24632
rect 29112 24572 29116 24628
rect 29116 24572 29172 24628
rect 29172 24572 29176 24628
rect 29112 24568 29176 24572
rect 29192 24628 29256 24632
rect 29192 24572 29196 24628
rect 29196 24572 29252 24628
rect 29252 24572 29256 24628
rect 29192 24568 29256 24572
rect 29272 24628 29336 24632
rect 29272 24572 29276 24628
rect 29276 24572 29332 24628
rect 29332 24572 29336 24628
rect 29272 24568 29336 24572
rect 29352 24628 29416 24632
rect 29352 24572 29356 24628
rect 29356 24572 29412 24628
rect 29412 24572 29416 24628
rect 29352 24568 29416 24572
rect 14112 24084 14176 24088
rect 14112 24028 14116 24084
rect 14116 24028 14172 24084
rect 14172 24028 14176 24084
rect 14112 24024 14176 24028
rect 14192 24084 14256 24088
rect 14192 24028 14196 24084
rect 14196 24028 14252 24084
rect 14252 24028 14256 24084
rect 14192 24024 14256 24028
rect 14272 24084 14336 24088
rect 14272 24028 14276 24084
rect 14276 24028 14332 24084
rect 14332 24028 14336 24084
rect 14272 24024 14336 24028
rect 14352 24084 14416 24088
rect 14352 24028 14356 24084
rect 14356 24028 14412 24084
rect 14412 24028 14416 24084
rect 14352 24024 14416 24028
rect 24112 24084 24176 24088
rect 24112 24028 24116 24084
rect 24116 24028 24172 24084
rect 24172 24028 24176 24084
rect 24112 24024 24176 24028
rect 24192 24084 24256 24088
rect 24192 24028 24196 24084
rect 24196 24028 24252 24084
rect 24252 24028 24256 24084
rect 24192 24024 24256 24028
rect 24272 24084 24336 24088
rect 24272 24028 24276 24084
rect 24276 24028 24332 24084
rect 24332 24028 24336 24084
rect 24272 24024 24336 24028
rect 24352 24084 24416 24088
rect 24352 24028 24356 24084
rect 24356 24028 24412 24084
rect 24412 24028 24416 24084
rect 24352 24024 24416 24028
rect 19112 23540 19176 23544
rect 19112 23484 19116 23540
rect 19116 23484 19172 23540
rect 19172 23484 19176 23540
rect 19112 23480 19176 23484
rect 19192 23540 19256 23544
rect 19192 23484 19196 23540
rect 19196 23484 19252 23540
rect 19252 23484 19256 23540
rect 19192 23480 19256 23484
rect 19272 23540 19336 23544
rect 19272 23484 19276 23540
rect 19276 23484 19332 23540
rect 19332 23484 19336 23540
rect 19272 23480 19336 23484
rect 19352 23540 19416 23544
rect 19352 23484 19356 23540
rect 19356 23484 19412 23540
rect 19412 23484 19416 23540
rect 19352 23480 19416 23484
rect 29112 23540 29176 23544
rect 29112 23484 29116 23540
rect 29116 23484 29172 23540
rect 29172 23484 29176 23540
rect 29112 23480 29176 23484
rect 29192 23540 29256 23544
rect 29192 23484 29196 23540
rect 29196 23484 29252 23540
rect 29252 23484 29256 23540
rect 29192 23480 29256 23484
rect 29272 23540 29336 23544
rect 29272 23484 29276 23540
rect 29276 23484 29332 23540
rect 29332 23484 29336 23540
rect 29272 23480 29336 23484
rect 29352 23540 29416 23544
rect 29352 23484 29356 23540
rect 29356 23484 29412 23540
rect 29412 23484 29416 23540
rect 29352 23480 29416 23484
rect 14112 22996 14176 23000
rect 14112 22940 14116 22996
rect 14116 22940 14172 22996
rect 14172 22940 14176 22996
rect 14112 22936 14176 22940
rect 14192 22996 14256 23000
rect 14192 22940 14196 22996
rect 14196 22940 14252 22996
rect 14252 22940 14256 22996
rect 14192 22936 14256 22940
rect 14272 22996 14336 23000
rect 14272 22940 14276 22996
rect 14276 22940 14332 22996
rect 14332 22940 14336 22996
rect 14272 22936 14336 22940
rect 14352 22996 14416 23000
rect 14352 22940 14356 22996
rect 14356 22940 14412 22996
rect 14412 22940 14416 22996
rect 14352 22936 14416 22940
rect 24112 22996 24176 23000
rect 24112 22940 24116 22996
rect 24116 22940 24172 22996
rect 24172 22940 24176 22996
rect 24112 22936 24176 22940
rect 24192 22996 24256 23000
rect 24192 22940 24196 22996
rect 24196 22940 24252 22996
rect 24252 22940 24256 22996
rect 24192 22936 24256 22940
rect 24272 22996 24336 23000
rect 24272 22940 24276 22996
rect 24276 22940 24332 22996
rect 24332 22940 24336 22996
rect 24272 22936 24336 22940
rect 24352 22996 24416 23000
rect 24352 22940 24356 22996
rect 24356 22940 24412 22996
rect 24412 22940 24416 22996
rect 24352 22936 24416 22940
rect 19112 22452 19176 22456
rect 19112 22396 19116 22452
rect 19116 22396 19172 22452
rect 19172 22396 19176 22452
rect 19112 22392 19176 22396
rect 19192 22452 19256 22456
rect 19192 22396 19196 22452
rect 19196 22396 19252 22452
rect 19252 22396 19256 22452
rect 19192 22392 19256 22396
rect 19272 22452 19336 22456
rect 19272 22396 19276 22452
rect 19276 22396 19332 22452
rect 19332 22396 19336 22452
rect 19272 22392 19336 22396
rect 19352 22452 19416 22456
rect 19352 22396 19356 22452
rect 19356 22396 19412 22452
rect 19412 22396 19416 22452
rect 19352 22392 19416 22396
rect 29112 22452 29176 22456
rect 29112 22396 29116 22452
rect 29116 22396 29172 22452
rect 29172 22396 29176 22452
rect 29112 22392 29176 22396
rect 29192 22452 29256 22456
rect 29192 22396 29196 22452
rect 29196 22396 29252 22452
rect 29252 22396 29256 22452
rect 29192 22392 29256 22396
rect 29272 22452 29336 22456
rect 29272 22396 29276 22452
rect 29276 22396 29332 22452
rect 29332 22396 29336 22452
rect 29272 22392 29336 22396
rect 29352 22452 29416 22456
rect 29352 22396 29356 22452
rect 29356 22396 29412 22452
rect 29412 22396 29416 22452
rect 29352 22392 29416 22396
rect 14112 21908 14176 21912
rect 14112 21852 14116 21908
rect 14116 21852 14172 21908
rect 14172 21852 14176 21908
rect 14112 21848 14176 21852
rect 14192 21908 14256 21912
rect 14192 21852 14196 21908
rect 14196 21852 14252 21908
rect 14252 21852 14256 21908
rect 14192 21848 14256 21852
rect 14272 21908 14336 21912
rect 14272 21852 14276 21908
rect 14276 21852 14332 21908
rect 14332 21852 14336 21908
rect 14272 21848 14336 21852
rect 14352 21908 14416 21912
rect 14352 21852 14356 21908
rect 14356 21852 14412 21908
rect 14412 21852 14416 21908
rect 14352 21848 14416 21852
rect 24112 21908 24176 21912
rect 24112 21852 24116 21908
rect 24116 21852 24172 21908
rect 24172 21852 24176 21908
rect 24112 21848 24176 21852
rect 24192 21908 24256 21912
rect 24192 21852 24196 21908
rect 24196 21852 24252 21908
rect 24252 21852 24256 21908
rect 24192 21848 24256 21852
rect 24272 21908 24336 21912
rect 24272 21852 24276 21908
rect 24276 21852 24332 21908
rect 24332 21852 24336 21908
rect 24272 21848 24336 21852
rect 24352 21908 24416 21912
rect 24352 21852 24356 21908
rect 24356 21852 24412 21908
rect 24412 21852 24416 21908
rect 24352 21848 24416 21852
rect 19112 21364 19176 21368
rect 19112 21308 19116 21364
rect 19116 21308 19172 21364
rect 19172 21308 19176 21364
rect 19112 21304 19176 21308
rect 19192 21364 19256 21368
rect 19192 21308 19196 21364
rect 19196 21308 19252 21364
rect 19252 21308 19256 21364
rect 19192 21304 19256 21308
rect 19272 21364 19336 21368
rect 19272 21308 19276 21364
rect 19276 21308 19332 21364
rect 19332 21308 19336 21364
rect 19272 21304 19336 21308
rect 19352 21364 19416 21368
rect 19352 21308 19356 21364
rect 19356 21308 19412 21364
rect 19412 21308 19416 21364
rect 19352 21304 19416 21308
rect 29112 21364 29176 21368
rect 29112 21308 29116 21364
rect 29116 21308 29172 21364
rect 29172 21308 29176 21364
rect 29112 21304 29176 21308
rect 29192 21364 29256 21368
rect 29192 21308 29196 21364
rect 29196 21308 29252 21364
rect 29252 21308 29256 21364
rect 29192 21304 29256 21308
rect 29272 21364 29336 21368
rect 29272 21308 29276 21364
rect 29276 21308 29332 21364
rect 29332 21308 29336 21364
rect 29272 21304 29336 21308
rect 29352 21364 29416 21368
rect 29352 21308 29356 21364
rect 29356 21308 29412 21364
rect 29412 21308 29416 21364
rect 29352 21304 29416 21308
rect 14112 20820 14176 20824
rect 14112 20764 14116 20820
rect 14116 20764 14172 20820
rect 14172 20764 14176 20820
rect 14112 20760 14176 20764
rect 14192 20820 14256 20824
rect 14192 20764 14196 20820
rect 14196 20764 14252 20820
rect 14252 20764 14256 20820
rect 14192 20760 14256 20764
rect 14272 20820 14336 20824
rect 14272 20764 14276 20820
rect 14276 20764 14332 20820
rect 14332 20764 14336 20820
rect 14272 20760 14336 20764
rect 14352 20820 14416 20824
rect 14352 20764 14356 20820
rect 14356 20764 14412 20820
rect 14412 20764 14416 20820
rect 14352 20760 14416 20764
rect 24112 20820 24176 20824
rect 24112 20764 24116 20820
rect 24116 20764 24172 20820
rect 24172 20764 24176 20820
rect 24112 20760 24176 20764
rect 24192 20820 24256 20824
rect 24192 20764 24196 20820
rect 24196 20764 24252 20820
rect 24252 20764 24256 20820
rect 24192 20760 24256 20764
rect 24272 20820 24336 20824
rect 24272 20764 24276 20820
rect 24276 20764 24332 20820
rect 24332 20764 24336 20820
rect 24272 20760 24336 20764
rect 24352 20820 24416 20824
rect 24352 20764 24356 20820
rect 24356 20764 24412 20820
rect 24412 20764 24416 20820
rect 24352 20760 24416 20764
rect 19112 20276 19176 20280
rect 19112 20220 19116 20276
rect 19116 20220 19172 20276
rect 19172 20220 19176 20276
rect 19112 20216 19176 20220
rect 19192 20276 19256 20280
rect 19192 20220 19196 20276
rect 19196 20220 19252 20276
rect 19252 20220 19256 20276
rect 19192 20216 19256 20220
rect 19272 20276 19336 20280
rect 19272 20220 19276 20276
rect 19276 20220 19332 20276
rect 19332 20220 19336 20276
rect 19272 20216 19336 20220
rect 19352 20276 19416 20280
rect 19352 20220 19356 20276
rect 19356 20220 19412 20276
rect 19412 20220 19416 20276
rect 19352 20216 19416 20220
rect 29112 20276 29176 20280
rect 29112 20220 29116 20276
rect 29116 20220 29172 20276
rect 29172 20220 29176 20276
rect 29112 20216 29176 20220
rect 29192 20276 29256 20280
rect 29192 20220 29196 20276
rect 29196 20220 29252 20276
rect 29252 20220 29256 20276
rect 29192 20216 29256 20220
rect 29272 20276 29336 20280
rect 29272 20220 29276 20276
rect 29276 20220 29332 20276
rect 29332 20220 29336 20276
rect 29272 20216 29336 20220
rect 29352 20276 29416 20280
rect 29352 20220 29356 20276
rect 29356 20220 29412 20276
rect 29412 20220 29416 20276
rect 29352 20216 29416 20220
rect 14112 19732 14176 19736
rect 14112 19676 14116 19732
rect 14116 19676 14172 19732
rect 14172 19676 14176 19732
rect 14112 19672 14176 19676
rect 14192 19732 14256 19736
rect 14192 19676 14196 19732
rect 14196 19676 14252 19732
rect 14252 19676 14256 19732
rect 14192 19672 14256 19676
rect 14272 19732 14336 19736
rect 14272 19676 14276 19732
rect 14276 19676 14332 19732
rect 14332 19676 14336 19732
rect 14272 19672 14336 19676
rect 14352 19732 14416 19736
rect 14352 19676 14356 19732
rect 14356 19676 14412 19732
rect 14412 19676 14416 19732
rect 14352 19672 14416 19676
rect 24112 19732 24176 19736
rect 24112 19676 24116 19732
rect 24116 19676 24172 19732
rect 24172 19676 24176 19732
rect 24112 19672 24176 19676
rect 24192 19732 24256 19736
rect 24192 19676 24196 19732
rect 24196 19676 24252 19732
rect 24252 19676 24256 19732
rect 24192 19672 24256 19676
rect 24272 19732 24336 19736
rect 24272 19676 24276 19732
rect 24276 19676 24332 19732
rect 24332 19676 24336 19732
rect 24272 19672 24336 19676
rect 24352 19732 24416 19736
rect 24352 19676 24356 19732
rect 24356 19676 24412 19732
rect 24412 19676 24416 19732
rect 24352 19672 24416 19676
rect 19112 19188 19176 19192
rect 19112 19132 19116 19188
rect 19116 19132 19172 19188
rect 19172 19132 19176 19188
rect 19112 19128 19176 19132
rect 19192 19188 19256 19192
rect 19192 19132 19196 19188
rect 19196 19132 19252 19188
rect 19252 19132 19256 19188
rect 19192 19128 19256 19132
rect 19272 19188 19336 19192
rect 19272 19132 19276 19188
rect 19276 19132 19332 19188
rect 19332 19132 19336 19188
rect 19272 19128 19336 19132
rect 19352 19188 19416 19192
rect 19352 19132 19356 19188
rect 19356 19132 19412 19188
rect 19412 19132 19416 19188
rect 19352 19128 19416 19132
rect 29112 19188 29176 19192
rect 29112 19132 29116 19188
rect 29116 19132 29172 19188
rect 29172 19132 29176 19188
rect 29112 19128 29176 19132
rect 29192 19188 29256 19192
rect 29192 19132 29196 19188
rect 29196 19132 29252 19188
rect 29252 19132 29256 19188
rect 29192 19128 29256 19132
rect 29272 19188 29336 19192
rect 29272 19132 29276 19188
rect 29276 19132 29332 19188
rect 29332 19132 29336 19188
rect 29272 19128 29336 19132
rect 29352 19188 29416 19192
rect 29352 19132 29356 19188
rect 29356 19132 29412 19188
rect 29412 19132 29416 19188
rect 29352 19128 29416 19132
rect 14112 18644 14176 18648
rect 14112 18588 14116 18644
rect 14116 18588 14172 18644
rect 14172 18588 14176 18644
rect 14112 18584 14176 18588
rect 14192 18644 14256 18648
rect 14192 18588 14196 18644
rect 14196 18588 14252 18644
rect 14252 18588 14256 18644
rect 14192 18584 14256 18588
rect 14272 18644 14336 18648
rect 14272 18588 14276 18644
rect 14276 18588 14332 18644
rect 14332 18588 14336 18644
rect 14272 18584 14336 18588
rect 14352 18644 14416 18648
rect 14352 18588 14356 18644
rect 14356 18588 14412 18644
rect 14412 18588 14416 18644
rect 14352 18584 14416 18588
rect 24112 18644 24176 18648
rect 24112 18588 24116 18644
rect 24116 18588 24172 18644
rect 24172 18588 24176 18644
rect 24112 18584 24176 18588
rect 24192 18644 24256 18648
rect 24192 18588 24196 18644
rect 24196 18588 24252 18644
rect 24252 18588 24256 18644
rect 24192 18584 24256 18588
rect 24272 18644 24336 18648
rect 24272 18588 24276 18644
rect 24276 18588 24332 18644
rect 24332 18588 24336 18644
rect 24272 18584 24336 18588
rect 24352 18644 24416 18648
rect 24352 18588 24356 18644
rect 24356 18588 24412 18644
rect 24412 18588 24416 18644
rect 24352 18584 24416 18588
rect 19112 18100 19176 18104
rect 19112 18044 19116 18100
rect 19116 18044 19172 18100
rect 19172 18044 19176 18100
rect 19112 18040 19176 18044
rect 19192 18100 19256 18104
rect 19192 18044 19196 18100
rect 19196 18044 19252 18100
rect 19252 18044 19256 18100
rect 19192 18040 19256 18044
rect 19272 18100 19336 18104
rect 19272 18044 19276 18100
rect 19276 18044 19332 18100
rect 19332 18044 19336 18100
rect 19272 18040 19336 18044
rect 19352 18100 19416 18104
rect 19352 18044 19356 18100
rect 19356 18044 19412 18100
rect 19412 18044 19416 18100
rect 19352 18040 19416 18044
rect 29112 18100 29176 18104
rect 29112 18044 29116 18100
rect 29116 18044 29172 18100
rect 29172 18044 29176 18100
rect 29112 18040 29176 18044
rect 29192 18100 29256 18104
rect 29192 18044 29196 18100
rect 29196 18044 29252 18100
rect 29252 18044 29256 18100
rect 29192 18040 29256 18044
rect 29272 18100 29336 18104
rect 29272 18044 29276 18100
rect 29276 18044 29332 18100
rect 29332 18044 29336 18100
rect 29272 18040 29336 18044
rect 29352 18100 29416 18104
rect 29352 18044 29356 18100
rect 29356 18044 29412 18100
rect 29412 18044 29416 18100
rect 29352 18040 29416 18044
rect 14112 17556 14176 17560
rect 14112 17500 14116 17556
rect 14116 17500 14172 17556
rect 14172 17500 14176 17556
rect 14112 17496 14176 17500
rect 14192 17556 14256 17560
rect 14192 17500 14196 17556
rect 14196 17500 14252 17556
rect 14252 17500 14256 17556
rect 14192 17496 14256 17500
rect 14272 17556 14336 17560
rect 14272 17500 14276 17556
rect 14276 17500 14332 17556
rect 14332 17500 14336 17556
rect 14272 17496 14336 17500
rect 14352 17556 14416 17560
rect 14352 17500 14356 17556
rect 14356 17500 14412 17556
rect 14412 17500 14416 17556
rect 14352 17496 14416 17500
rect 24112 17556 24176 17560
rect 24112 17500 24116 17556
rect 24116 17500 24172 17556
rect 24172 17500 24176 17556
rect 24112 17496 24176 17500
rect 24192 17556 24256 17560
rect 24192 17500 24196 17556
rect 24196 17500 24252 17556
rect 24252 17500 24256 17556
rect 24192 17496 24256 17500
rect 24272 17556 24336 17560
rect 24272 17500 24276 17556
rect 24276 17500 24332 17556
rect 24332 17500 24336 17556
rect 24272 17496 24336 17500
rect 24352 17556 24416 17560
rect 24352 17500 24356 17556
rect 24356 17500 24412 17556
rect 24412 17500 24416 17556
rect 24352 17496 24416 17500
rect 19112 17012 19176 17016
rect 19112 16956 19116 17012
rect 19116 16956 19172 17012
rect 19172 16956 19176 17012
rect 19112 16952 19176 16956
rect 19192 17012 19256 17016
rect 19192 16956 19196 17012
rect 19196 16956 19252 17012
rect 19252 16956 19256 17012
rect 19192 16952 19256 16956
rect 19272 17012 19336 17016
rect 19272 16956 19276 17012
rect 19276 16956 19332 17012
rect 19332 16956 19336 17012
rect 19272 16952 19336 16956
rect 19352 17012 19416 17016
rect 19352 16956 19356 17012
rect 19356 16956 19412 17012
rect 19412 16956 19416 17012
rect 19352 16952 19416 16956
rect 29112 17012 29176 17016
rect 29112 16956 29116 17012
rect 29116 16956 29172 17012
rect 29172 16956 29176 17012
rect 29112 16952 29176 16956
rect 29192 17012 29256 17016
rect 29192 16956 29196 17012
rect 29196 16956 29252 17012
rect 29252 16956 29256 17012
rect 29192 16952 29256 16956
rect 29272 17012 29336 17016
rect 29272 16956 29276 17012
rect 29276 16956 29332 17012
rect 29332 16956 29336 17012
rect 29272 16952 29336 16956
rect 29352 17012 29416 17016
rect 29352 16956 29356 17012
rect 29356 16956 29412 17012
rect 29412 16956 29416 17012
rect 29352 16952 29416 16956
rect 14112 16468 14176 16472
rect 14112 16412 14116 16468
rect 14116 16412 14172 16468
rect 14172 16412 14176 16468
rect 14112 16408 14176 16412
rect 14192 16468 14256 16472
rect 14192 16412 14196 16468
rect 14196 16412 14252 16468
rect 14252 16412 14256 16468
rect 14192 16408 14256 16412
rect 14272 16468 14336 16472
rect 14272 16412 14276 16468
rect 14276 16412 14332 16468
rect 14332 16412 14336 16468
rect 14272 16408 14336 16412
rect 14352 16468 14416 16472
rect 14352 16412 14356 16468
rect 14356 16412 14412 16468
rect 14412 16412 14416 16468
rect 14352 16408 14416 16412
rect 24112 16468 24176 16472
rect 24112 16412 24116 16468
rect 24116 16412 24172 16468
rect 24172 16412 24176 16468
rect 24112 16408 24176 16412
rect 24192 16468 24256 16472
rect 24192 16412 24196 16468
rect 24196 16412 24252 16468
rect 24252 16412 24256 16468
rect 24192 16408 24256 16412
rect 24272 16468 24336 16472
rect 24272 16412 24276 16468
rect 24276 16412 24332 16468
rect 24332 16412 24336 16468
rect 24272 16408 24336 16412
rect 24352 16468 24416 16472
rect 24352 16412 24356 16468
rect 24356 16412 24412 16468
rect 24412 16412 24416 16468
rect 24352 16408 24416 16412
rect 19112 15924 19176 15928
rect 19112 15868 19116 15924
rect 19116 15868 19172 15924
rect 19172 15868 19176 15924
rect 19112 15864 19176 15868
rect 19192 15924 19256 15928
rect 19192 15868 19196 15924
rect 19196 15868 19252 15924
rect 19252 15868 19256 15924
rect 19192 15864 19256 15868
rect 19272 15924 19336 15928
rect 19272 15868 19276 15924
rect 19276 15868 19332 15924
rect 19332 15868 19336 15924
rect 19272 15864 19336 15868
rect 19352 15924 19416 15928
rect 19352 15868 19356 15924
rect 19356 15868 19412 15924
rect 19412 15868 19416 15924
rect 19352 15864 19416 15868
rect 29112 15924 29176 15928
rect 29112 15868 29116 15924
rect 29116 15868 29172 15924
rect 29172 15868 29176 15924
rect 29112 15864 29176 15868
rect 29192 15924 29256 15928
rect 29192 15868 29196 15924
rect 29196 15868 29252 15924
rect 29252 15868 29256 15924
rect 29192 15864 29256 15868
rect 29272 15924 29336 15928
rect 29272 15868 29276 15924
rect 29276 15868 29332 15924
rect 29332 15868 29336 15924
rect 29272 15864 29336 15868
rect 29352 15924 29416 15928
rect 29352 15868 29356 15924
rect 29356 15868 29412 15924
rect 29412 15868 29416 15924
rect 29352 15864 29416 15868
rect 14112 15380 14176 15384
rect 14112 15324 14116 15380
rect 14116 15324 14172 15380
rect 14172 15324 14176 15380
rect 14112 15320 14176 15324
rect 14192 15380 14256 15384
rect 14192 15324 14196 15380
rect 14196 15324 14252 15380
rect 14252 15324 14256 15380
rect 14192 15320 14256 15324
rect 14272 15380 14336 15384
rect 14272 15324 14276 15380
rect 14276 15324 14332 15380
rect 14332 15324 14336 15380
rect 14272 15320 14336 15324
rect 14352 15380 14416 15384
rect 14352 15324 14356 15380
rect 14356 15324 14412 15380
rect 14412 15324 14416 15380
rect 14352 15320 14416 15324
rect 24112 15380 24176 15384
rect 24112 15324 24116 15380
rect 24116 15324 24172 15380
rect 24172 15324 24176 15380
rect 24112 15320 24176 15324
rect 24192 15380 24256 15384
rect 24192 15324 24196 15380
rect 24196 15324 24252 15380
rect 24252 15324 24256 15380
rect 24192 15320 24256 15324
rect 24272 15380 24336 15384
rect 24272 15324 24276 15380
rect 24276 15324 24332 15380
rect 24332 15324 24336 15380
rect 24272 15320 24336 15324
rect 24352 15380 24416 15384
rect 24352 15324 24356 15380
rect 24356 15324 24412 15380
rect 24412 15324 24416 15380
rect 24352 15320 24416 15324
rect 19112 14836 19176 14840
rect 19112 14780 19116 14836
rect 19116 14780 19172 14836
rect 19172 14780 19176 14836
rect 19112 14776 19176 14780
rect 19192 14836 19256 14840
rect 19192 14780 19196 14836
rect 19196 14780 19252 14836
rect 19252 14780 19256 14836
rect 19192 14776 19256 14780
rect 19272 14836 19336 14840
rect 19272 14780 19276 14836
rect 19276 14780 19332 14836
rect 19332 14780 19336 14836
rect 19272 14776 19336 14780
rect 19352 14836 19416 14840
rect 19352 14780 19356 14836
rect 19356 14780 19412 14836
rect 19412 14780 19416 14836
rect 19352 14776 19416 14780
rect 29112 14836 29176 14840
rect 29112 14780 29116 14836
rect 29116 14780 29172 14836
rect 29172 14780 29176 14836
rect 29112 14776 29176 14780
rect 29192 14836 29256 14840
rect 29192 14780 29196 14836
rect 29196 14780 29252 14836
rect 29252 14780 29256 14836
rect 29192 14776 29256 14780
rect 29272 14836 29336 14840
rect 29272 14780 29276 14836
rect 29276 14780 29332 14836
rect 29332 14780 29336 14836
rect 29272 14776 29336 14780
rect 29352 14836 29416 14840
rect 29352 14780 29356 14836
rect 29356 14780 29412 14836
rect 29412 14780 29416 14836
rect 29352 14776 29416 14780
rect 14112 14292 14176 14296
rect 14112 14236 14116 14292
rect 14116 14236 14172 14292
rect 14172 14236 14176 14292
rect 14112 14232 14176 14236
rect 14192 14292 14256 14296
rect 14192 14236 14196 14292
rect 14196 14236 14252 14292
rect 14252 14236 14256 14292
rect 14192 14232 14256 14236
rect 14272 14292 14336 14296
rect 14272 14236 14276 14292
rect 14276 14236 14332 14292
rect 14332 14236 14336 14292
rect 14272 14232 14336 14236
rect 14352 14292 14416 14296
rect 14352 14236 14356 14292
rect 14356 14236 14412 14292
rect 14412 14236 14416 14292
rect 14352 14232 14416 14236
rect 24112 14292 24176 14296
rect 24112 14236 24116 14292
rect 24116 14236 24172 14292
rect 24172 14236 24176 14292
rect 24112 14232 24176 14236
rect 24192 14292 24256 14296
rect 24192 14236 24196 14292
rect 24196 14236 24252 14292
rect 24252 14236 24256 14292
rect 24192 14232 24256 14236
rect 24272 14292 24336 14296
rect 24272 14236 24276 14292
rect 24276 14236 24332 14292
rect 24332 14236 24336 14292
rect 24272 14232 24336 14236
rect 24352 14292 24416 14296
rect 24352 14236 24356 14292
rect 24356 14236 24412 14292
rect 24412 14236 24416 14292
rect 24352 14232 24416 14236
rect 19112 13748 19176 13752
rect 19112 13692 19116 13748
rect 19116 13692 19172 13748
rect 19172 13692 19176 13748
rect 19112 13688 19176 13692
rect 19192 13748 19256 13752
rect 19192 13692 19196 13748
rect 19196 13692 19252 13748
rect 19252 13692 19256 13748
rect 19192 13688 19256 13692
rect 19272 13748 19336 13752
rect 19272 13692 19276 13748
rect 19276 13692 19332 13748
rect 19332 13692 19336 13748
rect 19272 13688 19336 13692
rect 19352 13748 19416 13752
rect 19352 13692 19356 13748
rect 19356 13692 19412 13748
rect 19412 13692 19416 13748
rect 19352 13688 19416 13692
rect 29112 13748 29176 13752
rect 29112 13692 29116 13748
rect 29116 13692 29172 13748
rect 29172 13692 29176 13748
rect 29112 13688 29176 13692
rect 29192 13748 29256 13752
rect 29192 13692 29196 13748
rect 29196 13692 29252 13748
rect 29252 13692 29256 13748
rect 29192 13688 29256 13692
rect 29272 13748 29336 13752
rect 29272 13692 29276 13748
rect 29276 13692 29332 13748
rect 29332 13692 29336 13748
rect 29272 13688 29336 13692
rect 29352 13748 29416 13752
rect 29352 13692 29356 13748
rect 29356 13692 29412 13748
rect 29412 13692 29416 13748
rect 29352 13688 29416 13692
rect 14112 13204 14176 13208
rect 14112 13148 14116 13204
rect 14116 13148 14172 13204
rect 14172 13148 14176 13204
rect 14112 13144 14176 13148
rect 14192 13204 14256 13208
rect 14192 13148 14196 13204
rect 14196 13148 14252 13204
rect 14252 13148 14256 13204
rect 14192 13144 14256 13148
rect 14272 13204 14336 13208
rect 14272 13148 14276 13204
rect 14276 13148 14332 13204
rect 14332 13148 14336 13204
rect 14272 13144 14336 13148
rect 14352 13204 14416 13208
rect 14352 13148 14356 13204
rect 14356 13148 14412 13204
rect 14412 13148 14416 13204
rect 14352 13144 14416 13148
rect 24112 13204 24176 13208
rect 24112 13148 24116 13204
rect 24116 13148 24172 13204
rect 24172 13148 24176 13204
rect 24112 13144 24176 13148
rect 24192 13204 24256 13208
rect 24192 13148 24196 13204
rect 24196 13148 24252 13204
rect 24252 13148 24256 13204
rect 24192 13144 24256 13148
rect 24272 13204 24336 13208
rect 24272 13148 24276 13204
rect 24276 13148 24332 13204
rect 24332 13148 24336 13204
rect 24272 13144 24336 13148
rect 24352 13204 24416 13208
rect 24352 13148 24356 13204
rect 24356 13148 24412 13204
rect 24412 13148 24416 13204
rect 24352 13144 24416 13148
rect 19112 12660 19176 12664
rect 19112 12604 19116 12660
rect 19116 12604 19172 12660
rect 19172 12604 19176 12660
rect 19112 12600 19176 12604
rect 19192 12660 19256 12664
rect 19192 12604 19196 12660
rect 19196 12604 19252 12660
rect 19252 12604 19256 12660
rect 19192 12600 19256 12604
rect 19272 12660 19336 12664
rect 19272 12604 19276 12660
rect 19276 12604 19332 12660
rect 19332 12604 19336 12660
rect 19272 12600 19336 12604
rect 19352 12660 19416 12664
rect 19352 12604 19356 12660
rect 19356 12604 19412 12660
rect 19412 12604 19416 12660
rect 19352 12600 19416 12604
rect 29112 12660 29176 12664
rect 29112 12604 29116 12660
rect 29116 12604 29172 12660
rect 29172 12604 29176 12660
rect 29112 12600 29176 12604
rect 29192 12660 29256 12664
rect 29192 12604 29196 12660
rect 29196 12604 29252 12660
rect 29252 12604 29256 12660
rect 29192 12600 29256 12604
rect 29272 12660 29336 12664
rect 29272 12604 29276 12660
rect 29276 12604 29332 12660
rect 29332 12604 29336 12660
rect 29272 12600 29336 12604
rect 29352 12660 29416 12664
rect 29352 12604 29356 12660
rect 29356 12604 29412 12660
rect 29412 12604 29416 12660
rect 29352 12600 29416 12604
rect 14112 12116 14176 12120
rect 14112 12060 14116 12116
rect 14116 12060 14172 12116
rect 14172 12060 14176 12116
rect 14112 12056 14176 12060
rect 14192 12116 14256 12120
rect 14192 12060 14196 12116
rect 14196 12060 14252 12116
rect 14252 12060 14256 12116
rect 14192 12056 14256 12060
rect 14272 12116 14336 12120
rect 14272 12060 14276 12116
rect 14276 12060 14332 12116
rect 14332 12060 14336 12116
rect 14272 12056 14336 12060
rect 14352 12116 14416 12120
rect 14352 12060 14356 12116
rect 14356 12060 14412 12116
rect 14412 12060 14416 12116
rect 14352 12056 14416 12060
rect 24112 12116 24176 12120
rect 24112 12060 24116 12116
rect 24116 12060 24172 12116
rect 24172 12060 24176 12116
rect 24112 12056 24176 12060
rect 24192 12116 24256 12120
rect 24192 12060 24196 12116
rect 24196 12060 24252 12116
rect 24252 12060 24256 12116
rect 24192 12056 24256 12060
rect 24272 12116 24336 12120
rect 24272 12060 24276 12116
rect 24276 12060 24332 12116
rect 24332 12060 24336 12116
rect 24272 12056 24336 12060
rect 24352 12116 24416 12120
rect 24352 12060 24356 12116
rect 24356 12060 24412 12116
rect 24412 12060 24416 12116
rect 24352 12056 24416 12060
rect 19112 11572 19176 11576
rect 19112 11516 19116 11572
rect 19116 11516 19172 11572
rect 19172 11516 19176 11572
rect 19112 11512 19176 11516
rect 19192 11572 19256 11576
rect 19192 11516 19196 11572
rect 19196 11516 19252 11572
rect 19252 11516 19256 11572
rect 19192 11512 19256 11516
rect 19272 11572 19336 11576
rect 19272 11516 19276 11572
rect 19276 11516 19332 11572
rect 19332 11516 19336 11572
rect 19272 11512 19336 11516
rect 19352 11572 19416 11576
rect 19352 11516 19356 11572
rect 19356 11516 19412 11572
rect 19412 11516 19416 11572
rect 19352 11512 19416 11516
rect 29112 11572 29176 11576
rect 29112 11516 29116 11572
rect 29116 11516 29172 11572
rect 29172 11516 29176 11572
rect 29112 11512 29176 11516
rect 29192 11572 29256 11576
rect 29192 11516 29196 11572
rect 29196 11516 29252 11572
rect 29252 11516 29256 11572
rect 29192 11512 29256 11516
rect 29272 11572 29336 11576
rect 29272 11516 29276 11572
rect 29276 11516 29332 11572
rect 29332 11516 29336 11572
rect 29272 11512 29336 11516
rect 29352 11572 29416 11576
rect 29352 11516 29356 11572
rect 29356 11516 29412 11572
rect 29412 11516 29416 11572
rect 29352 11512 29416 11516
rect 14112 11028 14176 11032
rect 14112 10972 14116 11028
rect 14116 10972 14172 11028
rect 14172 10972 14176 11028
rect 14112 10968 14176 10972
rect 14192 11028 14256 11032
rect 14192 10972 14196 11028
rect 14196 10972 14252 11028
rect 14252 10972 14256 11028
rect 14192 10968 14256 10972
rect 14272 11028 14336 11032
rect 14272 10972 14276 11028
rect 14276 10972 14332 11028
rect 14332 10972 14336 11028
rect 14272 10968 14336 10972
rect 14352 11028 14416 11032
rect 14352 10972 14356 11028
rect 14356 10972 14412 11028
rect 14412 10972 14416 11028
rect 14352 10968 14416 10972
rect 24112 11028 24176 11032
rect 24112 10972 24116 11028
rect 24116 10972 24172 11028
rect 24172 10972 24176 11028
rect 24112 10968 24176 10972
rect 24192 11028 24256 11032
rect 24192 10972 24196 11028
rect 24196 10972 24252 11028
rect 24252 10972 24256 11028
rect 24192 10968 24256 10972
rect 24272 11028 24336 11032
rect 24272 10972 24276 11028
rect 24276 10972 24332 11028
rect 24332 10972 24336 11028
rect 24272 10968 24336 10972
rect 24352 11028 24416 11032
rect 24352 10972 24356 11028
rect 24356 10972 24412 11028
rect 24412 10972 24416 11028
rect 24352 10968 24416 10972
rect 5008 5008 8992 8992
rect 14112 5008 14416 8992
rect 24112 5008 24416 8992
rect 32144 5008 36128 8992
rect 8 8 3992 3992
rect 19112 8 19416 3992
rect 29112 8 29416 3992
rect 37144 8 41128 3992
<< metal4 >>
rect 0 41032 4000 41040
rect 0 37048 8 41032
rect 3992 37048 4000 41032
rect 0 3992 4000 37048
rect 5000 36032 9000 36040
rect 5000 32048 5008 36032
rect 8992 32048 9000 36032
rect 5000 8992 9000 32048
rect 5000 5008 5008 8992
rect 8992 5008 9000 8992
rect 5000 5000 9000 5008
rect 14104 36032 14424 41040
rect 14104 32048 14112 36032
rect 14416 32048 14424 36032
rect 14104 29528 14424 32048
rect 14104 29464 14112 29528
rect 14176 29464 14192 29528
rect 14256 29464 14272 29528
rect 14336 29464 14352 29528
rect 14416 29464 14424 29528
rect 14104 28440 14424 29464
rect 14104 28376 14112 28440
rect 14176 28376 14192 28440
rect 14256 28376 14272 28440
rect 14336 28376 14352 28440
rect 14416 28376 14424 28440
rect 14104 27352 14424 28376
rect 14104 27288 14112 27352
rect 14176 27288 14192 27352
rect 14256 27288 14272 27352
rect 14336 27288 14352 27352
rect 14416 27288 14424 27352
rect 14104 26264 14424 27288
rect 14104 26200 14112 26264
rect 14176 26200 14192 26264
rect 14256 26200 14272 26264
rect 14336 26200 14352 26264
rect 14416 26200 14424 26264
rect 14104 25176 14424 26200
rect 14104 25112 14112 25176
rect 14176 25112 14192 25176
rect 14256 25112 14272 25176
rect 14336 25112 14352 25176
rect 14416 25112 14424 25176
rect 14104 24088 14424 25112
rect 14104 24024 14112 24088
rect 14176 24024 14192 24088
rect 14256 24024 14272 24088
rect 14336 24024 14352 24088
rect 14416 24024 14424 24088
rect 14104 23000 14424 24024
rect 14104 22936 14112 23000
rect 14176 22936 14192 23000
rect 14256 22936 14272 23000
rect 14336 22936 14352 23000
rect 14416 22936 14424 23000
rect 14104 21912 14424 22936
rect 14104 21848 14112 21912
rect 14176 21848 14192 21912
rect 14256 21848 14272 21912
rect 14336 21848 14352 21912
rect 14416 21848 14424 21912
rect 14104 20824 14424 21848
rect 14104 20760 14112 20824
rect 14176 20760 14192 20824
rect 14256 20760 14272 20824
rect 14336 20760 14352 20824
rect 14416 20760 14424 20824
rect 14104 19736 14424 20760
rect 14104 19672 14112 19736
rect 14176 19672 14192 19736
rect 14256 19672 14272 19736
rect 14336 19672 14352 19736
rect 14416 19672 14424 19736
rect 14104 18648 14424 19672
rect 14104 18584 14112 18648
rect 14176 18584 14192 18648
rect 14256 18584 14272 18648
rect 14336 18584 14352 18648
rect 14416 18584 14424 18648
rect 14104 17560 14424 18584
rect 14104 17496 14112 17560
rect 14176 17496 14192 17560
rect 14256 17496 14272 17560
rect 14336 17496 14352 17560
rect 14416 17496 14424 17560
rect 14104 16472 14424 17496
rect 14104 16408 14112 16472
rect 14176 16408 14192 16472
rect 14256 16408 14272 16472
rect 14336 16408 14352 16472
rect 14416 16408 14424 16472
rect 14104 15384 14424 16408
rect 14104 15320 14112 15384
rect 14176 15320 14192 15384
rect 14256 15320 14272 15384
rect 14336 15320 14352 15384
rect 14416 15320 14424 15384
rect 14104 14296 14424 15320
rect 14104 14232 14112 14296
rect 14176 14232 14192 14296
rect 14256 14232 14272 14296
rect 14336 14232 14352 14296
rect 14416 14232 14424 14296
rect 14104 13208 14424 14232
rect 14104 13144 14112 13208
rect 14176 13144 14192 13208
rect 14256 13144 14272 13208
rect 14336 13144 14352 13208
rect 14416 13144 14424 13208
rect 14104 12120 14424 13144
rect 14104 12056 14112 12120
rect 14176 12056 14192 12120
rect 14256 12056 14272 12120
rect 14336 12056 14352 12120
rect 14416 12056 14424 12120
rect 14104 11032 14424 12056
rect 14104 10968 14112 11032
rect 14176 10968 14192 11032
rect 14256 10968 14272 11032
rect 14336 10968 14352 11032
rect 14416 10968 14424 11032
rect 14104 8992 14424 10968
rect 14104 5008 14112 8992
rect 14416 5008 14424 8992
rect 0 8 8 3992
rect 3992 8 4000 3992
rect 0 0 4000 8
rect 14104 0 14424 5008
rect 19104 41032 19424 41040
rect 19104 37048 19112 41032
rect 19416 37048 19424 41032
rect 19104 30072 19424 37048
rect 19104 30008 19112 30072
rect 19176 30008 19192 30072
rect 19256 30008 19272 30072
rect 19336 30008 19352 30072
rect 19416 30008 19424 30072
rect 19104 28984 19424 30008
rect 19104 28920 19112 28984
rect 19176 28920 19192 28984
rect 19256 28920 19272 28984
rect 19336 28920 19352 28984
rect 19416 28920 19424 28984
rect 19104 27896 19424 28920
rect 19104 27832 19112 27896
rect 19176 27832 19192 27896
rect 19256 27832 19272 27896
rect 19336 27832 19352 27896
rect 19416 27832 19424 27896
rect 19104 26808 19424 27832
rect 19104 26744 19112 26808
rect 19176 26744 19192 26808
rect 19256 26744 19272 26808
rect 19336 26744 19352 26808
rect 19416 26744 19424 26808
rect 19104 25720 19424 26744
rect 19104 25656 19112 25720
rect 19176 25656 19192 25720
rect 19256 25656 19272 25720
rect 19336 25656 19352 25720
rect 19416 25656 19424 25720
rect 19104 24632 19424 25656
rect 19104 24568 19112 24632
rect 19176 24568 19192 24632
rect 19256 24568 19272 24632
rect 19336 24568 19352 24632
rect 19416 24568 19424 24632
rect 19104 23544 19424 24568
rect 19104 23480 19112 23544
rect 19176 23480 19192 23544
rect 19256 23480 19272 23544
rect 19336 23480 19352 23544
rect 19416 23480 19424 23544
rect 19104 22456 19424 23480
rect 19104 22392 19112 22456
rect 19176 22392 19192 22456
rect 19256 22392 19272 22456
rect 19336 22392 19352 22456
rect 19416 22392 19424 22456
rect 19104 21368 19424 22392
rect 19104 21304 19112 21368
rect 19176 21304 19192 21368
rect 19256 21304 19272 21368
rect 19336 21304 19352 21368
rect 19416 21304 19424 21368
rect 19104 20280 19424 21304
rect 19104 20216 19112 20280
rect 19176 20216 19192 20280
rect 19256 20216 19272 20280
rect 19336 20216 19352 20280
rect 19416 20216 19424 20280
rect 19104 19192 19424 20216
rect 19104 19128 19112 19192
rect 19176 19128 19192 19192
rect 19256 19128 19272 19192
rect 19336 19128 19352 19192
rect 19416 19128 19424 19192
rect 19104 18104 19424 19128
rect 19104 18040 19112 18104
rect 19176 18040 19192 18104
rect 19256 18040 19272 18104
rect 19336 18040 19352 18104
rect 19416 18040 19424 18104
rect 19104 17016 19424 18040
rect 19104 16952 19112 17016
rect 19176 16952 19192 17016
rect 19256 16952 19272 17016
rect 19336 16952 19352 17016
rect 19416 16952 19424 17016
rect 19104 15928 19424 16952
rect 19104 15864 19112 15928
rect 19176 15864 19192 15928
rect 19256 15864 19272 15928
rect 19336 15864 19352 15928
rect 19416 15864 19424 15928
rect 19104 14840 19424 15864
rect 19104 14776 19112 14840
rect 19176 14776 19192 14840
rect 19256 14776 19272 14840
rect 19336 14776 19352 14840
rect 19416 14776 19424 14840
rect 19104 13752 19424 14776
rect 19104 13688 19112 13752
rect 19176 13688 19192 13752
rect 19256 13688 19272 13752
rect 19336 13688 19352 13752
rect 19416 13688 19424 13752
rect 19104 12664 19424 13688
rect 19104 12600 19112 12664
rect 19176 12600 19192 12664
rect 19256 12600 19272 12664
rect 19336 12600 19352 12664
rect 19416 12600 19424 12664
rect 19104 11576 19424 12600
rect 19104 11512 19112 11576
rect 19176 11512 19192 11576
rect 19256 11512 19272 11576
rect 19336 11512 19352 11576
rect 19416 11512 19424 11576
rect 19104 3992 19424 11512
rect 19104 8 19112 3992
rect 19416 8 19424 3992
rect 19104 0 19424 8
rect 24104 36032 24424 41040
rect 24104 32048 24112 36032
rect 24416 32048 24424 36032
rect 24104 29528 24424 32048
rect 24104 29464 24112 29528
rect 24176 29464 24192 29528
rect 24256 29464 24272 29528
rect 24336 29464 24352 29528
rect 24416 29464 24424 29528
rect 24104 28440 24424 29464
rect 24104 28376 24112 28440
rect 24176 28376 24192 28440
rect 24256 28376 24272 28440
rect 24336 28376 24352 28440
rect 24416 28376 24424 28440
rect 24104 27352 24424 28376
rect 24104 27288 24112 27352
rect 24176 27288 24192 27352
rect 24256 27288 24272 27352
rect 24336 27288 24352 27352
rect 24416 27288 24424 27352
rect 24104 26264 24424 27288
rect 24104 26200 24112 26264
rect 24176 26200 24192 26264
rect 24256 26200 24272 26264
rect 24336 26200 24352 26264
rect 24416 26200 24424 26264
rect 24104 25176 24424 26200
rect 24104 25112 24112 25176
rect 24176 25112 24192 25176
rect 24256 25112 24272 25176
rect 24336 25112 24352 25176
rect 24416 25112 24424 25176
rect 24104 24088 24424 25112
rect 24104 24024 24112 24088
rect 24176 24024 24192 24088
rect 24256 24024 24272 24088
rect 24336 24024 24352 24088
rect 24416 24024 24424 24088
rect 24104 23000 24424 24024
rect 24104 22936 24112 23000
rect 24176 22936 24192 23000
rect 24256 22936 24272 23000
rect 24336 22936 24352 23000
rect 24416 22936 24424 23000
rect 24104 21912 24424 22936
rect 24104 21848 24112 21912
rect 24176 21848 24192 21912
rect 24256 21848 24272 21912
rect 24336 21848 24352 21912
rect 24416 21848 24424 21912
rect 24104 20824 24424 21848
rect 24104 20760 24112 20824
rect 24176 20760 24192 20824
rect 24256 20760 24272 20824
rect 24336 20760 24352 20824
rect 24416 20760 24424 20824
rect 24104 19736 24424 20760
rect 24104 19672 24112 19736
rect 24176 19672 24192 19736
rect 24256 19672 24272 19736
rect 24336 19672 24352 19736
rect 24416 19672 24424 19736
rect 24104 18648 24424 19672
rect 24104 18584 24112 18648
rect 24176 18584 24192 18648
rect 24256 18584 24272 18648
rect 24336 18584 24352 18648
rect 24416 18584 24424 18648
rect 24104 17560 24424 18584
rect 24104 17496 24112 17560
rect 24176 17496 24192 17560
rect 24256 17496 24272 17560
rect 24336 17496 24352 17560
rect 24416 17496 24424 17560
rect 24104 16472 24424 17496
rect 24104 16408 24112 16472
rect 24176 16408 24192 16472
rect 24256 16408 24272 16472
rect 24336 16408 24352 16472
rect 24416 16408 24424 16472
rect 24104 15384 24424 16408
rect 24104 15320 24112 15384
rect 24176 15320 24192 15384
rect 24256 15320 24272 15384
rect 24336 15320 24352 15384
rect 24416 15320 24424 15384
rect 24104 14296 24424 15320
rect 24104 14232 24112 14296
rect 24176 14232 24192 14296
rect 24256 14232 24272 14296
rect 24336 14232 24352 14296
rect 24416 14232 24424 14296
rect 24104 13208 24424 14232
rect 24104 13144 24112 13208
rect 24176 13144 24192 13208
rect 24256 13144 24272 13208
rect 24336 13144 24352 13208
rect 24416 13144 24424 13208
rect 24104 12120 24424 13144
rect 24104 12056 24112 12120
rect 24176 12056 24192 12120
rect 24256 12056 24272 12120
rect 24336 12056 24352 12120
rect 24416 12056 24424 12120
rect 24104 11032 24424 12056
rect 24104 10968 24112 11032
rect 24176 10968 24192 11032
rect 24256 10968 24272 11032
rect 24336 10968 24352 11032
rect 24416 10968 24424 11032
rect 24104 8992 24424 10968
rect 24104 5008 24112 8992
rect 24416 5008 24424 8992
rect 24104 0 24424 5008
rect 29104 41032 29424 41040
rect 29104 37048 29112 41032
rect 29416 37048 29424 41032
rect 29104 30072 29424 37048
rect 37136 41032 41136 41040
rect 37136 37048 37144 41032
rect 41128 37048 41136 41032
rect 29104 30008 29112 30072
rect 29176 30008 29192 30072
rect 29256 30008 29272 30072
rect 29336 30008 29352 30072
rect 29416 30008 29424 30072
rect 29104 28984 29424 30008
rect 29104 28920 29112 28984
rect 29176 28920 29192 28984
rect 29256 28920 29272 28984
rect 29336 28920 29352 28984
rect 29416 28920 29424 28984
rect 29104 27896 29424 28920
rect 29104 27832 29112 27896
rect 29176 27832 29192 27896
rect 29256 27832 29272 27896
rect 29336 27832 29352 27896
rect 29416 27832 29424 27896
rect 29104 26808 29424 27832
rect 29104 26744 29112 26808
rect 29176 26744 29192 26808
rect 29256 26744 29272 26808
rect 29336 26744 29352 26808
rect 29416 26744 29424 26808
rect 29104 25720 29424 26744
rect 29104 25656 29112 25720
rect 29176 25656 29192 25720
rect 29256 25656 29272 25720
rect 29336 25656 29352 25720
rect 29416 25656 29424 25720
rect 29104 24632 29424 25656
rect 29104 24568 29112 24632
rect 29176 24568 29192 24632
rect 29256 24568 29272 24632
rect 29336 24568 29352 24632
rect 29416 24568 29424 24632
rect 29104 23544 29424 24568
rect 29104 23480 29112 23544
rect 29176 23480 29192 23544
rect 29256 23480 29272 23544
rect 29336 23480 29352 23544
rect 29416 23480 29424 23544
rect 29104 22456 29424 23480
rect 29104 22392 29112 22456
rect 29176 22392 29192 22456
rect 29256 22392 29272 22456
rect 29336 22392 29352 22456
rect 29416 22392 29424 22456
rect 29104 21368 29424 22392
rect 29104 21304 29112 21368
rect 29176 21304 29192 21368
rect 29256 21304 29272 21368
rect 29336 21304 29352 21368
rect 29416 21304 29424 21368
rect 29104 20280 29424 21304
rect 29104 20216 29112 20280
rect 29176 20216 29192 20280
rect 29256 20216 29272 20280
rect 29336 20216 29352 20280
rect 29416 20216 29424 20280
rect 29104 19192 29424 20216
rect 29104 19128 29112 19192
rect 29176 19128 29192 19192
rect 29256 19128 29272 19192
rect 29336 19128 29352 19192
rect 29416 19128 29424 19192
rect 29104 18104 29424 19128
rect 29104 18040 29112 18104
rect 29176 18040 29192 18104
rect 29256 18040 29272 18104
rect 29336 18040 29352 18104
rect 29416 18040 29424 18104
rect 29104 17016 29424 18040
rect 29104 16952 29112 17016
rect 29176 16952 29192 17016
rect 29256 16952 29272 17016
rect 29336 16952 29352 17016
rect 29416 16952 29424 17016
rect 29104 15928 29424 16952
rect 29104 15864 29112 15928
rect 29176 15864 29192 15928
rect 29256 15864 29272 15928
rect 29336 15864 29352 15928
rect 29416 15864 29424 15928
rect 29104 14840 29424 15864
rect 29104 14776 29112 14840
rect 29176 14776 29192 14840
rect 29256 14776 29272 14840
rect 29336 14776 29352 14840
rect 29416 14776 29424 14840
rect 29104 13752 29424 14776
rect 29104 13688 29112 13752
rect 29176 13688 29192 13752
rect 29256 13688 29272 13752
rect 29336 13688 29352 13752
rect 29416 13688 29424 13752
rect 29104 12664 29424 13688
rect 29104 12600 29112 12664
rect 29176 12600 29192 12664
rect 29256 12600 29272 12664
rect 29336 12600 29352 12664
rect 29416 12600 29424 12664
rect 29104 11576 29424 12600
rect 29104 11512 29112 11576
rect 29176 11512 29192 11576
rect 29256 11512 29272 11576
rect 29336 11512 29352 11576
rect 29416 11512 29424 11576
rect 29104 3992 29424 11512
rect 32136 36032 36136 36040
rect 32136 32048 32144 36032
rect 36128 32048 36136 36032
rect 32136 8992 36136 32048
rect 32136 5008 32144 8992
rect 36128 5008 36136 8992
rect 32136 5000 36136 5008
rect 29104 8 29112 3992
rect 29416 8 29424 3992
rect 29104 0 29424 8
rect 37136 3992 41136 37048
rect 37136 8 37144 3992
rect 41128 8 41136 3992
rect 37136 0 41136 8
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[3\].id.delaybuf1
timestamp 1606789161
transform 1 0 29032 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[3\].id.delayint0
timestamp 1606789161
transform 1 0 28940 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_67
timestamp 1606789161
transform -1 0 30136 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_69
timestamp 1606789161
transform -1 0 30136 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_199
timestamp 1606789161
transform 1 0 29308 0 1 28952
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_34_198
timestamp 1606789161
transform 1 0 29216 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_34_204
timestamp 1606789161
transform 1 0 29768 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_33_184
timestamp 1606789161
transform 1 0 27928 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_168
timestamp 1606789161
transform 1 0 26456 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_174
timestamp 1606789161
transform 1 0 27836 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_180
timestamp 1606789161
transform 1 0 28112 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_182
timestamp 1606789161
transform 1 0 27744 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_180
timestamp 1606789161
transform 1 0 27560 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_34_187
timestamp 1606789161
transform 1 0 28204 0 -1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[4\].id.delayint0
timestamp 1606789161
transform 1 0 27100 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_33_168
timestamp 1606789161
transform 1 0 26456 0 1 28952
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_33_174
timestamp 1606789161
transform 1 0 27008 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_178
timestamp 1606789161
transform 1 0 27376 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[5\].id.delaybuf1
timestamp 1606789161
transform 1 0 26180 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[5\].id.delayenb1
timestamp 1606789161
transform 1 0 25444 0 1 28952
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_179
timestamp 1606789161
transform 1 0 25260 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_34_156
timestamp 1606789161
transform 1 0 25352 0 -1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_164
timestamp 1606789161
transform 1 0 26088 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[5\].id.delayint0
timestamp 1606789161
transform 1 0 24800 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_145
timestamp 1606789161
transform 1 0 24340 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_33_149
timestamp 1606789161
transform 1 0 24708 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_153
timestamp 1606789161
transform 1 0 25076 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_2  FILLER_34_153
timestamp 1606789161
transform 1 0 25076 0 -1 30040
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_34_129
timestamp 1606789161
transform 1 0 22868 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_141
timestamp 1606789161
transform 1 0 23972 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[6\].id.delaybuf1
timestamp 1606789161
transform 1 0 24064 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_138
timestamp 1606789161
transform 1 0 23696 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[6\].id.delayenb1
timestamp 1606789161
transform 1 0 22684 0 1 28952
box -38 -48 1050 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[6\].id.delayint0
timestamp 1606789161
transform 1 0 22592 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_173
timestamp 1606789161
transform 1 0 22224 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_178
timestamp 1606789161
transform 1 0 22408 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_33_121
timestamp 1606789161
transform 1 0 22132 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_123
timestamp 1606789161
transform 1 0 22316 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_123
timestamp 1606789161
transform 1 0 22316 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_34_125
timestamp 1606789161
transform 1 0 22500 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__a21bo_4  _439_
timestamp 1606789161
transform 1 0 20568 0 1 28952
box -38 -48 1234 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen0
timestamp 1606789161
transform 1 0 21120 0 -1 30040
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[7\].id.delaybuf0
timestamp 1606789161
transform 1 0 20292 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_100
timestamp 1606789161
transform 1 0 20200 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_33_117
timestamp 1606789161
transform 1 0 21764 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_97
timestamp 1606789161
transform 1 0 19924 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_105
timestamp 1606789161
transform 1 0 20660 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_34_109
timestamp 1606789161
transform 1 0 21028 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_34_117
timestamp 1606789161
transform 1 0 21764 0 -1 30040
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[7\].id.delaybuf1
timestamp 1606789161
transform 1 0 19648 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen1
timestamp 1606789161
transform 1 0 19556 0 1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[7\].id.delayint0
timestamp 1606789161
transform 1 0 18912 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_177
timestamp 1606789161
transform 1 0 19556 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_89
timestamp 1606789161
transform 1 0 19188 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_75
timestamp 1606789161
transform 1 0 17900 0 -1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_83
timestamp 1606789161
transform 1 0 18636 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_34_89
timestamp 1606789161
transform 1 0 19188 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[7\].id.delayenb0
timestamp 1606789161
transform 1 0 17532 0 1 28952
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_12  FILLER_34_63
timestamp 1606789161
transform 1 0 16796 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_172
timestamp 1606789161
transform 1 0 16612 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_176
timestamp 1606789161
transform 1 0 16704 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_33_62
timestamp 1606789161
transform 1 0 16704 0 1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_33_70
timestamp 1606789161
transform 1 0 17440 0 1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[8\].id.delayint0
timestamp 1606789161
transform 1 0 15416 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_33_57
timestamp 1606789161
transform 1 0 16244 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_51
timestamp 1606789161
transform 1 0 15692 0 -1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_34_59
timestamp 1606789161
transform 1 0 16428 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _449_
timestamp 1606789161
transform 1 0 15048 0 1 28952
box -38 -48 1234 592
use sky130_fd_sc_hd__a21bo_4  _511_
timestamp 1606789161
transform 1 0 13484 0 1 28952
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[8\].id.delaybuf1
timestamp 1606789161
transform 1 0 14772 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_175
timestamp 1606789161
transform 1 0 13852 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_33_40
timestamp 1606789161
transform 1 0 14680 0 1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_34_27
timestamp 1606789161
transform 1 0 13484 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_34_32
timestamp 1606789161
transform 1 0 13944 0 -1 30040
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_34_40
timestamp 1606789161
transform 1 0 14680 0 -1 30040
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_34_44
timestamp 1606789161
transform 1 0 15048 0 -1 30040
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_66
timestamp 1606789161
transform 1 0 11000 0 1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_68
timestamp 1606789161
transform 1 0 11000 0 -1 30040
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_33_3
timestamp 1606789161
transform 1 0 11276 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_33_15
timestamp 1606789161
transform 1 0 12380 0 1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_3
timestamp 1606789161
transform 1 0 11276 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_34_15
timestamp 1606789161
transform 1 0 12380 0 -1 30040
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _281_
timestamp 1606789161
transform 1 0 29124 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_65
timestamp 1606789161
transform -1 0 30136 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_32_196
timestamp 1606789161
transform 1 0 29032 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_200
timestamp 1606789161
transform 1 0 29400 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_204
timestamp 1606789161
transform 1 0 29768 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _545_
timestamp 1606789161
transform 1 0 27928 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen1
timestamp 1606789161
transform 1 0 26916 0 -1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_32_169
timestamp 1606789161
transform 1 0 26548 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_180
timestamp 1606789161
transform 1 0 27560 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_32_188
timestamp 1606789161
transform 1 0 28296 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__a21bo_4  _500_
timestamp 1606789161
transform 1 0 25352 0 -1 28952
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[6\].id.delaybuf0
timestamp 1606789161
transform 1 0 24248 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_171
timestamp 1606789161
transform 1 0 25076 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_148
timestamp 1606789161
transform 1 0 24616 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_32_152
timestamp 1606789161
transform 1 0 24984 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_32_154
timestamp 1606789161
transform 1 0 25168 0 -1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__a21bo_4  _503_
timestamp 1606789161
transform 1 0 22684 0 -1 28952
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_32_123
timestamp 1606789161
transform 1 0 22316 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_32_140
timestamp 1606789161
transform 1 0 23880 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[6\].id.delayenb0
timestamp 1606789161
transform 1 0 20660 0 -1 28952
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_32_101
timestamp 1606789161
transform 1 0 20292 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _428_
timestamp 1606789161
transform 1 0 19648 0 -1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[7\].id.delayen0
timestamp 1606789161
transform 1 0 17900 0 -1 28952
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_170
timestamp 1606789161
transform 1 0 19464 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_74
timestamp 1606789161
transform 1 0 17808 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_32_82
timestamp 1606789161
transform 1 0 18544 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_32_90
timestamp 1606789161
transform 1 0 19280 0 -1 28952
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_32_93
timestamp 1606789161
transform 1 0 19556 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[8\].id.delayenb0
timestamp 1606789161
transform 1 0 15416 0 -1 28952
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_8  FILLER_32_66
timestamp 1606789161
transform 1 0 17072 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[8\].id.delayenb1
timestamp 1606789161
transform 1 0 14036 0 -1 28952
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_169
timestamp 1606789161
transform 1 0 13852 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_30
timestamp 1606789161
transform 1 0 13760 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_32_32
timestamp 1606789161
transform 1 0 13944 0 -1 28952
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_32_44
timestamp 1606789161
transform 1 0 15048 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _280_
timestamp 1606789161
transform 1 0 11644 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_64
timestamp 1606789161
transform 1 0 11000 0 -1 28952
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_32_3
timestamp 1606789161
transform 1 0 11276 0 -1 28952
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_32_10
timestamp 1606789161
transform 1 0 11920 0 -1 28952
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_32_22
timestamp 1606789161
transform 1 0 13024 0 -1 28952
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[9\].id.delaybuf0
timestamp 1606789161
transform 1 0 28664 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_63
timestamp 1606789161
transform -1 0 30136 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_31_196
timestamp 1606789161
transform 1 0 29032 0 1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_31_204
timestamp 1606789161
transform 1 0 29768 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[5\].id.delaybuf0
timestamp 1606789161
transform 1 0 27928 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[5\].id.delayen0
timestamp 1606789161
transform 1 0 26456 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_168
timestamp 1606789161
transform 1 0 27836 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_175
timestamp 1606789161
transform 1 0 27100 0 1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_31_188
timestamp 1606789161
transform 1 0 28296 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[5\].id.delayenb0
timestamp 1606789161
transform 1 0 24432 0 1 27864
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_31_164
timestamp 1606789161
transform 1 0 26088 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[6\].id.delayen1
timestamp 1606789161
transform 1 0 22776 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_167
timestamp 1606789161
transform 1 0 22224 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_31_123
timestamp 1606789161
transform 1 0 22316 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_31_127
timestamp 1606789161
transform 1 0 22684 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_31_135
timestamp 1606789161
transform 1 0 23420 0 1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_143
timestamp 1606789161
transform 1 0 24156 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _427_
timestamp 1606789161
transform 1 0 20568 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_31_100
timestamp 1606789161
transform 1 0 20200 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_31_111
timestamp 1606789161
transform 1 0 21212 0 1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_31_119
timestamp 1606789161
transform 1 0 21948 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__a21bo_4  _435_
timestamp 1606789161
transform 1 0 17624 0 1 27864
box -38 -48 1234 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[7\].id.delayenb1
timestamp 1606789161
transform 1 0 19188 0 1 27864
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_31_85
timestamp 1606789161
transform 1 0 18820 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[8\].id.delaybuf0
timestamp 1606789161
transform 1 0 16888 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen0
timestamp 1606789161
transform 1 0 15416 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_166
timestamp 1606789161
transform 1 0 16612 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_55
timestamp 1606789161
transform 1 0 16060 0 1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_2  FILLER_31_62
timestamp 1606789161
transform 1 0 16704 0 1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_31_68
timestamp 1606789161
transform 1 0 17256 0 1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[8\].id.delayen1
timestamp 1606789161
transform 1 0 14128 0 1 27864
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_31_27
timestamp 1606789161
transform 1 0 13484 0 1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_33
timestamp 1606789161
transform 1 0 14036 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_31_41
timestamp 1606789161
transform 1 0 14772 0 1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_31_47
timestamp 1606789161
transform 1 0 15324 0 1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_62
timestamp 1606789161
transform 1 0 11000 0 1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_31_3
timestamp 1606789161
transform 1 0 11276 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_31_15
timestamp 1606789161
transform 1 0 12380 0 1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_61
timestamp 1606789161
transform -1 0 30136 0 -1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_201
timestamp 1606789161
transform 1 0 29492 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[3\].id.delayenb0
timestamp 1606789161
transform 1 0 27836 0 -1 27864
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_30_179
timestamp 1606789161
transform 1 0 27468 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[4\].id.delaybuf1
timestamp 1606789161
transform 1 0 25168 0 -1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[4\].id.delayenb0
timestamp 1606789161
transform 1 0 25812 0 -1 27864
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_165
timestamp 1606789161
transform 1 0 25076 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_30_146
timestamp 1606789161
transform 1 0 24432 0 -1 27864
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_30_152
timestamp 1606789161
transform 1 0 24984 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_157
timestamp 1606789161
transform 1 0 25444 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _453_
timestamp 1606789161
transform 1 0 23236 0 -1 27864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_30_129
timestamp 1606789161
transform 1 0 22868 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _404_
timestamp 1606789161
transform 1 0 21672 0 -1 27864
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_30_102
timestamp 1606789161
transform 1 0 20384 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_30_114
timestamp 1606789161
transform 1 0 21488 0 -1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__and4_4  _425_
timestamp 1606789161
transform 1 0 19556 0 -1 27864
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_164
timestamp 1606789161
transform 1 0 19464 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_30_82
timestamp 1606789161
transform 1 0 18544 0 -1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_90
timestamp 1606789161
transform 1 0 19280 0 -1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__o22a_4  _447_
timestamp 1606789161
transform 1 0 17256 0 -1 27864
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _448_
timestamp 1606789161
transform 1 0 16612 0 -1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_30_56
timestamp 1606789161
transform 1 0 16152 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_30_60
timestamp 1606789161
transform 1 0 16520 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_30_64
timestamp 1606789161
transform 1 0 16888 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _531_
timestamp 1606789161
transform 1 0 14680 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_163
timestamp 1606789161
transform 1 0 13852 0 -1 27864
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_30_29
timestamp 1606789161
transform 1 0 13668 0 -1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_30_32
timestamp 1606789161
transform 1 0 13944 0 -1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_30_44
timestamp 1606789161
transform 1 0 15048 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _530_
timestamp 1606789161
transform 1 0 12196 0 -1 27864
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_60
timestamp 1606789161
transform 1 0 11000 0 -1 27864
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_30_3
timestamp 1606789161
transform 1 0 11276 0 -1 27864
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_30_11
timestamp 1606789161
transform 1 0 12012 0 -1 27864
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_30_17
timestamp 1606789161
transform 1 0 12564 0 -1 27864
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_59
timestamp 1606789161
transform -1 0 30136 0 1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_196
timestamp 1606789161
transform 1 0 29032 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_29_204
timestamp 1606789161
transform 1 0 29768 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen0
timestamp 1606789161
transform 1 0 28388 0 1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen0
timestamp 1606789161
transform 1 0 26640 0 1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_162
timestamp 1606789161
transform 1 0 27836 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_29_169
timestamp 1606789161
transform 1 0 26548 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_29_177
timestamp 1606789161
transform 1 0 27284 0 1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_29_184
timestamp 1606789161
transform 1 0 27928 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_188
timestamp 1606789161
transform 1 0 28296 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _497_
timestamp 1606789161
transform 1 0 25536 0 1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_29_150
timestamp 1606789161
transform 1 0 24800 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_8  FILLER_29_161
timestamp 1606789161
transform 1 0 25812 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _419_
timestamp 1606789161
transform 1 0 22500 0 1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_4  _438_
timestamp 1606789161
transform 1 0 23604 0 1 26776
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_161
timestamp 1606789161
transform 1 0 22224 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_29_120
timestamp 1606789161
transform 1 0 22040 0 1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_29_123
timestamp 1606789161
transform 1 0 22316 0 1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_29_132
timestamp 1606789161
transform 1 0 23144 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_29_136
timestamp 1606789161
transform 1 0 23512 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _411_
timestamp 1606789161
transform 1 0 20108 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_29_108
timestamp 1606789161
transform 1 0 20936 0 1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _426_
timestamp 1606789161
transform 1 0 18912 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _434_
timestamp 1606789161
transform 1 0 17900 0 1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_29_82
timestamp 1606789161
transform 1 0 18544 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_29_95
timestamp 1606789161
transform 1 0 19740 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _433_
timestamp 1606789161
transform 1 0 16704 0 1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_160
timestamp 1606789161
transform 1 0 16612 0 1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_29_53
timestamp 1606789161
transform 1 0 15876 0 1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_29_71
timestamp 1606789161
transform 1 0 17532 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _558_
timestamp 1606789161
transform 1 0 13760 0 1 26776
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_29_26
timestamp 1606789161
transform 1 0 13392 0 1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _559_
timestamp 1606789161
transform 1 0 11276 0 1 26776
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_58
timestamp 1606789161
transform 1 0 11000 0 1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _284_
timestamp 1606789161
transform 1 0 29124 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_57
timestamp 1606789161
transform -1 0 30136 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_28_193
timestamp 1606789161
transform 1 0 28756 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_200
timestamp 1606789161
transform 1 0 29400 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_28_204
timestamp 1606789161
transform 1 0 29768 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[4\].id.delaybuf0
timestamp 1606789161
transform 1 0 28388 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[4\].id.delayenb1
timestamp 1606789161
transform 1 0 27008 0 -1 26776
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_4  FILLER_28_170
timestamp 1606789161
transform 1 0 26640 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_28_185
timestamp 1606789161
transform 1 0 28020 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _437_
timestamp 1606789161
transform 1 0 25168 0 -1 26776
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_159
timestamp 1606789161
transform 1 0 25076 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_28_145
timestamp 1606789161
transform 1 0 24340 0 -1 26776
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _418_
timestamp 1606789161
transform 1 0 22500 0 -1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _420_
timestamp 1606789161
transform 1 0 23696 0 -1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_28_121
timestamp 1606789161
transform 1 0 22132 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_28_132
timestamp 1606789161
transform 1 0 23144 0 -1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__and4_4  _410_
timestamp 1606789161
transform 1 0 20108 0 -1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _412_
timestamp 1606789161
transform 1 0 21488 0 -1 26776
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_28_108
timestamp 1606789161
transform 1 0 20936 0 -1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_158
timestamp 1606789161
transform 1 0 19464 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_28_79
timestamp 1606789161
transform 1 0 18268 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_28_91
timestamp 1606789161
transform 1 0 19372 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_28_93
timestamp 1606789161
transform 1 0 19556 0 -1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _270_
timestamp 1606789161
transform 1 0 15876 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _409_
timestamp 1606789161
transform 1 0 17440 0 -1 26776
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_28_49
timestamp 1606789161
transform 1 0 15508 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_56
timestamp 1606789161
transform 1 0 16152 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_68
timestamp 1606789161
transform 1 0 17256 0 -1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _271_
timestamp 1606789161
transform 1 0 15232 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_157
timestamp 1606789161
transform 1 0 13852 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_28_27
timestamp 1606789161
transform 1 0 13484 0 -1 26776
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_28_32
timestamp 1606789161
transform 1 0 13944 0 -1 26776
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_28_44
timestamp 1606789161
transform 1 0 15048 0 -1 26776
box -38 -48 222 592
use sky130_fd_sc_hd__a32o_4  _373_
timestamp 1606789161
transform 1 0 11920 0 -1 26776
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_56
timestamp 1606789161
transform 1 0 11000 0 -1 26776
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_28_3
timestamp 1606789161
transform 1 0 11276 0 -1 26776
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_28_9
timestamp 1606789161
transform 1 0 11828 0 -1 26776
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_53
timestamp 1606789161
transform -1 0 30136 0 -1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_55
timestamp 1606789161
transform -1 0 30136 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_199
timestamp 1606789161
transform 1 0 29308 0 -1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_27_196
timestamp 1606789161
transform 1 0 29032 0 1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_204
timestamp 1606789161
transform 1 0 29768 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _487_
timestamp 1606789161
transform 1 0 26548 0 -1 25688
box -38 -48 1326 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[3\].id.delayen1
timestamp 1606789161
transform 1 0 28388 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[3\].id.delayenb1
timestamp 1606789161
transform 1 0 28296 0 -1 25688
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_156
timestamp 1606789161
transform 1 0 27836 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_183
timestamp 1606789161
transform 1 0 27836 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_187
timestamp 1606789161
transform 1 0 28204 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_184
timestamp 1606789161
transform 1 0 27928 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_188
timestamp 1606789161
transform 1 0 28296 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[4\].id.delayen1
timestamp 1606789161
transform 1 0 26456 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_27_175
timestamp 1606789161
transform 1 0 27100 0 1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _496_
timestamp 1606789161
transform 1 0 24616 0 1 25688
box -38 -48 1326 592
use sky130_fd_sc_hd__or4_4  _499_
timestamp 1606789161
transform 1 0 25168 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_153
timestamp 1606789161
transform 1 0 25076 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_148
timestamp 1606789161
transform 1 0 24616 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_152
timestamp 1606789161
transform 1 0 24984 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_26_163
timestamp 1606789161
transform 1 0 25996 0 -1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_147
timestamp 1606789161
transform 1 0 24524 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_162
timestamp 1606789161
transform 1 0 25904 0 1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _423_
timestamp 1606789161
transform 1 0 23144 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _424_
timestamp 1606789161
transform 1 0 22316 0 -1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _495_
timestamp 1606789161
transform 1 0 23788 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_155
timestamp 1606789161
transform 1 0 22224 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_26_130
timestamp 1606789161
transform 1 0 22960 0 -1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_138
timestamp 1606789161
transform 1 0 23696 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_123
timestamp 1606789161
transform 1 0 22316 0 1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_27_131
timestamp 1606789161
transform 1 0 23052 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_27_139
timestamp 1606789161
transform 1 0 23788 0 1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _417_
timestamp 1606789161
transform 1 0 21304 0 -1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _464_
timestamp 1606789161
transform 1 0 21212 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _489_
timestamp 1606789161
transform 1 0 20108 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_26_103
timestamp 1606789161
transform 1 0 20476 0 -1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_26_111
timestamp 1606789161
transform 1 0 21212 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_119
timestamp 1606789161
transform 1 0 21948 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_106
timestamp 1606789161
transform 1 0 20752 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_27_110
timestamp 1606789161
transform 1 0 21120 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_118
timestamp 1606789161
transform 1 0 21856 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _493_
timestamp 1606789161
transform 1 0 19648 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_152
timestamp 1606789161
transform 1 0 19464 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_26_93
timestamp 1606789161
transform 1 0 19556 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_95
timestamp 1606789161
transform 1 0 19740 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _444_
timestamp 1606789161
transform 1 0 19096 0 1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_26_87
timestamp 1606789161
transform 1 0 19004 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_91
timestamp 1606789161
transform 1 0 19372 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_84
timestamp 1606789161
transform 1 0 18728 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _446_
timestamp 1606789161
transform 1 0 18176 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _462_
timestamp 1606789161
transform 1 0 17900 0 1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_26_74
timestamp 1606789161
transform 1 0 17808 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_71
timestamp 1606789161
transform 1 0 17532 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _445_
timestamp 1606789161
transform 1 0 16980 0 -1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _461_
timestamp 1606789161
transform 1 0 16704 0 1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_154
timestamp 1606789161
transform 1 0 16612 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_26_63
timestamp 1606789161
transform 1 0 16796 0 -1 25688
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_27_60
timestamp 1606789161
transform 1 0 16520 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _349_
timestamp 1606789161
transform 1 0 15876 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _374_
timestamp 1606789161
transform 1 0 15416 0 -1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_26_55
timestamp 1606789161
transform 1 0 16060 0 -1 25688
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_27_49
timestamp 1606789161
transform 1 0 15508 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_27_56
timestamp 1606789161
transform 1 0 16152 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _370_
timestamp 1606789161
transform 1 0 13944 0 -1 25688
box -38 -48 1142 592
use sky130_fd_sc_hd__a32o_4  _375_
timestamp 1606789161
transform 1 0 13944 0 1 25688
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_151
timestamp 1606789161
transform 1 0 13852 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_26
timestamp 1606789161
transform 1 0 13392 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_30
timestamp 1606789161
transform 1 0 13760 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_26_44
timestamp 1606789161
transform 1 0 15048 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_27_25
timestamp 1606789161
transform 1 0 13300 0 1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_27_31
timestamp 1606789161
transform 1 0 13852 0 1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _371_
timestamp 1606789161
transform 1 0 12472 0 1 25688
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _372_
timestamp 1606789161
transform 1 0 12748 0 -1 25688
box -38 -48 682 592
use sky130_fd_sc_hd__buf_2  _529_
timestamp 1606789161
transform 1 0 11920 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_26_14
timestamp 1606789161
transform 1 0 12288 0 -1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_26_18
timestamp 1606789161
transform 1 0 12656 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_27_10
timestamp 1606789161
transform 1 0 11920 0 1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _285_
timestamp 1606789161
transform 1 0 11644 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_52
timestamp 1606789161
transform 1 0 11000 0 -1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_54
timestamp 1606789161
transform 1 0 11000 0 1 25688
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_26_3
timestamp 1606789161
transform 1 0 11276 0 -1 25688
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_26_9
timestamp 1606789161
transform 1 0 11828 0 -1 25688
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_27_3
timestamp 1606789161
transform 1 0 11276 0 1 25688
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen1
timestamp 1606789161
transform 1 0 28572 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_51
timestamp 1606789161
transform -1 0 30136 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_25_198
timestamp 1606789161
transform 1 0 29216 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_204
timestamp 1606789161
transform 1 0 29768 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _488_
timestamp 1606789161
transform 1 0 27928 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[1\].id.delayint0
timestamp 1606789161
transform 1 0 26916 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_150
timestamp 1606789161
transform 1 0 27836 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_169
timestamp 1606789161
transform 1 0 26548 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_176
timestamp 1606789161
transform 1 0 27192 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_25_182
timestamp 1606789161
transform 1 0 27744 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_187
timestamp 1606789161
transform 1 0 28204 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _429_
timestamp 1606789161
transform 1 0 24892 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _450_
timestamp 1606789161
transform 1 0 25904 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_25_147
timestamp 1606789161
transform 1 0 24524 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_25_158
timestamp 1606789161
transform 1 0 25536 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _486_
timestamp 1606789161
transform 1 0 23696 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _498_
timestamp 1606789161
transform 1 0 22316 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_149
timestamp 1606789161
transform 1 0 22224 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_121
timestamp 1606789161
transform 1 0 22132 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_25_132
timestamp 1606789161
transform 1 0 23144 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__or4_4  _494_
timestamp 1606789161
transform 1 0 20568 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_25_100
timestamp 1606789161
transform 1 0 20200 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_25_113
timestamp 1606789161
transform 1 0 21396 0 1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _442_
timestamp 1606789161
transform 1 0 18176 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _490_
timestamp 1606789161
transform 1 0 19372 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_25_77
timestamp 1606789161
transform 1 0 18084 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_87
timestamp 1606789161
transform 1 0 19004 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _415_
timestamp 1606789161
transform 1 0 16704 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _501_
timestamp 1606789161
transform 1 0 15600 0 1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_148
timestamp 1606789161
transform 1 0 16612 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_25_49
timestamp 1606789161
transform 1 0 15508 0 1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_25_57
timestamp 1606789161
transform 1 0 16244 0 1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_25_71
timestamp 1606789161
transform 1 0 17532 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__nand2_4  _369_
timestamp 1606789161
transform 1 0 13944 0 1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_25_26
timestamp 1606789161
transform 1 0 13392 0 1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_25_41
timestamp 1606789161
transform 1 0 14772 0 1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _560_
timestamp 1606789161
transform 1 0 11276 0 1 24600
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_50
timestamp 1606789161
transform 1 0 11000 0 1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[3\].id.delaybuf0
timestamp 1606789161
transform 1 0 29124 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_49
timestamp 1606789161
transform -1 0 30136 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_24_193
timestamp 1606789161
transform 1 0 28756 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_201
timestamp 1606789161
transform 1 0 29492 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _451_
timestamp 1606789161
transform 1 0 27468 0 -1 24600
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_24_175
timestamp 1606789161
transform 1 0 27100 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _421_
timestamp 1606789161
transform 1 0 25812 0 -1 24600
box -38 -48 1326 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[9\].id.delaybuf1
timestamp 1606789161
transform 1 0 25168 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[9\].id.delayint0
timestamp 1606789161
transform 1 0 24432 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_147
timestamp 1606789161
transform 1 0 25076 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_145
timestamp 1606789161
transform 1 0 24340 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_24_149
timestamp 1606789161
transform 1 0 24708 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_157
timestamp 1606789161
transform 1 0 25444 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _521_
timestamp 1606789161
transform 1 0 23144 0 -1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_24_130
timestamp 1606789161
transform 1 0 22960 0 -1 24600
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_24_141
timestamp 1606789161
transform 1 0 23972 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _441_
timestamp 1606789161
transform 1 0 21212 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _484_
timestamp 1606789161
transform 1 0 20200 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_24_96
timestamp 1606789161
transform 1 0 19832 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_107
timestamp 1606789161
transform 1 0 20844 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_24_118
timestamp 1606789161
transform 1 0 21856 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _408_
timestamp 1606789161
transform 1 0 19556 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _520_
timestamp 1606789161
transform 1 0 18268 0 -1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_146
timestamp 1606789161
transform 1 0 19464 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_24_73
timestamp 1606789161
transform 1 0 17716 0 -1 24600
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_24_88
timestamp 1606789161
transform 1 0 19096 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _463_
timestamp 1606789161
transform 1 0 17072 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _491_
timestamp 1606789161
transform 1 0 15784 0 -1 24600
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_24_48
timestamp 1606789161
transform 1 0 15416 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_24_61
timestamp 1606789161
transform 1 0 16612 0 -1 24600
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_24_65
timestamp 1606789161
transform 1 0 16980 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _269_
timestamp 1606789161
transform 1 0 13944 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _492_
timestamp 1606789161
transform 1 0 15140 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_145
timestamp 1606789161
transform 1 0 13852 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_24_30
timestamp 1606789161
transform 1 0 13760 0 -1 24600
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_24_35
timestamp 1606789161
transform 1 0 14220 0 -1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_24_43
timestamp 1606789161
transform 1 0 14956 0 -1 24600
box -38 -48 222 592
use sky130_fd_sc_hd__or2_4  _366_
timestamp 1606789161
transform 1 0 12012 0 -1 24600
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_48
timestamp 1606789161
transform 1 0 11000 0 -1 24600
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_24_3
timestamp 1606789161
transform 1 0 11276 0 -1 24600
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_24_18
timestamp 1606789161
transform 1 0 12656 0 -1 24600
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _279_
timestamp 1606789161
transform 1 0 29124 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_47
timestamp 1606789161
transform -1 0 30136 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_23_191
timestamp 1606789161
transform 1 0 28572 0 1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_200
timestamp 1606789161
transform 1 0 29400 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_204
timestamp 1606789161
transform 1 0 29768 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _452_
timestamp 1606789161
transform 1 0 26916 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[9\].id.delayen0
timestamp 1606789161
transform 1 0 27928 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_144
timestamp 1606789161
transform 1 0 27836 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_167
timestamp 1606789161
transform 1 0 26364 0 1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_23_176
timestamp 1606789161
transform 1 0 27192 0 1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_23_182
timestamp 1606789161
transform 1 0 27744 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _422_
timestamp 1606789161
transform 1 0 26088 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__o21a_4  _436_
timestamp 1606789161
transform 1 0 24616 0 1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_23_147
timestamp 1606789161
transform 1 0 24524 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_160
timestamp 1606789161
transform 1 0 25720 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _460_
timestamp 1606789161
transform 1 0 22316 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__or2_4  _483_
timestamp 1606789161
transform 1 0 23328 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_143
timestamp 1606789161
transform 1 0 22224 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_23_130
timestamp 1606789161
transform 1 0 22960 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_23_141
timestamp 1606789161
transform 1 0 23972 0 1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _440_
timestamp 1606789161
transform 1 0 20016 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _510_
timestamp 1606789161
transform 1 0 21028 0 1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_23_105
timestamp 1606789161
transform 1 0 20660 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_118
timestamp 1606789161
transform 1 0 21856 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _443_
timestamp 1606789161
transform 1 0 18360 0 1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_23_75
timestamp 1606789161
transform 1 0 17900 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_23_79
timestamp 1606789161
transform 1 0 18268 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_23_87
timestamp 1606789161
transform 1 0 19004 0 1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_23_95
timestamp 1606789161
transform 1 0 19740 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _416_
timestamp 1606789161
transform 1 0 15968 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _478_
timestamp 1606789161
transform 1 0 17072 0 1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_142
timestamp 1606789161
transform 1 0 16612 0 1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_23_48
timestamp 1606789161
transform 1 0 15416 0 1 23512
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_23_57
timestamp 1606789161
transform 1 0 16244 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_23_62
timestamp 1606789161
transform 1 0 16704 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _361_
timestamp 1606789161
transform 1 0 14128 0 1 23512
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _363_
timestamp 1606789161
transform 1 0 13484 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_30
timestamp 1606789161
transform 1 0 13760 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _368_
timestamp 1606789161
transform 1 0 11552 0 1 23512
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_46
timestamp 1606789161
transform 1 0 11000 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_23_3
timestamp 1606789161
transform 1 0 11276 0 1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_23_23
timestamp 1606789161
transform 1 0 13116 0 1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_45
timestamp 1606789161
transform -1 0 30136 0 -1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_196
timestamp 1606789161
transform 1 0 29032 0 -1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_22_204
timestamp 1606789161
transform 1 0 29768 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[10\].id.delaybuf0
timestamp 1606789161
transform 1 0 26640 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[9\].id.delayenb0
timestamp 1606789161
transform 1 0 27376 0 -1 23512
box -38 -48 1694 592
use sky130_fd_sc_hd__fill_1  FILLER_22_169
timestamp 1606789161
transform 1 0 26548 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_174
timestamp 1606789161
transform 1 0 27008 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _504_
timestamp 1606789161
transform 1 0 25168 0 -1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_141
timestamp 1606789161
transform 1 0 25076 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_148
timestamp 1606789161
transform 1 0 24616 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_152
timestamp 1606789161
transform 1 0 24984 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_161
timestamp 1606789161
transform 1 0 25812 0 -1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _454_
timestamp 1606789161
transform 1 0 23972 0 -1 23512
box -38 -48 682 592
use sky130_fd_sc_hd__a211o_4  _516_
timestamp 1606789161
transform 1 0 22316 0 -1 23512
box -38 -48 1326 592
use sky130_fd_sc_hd__fill_2  FILLER_22_121
timestamp 1606789161
transform 1 0 22132 0 -1 23512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_22_137
timestamp 1606789161
transform 1 0 23604 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _509_
timestamp 1606789161
transform 1 0 20200 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_96
timestamp 1606789161
transform 1 0 19832 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_22_109
timestamp 1606789161
transform 1 0 21028 0 -1 23512
box -38 -48 1142 592
use sky130_fd_sc_hd__nor2_4  _414_
timestamp 1606789161
transform 1 0 17900 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__inv_2  _479_
timestamp 1606789161
transform 1 0 19556 0 -1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_140
timestamp 1606789161
transform 1 0 19464 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_22_74
timestamp 1606789161
transform 1 0 17808 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_22_84
timestamp 1606789161
transform 1 0 18728 0 -1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _335_
timestamp 1606789161
transform 1 0 17164 0 -1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _336_
timestamp 1606789161
transform 1 0 15968 0 -1 23512
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_22_49
timestamp 1606789161
transform 1 0 15508 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_22_53
timestamp 1606789161
transform 1 0 15876 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_63
timestamp 1606789161
transform 1 0 16796 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_22_70
timestamp 1606789161
transform 1 0 17440 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _364_
timestamp 1606789161
transform 1 0 13944 0 -1 23512
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_139
timestamp 1606789161
transform 1 0 13852 0 -1 23512
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_22_27
timestamp 1606789161
transform 1 0 13484 0 -1 23512
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _365_
timestamp 1606789161
transform 1 0 12196 0 -1 23512
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  PHY_44
timestamp 1606789161
transform 1 0 11000 0 -1 23512
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_22_3
timestamp 1606789161
transform 1 0 11276 0 -1 23512
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_22_11
timestamp 1606789161
transform 1 0 12012 0 -1 23512
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_43
timestamp 1606789161
transform -1 0 30136 0 1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_200
timestamp 1606789161
transform 1 0 29400 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_204
timestamp 1606789161
transform 1 0 29768 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen0
timestamp 1606789161
transform 1 0 26364 0 1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[9\].id.delayenb1
timestamp 1606789161
transform 1 0 28388 0 1 22424
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_138
timestamp 1606789161
transform 1 0 27836 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_174
timestamp 1606789161
transform 1 0 27008 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_21_182
timestamp 1606789161
transform 1 0 27744 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_21_184
timestamp 1606789161
transform 1 0 27928 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_21_188
timestamp 1606789161
transform 1 0 28296 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _430_
timestamp 1606789161
transform 1 0 25352 0 1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_21_152
timestamp 1606789161
transform 1 0 24984 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_21_163
timestamp 1606789161
transform 1 0 25996 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _455_
timestamp 1606789161
transform 1 0 23788 0 1 22424
box -38 -48 1234 592
use sky130_fd_sc_hd__or4_4  _517_
timestamp 1606789161
transform 1 0 22592 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_137
timestamp 1606789161
transform 1 0 22224 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_21_123
timestamp 1606789161
transform 1 0 22316 0 1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_21_135
timestamp 1606789161
transform 1 0 23420 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _480_
timestamp 1606789161
transform 1 0 20292 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_21_97
timestamp 1606789161
transform 1 0 19924 0 1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_21_110
timestamp 1606789161
transform 1 0 21120 0 1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__and4_4  _459_
timestamp 1606789161
transform 1 0 19096 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_21_80
timestamp 1606789161
transform 1 0 18360 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__o32a_4  _413_
timestamp 1606789161
transform 1 0 16704 0 1 22424
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_136
timestamp 1606789161
transform 1 0 16612 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_51
timestamp 1606789161
transform 1 0 15692 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_59
timestamp 1606789161
transform 1 0 16428 0 1 22424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _332_
timestamp 1606789161
transform 1 0 13852 0 1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _333_
timestamp 1606789161
transform 1 0 15048 0 1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_21_30
timestamp 1606789161
transform 1 0 13760 0 1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_21_34
timestamp 1606789161
transform 1 0 14128 0 1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_21_42
timestamp 1606789161
transform 1 0 14864 0 1 22424
box -38 -48 222 592
use sky130_fd_sc_hd__nand2_4  _367_
timestamp 1606789161
transform 1 0 11828 0 1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_42
timestamp 1606789161
transform 1 0 11000 0 1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_21_3
timestamp 1606789161
transform 1 0 11276 0 1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_21_18
timestamp 1606789161
transform 1 0 12656 0 1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[2\].id.delaybuf0
timestamp 1606789161
transform 1 0 28940 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_39
timestamp 1606789161
transform -1 0 30136 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_41
timestamp 1606789161
transform -1 0 30136 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_191
timestamp 1606789161
transform 1 0 28572 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_199
timestamp 1606789161
transform 1 0 29308 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_201
timestamp 1606789161
transform 1 0 29492 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _514_
timestamp 1606789161
transform 1 0 28296 0 -1 22424
box -38 -48 1234 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[1\].id.delaybuf0
timestamp 1606789161
transform 1 0 26916 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen1
timestamp 1606789161
transform 1 0 27928 0 1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_132
timestamp 1606789161
transform 1 0 27836 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_169
timestamp 1606789161
transform 1 0 26548 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_19_177
timestamp 1606789161
transform 1 0 27284 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_20_180
timestamp 1606789161
transform 1 0 27560 0 -1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[1\].id.delayenb0
timestamp 1606789161
transform 1 0 25904 0 -1 22424
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[1\].id.delayenb1
timestamp 1606789161
transform 1 0 25536 0 1 21336
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_2  FILLER_19_156
timestamp 1606789161
transform 1 0 25352 0 1 21336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_20_157
timestamp 1606789161
transform 1 0 25444 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_161
timestamp 1606789161
transform 1 0 25812 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _431_
timestamp 1606789161
transform 1 0 25168 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_135
timestamp 1606789161
transform 1 0 25076 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_19_148
timestamp 1606789161
transform 1 0 24616 0 1 21336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_20_148
timestamp 1606789161
transform 1 0 24616 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_152
timestamp 1606789161
transform 1 0 24984 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _502_
timestamp 1606789161
transform 1 0 23972 0 -1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__or4_4  _507_
timestamp 1606789161
transform 1 0 22592 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _513_
timestamp 1606789161
transform 1 0 22776 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _518_
timestamp 1606789161
transform 1 0 23788 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_131
timestamp 1606789161
transform 1 0 22224 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_123
timestamp 1606789161
transform 1 0 22316 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_19_135
timestamp 1606789161
transform 1 0 23420 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_124
timestamp 1606789161
transform 1 0 22408 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_137
timestamp 1606789161
transform 1 0 23604 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_118
timestamp 1606789161
transform 1 0 21856 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _465_
timestamp 1606789161
transform 1 0 21580 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__or4_4  _512_
timestamp 1606789161
transform 1 0 21028 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__decap_6  FILLER_20_108
timestamp 1606789161
transform 1 0 20936 0 -1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_20_114
timestamp 1606789161
transform 1 0 21488 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _356_
timestamp 1606789161
transform 1 0 20384 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _403_
timestamp 1606789161
transform 1 0 20292 0 -1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_19_98
timestamp 1606789161
transform 1 0 20016 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_19_105
timestamp 1606789161
transform 1 0 20660 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_96
timestamp 1606789161
transform 1 0 19832 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_20_100
timestamp 1606789161
transform 1 0 20200 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _358_
timestamp 1606789161
transform 1 0 19556 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_134
timestamp 1606789161
transform 1 0 19464 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _469_
timestamp 1606789161
transform 1 0 19188 0 1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__fill_1  FILLER_19_88
timestamp 1606789161
transform 1 0 19096 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_20_83
timestamp 1606789161
transform 1 0 18636 0 -1 22424
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_91
timestamp 1606789161
transform 1 0 19372 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _407_
timestamp 1606789161
transform 1 0 17716 0 1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _477_
timestamp 1606789161
transform 1 0 17808 0 -1 22424
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_19_80
timestamp 1606789161
transform 1 0 18360 0 1 21336
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_20_73
timestamp 1606789161
transform 1 0 17716 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_19_69
timestamp 1606789161
transform 1 0 17348 0 1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_20_69
timestamp 1606789161
transform 1 0 17348 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _357_
timestamp 1606789161
transform 1 0 16704 0 1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__and2_4  _359_
timestamp 1606789161
transform 1 0 16704 0 -1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_130
timestamp 1606789161
transform 1 0 16612 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_19_58
timestamp 1606789161
transform 1 0 16336 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_20_61
timestamp 1606789161
transform 1 0 16612 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _344_
timestamp 1606789161
transform 1 0 15416 0 -1 22424
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_19_50
timestamp 1606789161
transform 1 0 15600 0 1 21336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_6  FILLER_20_55
timestamp 1606789161
transform 1 0 16060 0 -1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__a32o_4  _360_
timestamp 1606789161
transform 1 0 14036 0 1 21336
box -38 -48 1602 592
use sky130_fd_sc_hd__o21a_4  _362_
timestamp 1606789161
transform 1 0 13944 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_133
timestamp 1606789161
transform 1 0 13852 0 -1 22424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_19_26
timestamp 1606789161
transform 1 0 13392 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_19_32
timestamp 1606789161
transform 1 0 13944 0 1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_20_25
timestamp 1606789161
transform 1 0 13300 0 -1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_20_44
timestamp 1606789161
transform 1 0 15048 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__a32o_4  _383_
timestamp 1606789161
transform 1 0 11828 0 1 21336
box -38 -48 1602 592
use sky130_fd_sc_hd__buf_2  _533_
timestamp 1606789161
transform 1 0 11828 0 -1 22424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_38
timestamp 1606789161
transform 1 0 11000 0 1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_40
timestamp 1606789161
transform 1 0 11000 0 -1 22424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_19_3
timestamp 1606789161
transform 1 0 11276 0 1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_20_3
timestamp 1606789161
transform 1 0 11276 0 -1 22424
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_20_13
timestamp 1606789161
transform 1 0 12196 0 -1 22424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_37
timestamp 1606789161
transform -1 0 30136 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_18_201
timestamp 1606789161
transform 1 0 29492 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[1\].id.delayen1
timestamp 1606789161
transform 1 0 26640 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[2\].id.delayenb0
timestamp 1606789161
transform 1 0 27836 0 -1 21336
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_6  FILLER_18_177
timestamp 1606789161
transform 1 0 27284 0 -1 21336
box -38 -48 590 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen0
timestamp 1606789161
transform 1 0 25628 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_129
timestamp 1606789161
transform 1 0 25076 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_149
timestamp 1606789161
transform 1 0 24708 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_18_154
timestamp 1606789161
transform 1 0 25168 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_158
timestamp 1606789161
transform 1 0 25536 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_166
timestamp 1606789161
transform 1 0 26272 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _508_
timestamp 1606789161
transform 1 0 23512 0 -1 21336
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_8  FILLER_18_125
timestamp 1606789161
transform 1 0 22500 0 -1 21336
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_18_133
timestamp 1606789161
transform 1 0 23236 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _475_
timestamp 1606789161
transform 1 0 21212 0 -1 21336
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_4  FILLER_18_107
timestamp 1606789161
transform 1 0 20844 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _470_
timestamp 1606789161
transform 1 0 19556 0 -1 21336
box -38 -48 1326 592
use sky130_fd_sc_hd__and4_4  _506_
timestamp 1606789161
transform 1 0 18268 0 -1 21336
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_128
timestamp 1606789161
transform 1 0 19464 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_74
timestamp 1606789161
transform 1 0 17808 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_78
timestamp 1606789161
transform 1 0 18176 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_88
timestamp 1606789161
transform 1 0 19096 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__o32a_4  _471_
timestamp 1606789161
transform 1 0 16152 0 -1 21336
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_18_52
timestamp 1606789161
transform 1 0 15784 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _273_
timestamp 1606789161
transform 1 0 14404 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _334_
timestamp 1606789161
transform 1 0 15140 0 -1 21336
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_127
timestamp 1606789161
transform 1 0 13852 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_26
timestamp 1606789161
transform 1 0 13392 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_30
timestamp 1606789161
transform 1 0 13760 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_32
timestamp 1606789161
transform 1 0 13944 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_36
timestamp 1606789161
transform 1 0 14312 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_18_40
timestamp 1606789161
transform 1 0 14680 0 -1 21336
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_18_44
timestamp 1606789161
transform 1 0 15048 0 -1 21336
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _556_
timestamp 1606789161
transform 1 0 11276 0 -1 21336
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_36
timestamp 1606789161
transform 1 0 11000 0 -1 21336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_35
timestamp 1606789161
transform -1 0 30136 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_195
timestamp 1606789161
transform 1 0 28940 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_203
timestamp 1606789161
transform 1 0 29676 0 1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[2\].id.delayenb1
timestamp 1606789161
transform 1 0 27928 0 1 20248
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_126
timestamp 1606789161
transform 1 0 27836 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_173
timestamp 1606789161
transform 1 0 26916 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_181
timestamp 1606789161
transform 1 0 27652 0 1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _476_
timestamp 1606789161
transform 1 0 24616 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[0\].id.delayenb0
timestamp 1606789161
transform 1 0 25260 0 1 20248
box -38 -48 1694 592
use sky130_fd_sc_hd__decap_4  FILLER_17_144
timestamp 1606789161
transform 1 0 24248 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_151
timestamp 1606789161
transform 1 0 24892 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _505_
timestamp 1606789161
transform 1 0 22316 0 1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[1\].id.delaybuf1
timestamp 1606789161
transform 1 0 23972 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_125
timestamp 1606789161
transform 1 0 22224 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_17_121
timestamp 1606789161
transform 1 0 22132 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_130
timestamp 1606789161
transform 1 0 22960 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_138
timestamp 1606789161
transform 1 0 23696 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__or4_4  _474_
timestamp 1606789161
transform 1 0 19924 0 1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__and2_4  _485_
timestamp 1606789161
transform 1 0 21120 0 1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_106
timestamp 1606789161
transform 1 0 20752 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_117
timestamp 1606789161
transform 1 0 21764 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _468_
timestamp 1606789161
transform 1 0 18912 0 1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__nor2_4  _472_
timestamp 1606789161
transform 1 0 17624 0 1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_4  FILLER_17_81
timestamp 1606789161
transform 1 0 18452 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_17_85
timestamp 1606789161
transform 1 0 18820 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_17_93
timestamp 1606789161
transform 1 0 19556 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_124
timestamp 1606789161
transform 1 0 16612 0 1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_17_50
timestamp 1606789161
transform 1 0 15600 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_17_58
timestamp 1606789161
transform 1 0 16336 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_17_62
timestamp 1606789161
transform 1 0 16704 0 1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_17_70
timestamp 1606789161
transform 1 0 17440 0 1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _354_
timestamp 1606789161
transform 1 0 15324 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _380_
timestamp 1606789161
transform 1 0 14312 0 1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_17_32
timestamp 1606789161
transform 1 0 13944 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_43
timestamp 1606789161
transform 1 0 14956 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _376_
timestamp 1606789161
transform 1 0 12656 0 1 20248
box -38 -48 1326 592
use sky130_fd_sc_hd__or2_4  _382_
timestamp 1606789161
transform 1 0 11644 0 1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_34
timestamp 1606789161
transform 1 0 11000 0 1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_17_3
timestamp 1606789161
transform 1 0 11276 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_17_14
timestamp 1606789161
transform 1 0 12288 0 1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[2\].id.delayen0
timestamp 1606789161
transform 1 0 28572 0 -1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1606789161
transform -1 0 30136 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_198
timestamp 1606789161
transform 1 0 29216 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_204
timestamp 1606789161
transform 1 0 29768 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _482_
timestamp 1606789161
transform 1 0 27100 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[0\].id.delaybuf1
timestamp 1606789161
transform 1 0 27744 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_16_168
timestamp 1606789161
transform 1 0 26456 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_174
timestamp 1606789161
transform 1 0 27008 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_16_178
timestamp 1606789161
transform 1 0 27376 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_16_185
timestamp 1606789161
transform 1 0 28020 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[0\].id.delayenb1
timestamp 1606789161
transform 1 0 25444 0 -1 20248
box -38 -48 1050 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_123
timestamp 1606789161
transform 1 0 25076 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_144
timestamp 1606789161
transform 1 0 24248 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_16_152
timestamp 1606789161
transform 1 0 24984 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_16_154
timestamp 1606789161
transform 1 0 25168 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _406_
timestamp 1606789161
transform 1 0 23972 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[0\].id.delayint0
timestamp 1606789161
transform 1 0 23328 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_16_124
timestamp 1606789161
transform 1 0 22408 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_16_132
timestamp 1606789161
transform 1 0 23144 0 -1 20248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_16_137
timestamp 1606789161
transform 1 0 23604 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__o22a_4  _481_
timestamp 1606789161
transform 1 0 21120 0 -1 20248
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_16_102
timestamp 1606789161
transform 1 0 20384 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__and4_4  _467_
timestamp 1606789161
transform 1 0 18176 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__and4_4  _473_
timestamp 1606789161
transform 1 0 19556 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_122
timestamp 1606789161
transform 1 0 19464 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_72
timestamp 1606789161
transform 1 0 17624 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_16_87
timestamp 1606789161
transform 1 0 19004 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_91
timestamp 1606789161
transform 1 0 19372 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _346_
timestamp 1606789161
transform 1 0 15784 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _355_
timestamp 1606789161
transform 1 0 16980 0 -1 20248
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  FILLER_16_49
timestamp 1606789161
transform 1 0 15508 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_61
timestamp 1606789161
transform 1 0 16612 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__nand2_4  _379_
timestamp 1606789161
transform 1 0 13944 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_121
timestamp 1606789161
transform 1 0 13852 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_16_24
timestamp 1606789161
transform 1 0 13208 0 -1 20248
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_16_30
timestamp 1606789161
transform 1 0 13760 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_41
timestamp 1606789161
transform 1 0 14772 0 -1 20248
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _282_
timestamp 1606789161
transform 1 0 11644 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _377_
timestamp 1606789161
transform 1 0 12380 0 -1 20248
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_32
timestamp 1606789161
transform 1 0 11000 0 -1 20248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_3
timestamp 1606789161
transform 1 0 11276 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_16_10
timestamp 1606789161
transform 1 0 11920 0 -1 20248
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_16_14
timestamp 1606789161
transform 1 0 12288 0 -1 20248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1606789161
transform -1 0 30136 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_15_201
timestamp 1606789161
transform 1 0 29492 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _432_
timestamp 1606789161
transform 1 0 28388 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[0\].id.delaybuf0
timestamp 1606789161
transform 1 0 26916 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_120
timestamp 1606789161
transform 1 0 27836 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_15_169
timestamp 1606789161
transform 1 0 26548 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_15_177
timestamp 1606789161
transform 1 0 27284 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_15_184
timestamp 1606789161
transform 1 0 27928 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_15_188
timestamp 1606789161
transform 1 0 28296 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _458_
timestamp 1606789161
transform 1 0 24984 0 1 19160
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_4  FILLER_15_148
timestamp 1606789161
transform 1 0 24616 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[10\].id.delayenb0
timestamp 1606789161
transform 1 0 22960 0 1 19160
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_119
timestamp 1606789161
transform 1 0 22224 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_15_120
timestamp 1606789161
transform 1 0 22040 0 1 19160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_15_123
timestamp 1606789161
transform 1 0 22316 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_129
timestamp 1606789161
transform 1 0 22868 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__or3_4  _405_
timestamp 1606789161
transform 1 0 20108 0 1 19160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_15_108
timestamp 1606789161
transform 1 0 20936 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _272_
timestamp 1606789161
transform 1 0 17716 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__and4_4  _466_
timestamp 1606789161
transform 1 0 18912 0 1 19160
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_15_76
timestamp 1606789161
transform 1 0 17992 0 1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_15_84
timestamp 1606789161
transform 1 0 18728 0 1 19160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_15_95
timestamp 1606789161
transform 1 0 19740 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _347_
timestamp 1606789161
transform 1 0 16704 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_118
timestamp 1606789161
transform 1 0 16612 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_15_54
timestamp 1606789161
transform 1 0 15968 0 1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_15_60
timestamp 1606789161
transform 1 0 16520 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_15_65
timestamp 1606789161
transform 1 0 16980 0 1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__o22a_4  _353_
timestamp 1606789161
transform 1 0 14680 0 1 19160
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_15_31
timestamp 1606789161
transform 1 0 13852 0 1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_15_39
timestamp 1606789161
transform 1 0 14588 0 1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__o21a_4  _378_
timestamp 1606789161
transform 1 0 12748 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1606789161
transform 1 0 11000 0 1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1606789161
transform 1 0 11276 0 1 19160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_15_15
timestamp 1606789161
transform 1 0 12380 0 1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[2\].id.delaybuf1
timestamp 1606789161
transform 1 0 29216 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[2\].id.delayint0
timestamp 1606789161
transform 1 0 28756 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1606789161
transform -1 0 30136 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1606789161
transform -1 0 30136 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_13_192
timestamp 1606789161
transform 1 0 28664 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_196
timestamp 1606789161
transform 1 0 29032 0 1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_13_204
timestamp 1606789161
transform 1 0 29768 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_194
timestamp 1606789161
transform 1 0 28848 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_201
timestamp 1606789161
transform 1 0 29492 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp01
timestamp 1606789161
transform 1 0 27652 0 -1 19160
box -38 -48 1234 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp00
timestamp 1606789161
transform 1 0 27928 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_114
timestamp 1606789161
transform 1 0 27836 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_179
timestamp 1606789161
transform 1 0 27468 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_188
timestamp 1606789161
transform 1 0 28296 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_14_180
timestamp 1606789161
transform 1 0 27560 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _278_
timestamp 1606789161
transform 1 0 27192 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_1  ringosc.iss.reseten0
timestamp 1606789161
transform 1 0 26548 0 -1 19160
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_13_171
timestamp 1606789161
transform 1 0 26732 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_175
timestamp 1606789161
transform 1 0 27100 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_14_174
timestamp 1606789161
transform 1 0 27008 0 -1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__conb_1  ringosc.iss.const1
timestamp 1606789161
transform 1 0 25628 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__or2_2  ringosc.iss.ctrlen0
timestamp 1606789161
transform 1 0 26272 0 1 18072
box -38 -48 498 592
use sky130_fd_sc_hd__decap_4  FILLER_13_162
timestamp 1606789161
transform 1 0 25904 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_165
timestamp 1606789161
transform 1 0 26180 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[0\].id.delayen1
timestamp 1606789161
transform 1 0 25536 0 -1 19160
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_117
timestamp 1606789161
transform 1 0 25076 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_13_153
timestamp 1606789161
transform 1 0 25076 0 1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_14_152
timestamp 1606789161
transform 1 0 24984 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_154
timestamp 1606789161
transform 1 0 25168 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[10\].id.delayint0
timestamp 1606789161
transform 1 0 24340 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[11\].id.delaybuf1
timestamp 1606789161
transform 1 0 24800 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_13_146
timestamp 1606789161
transform 1 0 24432 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_148
timestamp 1606789161
transform 1 0 24616 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_2  ringosc.dstage\[11\].id.delaybuf0
timestamp 1606789161
transform 1 0 24064 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_13_137
timestamp 1606789161
transform 1 0 23604 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_141
timestamp 1606789161
transform 1 0 23972 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_141
timestamp 1606789161
transform 1 0 23972 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.dstage\[10\].id.delaybuf1
timestamp 1606789161
transform 1 0 23328 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen0
timestamp 1606789161
transform 1 0 23328 0 -1 19160
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_13_130
timestamp 1606789161
transform 1 0 22960 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_14_130
timestamp 1606789161
transform 1 0 22960 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[10\].id.delayen1
timestamp 1606789161
transform 1 0 22316 0 1 18072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_113
timestamp 1606789161
transform 1 0 22224 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__inv_2  _283_
timestamp 1606789161
transform 1 0 21304 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__and3_4  _290_
timestamp 1606789161
transform 1 0 19924 0 1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[10\].id.delayenb1
timestamp 1606789161
transform 1 0 21948 0 -1 19160
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_13_96
timestamp 1606789161
transform 1 0 19832 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_106
timestamp 1606789161
transform 1 0 20752 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_13_118
timestamp 1606789161
transform 1 0 21856 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_14_103
timestamp 1606789161
transform 1 0 20476 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_111
timestamp 1606789161
transform 1 0 21212 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_14_115
timestamp 1606789161
transform 1 0 21580 0 -1 19160
box -38 -48 406 592
use sky130_fd_sc_hd__or4_4  _457_
timestamp 1606789161
transform 1 0 19648 0 -1 19160
box -38 -48 866 592
use sky130_fd_sc_hd__o22a_4  _515_
timestamp 1606789161
transform 1 0 17992 0 1 18072
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_116
timestamp 1606789161
transform 1 0 19464 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_72
timestamp 1606789161
transform 1 0 17624 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_90
timestamp 1606789161
transform 1 0 19280 0 1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_83
timestamp 1606789161
transform 1 0 18636 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_91
timestamp 1606789161
transform 1 0 19372 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_14_93
timestamp 1606789161
transform 1 0 19556 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__or4_4  _345_
timestamp 1606789161
transform 1 0 15416 0 1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _532_
timestamp 1606789161
transform 1 0 17256 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _557_
timestamp 1606789161
transform 1 0 16520 0 -1 19160
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_112
timestamp 1606789161
transform 1 0 16612 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_57
timestamp 1606789161
transform 1 0 16244 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_13_62
timestamp 1606789161
transform 1 0 16704 0 1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_14_52
timestamp 1606789161
transform 1 0 15784 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__a32o_4  _381_
timestamp 1606789161
transform 1 0 14220 0 -1 19160
box -38 -48 1602 592
use sky130_fd_sc_hd__inv_2  _387_
timestamp 1606789161
transform 1 0 14128 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_115
timestamp 1606789161
transform 1 0 13852 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_13_29
timestamp 1606789161
transform 1 0 13668 0 1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_13_33
timestamp 1606789161
transform 1 0 14036 0 1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_13_37
timestamp 1606789161
transform 1 0 14404 0 1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_13_45
timestamp 1606789161
transform 1 0 15140 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_14_25
timestamp 1606789161
transform 1 0 13300 0 -1 19160
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  FILLER_14_32
timestamp 1606789161
transform 1 0 13944 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _350_
timestamp 1606789161
transform 1 0 12380 0 1 18072
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ai_4  _352_
timestamp 1606789161
transform 1 0 12104 0 -1 19160
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1606789161
transform 1 0 11000 0 1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1606789161
transform 1 0 11000 0 -1 19160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1606789161
transform 1 0 11276 0 1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_14_3
timestamp 1606789161
transform 1 0 11276 0 -1 19160
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_14_11
timestamp 1606789161
transform 1 0 12012 0 -1 19160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1606789161
transform -1 0 30136 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_201
timestamp 1606789161
transform 1 0 29492 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__einvn_8  ringosc.iss.delayenb0
timestamp 1606789161
transform 1 0 26456 0 -1 18072
box -38 -48 1694 592
use sky130_fd_sc_hd__einvn_4  ringosc.iss.delayenb1
timestamp 1606789161
transform 1 0 28480 0 -1 18072
box -38 -48 1050 592
use sky130_fd_sc_hd__fill_1  FILLER_12_167
timestamp 1606789161
transform 1 0 26364 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_12_186
timestamp 1606789161
transform 1 0 28112 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen0
timestamp 1606789161
transform 1 0 25168 0 -1 18072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_111
timestamp 1606789161
transform 1 0 25076 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_146
timestamp 1606789161
transform 1 0 24432 0 -1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_152
timestamp 1606789161
transform 1 0 24984 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_161
timestamp 1606789161
transform 1 0 25812 0 -1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__einvn_4  ringosc.dstage\[11\].id.delayenb1
timestamp 1606789161
transform 1 0 23420 0 -1 18072
box -38 -48 1050 592
use sky130_fd_sc_hd__decap_8  FILLER_12_126
timestamp 1606789161
transform 1 0 22592 0 -1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_134
timestamp 1606789161
transform 1 0 23328 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _289_
timestamp 1606789161
transform 1 0 19924 0 -1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__buf_2  _539_
timestamp 1606789161
transform 1 0 21120 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_12_106
timestamp 1606789161
transform 1 0 20752 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_114
timestamp 1606789161
transform 1 0 21488 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_110
timestamp 1606789161
transform 1 0 19464 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_12_80
timestamp 1606789161
transform 1 0 18360 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_12_93
timestamp 1606789161
transform 1 0 19556 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__and4_4  _337_
timestamp 1606789161
transform 1 0 15416 0 -1 18072
box -38 -48 866 592
use sky130_fd_sc_hd__or2_4  _348_
timestamp 1606789161
transform 1 0 16612 0 -1 18072
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_12_57
timestamp 1606789161
transform 1 0 16244 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_12_68
timestamp 1606789161
transform 1 0 17256 0 -1 18072
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _384_
timestamp 1606789161
transform 1 0 13944 0 -1 18072
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_109
timestamp 1606789161
transform 1 0 13852 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_24
timestamp 1606789161
transform 1 0 13208 0 -1 18072
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_12_30
timestamp 1606789161
transform 1 0 13760 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_12_39
timestamp 1606789161
transform 1 0 14588 0 -1 18072
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_12_47
timestamp 1606789161
transform 1 0 15324 0 -1 18072
box -38 -48 130 592
use sky130_fd_sc_hd__a32o_4  _385_
timestamp 1606789161
transform 1 0 11644 0 -1 18072
box -38 -48 1602 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1606789161
transform 1 0 11000 0 -1 18072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_12_3
timestamp 1606789161
transform 1 0 11276 0 -1 18072
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1606789161
transform -1 0 30136 0 1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_11_201
timestamp 1606789161
transform 1 0 29492 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _522_
timestamp 1606789161
transform 1 0 28296 0 1 16984
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_108
timestamp 1606789161
transform 1 0 27836 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_11_177
timestamp 1606789161
transform 1 0 27284 0 1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_11_184
timestamp 1606789161
transform 1 0 27928 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _456_
timestamp 1606789161
transform 1 0 26088 0 1 16984
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_4  FILLER_11_160
timestamp 1606789161
transform 1 0 25720 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__a21bo_4  _519_
timestamp 1606789161
transform 1 0 22408 0 1 16984
box -38 -48 1234 592
use sky130_fd_sc_hd__einvn_8  ringosc.dstage\[11\].id.delayenb0
timestamp 1606789161
transform 1 0 24064 0 1 16984
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_107
timestamp 1606789161
transform 1 0 22224 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_121
timestamp 1606789161
transform 1 0 22132 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_123
timestamp 1606789161
transform 1 0 22316 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_137
timestamp 1606789161
transform 1 0 23604 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_11_141
timestamp 1606789161
transform 1 0 23972 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_113
timestamp 1606789161
transform 1 0 21396 0 1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _525_
timestamp 1606789161
transform 1 0 17900 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _550_
timestamp 1606789161
transform 1 0 19280 0 1 16984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_8  FILLER_11_79
timestamp 1606789161
transform 1 0 18268 0 1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_11_87
timestamp 1606789161
transform 1 0 19004 0 1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__or3_4  _343_
timestamp 1606789161
transform 1 0 16704 0 1 16984
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_106
timestamp 1606789161
transform 1 0 16612 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_11_52
timestamp 1606789161
transform 1 0 15784 0 1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_60
timestamp 1606789161
transform 1 0 16520 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_11_71
timestamp 1606789161
transform 1 0 17532 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _274_
timestamp 1606789161
transform 1 0 13392 0 1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _386_
timestamp 1606789161
transform 1 0 14496 0 1 16984
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_11_29
timestamp 1606789161
transform 1 0 13668 0 1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_11_37
timestamp 1606789161
transform 1 0 14404 0 1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__nand2_4  _351_
timestamp 1606789161
transform 1 0 12196 0 1 16984
box -38 -48 866 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1606789161
transform 1 0 11000 0 1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_11_3
timestamp 1606789161
transform 1 0 11276 0 1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_11_11
timestamp 1606789161
transform 1 0 12012 0 1 16984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_11_22
timestamp 1606789161
transform 1 0 13024 0 1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen1
timestamp 1606789161
transform 1 0 28572 0 -1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1606789161
transform -1 0 30136 0 -1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_10_198
timestamp 1606789161
transform 1 0 29216 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_204
timestamp 1606789161
transform 1 0 29768 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__einvp_2  ringosc.iss.delayen0
timestamp 1606789161
transform 1 0 27100 0 -1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__fill_2  FILLER_10_173
timestamp 1606789161
transform 1 0 26916 0 -1 16984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_10_182
timestamp 1606789161
transform 1 0 27744 0 -1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_10_190
timestamp 1606789161
transform 1 0 28480 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _523_
timestamp 1606789161
transform 1 0 25168 0 -1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__clkinv_1  ringosc.dstage\[11\].id.delayint0
timestamp 1606789161
transform 1 0 25904 0 -1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_105
timestamp 1606789161
transform 1 0 25076 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_10_151
timestamp 1606789161
transform 1 0 24892 0 -1 16984
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_10_158
timestamp 1606789161
transform 1 0 25536 0 -1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_10_165
timestamp 1606789161
transform 1 0 26180 0 -1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__einvp_2  ringosc.dstage\[11\].id.delayen1
timestamp 1606789161
transform 1 0 23512 0 -1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_10_130
timestamp 1606789161
transform 1 0 22960 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__decap_8  FILLER_10_143
timestamp 1606789161
transform 1 0 24156 0 -1 16984
box -38 -48 774 592
use sky130_fd_sc_hd__dfrtp_4  _551_
timestamp 1606789161
transform 1 0 20844 0 -1 16984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_10_101
timestamp 1606789161
transform 1 0 20292 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__or2_4  _401_
timestamp 1606789161
transform 1 0 19648 0 -1 16984
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_104
timestamp 1606789161
transform 1 0 19464 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_10_85
timestamp 1606789161
transform 1 0 18820 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_91
timestamp 1606789161
transform 1 0 19372 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_93
timestamp 1606789161
transform 1 0 19556 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _564_
timestamp 1606789161
transform 1 0 16704 0 -1 16984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_10_55
timestamp 1606789161
transform 1 0 16060 0 -1 16984
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_10_61
timestamp 1606789161
transform 1 0 16612 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _554_
timestamp 1606789161
transform 1 0 13944 0 -1 16984
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_103
timestamp 1606789161
transform 1 0 13852 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_10_26
timestamp 1606789161
transform 1 0 13392 0 -1 16984
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_10_30
timestamp 1606789161
transform 1 0 13760 0 -1 16984
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _555_
timestamp 1606789161
transform 1 0 11276 0 -1 16984
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1606789161
transform 1 0 11000 0 -1 16984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _527_
timestamp 1606789161
transform 1 0 28572 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1606789161
transform -1 0 30136 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_9_195
timestamp 1606789161
transform 1 0 28940 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_203
timestamp 1606789161
transform 1 0 29676 0 1 15896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _268_
timestamp 1606789161
transform 1 0 27928 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _342_
timestamp 1606789161
transform 1 0 27008 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_102
timestamp 1606789161
transform 1 0 27836 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_9_168
timestamp 1606789161
transform 1 0 26456 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_9_177
timestamp 1606789161
transform 1 0 27284 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_9_187
timestamp 1606789161
transform 1 0 28204 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _526_
timestamp 1606789161
transform 1 0 26088 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_160
timestamp 1606789161
transform 1 0 25720 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _538_
timestamp 1606789161
transform 1 0 22316 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _566_
timestamp 1606789161
transform 1 0 23604 0 1 15896
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_101
timestamp 1606789161
transform 1 0 22224 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_9_127
timestamp 1606789161
transform 1 0 22684 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_9_135
timestamp 1606789161
transform 1 0 23420 0 1 15896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _397_
timestamp 1606789161
transform 1 0 21396 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _398_
timestamp 1606789161
transform 1 0 20384 0 1 15896
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_9_97
timestamp 1606789161
transform 1 0 19924 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_101
timestamp 1606789161
transform 1 0 20292 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_109
timestamp 1606789161
transform 1 0 21028 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_9_116
timestamp 1606789161
transform 1 0 21672 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__and3_4  _400_
timestamp 1606789161
transform 1 0 19096 0 1 15896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_9_80
timestamp 1606789161
transform 1 0 18360 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__a2bb2o_4  _294_
timestamp 1606789161
transform 1 0 16888 0 1 15896
box -38 -48 1510 592
use sky130_fd_sc_hd__inv_2  _340_
timestamp 1606789161
transform 1 0 15876 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_100
timestamp 1606789161
transform 1 0 16612 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_9_49
timestamp 1606789161
transform 1 0 15508 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_9_56
timestamp 1606789161
transform 1 0 16152 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_60
timestamp 1606789161
transform 1 0 16520 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_9_62
timestamp 1606789161
transform 1 0 16704 0 1 15896
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _275_
timestamp 1606789161
transform 1 0 15232 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _535_
timestamp 1606789161
transform 1 0 14404 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_9_26
timestamp 1606789161
transform 1 0 13392 0 1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_9_34
timestamp 1606789161
transform 1 0 14128 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_9_41
timestamp 1606789161
transform 1 0 14772 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_9_45
timestamp 1606789161
transform 1 0 15140 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__buf_2  _534_
timestamp 1606789161
transform 1 0 11920 0 1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1606789161
transform 1 0 11000 0 1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_9_3
timestamp 1606789161
transform 1 0 11276 0 1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_9_9
timestamp 1606789161
transform 1 0 11828 0 1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_9_14
timestamp 1606789161
transform 1 0 12288 0 1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_17
timestamp 1606789161
transform -1 0 30136 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_201
timestamp 1606789161
transform 1 0 29492 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _562_
timestamp 1606789161
transform 1 0 27376 0 -1 15896
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_6  FILLER_8_171
timestamp 1606789161
transform 1 0 26732 0 -1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_8_177
timestamp 1606789161
transform 1 0 27284 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _295_
timestamp 1606789161
transform 1 0 25260 0 -1 15896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_99
timestamp 1606789161
transform 1 0 25076 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_8_145
timestamp 1606789161
transform 1 0 24340 0 -1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_8_154
timestamp 1606789161
transform 1 0 25168 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _292_
timestamp 1606789161
transform 1 0 22868 0 -1 15896
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_8_125
timestamp 1606789161
transform 1 0 22500 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__a21o_4  _313_
timestamp 1606789161
transform 1 0 21396 0 -1 15896
box -38 -48 1142 592
use sky130_fd_sc_hd__and3_4  _389_
timestamp 1606789161
transform 1 0 19832 0 -1 15896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_105
timestamp 1606789161
transform 1 0 20660 0 -1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _388_
timestamp 1606789161
transform 1 0 18360 0 -1 15896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_98
timestamp 1606789161
transform 1 0 19464 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_74
timestamp 1606789161
transform 1 0 17808 0 -1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_8_87
timestamp 1606789161
transform 1 0 19004 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_8_91
timestamp 1606789161
transform 1 0 19372 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_8_93
timestamp 1606789161
transform 1 0 19556 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__nand2_4  _299_
timestamp 1606789161
transform 1 0 16980 0 -1 15896
box -38 -48 866 592
use sky130_fd_sc_hd__decap_8  FILLER_8_54
timestamp 1606789161
transform 1 0 15968 0 -1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_8_62
timestamp 1606789161
transform 1 0 16704 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _293_
timestamp 1606789161
transform 1 0 14496 0 -1 15896
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_97
timestamp 1606789161
transform 1 0 13852 0 -1 15896
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_8_25
timestamp 1606789161
transform 1 0 13300 0 -1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_8_32
timestamp 1606789161
transform 1 0 13944 0 -1 15896
box -38 -48 590 592
use sky130_fd_sc_hd__and2_4  _301_
timestamp 1606789161
transform 1 0 11644 0 -1 15896
box -38 -48 682 592
use sky130_fd_sc_hd__inv_2  _328_
timestamp 1606789161
transform 1 0 13024 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1606789161
transform 1 0 11000 0 -1 15896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_8_3
timestamp 1606789161
transform 1 0 11276 0 -1 15896
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_8_14
timestamp 1606789161
transform 1 0 12288 0 -1 15896
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1606789161
transform -1 0 30136 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_15
timestamp 1606789161
transform -1 0 30136 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_201
timestamp 1606789161
transform 1 0 29492 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_200
timestamp 1606789161
transform 1 0 29400 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_204
timestamp 1606789161
transform 1 0 29768 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _296_
timestamp 1606789161
transform 1 0 27928 0 1 14808
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _561_
timestamp 1606789161
transform 1 0 27376 0 -1 14808
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_96
timestamp 1606789161
transform 1 0 27836 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_174
timestamp 1606789161
transform 1 0 27008 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_178
timestamp 1606789161
transform 1 0 27376 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_182
timestamp 1606789161
transform 1 0 27744 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__and2_4  _326_
timestamp 1606789161
transform 1 0 25168 0 -1 14808
box -38 -48 682 592
use sky130_fd_sc_hd__and4_4  _341_
timestamp 1606789161
transform 1 0 26180 0 -1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__dfrtp_4  _563_
timestamp 1606789161
transform 1 0 25260 0 1 14808
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_93
timestamp 1606789161
transform 1 0 25076 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_6_150
timestamp 1606789161
transform 1 0 24800 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_161
timestamp 1606789161
transform 1 0 25812 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_147
timestamp 1606789161
transform 1 0 24524 0 1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__inv_2  _264_
timestamp 1606789161
transform 1 0 23420 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__and2_4  _309_
timestamp 1606789161
transform 1 0 23880 0 1 14808
box -38 -48 682 592
use sky130_fd_sc_hd__a21bo_4  _315_
timestamp 1606789161
transform 1 0 22316 0 1 14808
box -38 -48 1234 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_95
timestamp 1606789161
transform 1 0 22224 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_131
timestamp 1606789161
transform 1 0 23052 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_6_138
timestamp 1606789161
transform 1 0 23696 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_121
timestamp 1606789161
transform 1 0 22132 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_136
timestamp 1606789161
transform 1 0 23512 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _263_
timestamp 1606789161
transform 1 0 21488 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _311_
timestamp 1606789161
transform 1 0 21764 0 -1 14808
box -38 -48 1326 592
use sky130_fd_sc_hd__a211o_4  _396_
timestamp 1606789161
transform 1 0 19832 0 1 14808
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_12  FILLER_6_101
timestamp 1606789161
transform 1 0 20292 0 -1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_6_113
timestamp 1606789161
transform 1 0 21396 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_110
timestamp 1606789161
transform 1 0 21120 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_117
timestamp 1606789161
transform 1 0 21764 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _390_
timestamp 1606789161
transform 1 0 19648 0 -1 14808
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_92
timestamp 1606789161
transform 1 0 19464 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_88
timestamp 1606789161
transform 1 0 19096 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_6_93
timestamp 1606789161
transform 1 0 19556 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_92
timestamp 1606789161
transform 1 0 19464 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _265_
timestamp 1606789161
transform 1 0 18820 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _399_
timestamp 1606789161
transform 1 0 18820 0 1 14808
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_6_81
timestamp 1606789161
transform 1 0 18452 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_7_81
timestamp 1606789161
transform 1 0 18452 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _267_
timestamp 1606789161
transform 1 0 18176 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_7_74
timestamp 1606789161
transform 1 0 17808 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _266_
timestamp 1606789161
transform 1 0 15416 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _300_
timestamp 1606789161
transform 1 0 16980 0 -1 14808
box -38 -48 1510 592
use sky130_fd_sc_hd__o21a_4  _303_
timestamp 1606789161
transform 1 0 16704 0 1 14808
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_94
timestamp 1606789161
transform 1 0 16612 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_6_61
timestamp 1606789161
transform 1 0 16612 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_7_51
timestamp 1606789161
transform 1 0 15692 0 1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_7_59
timestamp 1606789161
transform 1 0 16428 0 1 14808
box -38 -48 222 592
use sky130_fd_sc_hd__a2bb2o_4  _298_
timestamp 1606789161
transform 1 0 15140 0 -1 14808
box -38 -48 1510 592
use sky130_fd_sc_hd__buf_2  _524_
timestamp 1606789161
transform 1 0 13944 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_91
timestamp 1606789161
transform 1 0 13852 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_6_24
timestamp 1606789161
transform 1 0 13208 0 -1 14808
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_6_30
timestamp 1606789161
transform 1 0 13760 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_6_36
timestamp 1606789161
transform 1 0 14312 0 -1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_6_44
timestamp 1606789161
transform 1 0 15048 0 -1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_7_44
timestamp 1606789161
transform 1 0 15048 0 1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__nor2_4  _302_
timestamp 1606789161
transform 1 0 11368 0 1 14808
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _304_
timestamp 1606789161
transform 1 0 11276 0 -1 14808
box -38 -48 1326 592
use sky130_fd_sc_hd__inv_2  _305_
timestamp 1606789161
transform 1 0 12932 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _565_
timestamp 1606789161
transform 1 0 12932 0 1 14808
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1606789161
transform 1 0 11000 0 -1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1606789161
transform 1 0 11000 0 1 14808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_6_17
timestamp 1606789161
transform 1 0 12564 0 -1 14808
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_7_3
timestamp 1606789161
transform 1 0 11276 0 1 14808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_7_13
timestamp 1606789161
transform 1 0 12196 0 1 14808
box -38 -48 774 592
use sky130_fd_sc_hd__clkbuf_1  ringosc.iss.delaybuf0
timestamp 1606789161
transform 1 0 28940 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1606789161
transform -1 0 30136 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_191
timestamp 1606789161
transform 1 0 28572 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_5_198
timestamp 1606789161
transform 1 0 29216 0 1 13720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_5_204
timestamp 1606789161
transform 1 0 29768 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__or2_4  _297_
timestamp 1606789161
transform 1 0 27928 0 1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_90
timestamp 1606789161
transform 1 0 27836 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_172
timestamp 1606789161
transform 1 0 26824 0 1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_5_180
timestamp 1606789161
transform 1 0 27560 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_5_160
timestamp 1606789161
transform 1 0 25720 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__or2_4  _314_
timestamp 1606789161
transform 1 0 22316 0 1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__a22oi_4  _316_
timestamp 1606789161
transform 1 0 24156 0 1 13720
box -38 -48 1602 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_89
timestamp 1606789161
transform 1 0 22224 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_5_130
timestamp 1606789161
transform 1 0 22960 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_5_142
timestamp 1606789161
transform 1 0 24064 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__and4_4  _395_
timestamp 1606789161
transform 1 0 20016 0 1 13720
box -38 -48 866 592
use sky130_fd_sc_hd__decap_12  FILLER_5_107
timestamp 1606789161
transform 1 0 20844 0 1 13720
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_5_119
timestamp 1606789161
transform 1 0 21948 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_5_94
timestamp 1606789161
transform 1 0 19648 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _321_
timestamp 1606789161
transform 1 0 15600 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _540_
timestamp 1606789161
transform 1 0 16796 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _549_
timestamp 1606789161
transform 1 0 17532 0 1 13720
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_88
timestamp 1606789161
transform 1 0 16612 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_5_53
timestamp 1606789161
transform 1 0 15876 0 1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_5_62
timestamp 1606789161
transform 1 0 16704 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_67
timestamp 1606789161
transform 1 0 17164 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__or2_4  _331_
timestamp 1606789161
transform 1 0 14588 0 1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_4  FILLER_5_35
timestamp 1606789161
transform 1 0 14220 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_5_46
timestamp 1606789161
transform 1 0 15232 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _327_
timestamp 1606789161
transform 1 0 12932 0 1 13720
box -38 -48 1326 592
use sky130_fd_sc_hd__o21ai_4  _338_
timestamp 1606789161
transform 1 0 11368 0 1 13720
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1606789161
transform 1 0 11000 0 1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_5_3
timestamp 1606789161
transform 1 0 11276 0 1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_5_17
timestamp 1606789161
transform 1 0 12564 0 1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  _528_
timestamp 1606789161
transform 1 0 29032 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1606789161
transform -1 0 30136 0 -1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_4_192
timestamp 1606789161
transform 1 0 28664 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_4_200
timestamp 1606789161
transform 1 0 29400 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_204
timestamp 1606789161
transform 1 0 29768 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_4  _548_
timestamp 1606789161
transform 1 0 26548 0 -1 13720
box -38 -48 2154 592
use sky130_fd_sc_hd__and3_4  _320_
timestamp 1606789161
transform 1 0 25168 0 -1 13720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_87
timestamp 1606789161
transform 1 0 25076 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_149
timestamp 1606789161
transform 1 0 24708 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_4_163
timestamp 1606789161
transform 1 0 25996 0 -1 13720
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _317_
timestamp 1606789161
transform 1 0 23420 0 -1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _319_
timestamp 1606789161
transform 1 0 24064 0 -1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_8  FILLER_4_127
timestamp 1606789161
transform 1 0 22684 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_4_138
timestamp 1606789161
transform 1 0 23696 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _312_
timestamp 1606789161
transform 1 0 21212 0 -1 13720
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_8  FILLER_4_102
timestamp 1606789161
transform 1 0 20384 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_4_110
timestamp 1606789161
transform 1 0 21120 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__nor2_4  _392_
timestamp 1606789161
transform 1 0 19556 0 -1 13720
box -38 -48 866 592
use sky130_fd_sc_hd__a211o_4  _402_
timestamp 1606789161
transform 1 0 17716 0 -1 13720
box -38 -48 1326 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_86
timestamp 1606789161
transform 1 0 19464 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_4_87
timestamp 1606789161
transform 1 0 19004 0 -1 13720
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_4_91
timestamp 1606789161
transform 1 0 19372 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _310_
timestamp 1606789161
transform 1 0 15508 0 -1 13720
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_8  FILLER_4_63
timestamp 1606789161
transform 1 0 16796 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_4_71
timestamp 1606789161
transform 1 0 17532 0 -1 13720
box -38 -48 222 592
use sky130_fd_sc_hd__or4_4  _339_
timestamp 1606789161
transform 1 0 13944 0 -1 13720
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_85
timestamp 1606789161
transform 1 0 13852 0 -1 13720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_4_29
timestamp 1606789161
transform 1 0 13668 0 -1 13720
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_4_41
timestamp 1606789161
transform 1 0 14772 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__or2_4  _306_
timestamp 1606789161
transform 1 0 12288 0 -1 13720
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1606789161
transform 1 0 11000 0 -1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_3
timestamp 1606789161
transform 1 0 11276 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_4_11
timestamp 1606789161
transform 1 0 12012 0 -1 13720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_4_21
timestamp 1606789161
transform 1 0 12932 0 -1 13720
box -38 -48 774 592
use sky130_fd_sc_hd__clkinv_1  ringosc.iss.delayint0
timestamp 1606789161
transform 1 0 28664 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1606789161
transform -1 0 30136 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_3_195
timestamp 1606789161
transform 1 0 28940 0 1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_3_203
timestamp 1606789161
transform 1 0 29676 0 1 12632
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _541_
timestamp 1606789161
transform 1 0 27928 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_84
timestamp 1606789161
transform 1 0 27836 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_177
timestamp 1606789161
transform 1 0 27284 0 1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_3_188
timestamp 1606789161
transform 1 0 28296 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _287_
timestamp 1606789161
transform 1 0 25904 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__or2_4  _318_
timestamp 1606789161
transform 1 0 24892 0 1 12632
box -38 -48 682 592
use sky130_fd_sc_hd__fill_1  FILLER_3_150
timestamp 1606789161
transform 1 0 24800 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_3_158
timestamp 1606789161
transform 1 0 25536 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_3_165
timestamp 1606789161
transform 1 0 26180 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _261_
timestamp 1606789161
transform 1 0 22316 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__clkinv_2  ringosc.ibufp10
timestamp 1606789161
transform 1 0 23696 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_83
timestamp 1606789161
transform 1 0 22224 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_126
timestamp 1606789161
transform 1 0 22592 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_3_142
timestamp 1606789161
transform 1 0 24064 0 1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__a21o_4  _308_
timestamp 1606789161
transform 1 0 20752 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_118
timestamp 1606789161
transform 1 0 21856 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__a211o_4  _393_
timestamp 1606789161
transform 1 0 18360 0 1 12632
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_3_74
timestamp 1606789161
transform 1 0 17808 0 1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_94
timestamp 1606789161
transform 1 0 19648 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_82
timestamp 1606789161
transform 1 0 16612 0 1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_3_49
timestamp 1606789161
transform 1 0 15508 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_3_62
timestamp 1606789161
transform 1 0 16704 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__inv_2  _260_
timestamp 1606789161
transform 1 0 15232 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__a2bb2o_4  _324_
timestamp 1606789161
transform 1 0 13392 0 1 12632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_3_42
timestamp 1606789161
transform 1 0 14864 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__and2_4  _325_
timestamp 1606789161
transform 1 0 12380 0 1 12632
box -38 -48 682 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1606789161
transform 1 0 11000 0 1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_3_3
timestamp 1606789161
transform 1 0 11276 0 1 12632
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_3_22
timestamp 1606789161
transform 1 0 13024 0 1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1606789161
transform -1 0 30136 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_2_200
timestamp 1606789161
transform 1 0 29400 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_204
timestamp 1606789161
transform 1 0 29768 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _286_
timestamp 1606789161
transform 1 0 27928 0 -1 12632
box -38 -48 1510 592
use sky130_fd_sc_hd__decap_4  FILLER_2_180
timestamp 1606789161
transform 1 0 27560 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _547_
timestamp 1606789161
transform 1 0 25444 0 -1 12632
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_81
timestamp 1606789161
transform 1 0 25076 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_145
timestamp 1606789161
transform 1 0 24340 0 -1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_2_154
timestamp 1606789161
transform 1 0 25168 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_4  _567_
timestamp 1606789161
transform 1 0 22224 0 -1 12632
box -38 -48 2154 592
use sky130_fd_sc_hd__fill_1  FILLER_2_121
timestamp 1606789161
transform 1 0 22132 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__o22a_4  _323_
timestamp 1606789161
transform 1 0 20476 0 -1 12632
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_6  FILLER_2_96
timestamp 1606789161
transform 1 0 19832 0 -1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_102
timestamp 1606789161
transform 1 0 20384 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_117
timestamp 1606789161
transform 1 0 21764 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _394_
timestamp 1606789161
transform 1 0 19556 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_80
timestamp 1606789161
transform 1 0 19464 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_2_84
timestamp 1606789161
transform 1 0 18728 0 -1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _544_
timestamp 1606789161
transform 1 0 15876 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _553_
timestamp 1606789161
transform 1 0 16612 0 -1 12632
box -38 -48 2154 592
use sky130_fd_sc_hd__decap_4  FILLER_2_48
timestamp 1606789161
transform 1 0 15416 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_2_52
timestamp 1606789161
transform 1 0 15784 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_2_57
timestamp 1606789161
transform 1 0 16244 0 -1 12632
box -38 -48 406 592
use sky130_fd_sc_hd__a2bb2o_4  _322_
timestamp 1606789161
transform 1 0 13944 0 -1 12632
box -38 -48 1510 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_79
timestamp 1606789161
transform 1 0 13852 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_2_24
timestamp 1606789161
transform 1 0 13208 0 -1 12632
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_2_30
timestamp 1606789161
transform 1 0 13760 0 -1 12632
box -38 -48 130 592
use sky130_fd_sc_hd__o21ai_4  _330_
timestamp 1606789161
transform 1 0 12012 0 -1 12632
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1606789161
transform 1 0 11000 0 -1 12632
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_2_3
timestamp 1606789161
transform 1 0 11276 0 -1 12632
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1606789161
transform -1 0 30136 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1606789161
transform -1 0 30136 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_6  FILLER_0_199
timestamp 1606789161
transform 1 0 29308 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_6  FILLER_1_199
timestamp 1606789161
transform 1 0 29308 0 1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__inv_2  _276_
timestamp 1606789161
transform 1 0 27928 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _542_
timestamp 1606789161
transform 1 0 26364 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_75
timestamp 1606789161
transform 1 0 28112 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_78
timestamp 1606789161
transform 1 0 27836 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_172
timestamp 1606789161
transform 1 0 26824 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_184
timestamp 1606789161
transform 1 0 27928 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_12  FILLER_0_187
timestamp 1606789161
transform 1 0 28204 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_171
timestamp 1606789161
transform 1 0 26732 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_187
timestamp 1606789161
transform 1 0 28204 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _543_
timestamp 1606789161
transform 1 0 25352 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_74
timestamp 1606789161
transform 1 0 25260 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_0_160
timestamp 1606789161
transform 1 0 25720 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_163
timestamp 1606789161
transform 1 0 25996 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _546_
timestamp 1606789161
transform 1 0 23880 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__clkinv_8  ringosc.ibufp11
timestamp 1606789161
transform 1 0 22960 0 -1 11544
box -38 -48 1234 592
use sky130_fd_sc_hd__decap_12  FILLER_0_143
timestamp 1606789161
transform 1 0 24156 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_1_126
timestamp 1606789161
transform 1 0 22592 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_1_138
timestamp 1606789161
transform 1 0 23696 0 1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _262_
timestamp 1606789161
transform 1 0 22316 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_73
timestamp 1606789161
transform 1 0 22408 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_77
timestamp 1606789161
transform 1 0 22224 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_120
timestamp 1606789161
transform 1 0 22040 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_125
timestamp 1606789161
transform 1 0 22500 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_129
timestamp 1606789161
transform 1 0 22868 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _291_
timestamp 1606789161
transform 1 0 20568 0 -1 11544
box -38 -48 1510 592
use sky130_fd_sc_hd__and2_4  _307_
timestamp 1606789161
transform 1 0 21212 0 1 11544
box -38 -48 682 592
use sky130_fd_sc_hd__decap_6  FILLER_0_98
timestamp 1606789161
transform 1 0 20016 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_106
timestamp 1606789161
transform 1 0 20752 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_110
timestamp 1606789161
transform 1 0 21120 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_118
timestamp 1606789161
transform 1 0 21856 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _259_
timestamp 1606789161
transform 1 0 18636 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _537_
timestamp 1606789161
transform 1 0 19648 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__dfrtp_4  _552_
timestamp 1606789161
transform 1 0 18636 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_72
timestamp 1606789161
transform 1 0 19556 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_73
timestamp 1606789161
transform 1 0 17716 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_81
timestamp 1606789161
transform 1 0 18452 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_6  FILLER_0_86
timestamp 1606789161
transform 1 0 18912 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_92
timestamp 1606789161
transform 1 0 19464 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_1_79
timestamp 1606789161
transform 1 0 18268 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__o21a_4  _391_
timestamp 1606789161
transform 1 0 17164 0 1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__buf_2  _536_
timestamp 1606789161
transform 1 0 17348 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_71
timestamp 1606789161
transform 1 0 16704 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_76
timestamp 1606789161
transform 1 0 16612 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_58
timestamp 1606789161
transform 1 0 16336 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_0_63
timestamp 1606789161
transform 1 0 16796 0 -1 11544
box -38 -48 590 592
use sky130_fd_sc_hd__decap_4  FILLER_1_57
timestamp 1606789161
transform 1 0 16244 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_1_62
timestamp 1606789161
transform 1 0 16704 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_1_66
timestamp 1606789161
transform 1 0 17072 0 1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__a2bb2o_4  _288_
timestamp 1606789161
transform 1 0 14864 0 -1 11544
box -38 -48 1510 592
use sky130_fd_sc_hd__dfrtp_4  _568_
timestamp 1606789161
transform 1 0 14128 0 1 11544
box -38 -48 2154 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_70
timestamp 1606789161
transform 1 0 13852 0 -1 11544
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_27
timestamp 1606789161
transform 1 0 13484 0 -1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_32
timestamp 1606789161
transform 1 0 13944 0 -1 11544
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_40
timestamp 1606789161
transform 1 0 14680 0 -1 11544
box -38 -48 222 592
use sky130_fd_sc_hd__decap_4  FILLER_1_30
timestamp 1606789161
transform 1 0 13760 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__inv_2  _277_
timestamp 1606789161
transform 1 0 11644 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__o22a_4  _329_
timestamp 1606789161
transform 1 0 12472 0 1 11544
box -38 -48 1326 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1606789161
transform 1 0 11000 0 -1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1606789161
transform 1 0 11000 0 1 11544
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_0_3
timestamp 1606789161
transform 1 0 11276 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_0_15
timestamp 1606789161
transform 1 0 12380 0 -1 11544
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_1_3
timestamp 1606789161
transform 1 0 11276 0 1 11544
box -38 -48 406 592
use sky130_fd_sc_hd__decap_6  FILLER_1_10
timestamp 1606789161
transform 1 0 11920 0 1 11544
box -38 -48 590 592
<< labels >>
rlabel metal2 s 27762 31576 27818 32376 4 clockp[0]
port 1 nsew
rlabel metal2 s 21690 8824 21746 9624 4 clockp[1]
port 2 nsew
rlabel metal2 s 12306 8824 12362 9624 4 dco
port 3 nsew
rlabel metal2 s 10466 8824 10522 9624 4 div[0]
port 4 nsew
rlabel metal3 s 9896 17808 10696 17928 4 div[1]
port 5 nsew
rlabel metal2 s 27394 8824 27450 9624 4 div[2]
port 6 nsew
rlabel metal3 s 30504 10464 31304 10584 4 div[3]
port 7 nsew
rlabel metal3 s 9896 12368 10696 12488 4 div[4]
port 8 nsew
rlabel metal2 s 20218 31576 20274 32376 4 enable
port 9 nsew
rlabel metal2 s 14514 31576 14570 32376 4 ext_trim[0]
port 10 nsew
rlabel metal2 s 23898 31576 23954 32376 4 ext_trim[10]
port 11 nsew
rlabel metal3 s 9896 23520 10696 23640 4 ext_trim[11]
port 12 nsew
rlabel metal3 s 30504 13184 31304 13304 4 ext_trim[12]
port 13 nsew
rlabel metal2 s 29418 8824 29474 9624 4 ext_trim[13]
port 14 nsew
rlabel metal3 s 9896 20800 10696 20920 4 ext_trim[14]
port 15 nsew
rlabel metal2 s 14146 8824 14202 9624 4 ext_trim[15]
port 16 nsew
rlabel metal3 s 30504 27328 31304 27448 4 ext_trim[16]
port 17 nsew
rlabel metal3 s 9896 26240 10696 26360 4 ext_trim[17]
port 18 nsew
rlabel metal2 s 29602 31576 29658 32376 4 ext_trim[18]
port 19 nsew
rlabel metal2 s 18194 31576 18250 32376 4 ext_trim[19]
port 20 nsew
rlabel metal3 s 30504 24608 31304 24728 4 ext_trim[1]
port 21 nsew
rlabel metal2 s 25554 8824 25610 9624 4 ext_trim[20]
port 22 nsew
rlabel metal3 s 9896 29232 10696 29352 4 ext_trim[21]
port 23 nsew
rlabel metal3 s 30504 21616 31304 21736 4 ext_trim[22]
port 24 nsew
rlabel metal3 s 9896 15088 10696 15208 4 ext_trim[23]
port 25 nsew
rlabel metal2 s 19850 8824 19906 9624 4 ext_trim[24]
port 26 nsew
rlabel metal3 s 30504 16176 31304 16296 4 ext_trim[25]
port 27 nsew
rlabel metal3 s 30504 18896 31304 19016 4 ext_trim[2]
port 28 nsew
rlabel metal2 s 12490 31576 12546 32376 4 ext_trim[3]
port 29 nsew
rlabel metal2 s 25922 31576 25978 32376 4 ext_trim[4]
port 30 nsew
rlabel metal2 s 23714 8824 23770 9624 4 ext_trim[5]
port 31 nsew
rlabel metal2 s 22058 31576 22114 32376 4 ext_trim[6]
port 32 nsew
rlabel metal2 s 10650 31576 10706 32376 4 ext_trim[7]
port 33 nsew
rlabel metal2 s 16354 31576 16410 32376 4 ext_trim[8]
port 34 nsew
rlabel metal3 s 30504 30048 31304 30168 4 ext_trim[9]
port 35 nsew
rlabel metal2 s 18010 8824 18066 9624 4 osc
port 36 nsew
rlabel metal2 s 15986 8824 16042 9624 4 resetb
port 37 nsew
rlabel metal4 s 5000 5000 9000 36040 4 VPWR
port 38 nsew
rlabel metal4 s 0 0 4000 41040 4 VGND
port 39 nsew
<< properties >>
string FIXED_BBOX 0 0 41136 41040
string GDS_FILE digital_pll.gds
string GDS_END 2654930
string GDS_START 265824
<< end >>
