magic
tech sky130A
magscale 12 1
timestamp 1598787399
<< metal5 >>
rect 0 45 30 75
rect 0 0 30 30
<< properties >>
string FIXED_BBOX 0 -30 45 105
<< end >>
