*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* Simple testbench mainly to check SPICE model conversion from CDL
* Plots the transient response of the smallest inverter in the HD standard cell library

.lib "/home/tim/projects/efabless/tech/SW/sky130A/libs.tech/ngspice/sky130.lib.spice" tt
.include "/home/tim/projects/efabless/tech/SW/sky130A/libs.ref/sky130_fd_sc_hd/spice/sky130_fd_sc_hd.spice"

* .option TEMP=27

X0 in vss vss vdd vdd out sky130_fd_sc_hd__inv_1

V0 vdd vss PWL(0n 0.0 30n 1.8)
V1 vss 0 0.0

Vin in vss PWL(0n 0.0 100n 0.0 500n 1.8)

* Transient analysis
.control
tran 1n 1u
plot V(in) V(out)
.endc
.end
