magic
tech sky130A
timestamp 1619448499
<< metal2 >>
rect 9701 351760 9757 352480
rect 29159 351760 29215 352480
rect 48617 351760 48673 352480
rect 68075 351760 68131 352480
rect 87533 351760 87589 352480
rect 107037 351760 107093 352480
rect 126495 351760 126551 352480
rect 145953 351760 146009 352480
rect 165411 351760 165467 352480
rect 184869 351760 184925 352480
rect 204373 351760 204429 352480
rect 223831 351760 223887 352480
rect 243289 351760 243345 352480
rect 262747 351760 262803 352480
rect 282205 351760 282261 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4365 -480 4421 240
rect 4963 -480 5019 240
rect 5561 -480 5617 240
rect 6159 -480 6215 240
rect 6757 -480 6813 240
rect 7355 -480 7411 240
rect 7953 -480 8009 240
rect 8505 -480 8561 240
rect 9103 -480 9159 240
rect 9701 -480 9757 240
rect 10299 -480 10355 240
rect 10897 -480 10953 240
rect 11495 -480 11551 240
rect 12093 -480 12149 240
rect 12645 -480 12701 240
rect 13243 -480 13299 240
rect 13841 -480 13897 240
rect 14439 -480 14495 240
rect 15037 -480 15093 240
rect 15635 -480 15691 240
rect 16187 -480 16243 240
rect 16785 -480 16841 240
rect 17383 -480 17439 240
rect 17981 -480 18037 240
rect 18579 -480 18635 240
rect 19177 -480 19233 240
rect 19775 -480 19831 240
rect 20327 -480 20383 240
rect 20925 -480 20981 240
rect 21523 -480 21579 240
rect 22121 -480 22177 240
rect 22719 -480 22775 240
rect 23317 -480 23373 240
rect 23915 -480 23971 240
rect 24467 -480 24523 240
rect 25065 -480 25121 240
rect 25663 -480 25719 240
rect 26261 -480 26317 240
rect 26859 -480 26915 240
rect 27457 -480 27513 240
rect 28009 -480 28065 240
rect 28607 -480 28663 240
rect 29205 -480 29261 240
rect 29803 -480 29859 240
rect 30401 -480 30457 240
rect 30999 -480 31055 240
rect 31597 -480 31653 240
rect 32149 -480 32205 240
rect 32747 -480 32803 240
rect 33345 -480 33401 240
rect 33943 -480 33999 240
rect 34541 -480 34597 240
rect 35139 -480 35195 240
rect 35737 -480 35793 240
rect 36289 -480 36345 240
rect 36887 -480 36943 240
rect 37485 -480 37541 240
rect 38083 -480 38139 240
rect 38681 -480 38737 240
rect 39279 -480 39335 240
rect 39831 -480 39887 240
rect 40429 -480 40485 240
rect 41027 -480 41083 240
rect 41625 -480 41681 240
rect 42223 -480 42279 240
rect 42821 -480 42877 240
rect 43419 -480 43475 240
rect 43971 -480 44027 240
rect 44569 -480 44625 240
rect 45167 -480 45223 240
rect 45765 -480 45821 240
rect 46363 -480 46419 240
rect 46961 -480 47017 240
rect 47559 -480 47615 240
rect 48111 -480 48167 240
rect 48709 -480 48765 240
rect 49307 -480 49363 240
rect 49905 -480 49961 240
rect 50503 -480 50559 240
rect 51101 -480 51157 240
rect 51653 -480 51709 240
rect 52251 -480 52307 240
rect 52849 -480 52905 240
rect 53447 -480 53503 240
rect 54045 -480 54101 240
rect 54643 -480 54699 240
rect 55241 -480 55297 240
rect 55793 -480 55849 240
rect 56391 -480 56447 240
rect 56989 -480 57045 240
rect 57587 -480 57643 240
rect 58185 -480 58241 240
rect 58783 -480 58839 240
rect 59381 -480 59437 240
rect 59933 -480 59989 240
rect 60531 -480 60587 240
rect 61129 -480 61185 240
rect 61727 -480 61783 240
rect 62325 -480 62381 240
rect 62923 -480 62979 240
rect 63475 -480 63531 240
rect 64073 -480 64129 240
rect 64671 -480 64727 240
rect 65269 -480 65325 240
rect 65867 -480 65923 240
rect 66465 -480 66521 240
rect 67063 -480 67119 240
rect 67615 -480 67671 240
rect 68213 -480 68269 240
rect 68811 -480 68867 240
rect 69409 -480 69465 240
rect 70007 -480 70063 240
rect 70605 -480 70661 240
rect 71203 -480 71259 240
rect 71755 -480 71811 240
rect 72353 -480 72409 240
rect 72951 -480 73007 240
rect 73549 -480 73605 240
rect 74147 -480 74203 240
rect 74745 -480 74801 240
rect 75297 -480 75353 240
rect 75895 -480 75951 240
rect 76493 -480 76549 240
rect 77091 -480 77147 240
rect 77689 -480 77745 240
rect 78287 -480 78343 240
rect 78885 -480 78941 240
rect 79437 -480 79493 240
rect 80035 -480 80091 240
rect 80633 -480 80689 240
rect 81231 -480 81287 240
rect 81829 -480 81885 240
rect 82427 -480 82483 240
rect 83025 -480 83081 240
rect 83577 -480 83633 240
rect 84175 -480 84231 240
rect 84773 -480 84829 240
rect 85371 -480 85427 240
rect 85969 -480 86025 240
rect 86567 -480 86623 240
rect 87119 -480 87175 240
rect 87717 -480 87773 240
rect 88315 -480 88371 240
rect 88913 -480 88969 240
rect 89511 -480 89567 240
rect 90109 -480 90165 240
rect 90707 -480 90763 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92455 -480 92511 240
rect 93053 -480 93109 240
rect 93651 -480 93707 240
rect 94249 -480 94305 240
rect 94847 -480 94903 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98941 -480 98997 240
rect 99539 -480 99595 240
rect 100137 -480 100193 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103081 -480 103137 240
rect 103679 -480 103735 240
rect 104277 -480 104333 240
rect 104875 -480 104931 240
rect 105473 -480 105529 240
rect 106071 -480 106127 240
rect 106669 -480 106725 240
rect 107221 -480 107277 240
rect 107819 -480 107875 240
rect 108417 -480 108473 240
rect 109015 -480 109071 240
rect 109613 -480 109669 240
rect 110211 -480 110267 240
rect 110763 -480 110819 240
rect 111361 -480 111417 240
rect 111959 -480 112015 240
rect 112557 -480 112613 240
rect 113155 -480 113211 240
rect 113753 -480 113809 240
rect 114351 -480 114407 240
rect 114903 -480 114959 240
rect 115501 -480 115557 240
rect 116099 -480 116155 240
rect 116697 -480 116753 240
rect 117295 -480 117351 240
rect 117893 -480 117949 240
rect 118491 -480 118547 240
rect 119043 -480 119099 240
rect 119641 -480 119697 240
rect 120239 -480 120295 240
rect 120837 -480 120893 240
rect 121435 -480 121491 240
rect 122033 -480 122089 240
rect 122585 -480 122641 240
rect 123183 -480 123239 240
rect 123781 -480 123837 240
rect 124379 -480 124435 240
rect 124977 -480 125033 240
rect 125575 -480 125631 240
rect 126173 -480 126229 240
rect 126725 -480 126781 240
rect 127323 -480 127379 240
rect 127921 -480 127977 240
rect 128519 -480 128575 240
rect 129117 -480 129173 240
rect 129715 -480 129771 240
rect 130313 -480 130369 240
rect 130865 -480 130921 240
rect 131463 -480 131519 240
rect 132061 -480 132117 240
rect 132659 -480 132715 240
rect 133257 -480 133313 240
rect 133855 -480 133911 240
rect 134407 -480 134463 240
rect 135005 -480 135061 240
rect 135603 -480 135659 240
rect 136201 -480 136257 240
rect 136799 -480 136855 240
rect 137397 -480 137453 240
rect 137995 -480 138051 240
rect 138547 -480 138603 240
rect 139145 -480 139201 240
rect 139743 -480 139799 240
rect 140341 -480 140397 240
rect 140939 -480 140995 240
rect 141537 -480 141593 240
rect 142135 -480 142191 240
rect 142687 -480 142743 240
rect 143285 -480 143341 240
rect 143883 -480 143939 240
rect 144481 -480 144537 240
rect 145079 -480 145135 240
rect 145677 -480 145733 240
rect 146275 -480 146331 240
rect 146827 -480 146883 240
rect 147425 -480 147481 240
rect 148023 -480 148079 240
rect 148621 -480 148677 240
rect 149219 -480 149275 240
rect 149817 -480 149873 240
rect 150369 -480 150425 240
rect 150967 -480 151023 240
rect 151565 -480 151621 240
rect 152163 -480 152219 240
rect 152761 -480 152817 240
rect 153359 -480 153415 240
rect 153957 -480 154013 240
rect 154509 -480 154565 240
rect 155107 -480 155163 240
rect 155705 -480 155761 240
rect 156303 -480 156359 240
rect 156901 -480 156957 240
rect 157499 -480 157555 240
rect 158097 -480 158153 240
rect 158649 -480 158705 240
rect 159247 -480 159303 240
rect 159845 -480 159901 240
rect 160443 -480 160499 240
rect 161041 -480 161097 240
rect 161639 -480 161695 240
rect 162191 -480 162247 240
rect 162789 -480 162845 240
rect 163387 -480 163443 240
rect 163985 -480 164041 240
rect 164583 -480 164639 240
rect 165181 -480 165237 240
rect 165779 -480 165835 240
rect 166331 -480 166387 240
rect 166929 -480 166985 240
rect 167527 -480 167583 240
rect 168125 -480 168181 240
rect 168723 -480 168779 240
rect 169321 -480 169377 240
rect 169919 -480 169975 240
rect 170471 -480 170527 240
rect 171069 -480 171125 240
rect 171667 -480 171723 240
rect 172265 -480 172321 240
rect 172863 -480 172919 240
rect 173461 -480 173517 240
rect 174013 -480 174069 240
rect 174611 -480 174667 240
rect 175209 -480 175265 240
rect 175807 -480 175863 240
rect 176405 -480 176461 240
rect 177003 -480 177059 240
rect 177601 -480 177657 240
rect 178153 -480 178209 240
rect 178751 -480 178807 240
rect 179349 -480 179405 240
rect 179947 -480 180003 240
rect 180545 -480 180601 240
rect 181143 -480 181199 240
rect 181741 -480 181797 240
rect 182293 -480 182349 240
rect 182891 -480 182947 240
rect 183489 -480 183545 240
rect 184087 -480 184143 240
rect 184685 -480 184741 240
rect 185283 -480 185339 240
rect 185835 -480 185891 240
rect 186433 -480 186489 240
rect 187031 -480 187087 240
rect 187629 -480 187685 240
rect 188227 -480 188283 240
rect 188825 -480 188881 240
rect 189423 -480 189479 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192367 -480 192423 240
rect 192965 -480 193021 240
rect 193563 -480 193619 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197657 -480 197713 240
rect 198255 -480 198311 240
rect 198853 -480 198909 240
rect 199451 -480 199507 240
rect 200049 -480 200105 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201797 -480 201853 240
rect 202395 -480 202451 240
rect 202993 -480 203049 240
rect 203591 -480 203647 240
rect 204189 -480 204245 240
rect 204787 -480 204843 240
rect 205385 -480 205441 240
rect 205937 -480 205993 240
rect 206535 -480 206591 240
rect 207133 -480 207189 240
rect 207731 -480 207787 240
rect 208329 -480 208385 240
rect 208927 -480 208983 240
rect 209479 -480 209535 240
rect 210077 -480 210133 240
rect 210675 -480 210731 240
rect 211273 -480 211329 240
rect 211871 -480 211927 240
rect 212469 -480 212525 240
rect 213067 -480 213123 240
rect 213619 -480 213675 240
rect 214217 -480 214273 240
rect 214815 -480 214871 240
rect 215413 -480 215469 240
rect 216011 -480 216067 240
rect 216609 -480 216665 240
rect 217207 -480 217263 240
rect 217759 -480 217815 240
rect 218357 -480 218413 240
rect 218955 -480 219011 240
rect 219553 -480 219609 240
rect 220151 -480 220207 240
rect 220749 -480 220805 240
rect 221301 -480 221357 240
rect 221899 -480 221955 240
rect 222497 -480 222553 240
rect 223095 -480 223151 240
rect 223693 -480 223749 240
rect 224291 -480 224347 240
rect 224889 -480 224945 240
rect 225441 -480 225497 240
rect 226039 -480 226095 240
rect 226637 -480 226693 240
rect 227235 -480 227291 240
rect 227833 -480 227889 240
rect 228431 -480 228487 240
rect 229029 -480 229085 240
rect 229581 -480 229637 240
rect 230179 -480 230235 240
rect 230777 -480 230833 240
rect 231375 -480 231431 240
rect 231973 -480 232029 240
rect 232571 -480 232627 240
rect 233123 -480 233179 240
rect 233721 -480 233777 240
rect 234319 -480 234375 240
rect 234917 -480 234973 240
rect 235515 -480 235571 240
rect 236113 -480 236169 240
rect 236711 -480 236767 240
rect 237263 -480 237319 240
rect 237861 -480 237917 240
rect 238459 -480 238515 240
rect 239057 -480 239113 240
rect 239655 -480 239711 240
rect 240253 -480 240309 240
rect 240851 -480 240907 240
rect 241403 -480 241459 240
rect 242001 -480 242057 240
rect 242599 -480 242655 240
rect 243197 -480 243253 240
rect 243795 -480 243851 240
rect 244393 -480 244449 240
rect 244945 -480 245001 240
rect 245543 -480 245599 240
rect 246141 -480 246197 240
rect 246739 -480 246795 240
rect 247337 -480 247393 240
rect 247935 -480 247991 240
rect 248533 -480 248589 240
rect 249085 -480 249141 240
rect 249683 -480 249739 240
rect 250281 -480 250337 240
rect 250879 -480 250935 240
rect 251477 -480 251533 240
rect 252075 -480 252131 240
rect 252673 -480 252729 240
rect 253225 -480 253281 240
rect 253823 -480 253879 240
rect 254421 -480 254477 240
rect 255019 -480 255075 240
rect 255617 -480 255673 240
rect 256215 -480 256271 240
rect 256767 -480 256823 240
rect 257365 -480 257421 240
rect 257963 -480 258019 240
rect 258561 -480 258617 240
rect 259159 -480 259215 240
rect 259757 -480 259813 240
rect 260355 -480 260411 240
rect 260907 -480 260963 240
rect 261505 -480 261561 240
rect 262103 -480 262159 240
rect 262701 -480 262757 240
rect 263299 -480 263355 240
rect 263897 -480 263953 240
rect 264495 -480 264551 240
rect 265047 -480 265103 240
rect 265645 -480 265701 240
rect 266243 -480 266299 240
rect 266841 -480 266897 240
rect 267439 -480 267495 240
rect 268037 -480 268093 240
rect 268589 -480 268645 240
rect 269187 -480 269243 240
rect 269785 -480 269841 240
rect 270383 -480 270439 240
rect 270981 -480 271037 240
rect 271579 -480 271635 240
rect 272177 -480 272233 240
rect 272729 -480 272785 240
rect 273327 -480 273383 240
rect 273925 -480 273981 240
rect 274523 -480 274579 240
rect 275121 -480 275177 240
rect 275719 -480 275775 240
rect 276317 -480 276373 240
rect 276869 -480 276925 240
rect 277467 -480 277523 240
rect 278065 -480 278121 240
rect 278663 -480 278719 240
rect 279261 -480 279317 240
rect 279859 -480 279915 240
rect 280411 -480 280467 240
rect 281009 -480 281065 240
rect 281607 -480 281663 240
rect 282205 -480 282261 240
rect 282803 -480 282859 240
rect 283401 -480 283457 240
rect 283999 -480 284055 240
rect 284551 -480 284607 240
rect 285149 -480 285205 240
rect 285747 -480 285803 240
rect 286345 -480 286401 240
rect 286943 -480 286999 240
rect 287541 -480 287597 240
rect 288139 -480 288195 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect -480 349494 240 349614
rect 291760 349426 292480 349546
rect -480 344802 240 344922
rect 291760 344462 292480 344582
rect -480 340110 240 340230
rect 291760 339498 292480 339618
rect -480 335418 240 335538
rect 291760 334534 292480 334654
rect -480 330726 240 330846
rect 291760 329570 292480 329690
rect -480 326034 240 326154
rect 291760 324606 292480 324726
rect -480 321342 240 321462
rect 291760 319642 292480 319762
rect -480 316650 240 316770
rect 291760 314678 292480 314798
rect -480 311958 240 312078
rect 291760 309714 292480 309834
rect -480 307266 240 307386
rect 291760 304750 292480 304870
rect -480 302574 240 302694
rect 291760 299854 292480 299974
rect -480 297882 240 298002
rect 291760 294890 292480 295010
rect -480 293190 240 293310
rect 291760 289926 292480 290046
rect -480 288498 240 288618
rect 291760 284962 292480 285082
rect -480 283806 240 283926
rect 291760 279998 292480 280118
rect -480 279114 240 279234
rect 291760 275034 292480 275154
rect -480 274422 240 274542
rect 291760 270070 292480 270190
rect -480 269730 240 269850
rect -480 265038 240 265158
rect 291760 265106 292480 265226
rect -480 260346 240 260466
rect 291760 260142 292480 260262
rect -480 255654 240 255774
rect 291760 255178 292480 255298
rect -480 250962 240 251082
rect 291760 250282 292480 250402
rect -480 246270 240 246390
rect 291760 245318 292480 245438
rect -480 241578 240 241698
rect 291760 240354 292480 240474
rect -480 236886 240 237006
rect 291760 235390 292480 235510
rect -480 232194 240 232314
rect 291760 230426 292480 230546
rect -480 227502 240 227622
rect 291760 225462 292480 225582
rect -480 222810 240 222930
rect 291760 220498 292480 220618
rect -480 218118 240 218238
rect 291760 215534 292480 215654
rect -480 213426 240 213546
rect 291760 210570 292480 210690
rect -480 208734 240 208854
rect 291760 205606 292480 205726
rect -480 204042 240 204162
rect 291760 200710 292480 200830
rect -480 199350 240 199470
rect 291760 195746 292480 195866
rect -480 194658 240 194778
rect 291760 190782 292480 190902
rect -480 189966 240 190086
rect 291760 185818 292480 185938
rect -480 185274 240 185394
rect 291760 180854 292480 180974
rect -480 180582 240 180702
rect -480 175890 240 176010
rect 291760 175890 292480 176010
rect -480 171198 240 171318
rect 291760 170926 292480 171046
rect -480 166506 240 166626
rect 291760 165962 292480 166082
rect -480 161814 240 161934
rect 291760 160998 292480 161118
rect -480 157122 240 157242
rect 291760 156034 292480 156154
rect -480 152430 240 152550
rect 291760 151138 292480 151258
rect -480 147738 240 147858
rect 291760 146174 292480 146294
rect -480 143046 240 143166
rect 291760 141210 292480 141330
rect -480 138354 240 138474
rect 291760 136246 292480 136366
rect -480 133662 240 133782
rect 291760 131282 292480 131402
rect -480 128970 240 129090
rect 291760 126318 292480 126438
rect -480 124278 240 124398
rect 291760 121354 292480 121474
rect -480 119586 240 119706
rect 291760 116390 292480 116510
rect -480 114894 240 115014
rect 291760 111426 292480 111546
rect -480 110202 240 110322
rect 291760 106462 292480 106582
rect -480 105510 240 105630
rect 291760 101566 292480 101686
rect -480 100818 240 100938
rect 291760 96602 292480 96722
rect -480 96126 240 96246
rect 291760 91638 292480 91758
rect -480 91434 240 91554
rect -480 86742 240 86862
rect 291760 86674 292480 86794
rect -480 82050 240 82170
rect 291760 81710 292480 81830
rect -480 77358 240 77478
rect 291760 76746 292480 76866
rect -480 72666 240 72786
rect 291760 71782 292480 71902
rect -480 67974 240 68094
rect 291760 66818 292480 66938
rect -480 63282 240 63402
rect 291760 61854 292480 61974
rect -480 58590 240 58710
rect 291760 56890 292480 57010
rect -480 53898 240 54018
rect 291760 51994 292480 52114
rect -480 49206 240 49326
rect 291760 47030 292480 47150
rect -480 44514 240 44634
rect 291760 42066 292480 42186
rect -480 39822 240 39942
rect 291760 37102 292480 37222
rect -480 35130 240 35250
rect 291760 32138 292480 32258
rect -480 30438 240 30558
rect 291760 27174 292480 27294
rect -480 25746 240 25866
rect 291760 22210 292480 22330
rect -480 21054 240 21174
rect 291760 17246 292480 17366
rect -480 16362 240 16482
rect 291760 12282 292480 12402
rect -480 11670 240 11790
rect 291760 7318 292480 7438
rect -480 6978 240 7098
rect 291760 2422 292480 2542
rect -480 2286 240 2406
<< metal4 >>
rect -4288 355709 -3988 355720
rect -4288 355591 -4197 355709
rect -4079 355591 -3988 355709
rect -4288 355549 -3988 355591
rect -4288 355431 -4197 355549
rect -4079 355431 -3988 355549
rect -4288 -3463 -3988 355431
rect 295950 355709 296250 355720
rect 295950 355591 296041 355709
rect 296159 355591 296250 355709
rect 295950 355549 296250 355591
rect 295950 355431 296041 355549
rect 296159 355431 296250 355549
rect -3818 355239 -3518 355250
rect -3818 355121 -3727 355239
rect -3609 355121 -3518 355239
rect -3818 355079 -3518 355121
rect -3818 354961 -3727 355079
rect -3609 354961 -3518 355079
rect -3818 -2993 -3518 354961
rect 295480 355239 295780 355250
rect 295480 355121 295571 355239
rect 295689 355121 295780 355239
rect 295480 355079 295780 355121
rect 295480 354961 295571 355079
rect 295689 354961 295780 355079
rect -3348 354769 -3048 354780
rect -3348 354651 -3257 354769
rect -3139 354651 -3048 354769
rect -3348 354609 -3048 354651
rect -3348 354491 -3257 354609
rect -3139 354491 -3048 354609
rect -3348 -2523 -3048 354491
rect 295010 354769 295310 354780
rect 295010 354651 295101 354769
rect 295219 354651 295310 354769
rect 295010 354609 295310 354651
rect 295010 354491 295101 354609
rect 295219 354491 295310 354609
rect -2878 354299 -2578 354310
rect -2878 354181 -2787 354299
rect -2669 354181 -2578 354299
rect -2878 354139 -2578 354181
rect -2878 354021 -2787 354139
rect -2669 354021 -2578 354139
rect -2878 -2053 -2578 354021
rect 294540 354299 294840 354310
rect 294540 354181 294631 354299
rect 294749 354181 294840 354299
rect 294540 354139 294840 354181
rect 294540 354021 294631 354139
rect 294749 354021 294840 354139
rect -2408 353829 -2108 353840
rect -2408 353711 -2317 353829
rect -2199 353711 -2108 353829
rect -2408 353669 -2108 353711
rect -2408 353551 -2317 353669
rect -2199 353551 -2108 353669
rect -2408 -1583 -2108 353551
rect 294070 353829 294370 353840
rect 294070 353711 294161 353829
rect 294279 353711 294370 353829
rect 294070 353669 294370 353711
rect 294070 353551 294161 353669
rect 294279 353551 294370 353669
rect -1938 353359 -1638 353370
rect -1938 353241 -1847 353359
rect -1729 353241 -1638 353359
rect -1938 353199 -1638 353241
rect -1938 353081 -1847 353199
rect -1729 353081 -1638 353199
rect -1938 -1113 -1638 353081
rect 293600 353359 293900 353370
rect 293600 353241 293691 353359
rect 293809 353241 293900 353359
rect 293600 353199 293900 353241
rect 293600 353081 293691 353199
rect 293809 353081 293900 353199
rect -1468 352889 -1168 352900
rect -1468 352771 -1377 352889
rect -1259 352771 -1168 352889
rect -1468 352729 -1168 352771
rect -1468 352611 -1377 352729
rect -1259 352611 -1168 352729
rect -1468 -643 -1168 352611
rect 293130 352889 293430 352900
rect 293130 352771 293221 352889
rect 293339 352771 293430 352889
rect 293130 352729 293430 352771
rect 293130 352611 293221 352729
rect 293339 352611 293430 352729
rect -998 352419 -698 352430
rect -998 352301 -907 352419
rect -789 352301 -698 352419
rect -998 352259 -698 352301
rect -998 352141 -907 352259
rect -789 352141 -698 352259
rect -998 -173 -698 352141
rect -998 -291 -907 -173
rect -789 -291 -698 -173
rect -998 -333 -698 -291
rect -998 -451 -907 -333
rect -789 -451 -698 -333
rect -998 -462 -698 -451
rect 292660 352419 292960 352430
rect 292660 352301 292751 352419
rect 292869 352301 292960 352419
rect 292660 352259 292960 352301
rect 292660 352141 292751 352259
rect 292869 352141 292960 352259
rect 292660 -173 292960 352141
rect 292660 -291 292751 -173
rect 292869 -291 292960 -173
rect 292660 -333 292960 -291
rect 292660 -451 292751 -333
rect 292869 -451 292960 -333
rect 292660 -462 292960 -451
rect -1468 -761 -1377 -643
rect -1259 -761 -1168 -643
rect -1468 -803 -1168 -761
rect -1468 -921 -1377 -803
rect -1259 -921 -1168 -803
rect -1468 -932 -1168 -921
rect 293130 -643 293430 352611
rect 293130 -761 293221 -643
rect 293339 -761 293430 -643
rect 293130 -803 293430 -761
rect 293130 -921 293221 -803
rect 293339 -921 293430 -803
rect 293130 -932 293430 -921
rect -1938 -1231 -1847 -1113
rect -1729 -1231 -1638 -1113
rect -1938 -1273 -1638 -1231
rect -1938 -1391 -1847 -1273
rect -1729 -1391 -1638 -1273
rect -1938 -1402 -1638 -1391
rect 293600 -1113 293900 353081
rect 293600 -1231 293691 -1113
rect 293809 -1231 293900 -1113
rect 293600 -1273 293900 -1231
rect 293600 -1391 293691 -1273
rect 293809 -1391 293900 -1273
rect 293600 -1402 293900 -1391
rect -2408 -1701 -2317 -1583
rect -2199 -1701 -2108 -1583
rect -2408 -1743 -2108 -1701
rect -2408 -1861 -2317 -1743
rect -2199 -1861 -2108 -1743
rect -2408 -1872 -2108 -1861
rect 294070 -1583 294370 353551
rect 294070 -1701 294161 -1583
rect 294279 -1701 294370 -1583
rect 294070 -1743 294370 -1701
rect 294070 -1861 294161 -1743
rect 294279 -1861 294370 -1743
rect 294070 -1872 294370 -1861
rect -2878 -2171 -2787 -2053
rect -2669 -2171 -2578 -2053
rect -2878 -2213 -2578 -2171
rect -2878 -2331 -2787 -2213
rect -2669 -2331 -2578 -2213
rect -2878 -2342 -2578 -2331
rect 294540 -2053 294840 354021
rect 294540 -2171 294631 -2053
rect 294749 -2171 294840 -2053
rect 294540 -2213 294840 -2171
rect 294540 -2331 294631 -2213
rect 294749 -2331 294840 -2213
rect 294540 -2342 294840 -2331
rect -3348 -2641 -3257 -2523
rect -3139 -2641 -3048 -2523
rect -3348 -2683 -3048 -2641
rect -3348 -2801 -3257 -2683
rect -3139 -2801 -3048 -2683
rect -3348 -2812 -3048 -2801
rect 295010 -2523 295310 354491
rect 295010 -2641 295101 -2523
rect 295219 -2641 295310 -2523
rect 295010 -2683 295310 -2641
rect 295010 -2801 295101 -2683
rect 295219 -2801 295310 -2683
rect 295010 -2812 295310 -2801
rect -3818 -3111 -3727 -2993
rect -3609 -3111 -3518 -2993
rect -3818 -3153 -3518 -3111
rect -3818 -3271 -3727 -3153
rect -3609 -3271 -3518 -3153
rect -3818 -3282 -3518 -3271
rect 295480 -2993 295780 354961
rect 295480 -3111 295571 -2993
rect 295689 -3111 295780 -2993
rect 295480 -3153 295780 -3111
rect 295480 -3271 295571 -3153
rect 295689 -3271 295780 -3153
rect 295480 -3282 295780 -3271
rect -4288 -3581 -4197 -3463
rect -4079 -3581 -3988 -3463
rect -4288 -3623 -3988 -3581
rect -4288 -3741 -4197 -3623
rect -4079 -3741 -3988 -3623
rect -4288 -3752 -3988 -3741
rect 295950 -3463 296250 355431
rect 295950 -3581 296041 -3463
rect 296159 -3581 296250 -3463
rect 295950 -3623 296250 -3581
rect 295950 -3741 296041 -3623
rect 296159 -3741 296250 -3623
rect 295950 -3752 296250 -3741
<< via4 >>
rect -4197 355591 -4079 355709
rect -4197 355431 -4079 355549
rect 296041 355591 296159 355709
rect 296041 355431 296159 355549
rect -3727 355121 -3609 355239
rect -3727 354961 -3609 355079
rect 295571 355121 295689 355239
rect 295571 354961 295689 355079
rect -3257 354651 -3139 354769
rect -3257 354491 -3139 354609
rect 295101 354651 295219 354769
rect 295101 354491 295219 354609
rect -2787 354181 -2669 354299
rect -2787 354021 -2669 354139
rect 294631 354181 294749 354299
rect 294631 354021 294749 354139
rect -2317 353711 -2199 353829
rect -2317 353551 -2199 353669
rect 294161 353711 294279 353829
rect 294161 353551 294279 353669
rect -1847 353241 -1729 353359
rect -1847 353081 -1729 353199
rect 293691 353241 293809 353359
rect 293691 353081 293809 353199
rect -1377 352771 -1259 352889
rect -1377 352611 -1259 352729
rect 293221 352771 293339 352889
rect 293221 352611 293339 352729
rect -907 352301 -789 352419
rect -907 352141 -789 352259
rect -907 -291 -789 -173
rect -907 -451 -789 -333
rect 292751 352301 292869 352419
rect 292751 352141 292869 352259
rect 292751 -291 292869 -173
rect 292751 -451 292869 -333
rect -1377 -761 -1259 -643
rect -1377 -921 -1259 -803
rect 293221 -761 293339 -643
rect 293221 -921 293339 -803
rect -1847 -1231 -1729 -1113
rect -1847 -1391 -1729 -1273
rect 293691 -1231 293809 -1113
rect 293691 -1391 293809 -1273
rect -2317 -1701 -2199 -1583
rect -2317 -1861 -2199 -1743
rect 294161 -1701 294279 -1583
rect 294161 -1861 294279 -1743
rect -2787 -2171 -2669 -2053
rect -2787 -2331 -2669 -2213
rect 294631 -2171 294749 -2053
rect 294631 -2331 294749 -2213
rect -3257 -2641 -3139 -2523
rect -3257 -2801 -3139 -2683
rect 295101 -2641 295219 -2523
rect 295101 -2801 295219 -2683
rect -3727 -3111 -3609 -2993
rect -3727 -3271 -3609 -3153
rect 295571 -3111 295689 -2993
rect 295571 -3271 295689 -3153
rect -4197 -3581 -4079 -3463
rect -4197 -3741 -4079 -3623
rect 296041 -3581 296159 -3463
rect 296041 -3741 296159 -3623
<< metal5 >>
rect -4288 355720 -3988 355721
rect 295950 355720 296250 355721
rect -4288 355709 296250 355720
rect -4288 355591 -4197 355709
rect -4079 355591 296041 355709
rect 296159 355591 296250 355709
rect -4288 355549 296250 355591
rect -4288 355431 -4197 355549
rect -4079 355431 296041 355549
rect 296159 355431 296250 355549
rect -4288 355420 296250 355431
rect -4288 355419 -3988 355420
rect 295950 355419 296250 355420
rect -3818 355250 -3518 355251
rect 295480 355250 295780 355251
rect -3818 355239 295780 355250
rect -3818 355121 -3727 355239
rect -3609 355121 295571 355239
rect 295689 355121 295780 355239
rect -3818 355079 295780 355121
rect -3818 354961 -3727 355079
rect -3609 354961 295571 355079
rect 295689 354961 295780 355079
rect -3818 354950 295780 354961
rect -3818 354949 -3518 354950
rect 295480 354949 295780 354950
rect -3348 354780 -3048 354781
rect 295010 354780 295310 354781
rect -3348 354769 295310 354780
rect -3348 354651 -3257 354769
rect -3139 354651 295101 354769
rect 295219 354651 295310 354769
rect -3348 354609 295310 354651
rect -3348 354491 -3257 354609
rect -3139 354491 295101 354609
rect 295219 354491 295310 354609
rect -3348 354480 295310 354491
rect -3348 354479 -3048 354480
rect 295010 354479 295310 354480
rect -2878 354310 -2578 354311
rect 294540 354310 294840 354311
rect -2878 354299 294840 354310
rect -2878 354181 -2787 354299
rect -2669 354181 294631 354299
rect 294749 354181 294840 354299
rect -2878 354139 294840 354181
rect -2878 354021 -2787 354139
rect -2669 354021 294631 354139
rect 294749 354021 294840 354139
rect -2878 354010 294840 354021
rect -2878 354009 -2578 354010
rect 294540 354009 294840 354010
rect -2408 353840 -2108 353841
rect 294070 353840 294370 353841
rect -2408 353829 294370 353840
rect -2408 353711 -2317 353829
rect -2199 353711 294161 353829
rect 294279 353711 294370 353829
rect -2408 353669 294370 353711
rect -2408 353551 -2317 353669
rect -2199 353551 294161 353669
rect 294279 353551 294370 353669
rect -2408 353540 294370 353551
rect -2408 353539 -2108 353540
rect 294070 353539 294370 353540
rect -1938 353370 -1638 353371
rect 293600 353370 293900 353371
rect -1938 353359 293900 353370
rect -1938 353241 -1847 353359
rect -1729 353241 293691 353359
rect 293809 353241 293900 353359
rect -1938 353199 293900 353241
rect -1938 353081 -1847 353199
rect -1729 353081 293691 353199
rect 293809 353081 293900 353199
rect -1938 353070 293900 353081
rect -1938 353069 -1638 353070
rect 293600 353069 293900 353070
rect -1468 352900 -1168 352901
rect 293130 352900 293430 352901
rect -1468 352889 293430 352900
rect -1468 352771 -1377 352889
rect -1259 352771 293221 352889
rect 293339 352771 293430 352889
rect -1468 352729 293430 352771
rect -1468 352611 -1377 352729
rect -1259 352611 293221 352729
rect 293339 352611 293430 352729
rect -1468 352600 293430 352611
rect -1468 352599 -1168 352600
rect 293130 352599 293430 352600
rect -998 352430 -698 352431
rect 292660 352430 292960 352431
rect -998 352419 292960 352430
rect -998 352301 -907 352419
rect -789 352301 292751 352419
rect 292869 352301 292960 352419
rect -998 352259 292960 352301
rect -998 352141 -907 352259
rect -789 352141 292751 352259
rect 292869 352141 292960 352259
rect -998 352130 292960 352141
rect -998 352129 -698 352130
rect 292660 352129 292960 352130
rect -998 -162 -698 -161
rect 292660 -162 292960 -161
rect -998 -173 292960 -162
rect -998 -291 -907 -173
rect -789 -291 292751 -173
rect 292869 -291 292960 -173
rect -998 -333 292960 -291
rect -998 -451 -907 -333
rect -789 -451 292751 -333
rect 292869 -451 292960 -333
rect -998 -462 292960 -451
rect -998 -463 -698 -462
rect 292660 -463 292960 -462
rect -1468 -632 -1168 -631
rect 293130 -632 293430 -631
rect -1468 -643 293430 -632
rect -1468 -761 -1377 -643
rect -1259 -761 293221 -643
rect 293339 -761 293430 -643
rect -1468 -803 293430 -761
rect -1468 -921 -1377 -803
rect -1259 -921 293221 -803
rect 293339 -921 293430 -803
rect -1468 -932 293430 -921
rect -1468 -933 -1168 -932
rect 293130 -933 293430 -932
rect -1938 -1102 -1638 -1101
rect 293600 -1102 293900 -1101
rect -1938 -1113 293900 -1102
rect -1938 -1231 -1847 -1113
rect -1729 -1231 293691 -1113
rect 293809 -1231 293900 -1113
rect -1938 -1273 293900 -1231
rect -1938 -1391 -1847 -1273
rect -1729 -1391 293691 -1273
rect 293809 -1391 293900 -1273
rect -1938 -1402 293900 -1391
rect -1938 -1403 -1638 -1402
rect 293600 -1403 293900 -1402
rect -2408 -1572 -2108 -1571
rect 294070 -1572 294370 -1571
rect -2408 -1583 294370 -1572
rect -2408 -1701 -2317 -1583
rect -2199 -1701 294161 -1583
rect 294279 -1701 294370 -1583
rect -2408 -1743 294370 -1701
rect -2408 -1861 -2317 -1743
rect -2199 -1861 294161 -1743
rect 294279 -1861 294370 -1743
rect -2408 -1872 294370 -1861
rect -2408 -1873 -2108 -1872
rect 294070 -1873 294370 -1872
rect -2878 -2042 -2578 -2041
rect 294540 -2042 294840 -2041
rect -2878 -2053 294840 -2042
rect -2878 -2171 -2787 -2053
rect -2669 -2171 294631 -2053
rect 294749 -2171 294840 -2053
rect -2878 -2213 294840 -2171
rect -2878 -2331 -2787 -2213
rect -2669 -2331 294631 -2213
rect 294749 -2331 294840 -2213
rect -2878 -2342 294840 -2331
rect -2878 -2343 -2578 -2342
rect 294540 -2343 294840 -2342
rect -3348 -2512 -3048 -2511
rect 295010 -2512 295310 -2511
rect -3348 -2523 295310 -2512
rect -3348 -2641 -3257 -2523
rect -3139 -2641 295101 -2523
rect 295219 -2641 295310 -2523
rect -3348 -2683 295310 -2641
rect -3348 -2801 -3257 -2683
rect -3139 -2801 295101 -2683
rect 295219 -2801 295310 -2683
rect -3348 -2812 295310 -2801
rect -3348 -2813 -3048 -2812
rect 295010 -2813 295310 -2812
rect -3818 -2982 -3518 -2981
rect 295480 -2982 295780 -2981
rect -3818 -2993 295780 -2982
rect -3818 -3111 -3727 -2993
rect -3609 -3111 295571 -2993
rect 295689 -3111 295780 -2993
rect -3818 -3153 295780 -3111
rect -3818 -3271 -3727 -3153
rect -3609 -3271 295571 -3153
rect 295689 -3271 295780 -3153
rect -3818 -3282 295780 -3271
rect -3818 -3283 -3518 -3282
rect 295480 -3283 295780 -3282
rect -4288 -3452 -3988 -3451
rect 295950 -3452 296250 -3451
rect -4288 -3463 296250 -3452
rect -4288 -3581 -4197 -3463
rect -4079 -3581 296041 -3463
rect 296159 -3581 296250 -3463
rect -4288 -3623 296250 -3581
rect -4288 -3741 -4197 -3623
rect -4079 -3741 296041 -3623
rect 296159 -3741 296250 -3623
rect -4288 -3752 296250 -3741
rect -4288 -3753 -3988 -3752
rect 295950 -3753 296250 -3752
<< labels >>
rlabel metal3 s 291760 141210 292480 141330 6 gpio_analog[0]
port 0 nsew signal bidirectional
rlabel metal3 s -480 279114 240 279234 4 gpio_analog[10]
port 1 nsew signal bidirectional
rlabel metal3 s -480 250962 240 251082 4 gpio_analog[11]
port 2 nsew signal bidirectional
rlabel metal3 s -480 222810 240 222930 4 gpio_analog[12]
port 3 nsew signal bidirectional
rlabel metal3 s -480 194658 240 194778 4 gpio_analog[13]
port 4 nsew signal bidirectional
rlabel metal3 s -480 166506 240 166626 4 gpio_analog[14]
port 5 nsew signal bidirectional
rlabel metal3 s -480 138354 240 138474 4 gpio_analog[15]
port 6 nsew signal bidirectional
rlabel metal3 s -480 110202 240 110322 4 gpio_analog[16]
port 7 nsew signal bidirectional
rlabel metal3 s -480 82050 240 82170 4 gpio_analog[17]
port 8 nsew signal bidirectional
rlabel metal3 s 291760 170926 292480 171046 6 gpio_analog[1]
port 9 nsew signal bidirectional
rlabel metal3 s 291760 200710 292480 200830 6 gpio_analog[2]
port 10 nsew signal bidirectional
rlabel metal3 s 291760 230426 292480 230546 6 gpio_analog[3]
port 11 nsew signal bidirectional
rlabel metal3 s 291760 260142 292480 260262 6 gpio_analog[4]
port 12 nsew signal bidirectional
rlabel metal3 s 291760 289926 292480 290046 6 gpio_analog[5]
port 13 nsew signal bidirectional
rlabel metal3 s 291760 319642 292480 319762 6 gpio_analog[6]
port 14 nsew signal bidirectional
rlabel metal3 s -480 344802 240 344922 4 gpio_analog[7]
port 15 nsew signal bidirectional
rlabel metal3 s -480 335418 240 335538 4 gpio_analog[8]
port 16 nsew signal bidirectional
rlabel metal3 s -480 307266 240 307386 4 gpio_analog[9]
port 17 nsew signal bidirectional
rlabel metal3 s 291760 146174 292480 146294 6 gpio_noesd[0]
port 18 nsew signal bidirectional
rlabel metal3 s -480 274422 240 274542 4 gpio_noesd[10]
port 19 nsew signal bidirectional
rlabel metal3 s -480 246270 240 246390 4 gpio_noesd[11]
port 20 nsew signal bidirectional
rlabel metal3 s -480 218118 240 218238 4 gpio_noesd[12]
port 21 nsew signal bidirectional
rlabel metal3 s -480 189966 240 190086 4 gpio_noesd[13]
port 22 nsew signal bidirectional
rlabel metal3 s -480 161814 240 161934 4 gpio_noesd[14]
port 23 nsew signal bidirectional
rlabel metal3 s -480 133662 240 133782 4 gpio_noesd[15]
port 24 nsew signal bidirectional
rlabel metal3 s -480 105510 240 105630 4 gpio_noesd[16]
port 25 nsew signal bidirectional
rlabel metal3 s -480 77358 240 77478 4 gpio_noesd[17]
port 26 nsew signal bidirectional
rlabel metal3 s 291760 175890 292480 176010 6 gpio_noesd[1]
port 27 nsew signal bidirectional
rlabel metal3 s 291760 205606 292480 205726 6 gpio_noesd[2]
port 28 nsew signal bidirectional
rlabel metal3 s 291760 235390 292480 235510 6 gpio_noesd[3]
port 29 nsew signal bidirectional
rlabel metal3 s 291760 265106 292480 265226 6 gpio_noesd[4]
port 30 nsew signal bidirectional
rlabel metal3 s 291760 294890 292480 295010 6 gpio_noesd[5]
port 31 nsew signal bidirectional
rlabel metal3 s 291760 324606 292480 324726 6 gpio_noesd[6]
port 32 nsew signal bidirectional
rlabel metal3 s -480 340110 240 340230 4 gpio_noesd[7]
port 33 nsew signal bidirectional
rlabel metal3 s -480 330726 240 330846 4 gpio_noesd[8]
port 34 nsew signal bidirectional
rlabel metal3 s -480 302574 240 302694 4 gpio_noesd[9]
port 35 nsew signal bidirectional
rlabel metal3 s 291760 349426 292480 349546 6 io_analog[0]
port 36 nsew signal bidirectional
rlabel metal3 s -480 349494 240 349614 4 io_analog[10]
port 37 nsew signal bidirectional
rlabel metal2 s 282205 351760 282261 352480 6 io_analog[1]
port 38 nsew signal bidirectional
rlabel metal2 s 262747 351760 262803 352480 6 io_analog[2]
port 39 nsew signal bidirectional
rlabel metal2 s 243289 351760 243345 352480 6 io_analog[3]
port 40 nsew signal bidirectional
rlabel metal2 s 184869 351760 184925 352480 6 io_analog[4]
port 41 nsew signal bidirectional
rlabel metal2 s 126495 351760 126551 352480 6 io_analog[5]
port 42 nsew signal bidirectional
rlabel metal2 s 68075 351760 68131 352480 6 io_analog[6]
port 43 nsew signal bidirectional
rlabel metal2 s 48617 351760 48673 352480 6 io_analog[7]
port 44 nsew signal bidirectional
rlabel metal2 s 29159 351760 29215 352480 6 io_analog[8]
port 45 nsew signal bidirectional
rlabel metal2 s 9701 351760 9757 352480 6 io_analog[9]
port 46 nsew signal bidirectional
rlabel metal2 s 223831 351760 223887 352480 6 io_clamp_high[0]
port 47 nsew signal bidirectional
rlabel metal2 s 165411 351760 165467 352480 6 io_clamp_high[1]
port 48 nsew signal bidirectional
rlabel metal2 s 107037 351760 107093 352480 6 io_clamp_high[2]
port 49 nsew signal bidirectional
rlabel metal2 s 204373 351760 204429 352480 6 io_clamp_low[0]
port 50 nsew signal bidirectional
rlabel metal2 s 145953 351760 146009 352480 6 io_clamp_low[1]
port 51 nsew signal bidirectional
rlabel metal2 s 87533 351760 87589 352480 6 io_clamp_low[2]
port 52 nsew signal bidirectional
rlabel metal3 s 291760 7318 292480 7438 6 io_in[0]
port 53 nsew signal input
rlabel metal3 s 291760 12282 292480 12402 6 io_out[0]
port 54 nsew signal tristate
rlabel metal3 s 291760 245318 292480 245438 6 io_in[10]
port 55 nsew signal input
rlabel metal3 s 291760 250282 292480 250402 6 io_out[10]
port 56 nsew signal tristate
rlabel metal3 s 291760 275034 292480 275154 6 io_in[11]
port 57 nsew signal input
rlabel metal3 s 291760 279998 292480 280118 6 io_out[11]
port 58 nsew signal tristate
rlabel metal3 s 291760 304750 292480 304870 6 io_in[12]
port 59 nsew signal input
rlabel metal3 s 291760 309714 292480 309834 6 io_out[12]
port 60 nsew signal tristate
rlabel metal3 s 291760 334534 292480 334654 6 io_in[13]
port 61 nsew signal input
rlabel metal3 s 291760 339498 292480 339618 6 io_out[13]
port 62 nsew signal tristate
rlabel metal3 s -480 321342 240 321462 4 io_in[14]
port 63 nsew signal input
rlabel metal3 s -480 316650 240 316770 4 io_out[14]
port 64 nsew signal tristate
rlabel metal3 s -480 293190 240 293310 4 io_in[15]
port 65 nsew signal input
rlabel metal3 s -480 288498 240 288618 4 io_out[15]
port 66 nsew signal tristate
rlabel metal3 s -480 265038 240 265158 4 io_in[16]
port 67 nsew signal input
rlabel metal3 s -480 260346 240 260466 4 io_out[16]
port 68 nsew signal tristate
rlabel metal3 s -480 236886 240 237006 4 io_in[17]
port 69 nsew signal input
rlabel metal3 s -480 232194 240 232314 4 io_out[17]
port 70 nsew signal tristate
rlabel metal3 s -480 208734 240 208854 4 io_in[18]
port 71 nsew signal input
rlabel metal3 s -480 204042 240 204162 4 io_out[18]
port 72 nsew signal tristate
rlabel metal3 s -480 180582 240 180702 4 io_in[19]
port 73 nsew signal input
rlabel metal3 s -480 175890 240 176010 4 io_out[19]
port 74 nsew signal tristate
rlabel metal3 s 291760 27174 292480 27294 6 io_in[1]
port 75 nsew signal input
rlabel metal3 s 291760 32138 292480 32258 6 io_out[1]
port 76 nsew signal tristate
rlabel metal3 s -480 152430 240 152550 4 io_in[20]
port 77 nsew signal input
rlabel metal3 s -480 147738 240 147858 4 io_out[20]
port 78 nsew signal tristate
rlabel metal3 s -480 124278 240 124398 4 io_in[21]
port 79 nsew signal input
rlabel metal3 s -480 119586 240 119706 4 io_out[21]
port 80 nsew signal tristate
rlabel metal3 s -480 96126 240 96246 4 io_in[22]
port 81 nsew signal input
rlabel metal3 s -480 91434 240 91554 4 io_out[22]
port 82 nsew signal tristate
rlabel metal3 s -480 67974 240 68094 4 io_in[23]
port 83 nsew signal input
rlabel metal3 s -480 63282 240 63402 4 io_out[23]
port 84 nsew signal tristate
rlabel metal3 s -480 49206 240 49326 4 io_in[24]
port 85 nsew signal input
rlabel metal3 s -480 44514 240 44634 4 io_out[24]
port 86 nsew signal tristate
rlabel metal3 s -480 30438 240 30558 4 io_in[25]
port 87 nsew signal input
rlabel metal3 s -480 25746 240 25866 4 io_out[25]
port 88 nsew signal tristate
rlabel metal3 s -480 11670 240 11790 4 io_in[26]
port 89 nsew signal input
rlabel metal3 s -480 6978 240 7098 4 io_out[26]
port 90 nsew signal tristate
rlabel metal3 s 291760 47030 292480 47150 6 io_in[2]
port 91 nsew signal input
rlabel metal3 s 291760 51994 292480 52114 6 io_out[2]
port 92 nsew signal tristate
rlabel metal3 s 291760 66818 292480 66938 6 io_in[3]
port 93 nsew signal input
rlabel metal3 s 291760 71782 292480 71902 6 io_out[3]
port 94 nsew signal tristate
rlabel metal3 s 291760 86674 292480 86794 6 io_in[4]
port 95 nsew signal input
rlabel metal3 s 291760 91638 292480 91758 6 io_out[4]
port 96 nsew signal tristate
rlabel metal3 s 291760 106462 292480 106582 6 io_in[5]
port 97 nsew signal input
rlabel metal3 s 291760 111426 292480 111546 6 io_out[5]
port 98 nsew signal tristate
rlabel metal3 s 291760 126318 292480 126438 6 io_in[6]
port 99 nsew signal input
rlabel metal3 s 291760 131282 292480 131402 6 io_out[6]
port 100 nsew signal tristate
rlabel metal3 s 291760 156034 292480 156154 6 io_in[7]
port 101 nsew signal input
rlabel metal3 s 291760 160998 292480 161118 6 io_out[7]
port 102 nsew signal tristate
rlabel metal3 s 291760 185818 292480 185938 6 io_in[8]
port 103 nsew signal input
rlabel metal3 s 291760 190782 292480 190902 6 io_out[8]
port 104 nsew signal tristate
rlabel metal3 s 291760 215534 292480 215654 6 io_in[9]
port 105 nsew signal input
rlabel metal3 s 291760 220498 292480 220618 6 io_out[9]
port 106 nsew signal tristate
rlabel metal3 s 291760 2422 292480 2542 6 io_in_3v3[0]
port 107 nsew signal input
rlabel metal3 s 291760 240354 292480 240474 6 io_in_3v3[10]
port 108 nsew signal input
rlabel metal3 s 291760 270070 292480 270190 6 io_in_3v3[11]
port 109 nsew signal input
rlabel metal3 s 291760 299854 292480 299974 6 io_in_3v3[12]
port 110 nsew signal input
rlabel metal3 s 291760 329570 292480 329690 6 io_in_3v3[13]
port 111 nsew signal input
rlabel metal3 s -480 326034 240 326154 4 io_in_3v3[14]
port 112 nsew signal input
rlabel metal3 s -480 297882 240 298002 4 io_in_3v3[15]
port 113 nsew signal input
rlabel metal3 s -480 269730 240 269850 4 io_in_3v3[16]
port 114 nsew signal input
rlabel metal3 s -480 241578 240 241698 4 io_in_3v3[17]
port 115 nsew signal input
rlabel metal3 s -480 213426 240 213546 4 io_in_3v3[18]
port 116 nsew signal input
rlabel metal3 s -480 185274 240 185394 4 io_in_3v3[19]
port 117 nsew signal input
rlabel metal3 s 291760 22210 292480 22330 6 io_in_3v3[1]
port 118 nsew signal input
rlabel metal3 s -480 157122 240 157242 4 io_in_3v3[20]
port 119 nsew signal input
rlabel metal3 s -480 128970 240 129090 4 io_in_3v3[21]
port 120 nsew signal input
rlabel metal3 s -480 100818 240 100938 4 io_in_3v3[22]
port 121 nsew signal input
rlabel metal3 s -480 72666 240 72786 4 io_in_3v3[23]
port 122 nsew signal input
rlabel metal3 s -480 53898 240 54018 4 io_in_3v3[24]
port 123 nsew signal input
rlabel metal3 s -480 35130 240 35250 4 io_in_3v3[25]
port 124 nsew signal input
rlabel metal3 s -480 16362 240 16482 4 io_in_3v3[26]
port 125 nsew signal input
rlabel metal3 s 291760 42066 292480 42186 6 io_in_3v3[2]
port 126 nsew signal input
rlabel metal3 s 291760 61854 292480 61974 6 io_in_3v3[3]
port 127 nsew signal input
rlabel metal3 s 291760 81710 292480 81830 6 io_in_3v3[4]
port 128 nsew signal input
rlabel metal3 s 291760 101566 292480 101686 6 io_in_3v3[5]
port 129 nsew signal input
rlabel metal3 s 291760 121354 292480 121474 6 io_in_3v3[6]
port 130 nsew signal input
rlabel metal3 s 291760 151138 292480 151258 6 io_in_3v3[7]
port 131 nsew signal input
rlabel metal3 s 291760 180854 292480 180974 6 io_in_3v3[8]
port 132 nsew signal input
rlabel metal3 s 291760 210570 292480 210690 6 io_in_3v3[9]
port 133 nsew signal input
rlabel metal3 s 291760 17246 292480 17366 6 io_oeb[0]
port 134 nsew signal tristate
rlabel metal3 s 291760 255178 292480 255298 6 io_oeb[10]
port 135 nsew signal tristate
rlabel metal3 s 291760 284962 292480 285082 6 io_oeb[11]
port 136 nsew signal tristate
rlabel metal3 s 291760 314678 292480 314798 6 io_oeb[12]
port 137 nsew signal tristate
rlabel metal3 s 291760 344462 292480 344582 6 io_oeb[13]
port 138 nsew signal tristate
rlabel metal3 s -480 311958 240 312078 4 io_oeb[14]
port 139 nsew signal tristate
rlabel metal3 s -480 283806 240 283926 4 io_oeb[15]
port 140 nsew signal tristate
rlabel metal3 s -480 255654 240 255774 4 io_oeb[16]
port 141 nsew signal tristate
rlabel metal3 s -480 227502 240 227622 4 io_oeb[17]
port 142 nsew signal tristate
rlabel metal3 s -480 199350 240 199470 4 io_oeb[18]
port 143 nsew signal tristate
rlabel metal3 s -480 171198 240 171318 4 io_oeb[19]
port 144 nsew signal tristate
rlabel metal3 s 291760 37102 292480 37222 6 io_oeb[1]
port 145 nsew signal tristate
rlabel metal3 s -480 143046 240 143166 4 io_oeb[20]
port 146 nsew signal tristate
rlabel metal3 s -480 114894 240 115014 4 io_oeb[21]
port 147 nsew signal tristate
rlabel metal3 s -480 86742 240 86862 4 io_oeb[22]
port 148 nsew signal tristate
rlabel metal3 s -480 58590 240 58710 4 io_oeb[23]
port 149 nsew signal tristate
rlabel metal3 s -480 39822 240 39942 4 io_oeb[24]
port 150 nsew signal tristate
rlabel metal3 s -480 21054 240 21174 4 io_oeb[25]
port 151 nsew signal tristate
rlabel metal3 s -480 2286 240 2406 4 io_oeb[26]
port 152 nsew signal tristate
rlabel metal3 s 291760 56890 292480 57010 6 io_oeb[2]
port 153 nsew signal tristate
rlabel metal3 s 291760 76746 292480 76866 6 io_oeb[3]
port 154 nsew signal tristate
rlabel metal3 s 291760 96602 292480 96722 6 io_oeb[4]
port 155 nsew signal tristate
rlabel metal3 s 291760 116390 292480 116510 6 io_oeb[5]
port 156 nsew signal tristate
rlabel metal3 s 291760 136246 292480 136366 6 io_oeb[6]
port 157 nsew signal tristate
rlabel metal3 s 291760 165962 292480 166082 6 io_oeb[7]
port 158 nsew signal tristate
rlabel metal3 s 291760 195746 292480 195866 6 io_oeb[8]
port 159 nsew signal tristate
rlabel metal3 s 291760 225462 292480 225582 6 io_oeb[9]
port 160 nsew signal tristate
rlabel metal2 s 62923 -480 62979 240 8 la_data_in[0]
port 161 nsew signal input
rlabel metal2 s 240253 -480 240309 240 8 la_data_in[100]
port 162 nsew signal input
rlabel metal2 s 242001 -480 242057 240 8 la_data_in[101]
port 163 nsew signal input
rlabel metal2 s 243795 -480 243851 240 8 la_data_in[102]
port 164 nsew signal input
rlabel metal2 s 245543 -480 245599 240 8 la_data_in[103]
port 165 nsew signal input
rlabel metal2 s 247337 -480 247393 240 8 la_data_in[104]
port 166 nsew signal input
rlabel metal2 s 249085 -480 249141 240 8 la_data_in[105]
port 167 nsew signal input
rlabel metal2 s 250879 -480 250935 240 8 la_data_in[106]
port 168 nsew signal input
rlabel metal2 s 252673 -480 252729 240 8 la_data_in[107]
port 169 nsew signal input
rlabel metal2 s 254421 -480 254477 240 8 la_data_in[108]
port 170 nsew signal input
rlabel metal2 s 256215 -480 256271 240 8 la_data_in[109]
port 171 nsew signal input
rlabel metal2 s 80633 -480 80689 240 8 la_data_in[10]
port 172 nsew signal input
rlabel metal2 s 257963 -480 258019 240 8 la_data_in[110]
port 173 nsew signal input
rlabel metal2 s 259757 -480 259813 240 8 la_data_in[111]
port 174 nsew signal input
rlabel metal2 s 261505 -480 261561 240 8 la_data_in[112]
port 175 nsew signal input
rlabel metal2 s 263299 -480 263355 240 8 la_data_in[113]
port 176 nsew signal input
rlabel metal2 s 265047 -480 265103 240 8 la_data_in[114]
port 177 nsew signal input
rlabel metal2 s 266841 -480 266897 240 8 la_data_in[115]
port 178 nsew signal input
rlabel metal2 s 268589 -480 268645 240 8 la_data_in[116]
port 179 nsew signal input
rlabel metal2 s 270383 -480 270439 240 8 la_data_in[117]
port 180 nsew signal input
rlabel metal2 s 272177 -480 272233 240 8 la_data_in[118]
port 181 nsew signal input
rlabel metal2 s 273925 -480 273981 240 8 la_data_in[119]
port 182 nsew signal input
rlabel metal2 s 82427 -480 82483 240 8 la_data_in[11]
port 183 nsew signal input
rlabel metal2 s 275719 -480 275775 240 8 la_data_in[120]
port 184 nsew signal input
rlabel metal2 s 277467 -480 277523 240 8 la_data_in[121]
port 185 nsew signal input
rlabel metal2 s 279261 -480 279317 240 8 la_data_in[122]
port 186 nsew signal input
rlabel metal2 s 281009 -480 281065 240 8 la_data_in[123]
port 187 nsew signal input
rlabel metal2 s 282803 -480 282859 240 8 la_data_in[124]
port 188 nsew signal input
rlabel metal2 s 284551 -480 284607 240 8 la_data_in[125]
port 189 nsew signal input
rlabel metal2 s 286345 -480 286401 240 8 la_data_in[126]
port 190 nsew signal input
rlabel metal2 s 288139 -480 288195 240 8 la_data_in[127]
port 191 nsew signal input
rlabel metal2 s 84175 -480 84231 240 8 la_data_in[12]
port 192 nsew signal input
rlabel metal2 s 85969 -480 86025 240 8 la_data_in[13]
port 193 nsew signal input
rlabel metal2 s 87717 -480 87773 240 8 la_data_in[14]
port 194 nsew signal input
rlabel metal2 s 89511 -480 89567 240 8 la_data_in[15]
port 195 nsew signal input
rlabel metal2 s 91259 -480 91315 240 8 la_data_in[16]
port 196 nsew signal input
rlabel metal2 s 93053 -480 93109 240 8 la_data_in[17]
port 197 nsew signal input
rlabel metal2 s 94847 -480 94903 240 8 la_data_in[18]
port 198 nsew signal input
rlabel metal2 s 96595 -480 96651 240 8 la_data_in[19]
port 199 nsew signal input
rlabel metal2 s 64671 -480 64727 240 8 la_data_in[1]
port 200 nsew signal input
rlabel metal2 s 98389 -480 98445 240 8 la_data_in[20]
port 201 nsew signal input
rlabel metal2 s 100137 -480 100193 240 8 la_data_in[21]
port 202 nsew signal input
rlabel metal2 s 101931 -480 101987 240 8 la_data_in[22]
port 203 nsew signal input
rlabel metal2 s 103679 -480 103735 240 8 la_data_in[23]
port 204 nsew signal input
rlabel metal2 s 105473 -480 105529 240 8 la_data_in[24]
port 205 nsew signal input
rlabel metal2 s 107221 -480 107277 240 8 la_data_in[25]
port 206 nsew signal input
rlabel metal2 s 109015 -480 109071 240 8 la_data_in[26]
port 207 nsew signal input
rlabel metal2 s 110763 -480 110819 240 8 la_data_in[27]
port 208 nsew signal input
rlabel metal2 s 112557 -480 112613 240 8 la_data_in[28]
port 209 nsew signal input
rlabel metal2 s 114351 -480 114407 240 8 la_data_in[29]
port 210 nsew signal input
rlabel metal2 s 66465 -480 66521 240 8 la_data_in[2]
port 211 nsew signal input
rlabel metal2 s 116099 -480 116155 240 8 la_data_in[30]
port 212 nsew signal input
rlabel metal2 s 117893 -480 117949 240 8 la_data_in[31]
port 213 nsew signal input
rlabel metal2 s 119641 -480 119697 240 8 la_data_in[32]
port 214 nsew signal input
rlabel metal2 s 121435 -480 121491 240 8 la_data_in[33]
port 215 nsew signal input
rlabel metal2 s 123183 -480 123239 240 8 la_data_in[34]
port 216 nsew signal input
rlabel metal2 s 124977 -480 125033 240 8 la_data_in[35]
port 217 nsew signal input
rlabel metal2 s 126725 -480 126781 240 8 la_data_in[36]
port 218 nsew signal input
rlabel metal2 s 128519 -480 128575 240 8 la_data_in[37]
port 219 nsew signal input
rlabel metal2 s 130313 -480 130369 240 8 la_data_in[38]
port 220 nsew signal input
rlabel metal2 s 132061 -480 132117 240 8 la_data_in[39]
port 221 nsew signal input
rlabel metal2 s 68213 -480 68269 240 8 la_data_in[3]
port 222 nsew signal input
rlabel metal2 s 133855 -480 133911 240 8 la_data_in[40]
port 223 nsew signal input
rlabel metal2 s 135603 -480 135659 240 8 la_data_in[41]
port 224 nsew signal input
rlabel metal2 s 137397 -480 137453 240 8 la_data_in[42]
port 225 nsew signal input
rlabel metal2 s 139145 -480 139201 240 8 la_data_in[43]
port 226 nsew signal input
rlabel metal2 s 140939 -480 140995 240 8 la_data_in[44]
port 227 nsew signal input
rlabel metal2 s 142687 -480 142743 240 8 la_data_in[45]
port 228 nsew signal input
rlabel metal2 s 144481 -480 144537 240 8 la_data_in[46]
port 229 nsew signal input
rlabel metal2 s 146275 -480 146331 240 8 la_data_in[47]
port 230 nsew signal input
rlabel metal2 s 148023 -480 148079 240 8 la_data_in[48]
port 231 nsew signal input
rlabel metal2 s 149817 -480 149873 240 8 la_data_in[49]
port 232 nsew signal input
rlabel metal2 s 70007 -480 70063 240 8 la_data_in[4]
port 233 nsew signal input
rlabel metal2 s 151565 -480 151621 240 8 la_data_in[50]
port 234 nsew signal input
rlabel metal2 s 153359 -480 153415 240 8 la_data_in[51]
port 235 nsew signal input
rlabel metal2 s 155107 -480 155163 240 8 la_data_in[52]
port 236 nsew signal input
rlabel metal2 s 156901 -480 156957 240 8 la_data_in[53]
port 237 nsew signal input
rlabel metal2 s 158649 -480 158705 240 8 la_data_in[54]
port 238 nsew signal input
rlabel metal2 s 160443 -480 160499 240 8 la_data_in[55]
port 239 nsew signal input
rlabel metal2 s 162191 -480 162247 240 8 la_data_in[56]
port 240 nsew signal input
rlabel metal2 s 163985 -480 164041 240 8 la_data_in[57]
port 241 nsew signal input
rlabel metal2 s 165779 -480 165835 240 8 la_data_in[58]
port 242 nsew signal input
rlabel metal2 s 167527 -480 167583 240 8 la_data_in[59]
port 243 nsew signal input
rlabel metal2 s 71755 -480 71811 240 8 la_data_in[5]
port 244 nsew signal input
rlabel metal2 s 169321 -480 169377 240 8 la_data_in[60]
port 245 nsew signal input
rlabel metal2 s 171069 -480 171125 240 8 la_data_in[61]
port 246 nsew signal input
rlabel metal2 s 172863 -480 172919 240 8 la_data_in[62]
port 247 nsew signal input
rlabel metal2 s 174611 -480 174667 240 8 la_data_in[63]
port 248 nsew signal input
rlabel metal2 s 176405 -480 176461 240 8 la_data_in[64]
port 249 nsew signal input
rlabel metal2 s 178153 -480 178209 240 8 la_data_in[65]
port 250 nsew signal input
rlabel metal2 s 179947 -480 180003 240 8 la_data_in[66]
port 251 nsew signal input
rlabel metal2 s 181741 -480 181797 240 8 la_data_in[67]
port 252 nsew signal input
rlabel metal2 s 183489 -480 183545 240 8 la_data_in[68]
port 253 nsew signal input
rlabel metal2 s 185283 -480 185339 240 8 la_data_in[69]
port 254 nsew signal input
rlabel metal2 s 73549 -480 73605 240 8 la_data_in[6]
port 255 nsew signal input
rlabel metal2 s 187031 -480 187087 240 8 la_data_in[70]
port 256 nsew signal input
rlabel metal2 s 188825 -480 188881 240 8 la_data_in[71]
port 257 nsew signal input
rlabel metal2 s 190573 -480 190629 240 8 la_data_in[72]
port 258 nsew signal input
rlabel metal2 s 192367 -480 192423 240 8 la_data_in[73]
port 259 nsew signal input
rlabel metal2 s 194115 -480 194171 240 8 la_data_in[74]
port 260 nsew signal input
rlabel metal2 s 195909 -480 195965 240 8 la_data_in[75]
port 261 nsew signal input
rlabel metal2 s 197657 -480 197713 240 8 la_data_in[76]
port 262 nsew signal input
rlabel metal2 s 199451 -480 199507 240 8 la_data_in[77]
port 263 nsew signal input
rlabel metal2 s 201245 -480 201301 240 8 la_data_in[78]
port 264 nsew signal input
rlabel metal2 s 202993 -480 203049 240 8 la_data_in[79]
port 265 nsew signal input
rlabel metal2 s 75297 -480 75353 240 8 la_data_in[7]
port 266 nsew signal input
rlabel metal2 s 204787 -480 204843 240 8 la_data_in[80]
port 267 nsew signal input
rlabel metal2 s 206535 -480 206591 240 8 la_data_in[81]
port 268 nsew signal input
rlabel metal2 s 208329 -480 208385 240 8 la_data_in[82]
port 269 nsew signal input
rlabel metal2 s 210077 -480 210133 240 8 la_data_in[83]
port 270 nsew signal input
rlabel metal2 s 211871 -480 211927 240 8 la_data_in[84]
port 271 nsew signal input
rlabel metal2 s 213619 -480 213675 240 8 la_data_in[85]
port 272 nsew signal input
rlabel metal2 s 215413 -480 215469 240 8 la_data_in[86]
port 273 nsew signal input
rlabel metal2 s 217207 -480 217263 240 8 la_data_in[87]
port 274 nsew signal input
rlabel metal2 s 218955 -480 219011 240 8 la_data_in[88]
port 275 nsew signal input
rlabel metal2 s 220749 -480 220805 240 8 la_data_in[89]
port 276 nsew signal input
rlabel metal2 s 77091 -480 77147 240 8 la_data_in[8]
port 277 nsew signal input
rlabel metal2 s 222497 -480 222553 240 8 la_data_in[90]
port 278 nsew signal input
rlabel metal2 s 224291 -480 224347 240 8 la_data_in[91]
port 279 nsew signal input
rlabel metal2 s 226039 -480 226095 240 8 la_data_in[92]
port 280 nsew signal input
rlabel metal2 s 227833 -480 227889 240 8 la_data_in[93]
port 281 nsew signal input
rlabel metal2 s 229581 -480 229637 240 8 la_data_in[94]
port 282 nsew signal input
rlabel metal2 s 231375 -480 231431 240 8 la_data_in[95]
port 283 nsew signal input
rlabel metal2 s 233123 -480 233179 240 8 la_data_in[96]
port 284 nsew signal input
rlabel metal2 s 234917 -480 234973 240 8 la_data_in[97]
port 285 nsew signal input
rlabel metal2 s 236711 -480 236767 240 8 la_data_in[98]
port 286 nsew signal input
rlabel metal2 s 238459 -480 238515 240 8 la_data_in[99]
port 287 nsew signal input
rlabel metal2 s 78885 -480 78941 240 8 la_data_in[9]
port 288 nsew signal input
rlabel metal2 s 63475 -480 63531 240 8 la_data_out[0]
port 289 nsew signal tristate
rlabel metal2 s 240851 -480 240907 240 8 la_data_out[100]
port 290 nsew signal tristate
rlabel metal2 s 242599 -480 242655 240 8 la_data_out[101]
port 291 nsew signal tristate
rlabel metal2 s 244393 -480 244449 240 8 la_data_out[102]
port 292 nsew signal tristate
rlabel metal2 s 246141 -480 246197 240 8 la_data_out[103]
port 293 nsew signal tristate
rlabel metal2 s 247935 -480 247991 240 8 la_data_out[104]
port 294 nsew signal tristate
rlabel metal2 s 249683 -480 249739 240 8 la_data_out[105]
port 295 nsew signal tristate
rlabel metal2 s 251477 -480 251533 240 8 la_data_out[106]
port 296 nsew signal tristate
rlabel metal2 s 253225 -480 253281 240 8 la_data_out[107]
port 297 nsew signal tristate
rlabel metal2 s 255019 -480 255075 240 8 la_data_out[108]
port 298 nsew signal tristate
rlabel metal2 s 256767 -480 256823 240 8 la_data_out[109]
port 299 nsew signal tristate
rlabel metal2 s 81231 -480 81287 240 8 la_data_out[10]
port 300 nsew signal tristate
rlabel metal2 s 258561 -480 258617 240 8 la_data_out[110]
port 301 nsew signal tristate
rlabel metal2 s 260355 -480 260411 240 8 la_data_out[111]
port 302 nsew signal tristate
rlabel metal2 s 262103 -480 262159 240 8 la_data_out[112]
port 303 nsew signal tristate
rlabel metal2 s 263897 -480 263953 240 8 la_data_out[113]
port 304 nsew signal tristate
rlabel metal2 s 265645 -480 265701 240 8 la_data_out[114]
port 305 nsew signal tristate
rlabel metal2 s 267439 -480 267495 240 8 la_data_out[115]
port 306 nsew signal tristate
rlabel metal2 s 269187 -480 269243 240 8 la_data_out[116]
port 307 nsew signal tristate
rlabel metal2 s 270981 -480 271037 240 8 la_data_out[117]
port 308 nsew signal tristate
rlabel metal2 s 272729 -480 272785 240 8 la_data_out[118]
port 309 nsew signal tristate
rlabel metal2 s 274523 -480 274579 240 8 la_data_out[119]
port 310 nsew signal tristate
rlabel metal2 s 83025 -480 83081 240 8 la_data_out[11]
port 311 nsew signal tristate
rlabel metal2 s 276317 -480 276373 240 8 la_data_out[120]
port 312 nsew signal tristate
rlabel metal2 s 278065 -480 278121 240 8 la_data_out[121]
port 313 nsew signal tristate
rlabel metal2 s 279859 -480 279915 240 8 la_data_out[122]
port 314 nsew signal tristate
rlabel metal2 s 281607 -480 281663 240 8 la_data_out[123]
port 315 nsew signal tristate
rlabel metal2 s 283401 -480 283457 240 8 la_data_out[124]
port 316 nsew signal tristate
rlabel metal2 s 285149 -480 285205 240 8 la_data_out[125]
port 317 nsew signal tristate
rlabel metal2 s 286943 -480 286999 240 8 la_data_out[126]
port 318 nsew signal tristate
rlabel metal2 s 288691 -480 288747 240 8 la_data_out[127]
port 319 nsew signal tristate
rlabel metal2 s 84773 -480 84829 240 8 la_data_out[12]
port 320 nsew signal tristate
rlabel metal2 s 86567 -480 86623 240 8 la_data_out[13]
port 321 nsew signal tristate
rlabel metal2 s 88315 -480 88371 240 8 la_data_out[14]
port 322 nsew signal tristate
rlabel metal2 s 90109 -480 90165 240 8 la_data_out[15]
port 323 nsew signal tristate
rlabel metal2 s 91857 -480 91913 240 8 la_data_out[16]
port 324 nsew signal tristate
rlabel metal2 s 93651 -480 93707 240 8 la_data_out[17]
port 325 nsew signal tristate
rlabel metal2 s 95399 -480 95455 240 8 la_data_out[18]
port 326 nsew signal tristate
rlabel metal2 s 97193 -480 97249 240 8 la_data_out[19]
port 327 nsew signal tristate
rlabel metal2 s 65269 -480 65325 240 8 la_data_out[1]
port 328 nsew signal tristate
rlabel metal2 s 98941 -480 98997 240 8 la_data_out[20]
port 329 nsew signal tristate
rlabel metal2 s 100735 -480 100791 240 8 la_data_out[21]
port 330 nsew signal tristate
rlabel metal2 s 102529 -480 102585 240 8 la_data_out[22]
port 331 nsew signal tristate
rlabel metal2 s 104277 -480 104333 240 8 la_data_out[23]
port 332 nsew signal tristate
rlabel metal2 s 106071 -480 106127 240 8 la_data_out[24]
port 333 nsew signal tristate
rlabel metal2 s 107819 -480 107875 240 8 la_data_out[25]
port 334 nsew signal tristate
rlabel metal2 s 109613 -480 109669 240 8 la_data_out[26]
port 335 nsew signal tristate
rlabel metal2 s 111361 -480 111417 240 8 la_data_out[27]
port 336 nsew signal tristate
rlabel metal2 s 113155 -480 113211 240 8 la_data_out[28]
port 337 nsew signal tristate
rlabel metal2 s 114903 -480 114959 240 8 la_data_out[29]
port 338 nsew signal tristate
rlabel metal2 s 67063 -480 67119 240 8 la_data_out[2]
port 339 nsew signal tristate
rlabel metal2 s 116697 -480 116753 240 8 la_data_out[30]
port 340 nsew signal tristate
rlabel metal2 s 118491 -480 118547 240 8 la_data_out[31]
port 341 nsew signal tristate
rlabel metal2 s 120239 -480 120295 240 8 la_data_out[32]
port 342 nsew signal tristate
rlabel metal2 s 122033 -480 122089 240 8 la_data_out[33]
port 343 nsew signal tristate
rlabel metal2 s 123781 -480 123837 240 8 la_data_out[34]
port 344 nsew signal tristate
rlabel metal2 s 125575 -480 125631 240 8 la_data_out[35]
port 345 nsew signal tristate
rlabel metal2 s 127323 -480 127379 240 8 la_data_out[36]
port 346 nsew signal tristate
rlabel metal2 s 129117 -480 129173 240 8 la_data_out[37]
port 347 nsew signal tristate
rlabel metal2 s 130865 -480 130921 240 8 la_data_out[38]
port 348 nsew signal tristate
rlabel metal2 s 132659 -480 132715 240 8 la_data_out[39]
port 349 nsew signal tristate
rlabel metal2 s 68811 -480 68867 240 8 la_data_out[3]
port 350 nsew signal tristate
rlabel metal2 s 134407 -480 134463 240 8 la_data_out[40]
port 351 nsew signal tristate
rlabel metal2 s 136201 -480 136257 240 8 la_data_out[41]
port 352 nsew signal tristate
rlabel metal2 s 137995 -480 138051 240 8 la_data_out[42]
port 353 nsew signal tristate
rlabel metal2 s 139743 -480 139799 240 8 la_data_out[43]
port 354 nsew signal tristate
rlabel metal2 s 141537 -480 141593 240 8 la_data_out[44]
port 355 nsew signal tristate
rlabel metal2 s 143285 -480 143341 240 8 la_data_out[45]
port 356 nsew signal tristate
rlabel metal2 s 145079 -480 145135 240 8 la_data_out[46]
port 357 nsew signal tristate
rlabel metal2 s 146827 -480 146883 240 8 la_data_out[47]
port 358 nsew signal tristate
rlabel metal2 s 148621 -480 148677 240 8 la_data_out[48]
port 359 nsew signal tristate
rlabel metal2 s 150369 -480 150425 240 8 la_data_out[49]
port 360 nsew signal tristate
rlabel metal2 s 70605 -480 70661 240 8 la_data_out[4]
port 361 nsew signal tristate
rlabel metal2 s 152163 -480 152219 240 8 la_data_out[50]
port 362 nsew signal tristate
rlabel metal2 s 153957 -480 154013 240 8 la_data_out[51]
port 363 nsew signal tristate
rlabel metal2 s 155705 -480 155761 240 8 la_data_out[52]
port 364 nsew signal tristate
rlabel metal2 s 157499 -480 157555 240 8 la_data_out[53]
port 365 nsew signal tristate
rlabel metal2 s 159247 -480 159303 240 8 la_data_out[54]
port 366 nsew signal tristate
rlabel metal2 s 161041 -480 161097 240 8 la_data_out[55]
port 367 nsew signal tristate
rlabel metal2 s 162789 -480 162845 240 8 la_data_out[56]
port 368 nsew signal tristate
rlabel metal2 s 164583 -480 164639 240 8 la_data_out[57]
port 369 nsew signal tristate
rlabel metal2 s 166331 -480 166387 240 8 la_data_out[58]
port 370 nsew signal tristate
rlabel metal2 s 168125 -480 168181 240 8 la_data_out[59]
port 371 nsew signal tristate
rlabel metal2 s 72353 -480 72409 240 8 la_data_out[5]
port 372 nsew signal tristate
rlabel metal2 s 169919 -480 169975 240 8 la_data_out[60]
port 373 nsew signal tristate
rlabel metal2 s 171667 -480 171723 240 8 la_data_out[61]
port 374 nsew signal tristate
rlabel metal2 s 173461 -480 173517 240 8 la_data_out[62]
port 375 nsew signal tristate
rlabel metal2 s 175209 -480 175265 240 8 la_data_out[63]
port 376 nsew signal tristate
rlabel metal2 s 177003 -480 177059 240 8 la_data_out[64]
port 377 nsew signal tristate
rlabel metal2 s 178751 -480 178807 240 8 la_data_out[65]
port 378 nsew signal tristate
rlabel metal2 s 180545 -480 180601 240 8 la_data_out[66]
port 379 nsew signal tristate
rlabel metal2 s 182293 -480 182349 240 8 la_data_out[67]
port 380 nsew signal tristate
rlabel metal2 s 184087 -480 184143 240 8 la_data_out[68]
port 381 nsew signal tristate
rlabel metal2 s 185835 -480 185891 240 8 la_data_out[69]
port 382 nsew signal tristate
rlabel metal2 s 74147 -480 74203 240 8 la_data_out[6]
port 383 nsew signal tristate
rlabel metal2 s 187629 -480 187685 240 8 la_data_out[70]
port 384 nsew signal tristate
rlabel metal2 s 189423 -480 189479 240 8 la_data_out[71]
port 385 nsew signal tristate
rlabel metal2 s 191171 -480 191227 240 8 la_data_out[72]
port 386 nsew signal tristate
rlabel metal2 s 192965 -480 193021 240 8 la_data_out[73]
port 387 nsew signal tristate
rlabel metal2 s 194713 -480 194769 240 8 la_data_out[74]
port 388 nsew signal tristate
rlabel metal2 s 196507 -480 196563 240 8 la_data_out[75]
port 389 nsew signal tristate
rlabel metal2 s 198255 -480 198311 240 8 la_data_out[76]
port 390 nsew signal tristate
rlabel metal2 s 200049 -480 200105 240 8 la_data_out[77]
port 391 nsew signal tristate
rlabel metal2 s 201797 -480 201853 240 8 la_data_out[78]
port 392 nsew signal tristate
rlabel metal2 s 203591 -480 203647 240 8 la_data_out[79]
port 393 nsew signal tristate
rlabel metal2 s 75895 -480 75951 240 8 la_data_out[7]
port 394 nsew signal tristate
rlabel metal2 s 205385 -480 205441 240 8 la_data_out[80]
port 395 nsew signal tristate
rlabel metal2 s 207133 -480 207189 240 8 la_data_out[81]
port 396 nsew signal tristate
rlabel metal2 s 208927 -480 208983 240 8 la_data_out[82]
port 397 nsew signal tristate
rlabel metal2 s 210675 -480 210731 240 8 la_data_out[83]
port 398 nsew signal tristate
rlabel metal2 s 212469 -480 212525 240 8 la_data_out[84]
port 399 nsew signal tristate
rlabel metal2 s 214217 -480 214273 240 8 la_data_out[85]
port 400 nsew signal tristate
rlabel metal2 s 216011 -480 216067 240 8 la_data_out[86]
port 401 nsew signal tristate
rlabel metal2 s 217759 -480 217815 240 8 la_data_out[87]
port 402 nsew signal tristate
rlabel metal2 s 219553 -480 219609 240 8 la_data_out[88]
port 403 nsew signal tristate
rlabel metal2 s 221301 -480 221357 240 8 la_data_out[89]
port 404 nsew signal tristate
rlabel metal2 s 77689 -480 77745 240 8 la_data_out[8]
port 405 nsew signal tristate
rlabel metal2 s 223095 -480 223151 240 8 la_data_out[90]
port 406 nsew signal tristate
rlabel metal2 s 224889 -480 224945 240 8 la_data_out[91]
port 407 nsew signal tristate
rlabel metal2 s 226637 -480 226693 240 8 la_data_out[92]
port 408 nsew signal tristate
rlabel metal2 s 228431 -480 228487 240 8 la_data_out[93]
port 409 nsew signal tristate
rlabel metal2 s 230179 -480 230235 240 8 la_data_out[94]
port 410 nsew signal tristate
rlabel metal2 s 231973 -480 232029 240 8 la_data_out[95]
port 411 nsew signal tristate
rlabel metal2 s 233721 -480 233777 240 8 la_data_out[96]
port 412 nsew signal tristate
rlabel metal2 s 235515 -480 235571 240 8 la_data_out[97]
port 413 nsew signal tristate
rlabel metal2 s 237263 -480 237319 240 8 la_data_out[98]
port 414 nsew signal tristate
rlabel metal2 s 239057 -480 239113 240 8 la_data_out[99]
port 415 nsew signal tristate
rlabel metal2 s 79437 -480 79493 240 8 la_data_out[9]
port 416 nsew signal tristate
rlabel metal2 s 64073 -480 64129 240 8 la_oenb[0]
port 417 nsew signal input
rlabel metal2 s 241403 -480 241459 240 8 la_oenb[100]
port 418 nsew signal input
rlabel metal2 s 243197 -480 243253 240 8 la_oenb[101]
port 419 nsew signal input
rlabel metal2 s 244945 -480 245001 240 8 la_oenb[102]
port 420 nsew signal input
rlabel metal2 s 246739 -480 246795 240 8 la_oenb[103]
port 421 nsew signal input
rlabel metal2 s 248533 -480 248589 240 8 la_oenb[104]
port 422 nsew signal input
rlabel metal2 s 250281 -480 250337 240 8 la_oenb[105]
port 423 nsew signal input
rlabel metal2 s 252075 -480 252131 240 8 la_oenb[106]
port 424 nsew signal input
rlabel metal2 s 253823 -480 253879 240 8 la_oenb[107]
port 425 nsew signal input
rlabel metal2 s 255617 -480 255673 240 8 la_oenb[108]
port 426 nsew signal input
rlabel metal2 s 257365 -480 257421 240 8 la_oenb[109]
port 427 nsew signal input
rlabel metal2 s 81829 -480 81885 240 8 la_oenb[10]
port 428 nsew signal input
rlabel metal2 s 259159 -480 259215 240 8 la_oenb[110]
port 429 nsew signal input
rlabel metal2 s 260907 -480 260963 240 8 la_oenb[111]
port 430 nsew signal input
rlabel metal2 s 262701 -480 262757 240 8 la_oenb[112]
port 431 nsew signal input
rlabel metal2 s 264495 -480 264551 240 8 la_oenb[113]
port 432 nsew signal input
rlabel metal2 s 266243 -480 266299 240 8 la_oenb[114]
port 433 nsew signal input
rlabel metal2 s 268037 -480 268093 240 8 la_oenb[115]
port 434 nsew signal input
rlabel metal2 s 269785 -480 269841 240 8 la_oenb[116]
port 435 nsew signal input
rlabel metal2 s 271579 -480 271635 240 8 la_oenb[117]
port 436 nsew signal input
rlabel metal2 s 273327 -480 273383 240 8 la_oenb[118]
port 437 nsew signal input
rlabel metal2 s 275121 -480 275177 240 8 la_oenb[119]
port 438 nsew signal input
rlabel metal2 s 83577 -480 83633 240 8 la_oenb[11]
port 439 nsew signal input
rlabel metal2 s 276869 -480 276925 240 8 la_oenb[120]
port 440 nsew signal input
rlabel metal2 s 278663 -480 278719 240 8 la_oenb[121]
port 441 nsew signal input
rlabel metal2 s 280411 -480 280467 240 8 la_oenb[122]
port 442 nsew signal input
rlabel metal2 s 282205 -480 282261 240 8 la_oenb[123]
port 443 nsew signal input
rlabel metal2 s 283999 -480 284055 240 8 la_oenb[124]
port 444 nsew signal input
rlabel metal2 s 285747 -480 285803 240 8 la_oenb[125]
port 445 nsew signal input
rlabel metal2 s 287541 -480 287597 240 8 la_oenb[126]
port 446 nsew signal input
rlabel metal2 s 289289 -480 289345 240 8 la_oenb[127]
port 447 nsew signal input
rlabel metal2 s 85371 -480 85427 240 8 la_oenb[12]
port 448 nsew signal input
rlabel metal2 s 87119 -480 87175 240 8 la_oenb[13]
port 449 nsew signal input
rlabel metal2 s 88913 -480 88969 240 8 la_oenb[14]
port 450 nsew signal input
rlabel metal2 s 90707 -480 90763 240 8 la_oenb[15]
port 451 nsew signal input
rlabel metal2 s 92455 -480 92511 240 8 la_oenb[16]
port 452 nsew signal input
rlabel metal2 s 94249 -480 94305 240 8 la_oenb[17]
port 453 nsew signal input
rlabel metal2 s 95997 -480 96053 240 8 la_oenb[18]
port 454 nsew signal input
rlabel metal2 s 97791 -480 97847 240 8 la_oenb[19]
port 455 nsew signal input
rlabel metal2 s 65867 -480 65923 240 8 la_oenb[1]
port 456 nsew signal input
rlabel metal2 s 99539 -480 99595 240 8 la_oenb[20]
port 457 nsew signal input
rlabel metal2 s 101333 -480 101389 240 8 la_oenb[21]
port 458 nsew signal input
rlabel metal2 s 103081 -480 103137 240 8 la_oenb[22]
port 459 nsew signal input
rlabel metal2 s 104875 -480 104931 240 8 la_oenb[23]
port 460 nsew signal input
rlabel metal2 s 106669 -480 106725 240 8 la_oenb[24]
port 461 nsew signal input
rlabel metal2 s 108417 -480 108473 240 8 la_oenb[25]
port 462 nsew signal input
rlabel metal2 s 110211 -480 110267 240 8 la_oenb[26]
port 463 nsew signal input
rlabel metal2 s 111959 -480 112015 240 8 la_oenb[27]
port 464 nsew signal input
rlabel metal2 s 113753 -480 113809 240 8 la_oenb[28]
port 465 nsew signal input
rlabel metal2 s 115501 -480 115557 240 8 la_oenb[29]
port 466 nsew signal input
rlabel metal2 s 67615 -480 67671 240 8 la_oenb[2]
port 467 nsew signal input
rlabel metal2 s 117295 -480 117351 240 8 la_oenb[30]
port 468 nsew signal input
rlabel metal2 s 119043 -480 119099 240 8 la_oenb[31]
port 469 nsew signal input
rlabel metal2 s 120837 -480 120893 240 8 la_oenb[32]
port 470 nsew signal input
rlabel metal2 s 122585 -480 122641 240 8 la_oenb[33]
port 471 nsew signal input
rlabel metal2 s 124379 -480 124435 240 8 la_oenb[34]
port 472 nsew signal input
rlabel metal2 s 126173 -480 126229 240 8 la_oenb[35]
port 473 nsew signal input
rlabel metal2 s 127921 -480 127977 240 8 la_oenb[36]
port 474 nsew signal input
rlabel metal2 s 129715 -480 129771 240 8 la_oenb[37]
port 475 nsew signal input
rlabel metal2 s 131463 -480 131519 240 8 la_oenb[38]
port 476 nsew signal input
rlabel metal2 s 133257 -480 133313 240 8 la_oenb[39]
port 477 nsew signal input
rlabel metal2 s 69409 -480 69465 240 8 la_oenb[3]
port 478 nsew signal input
rlabel metal2 s 135005 -480 135061 240 8 la_oenb[40]
port 479 nsew signal input
rlabel metal2 s 136799 -480 136855 240 8 la_oenb[41]
port 480 nsew signal input
rlabel metal2 s 138547 -480 138603 240 8 la_oenb[42]
port 481 nsew signal input
rlabel metal2 s 140341 -480 140397 240 8 la_oenb[43]
port 482 nsew signal input
rlabel metal2 s 142135 -480 142191 240 8 la_oenb[44]
port 483 nsew signal input
rlabel metal2 s 143883 -480 143939 240 8 la_oenb[45]
port 484 nsew signal input
rlabel metal2 s 145677 -480 145733 240 8 la_oenb[46]
port 485 nsew signal input
rlabel metal2 s 147425 -480 147481 240 8 la_oenb[47]
port 486 nsew signal input
rlabel metal2 s 149219 -480 149275 240 8 la_oenb[48]
port 487 nsew signal input
rlabel metal2 s 150967 -480 151023 240 8 la_oenb[49]
port 488 nsew signal input
rlabel metal2 s 71203 -480 71259 240 8 la_oenb[4]
port 489 nsew signal input
rlabel metal2 s 152761 -480 152817 240 8 la_oenb[50]
port 490 nsew signal input
rlabel metal2 s 154509 -480 154565 240 8 la_oenb[51]
port 491 nsew signal input
rlabel metal2 s 156303 -480 156359 240 8 la_oenb[52]
port 492 nsew signal input
rlabel metal2 s 158097 -480 158153 240 8 la_oenb[53]
port 493 nsew signal input
rlabel metal2 s 159845 -480 159901 240 8 la_oenb[54]
port 494 nsew signal input
rlabel metal2 s 161639 -480 161695 240 8 la_oenb[55]
port 495 nsew signal input
rlabel metal2 s 163387 -480 163443 240 8 la_oenb[56]
port 496 nsew signal input
rlabel metal2 s 165181 -480 165237 240 8 la_oenb[57]
port 497 nsew signal input
rlabel metal2 s 166929 -480 166985 240 8 la_oenb[58]
port 498 nsew signal input
rlabel metal2 s 168723 -480 168779 240 8 la_oenb[59]
port 499 nsew signal input
rlabel metal2 s 72951 -480 73007 240 8 la_oenb[5]
port 500 nsew signal input
rlabel metal2 s 170471 -480 170527 240 8 la_oenb[60]
port 501 nsew signal input
rlabel metal2 s 172265 -480 172321 240 8 la_oenb[61]
port 502 nsew signal input
rlabel metal2 s 174013 -480 174069 240 8 la_oenb[62]
port 503 nsew signal input
rlabel metal2 s 175807 -480 175863 240 8 la_oenb[63]
port 504 nsew signal input
rlabel metal2 s 177601 -480 177657 240 8 la_oenb[64]
port 505 nsew signal input
rlabel metal2 s 179349 -480 179405 240 8 la_oenb[65]
port 506 nsew signal input
rlabel metal2 s 181143 -480 181199 240 8 la_oenb[66]
port 507 nsew signal input
rlabel metal2 s 182891 -480 182947 240 8 la_oenb[67]
port 508 nsew signal input
rlabel metal2 s 184685 -480 184741 240 8 la_oenb[68]
port 509 nsew signal input
rlabel metal2 s 186433 -480 186489 240 8 la_oenb[69]
port 510 nsew signal input
rlabel metal2 s 74745 -480 74801 240 8 la_oenb[6]
port 511 nsew signal input
rlabel metal2 s 188227 -480 188283 240 8 la_oenb[70]
port 512 nsew signal input
rlabel metal2 s 189975 -480 190031 240 8 la_oenb[71]
port 513 nsew signal input
rlabel metal2 s 191769 -480 191825 240 8 la_oenb[72]
port 514 nsew signal input
rlabel metal2 s 193563 -480 193619 240 8 la_oenb[73]
port 515 nsew signal input
rlabel metal2 s 195311 -480 195367 240 8 la_oenb[74]
port 516 nsew signal input
rlabel metal2 s 197105 -480 197161 240 8 la_oenb[75]
port 517 nsew signal input
rlabel metal2 s 198853 -480 198909 240 8 la_oenb[76]
port 518 nsew signal input
rlabel metal2 s 200647 -480 200703 240 8 la_oenb[77]
port 519 nsew signal input
rlabel metal2 s 202395 -480 202451 240 8 la_oenb[78]
port 520 nsew signal input
rlabel metal2 s 204189 -480 204245 240 8 la_oenb[79]
port 521 nsew signal input
rlabel metal2 s 76493 -480 76549 240 8 la_oenb[7]
port 522 nsew signal input
rlabel metal2 s 205937 -480 205993 240 8 la_oenb[80]
port 523 nsew signal input
rlabel metal2 s 207731 -480 207787 240 8 la_oenb[81]
port 524 nsew signal input
rlabel metal2 s 209479 -480 209535 240 8 la_oenb[82]
port 525 nsew signal input
rlabel metal2 s 211273 -480 211329 240 8 la_oenb[83]
port 526 nsew signal input
rlabel metal2 s 213067 -480 213123 240 8 la_oenb[84]
port 527 nsew signal input
rlabel metal2 s 214815 -480 214871 240 8 la_oenb[85]
port 528 nsew signal input
rlabel metal2 s 216609 -480 216665 240 8 la_oenb[86]
port 529 nsew signal input
rlabel metal2 s 218357 -480 218413 240 8 la_oenb[87]
port 530 nsew signal input
rlabel metal2 s 220151 -480 220207 240 8 la_oenb[88]
port 531 nsew signal input
rlabel metal2 s 221899 -480 221955 240 8 la_oenb[89]
port 532 nsew signal input
rlabel metal2 s 78287 -480 78343 240 8 la_oenb[8]
port 533 nsew signal input
rlabel metal2 s 223693 -480 223749 240 8 la_oenb[90]
port 534 nsew signal input
rlabel metal2 s 225441 -480 225497 240 8 la_oenb[91]
port 535 nsew signal input
rlabel metal2 s 227235 -480 227291 240 8 la_oenb[92]
port 536 nsew signal input
rlabel metal2 s 229029 -480 229085 240 8 la_oenb[93]
port 537 nsew signal input
rlabel metal2 s 230777 -480 230833 240 8 la_oenb[94]
port 538 nsew signal input
rlabel metal2 s 232571 -480 232627 240 8 la_oenb[95]
port 539 nsew signal input
rlabel metal2 s 234319 -480 234375 240 8 la_oenb[96]
port 540 nsew signal input
rlabel metal2 s 236113 -480 236169 240 8 la_oenb[97]
port 541 nsew signal input
rlabel metal2 s 237861 -480 237917 240 8 la_oenb[98]
port 542 nsew signal input
rlabel metal2 s 239655 -480 239711 240 8 la_oenb[99]
port 543 nsew signal input
rlabel metal2 s 80035 -480 80091 240 8 la_oenb[9]
port 544 nsew signal input
rlabel metal2 s 289887 -480 289943 240 8 user_clock2
port 545 nsew signal input
rlabel metal2 s 290485 -480 290541 240 8 user_irq[0]
port 546 nsew signal tristate
rlabel metal2 s 291083 -480 291139 240 8 user_irq[1]
port 547 nsew signal tristate
rlabel metal2 s 291681 -480 291737 240 8 user_irq[2]
port 548 nsew signal tristate
rlabel metal2 s 271 -480 327 240 8 wb_clk_i
port 549 nsew signal input
rlabel metal2 s 823 -480 879 240 8 wb_rst_i
port 550 nsew signal input
rlabel metal2 s 1421 -480 1477 240 8 wbs_ack_o
port 551 nsew signal tristate
rlabel metal2 s 3813 -480 3869 240 8 wbs_adr_i[0]
port 552 nsew signal input
rlabel metal2 s 23915 -480 23971 240 8 wbs_adr_i[10]
port 553 nsew signal input
rlabel metal2 s 25663 -480 25719 240 8 wbs_adr_i[11]
port 554 nsew signal input
rlabel metal2 s 27457 -480 27513 240 8 wbs_adr_i[12]
port 555 nsew signal input
rlabel metal2 s 29205 -480 29261 240 8 wbs_adr_i[13]
port 556 nsew signal input
rlabel metal2 s 30999 -480 31055 240 8 wbs_adr_i[14]
port 557 nsew signal input
rlabel metal2 s 32747 -480 32803 240 8 wbs_adr_i[15]
port 558 nsew signal input
rlabel metal2 s 34541 -480 34597 240 8 wbs_adr_i[16]
port 559 nsew signal input
rlabel metal2 s 36289 -480 36345 240 8 wbs_adr_i[17]
port 560 nsew signal input
rlabel metal2 s 38083 -480 38139 240 8 wbs_adr_i[18]
port 561 nsew signal input
rlabel metal2 s 39831 -480 39887 240 8 wbs_adr_i[19]
port 562 nsew signal input
rlabel metal2 s 6159 -480 6215 240 8 wbs_adr_i[1]
port 563 nsew signal input
rlabel metal2 s 41625 -480 41681 240 8 wbs_adr_i[20]
port 564 nsew signal input
rlabel metal2 s 43419 -480 43475 240 8 wbs_adr_i[21]
port 565 nsew signal input
rlabel metal2 s 45167 -480 45223 240 8 wbs_adr_i[22]
port 566 nsew signal input
rlabel metal2 s 46961 -480 47017 240 8 wbs_adr_i[23]
port 567 nsew signal input
rlabel metal2 s 48709 -480 48765 240 8 wbs_adr_i[24]
port 568 nsew signal input
rlabel metal2 s 50503 -480 50559 240 8 wbs_adr_i[25]
port 569 nsew signal input
rlabel metal2 s 52251 -480 52307 240 8 wbs_adr_i[26]
port 570 nsew signal input
rlabel metal2 s 54045 -480 54101 240 8 wbs_adr_i[27]
port 571 nsew signal input
rlabel metal2 s 55793 -480 55849 240 8 wbs_adr_i[28]
port 572 nsew signal input
rlabel metal2 s 57587 -480 57643 240 8 wbs_adr_i[29]
port 573 nsew signal input
rlabel metal2 s 8505 -480 8561 240 8 wbs_adr_i[2]
port 574 nsew signal input
rlabel metal2 s 59381 -480 59437 240 8 wbs_adr_i[30]
port 575 nsew signal input
rlabel metal2 s 61129 -480 61185 240 8 wbs_adr_i[31]
port 576 nsew signal input
rlabel metal2 s 10897 -480 10953 240 8 wbs_adr_i[3]
port 577 nsew signal input
rlabel metal2 s 13243 -480 13299 240 8 wbs_adr_i[4]
port 578 nsew signal input
rlabel metal2 s 15037 -480 15093 240 8 wbs_adr_i[5]
port 579 nsew signal input
rlabel metal2 s 16785 -480 16841 240 8 wbs_adr_i[6]
port 580 nsew signal input
rlabel metal2 s 18579 -480 18635 240 8 wbs_adr_i[7]
port 581 nsew signal input
rlabel metal2 s 20327 -480 20383 240 8 wbs_adr_i[8]
port 582 nsew signal input
rlabel metal2 s 22121 -480 22177 240 8 wbs_adr_i[9]
port 583 nsew signal input
rlabel metal2 s 2019 -480 2075 240 8 wbs_cyc_i
port 584 nsew signal input
rlabel metal2 s 4365 -480 4421 240 8 wbs_dat_i[0]
port 585 nsew signal input
rlabel metal2 s 24467 -480 24523 240 8 wbs_dat_i[10]
port 586 nsew signal input
rlabel metal2 s 26261 -480 26317 240 8 wbs_dat_i[11]
port 587 nsew signal input
rlabel metal2 s 28009 -480 28065 240 8 wbs_dat_i[12]
port 588 nsew signal input
rlabel metal2 s 29803 -480 29859 240 8 wbs_dat_i[13]
port 589 nsew signal input
rlabel metal2 s 31597 -480 31653 240 8 wbs_dat_i[14]
port 590 nsew signal input
rlabel metal2 s 33345 -480 33401 240 8 wbs_dat_i[15]
port 591 nsew signal input
rlabel metal2 s 35139 -480 35195 240 8 wbs_dat_i[16]
port 592 nsew signal input
rlabel metal2 s 36887 -480 36943 240 8 wbs_dat_i[17]
port 593 nsew signal input
rlabel metal2 s 38681 -480 38737 240 8 wbs_dat_i[18]
port 594 nsew signal input
rlabel metal2 s 40429 -480 40485 240 8 wbs_dat_i[19]
port 595 nsew signal input
rlabel metal2 s 6757 -480 6813 240 8 wbs_dat_i[1]
port 596 nsew signal input
rlabel metal2 s 42223 -480 42279 240 8 wbs_dat_i[20]
port 597 nsew signal input
rlabel metal2 s 43971 -480 44027 240 8 wbs_dat_i[21]
port 598 nsew signal input
rlabel metal2 s 45765 -480 45821 240 8 wbs_dat_i[22]
port 599 nsew signal input
rlabel metal2 s 47559 -480 47615 240 8 wbs_dat_i[23]
port 600 nsew signal input
rlabel metal2 s 49307 -480 49363 240 8 wbs_dat_i[24]
port 601 nsew signal input
rlabel metal2 s 51101 -480 51157 240 8 wbs_dat_i[25]
port 602 nsew signal input
rlabel metal2 s 52849 -480 52905 240 8 wbs_dat_i[26]
port 603 nsew signal input
rlabel metal2 s 54643 -480 54699 240 8 wbs_dat_i[27]
port 604 nsew signal input
rlabel metal2 s 56391 -480 56447 240 8 wbs_dat_i[28]
port 605 nsew signal input
rlabel metal2 s 58185 -480 58241 240 8 wbs_dat_i[29]
port 606 nsew signal input
rlabel metal2 s 9103 -480 9159 240 8 wbs_dat_i[2]
port 607 nsew signal input
rlabel metal2 s 59933 -480 59989 240 8 wbs_dat_i[30]
port 608 nsew signal input
rlabel metal2 s 61727 -480 61783 240 8 wbs_dat_i[31]
port 609 nsew signal input
rlabel metal2 s 11495 -480 11551 240 8 wbs_dat_i[3]
port 610 nsew signal input
rlabel metal2 s 13841 -480 13897 240 8 wbs_dat_i[4]
port 611 nsew signal input
rlabel metal2 s 15635 -480 15691 240 8 wbs_dat_i[5]
port 612 nsew signal input
rlabel metal2 s 17383 -480 17439 240 8 wbs_dat_i[6]
port 613 nsew signal input
rlabel metal2 s 19177 -480 19233 240 8 wbs_dat_i[7]
port 614 nsew signal input
rlabel metal2 s 20925 -480 20981 240 8 wbs_dat_i[8]
port 615 nsew signal input
rlabel metal2 s 22719 -480 22775 240 8 wbs_dat_i[9]
port 616 nsew signal input
rlabel metal2 s 4963 -480 5019 240 8 wbs_dat_o[0]
port 617 nsew signal tristate
rlabel metal2 s 25065 -480 25121 240 8 wbs_dat_o[10]
port 618 nsew signal tristate
rlabel metal2 s 26859 -480 26915 240 8 wbs_dat_o[11]
port 619 nsew signal tristate
rlabel metal2 s 28607 -480 28663 240 8 wbs_dat_o[12]
port 620 nsew signal tristate
rlabel metal2 s 30401 -480 30457 240 8 wbs_dat_o[13]
port 621 nsew signal tristate
rlabel metal2 s 32149 -480 32205 240 8 wbs_dat_o[14]
port 622 nsew signal tristate
rlabel metal2 s 33943 -480 33999 240 8 wbs_dat_o[15]
port 623 nsew signal tristate
rlabel metal2 s 35737 -480 35793 240 8 wbs_dat_o[16]
port 624 nsew signal tristate
rlabel metal2 s 37485 -480 37541 240 8 wbs_dat_o[17]
port 625 nsew signal tristate
rlabel metal2 s 39279 -480 39335 240 8 wbs_dat_o[18]
port 626 nsew signal tristate
rlabel metal2 s 41027 -480 41083 240 8 wbs_dat_o[19]
port 627 nsew signal tristate
rlabel metal2 s 7355 -480 7411 240 8 wbs_dat_o[1]
port 628 nsew signal tristate
rlabel metal2 s 42821 -480 42877 240 8 wbs_dat_o[20]
port 629 nsew signal tristate
rlabel metal2 s 44569 -480 44625 240 8 wbs_dat_o[21]
port 630 nsew signal tristate
rlabel metal2 s 46363 -480 46419 240 8 wbs_dat_o[22]
port 631 nsew signal tristate
rlabel metal2 s 48111 -480 48167 240 8 wbs_dat_o[23]
port 632 nsew signal tristate
rlabel metal2 s 49905 -480 49961 240 8 wbs_dat_o[24]
port 633 nsew signal tristate
rlabel metal2 s 51653 -480 51709 240 8 wbs_dat_o[25]
port 634 nsew signal tristate
rlabel metal2 s 53447 -480 53503 240 8 wbs_dat_o[26]
port 635 nsew signal tristate
rlabel metal2 s 55241 -480 55297 240 8 wbs_dat_o[27]
port 636 nsew signal tristate
rlabel metal2 s 56989 -480 57045 240 8 wbs_dat_o[28]
port 637 nsew signal tristate
rlabel metal2 s 58783 -480 58839 240 8 wbs_dat_o[29]
port 638 nsew signal tristate
rlabel metal2 s 9701 -480 9757 240 8 wbs_dat_o[2]
port 639 nsew signal tristate
rlabel metal2 s 60531 -480 60587 240 8 wbs_dat_o[30]
port 640 nsew signal tristate
rlabel metal2 s 62325 -480 62381 240 8 wbs_dat_o[31]
port 641 nsew signal tristate
rlabel metal2 s 12093 -480 12149 240 8 wbs_dat_o[3]
port 642 nsew signal tristate
rlabel metal2 s 14439 -480 14495 240 8 wbs_dat_o[4]
port 643 nsew signal tristate
rlabel metal2 s 16187 -480 16243 240 8 wbs_dat_o[5]
port 644 nsew signal tristate
rlabel metal2 s 17981 -480 18037 240 8 wbs_dat_o[6]
port 645 nsew signal tristate
rlabel metal2 s 19775 -480 19831 240 8 wbs_dat_o[7]
port 646 nsew signal tristate
rlabel metal2 s 21523 -480 21579 240 8 wbs_dat_o[8]
port 647 nsew signal tristate
rlabel metal2 s 23317 -480 23373 240 8 wbs_dat_o[9]
port 648 nsew signal tristate
rlabel metal2 s 5561 -480 5617 240 8 wbs_sel_i[0]
port 649 nsew signal input
rlabel metal2 s 7953 -480 8009 240 8 wbs_sel_i[1]
port 650 nsew signal input
rlabel metal2 s 10299 -480 10355 240 8 wbs_sel_i[2]
port 651 nsew signal input
rlabel metal2 s 12645 -480 12701 240 8 wbs_sel_i[3]
port 652 nsew signal input
rlabel metal2 s 2617 -480 2673 240 8 wbs_stb_i
port 653 nsew signal input
rlabel metal2 s 3215 -480 3271 240 8 wbs_we_i
port 654 nsew signal input
rlabel metal4 s 292660 -462 292960 352430 6 vccd1
port 655 nsew power bidirectional
rlabel metal4 s -998 -462 -698 352430 4 vccd1.extra1
port 656 nsew power bidirectional
rlabel metal5 s -998 352130 292960 352430 6 vccd1.extra2
port 657 nsew power bidirectional
rlabel metal5 s -998 -462 292960 -162 8 vccd1.extra3
port 658 nsew power bidirectional
rlabel metal4 s 293130 -932 293430 352900 6 vssd1
port 659 nsew ground bidirectional
rlabel metal4 s -1468 -932 -1168 352900 4 vssd1.extra1
port 660 nsew ground bidirectional
rlabel metal5 s -1468 352600 293430 352900 6 vssd1.extra2
port 661 nsew ground bidirectional
rlabel metal5 s -1468 -932 293430 -632 8 vssd1.extra3
port 662 nsew ground bidirectional
rlabel metal4 s 293600 -1402 293900 353370 6 vccd2
port 663 nsew power bidirectional
rlabel metal4 s -1938 -1402 -1638 353370 4 vccd2.extra1
port 664 nsew power bidirectional
rlabel metal5 s -1938 353070 293900 353370 6 vccd2.extra2
port 665 nsew power bidirectional
rlabel metal5 s -1938 -1402 293900 -1102 8 vccd2.extra3
port 666 nsew power bidirectional
rlabel metal4 s 294070 -1872 294370 353840 6 vssd2
port 667 nsew ground bidirectional
rlabel metal4 s -2408 -1872 -2108 353840 4 vssd2.extra1
port 668 nsew ground bidirectional
rlabel metal5 s -2408 353540 294370 353840 6 vssd2.extra2
port 669 nsew ground bidirectional
rlabel metal5 s -2408 -1872 294370 -1572 8 vssd2.extra3
port 670 nsew ground bidirectional
rlabel metal4 s 294540 -2342 294840 354310 6 vdda1
port 671 nsew power bidirectional
rlabel metal4 s -2878 -2342 -2578 354310 4 vdda1.extra1
port 672 nsew power bidirectional
rlabel metal5 s -2878 354010 294840 354310 6 vdda1.extra2
port 673 nsew power bidirectional
rlabel metal5 s -2878 -2342 294840 -2042 8 vdda1.extra3
port 674 nsew power bidirectional
rlabel metal4 s 295010 -2812 295310 354780 6 vssa1
port 675 nsew ground bidirectional
rlabel metal4 s -3348 -2812 -3048 354780 4 vssa1.extra1
port 676 nsew ground bidirectional
rlabel metal5 s -3348 354480 295310 354780 6 vssa1.extra2
port 677 nsew ground bidirectional
rlabel metal5 s -3348 -2812 295310 -2512 8 vssa1.extra3
port 678 nsew ground bidirectional
rlabel metal4 s 295480 -3282 295780 355250 6 vdda2
port 679 nsew power bidirectional
rlabel metal4 s -3818 -3282 -3518 355250 4 vdda2.extra1
port 680 nsew power bidirectional
rlabel metal5 s -3818 354950 295780 355250 6 vdda2.extra2
port 681 nsew power bidirectional
rlabel metal5 s -3818 -3282 295780 -2982 8 vdda2.extra3
port 682 nsew power bidirectional
rlabel metal4 s 295950 -3752 296250 355720 6 vssa2
port 683 nsew ground bidirectional
rlabel metal4 s -4288 -3752 -3988 355720 4 vssa2.extra1
port 684 nsew ground bidirectional
rlabel metal5 s -4288 355420 296250 355720 6 vssa2.extra2
port 685 nsew ground bidirectional
rlabel metal5 s -4288 -3752 296250 -3452 8 vssa2.extra3
port 686 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
