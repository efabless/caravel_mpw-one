magic
tech sky130A
magscale 1 2
timestamp 1623348570
<< checkpaint >>
rect -1288 -1260 11504 1935
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_10
timestamp 1623348570
transform 1 0 9360 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_9
timestamp 1623348570
transform 1 0 8504 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_8
timestamp 1623348570
transform 1 0 7648 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_7
timestamp 1623348570
transform 1 0 6792 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_6
timestamp 1623348570
transform 1 0 5936 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_5
timestamp 1623348570
transform 1 0 5080 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_4
timestamp 1623348570
transform 1 0 4224 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_3
timestamp 1623348570
transform 1 0 3368 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_2
timestamp 1623348570
transform 1 0 2512 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_1
timestamp 1623348570
transform 1 0 1656 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd2__example_55959141808559  sky130_fd_pr__hvdfl1sd2__example_55959141808559_0
timestamp 1623348570
transform 1 0 800 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808700  sky130_fd_pr__hvdfl1sd__example_55959141808700_0
timestamp 1623348570
transform -1 0 0 0 1 0
box 0 0 1 1
use sky130_fd_pr__hvdfl1sd__example_55959141808700  sky130_fd_pr__hvdfl1sd__example_55959141808700_1
timestamp 1623348570
transform 1 0 10216 0 1 0
box 0 0 1 1
<< labels >>
flabel comment s 10244 675 10244 675 0 FreeSans 300 0 0 0 S
flabel comment s 9388 675 9388 675 0 FreeSans 300 0 0 0 D
flabel comment s 8532 675 8532 675 0 FreeSans 300 0 0 0 S
flabel comment s 7676 675 7676 675 0 FreeSans 300 0 0 0 D
flabel comment s 6820 675 6820 675 0 FreeSans 300 0 0 0 S
flabel comment s 5964 675 5964 675 0 FreeSans 300 0 0 0 D
flabel comment s 5108 675 5108 675 0 FreeSans 300 0 0 0 S
flabel comment s 4252 675 4252 675 0 FreeSans 300 0 0 0 D
flabel comment s 3396 675 3396 675 0 FreeSans 300 0 0 0 S
flabel comment s 2540 675 2540 675 0 FreeSans 300 0 0 0 D
flabel comment s 1684 675 1684 675 0 FreeSans 300 0 0 0 S
flabel comment s 828 675 828 675 0 FreeSans 300 0 0 0 D
flabel comment s -28 675 -28 675 0 FreeSans 300 0 0 0 S
<< properties >>
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_io/gds/sky130_fd_io.gds
string GDS_END 15473678
string GDS_START 15467054
<< end >>
