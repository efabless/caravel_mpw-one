magic
tech sky130A
magscale 1 2
timestamp 1606852874
<< obsli1 >>
rect 76168 997646 92232 1037541
rect 127568 997646 143632 1037541
rect 178968 997646 195032 1037541
rect 230368 997646 246432 1037541
rect 281968 997646 298032 1037541
rect 333614 998007 347955 1037539
rect 383768 997646 399832 1037541
rect 472768 997646 488832 1037541
rect 524168 997646 540232 1037541
rect 575814 998007 590155 1037539
rect 625968 997646 642032 1037541
rect 59 954168 39954 970232
rect 677646 951568 717541 967632
rect 44 912048 39396 926951
rect 678204 907649 717556 922552
rect 61 869922 39593 884371
rect 677646 862368 717541 878432
rect 61 827814 39593 842155
rect 678007 818829 717539 833278
rect 59 784368 39954 800432
rect 677646 773168 717541 789232
rect 59 741168 39954 757232
rect 677646 728168 717541 744232
rect 59 697968 39954 714032
rect 677646 683168 717541 699232
rect 59 654768 39954 670832
rect 677646 637968 717541 654032
rect 59 611568 39954 627632
rect 677646 592968 717541 609032
rect 59 568368 39954 584432
rect 677646 547768 717541 563832
rect 59 525168 39954 541232
rect 678007 504229 717539 518678
rect 61 483122 39593 497571
rect 678204 459849 717556 474752
rect 44 440848 39396 455751
rect 678007 416045 717539 430386
rect 59 397568 39954 413632
rect 677646 370568 717541 386632
rect 59 354368 39954 370432
rect 59 311168 39954 327232
rect 677646 325368 717541 341432
rect 59 267968 39954 284032
rect 677646 280368 717541 296432
rect 59 224768 39954 240832
rect 677646 235368 717541 251432
rect 59 181568 39954 197632
rect 677646 190168 717541 206232
rect 677646 145168 717541 161232
rect 61 110322 39593 124771
rect 677646 99968 717541 116032
rect 44 68048 39396 82951
rect 79245 61 93586 39593
rect 132600 156 147600 39963
rect 186368 59 202432 39954
rect 241249 44 256152 39396
rect 294968 59 311032 39954
rect 349768 59 365832 39954
rect 404568 59 420632 39954
rect 459368 59 475432 39954
rect 514168 59 530232 39954
rect 569445 61 583786 39593
rect 623229 61 637678 39593
<< metal1 >>
rect 84016 995596 84068 995648
rect 91744 995596 91796 995648
rect 238208 995596 238260 995648
rect 245936 995596 245988 995648
rect 531964 995596 532016 995648
rect 539692 995596 539744 995648
rect 135352 995460 135404 995512
rect 143172 995460 143224 995512
rect 633808 995460 633860 995512
rect 641536 995460 641588 995512
rect 289636 995256 289688 995308
rect 297640 995256 297692 995308
rect 391480 995256 391532 995308
rect 399484 995256 399536 995308
rect 480444 995256 480496 995308
rect 488448 995256 488500 995308
rect 231860 995052 231912 995104
rect 244188 995052 244240 995104
rect 463786 992264 463792 992316
rect 463844 992304 463850 992316
rect 475470 992304 475476 992316
rect 463844 992276 475476 992304
rect 463844 992264 463850 992276
rect 475470 992264 475476 992276
rect 475528 992304 475534 992316
rect 482922 992304 482928 992316
rect 475528 992276 482928 992304
rect 475528 992264 475534 992276
rect 482922 992264 482928 992276
rect 482980 992264 482986 992316
rect 141424 992060 141476 992112
rect 154396 992060 154448 992112
rect 130286 990876 130292 990888
rect 130120 990848 130292 990876
rect 130120 990820 130148 990848
rect 130286 990836 130292 990848
rect 130344 990876 130350 990888
rect 130344 990848 130424 990876
rect 130344 990836 130350 990848
rect 79042 990768 79048 990820
rect 79100 990808 79106 990820
rect 110414 990808 110420 990820
rect 79100 990780 110420 990808
rect 79100 990768 79106 990780
rect 110414 990768 110420 990780
rect 110472 990768 110478 990820
rect 130102 990768 130108 990820
rect 130160 990768 130166 990820
rect 130396 990808 130424 990848
rect 419534 990836 419540 990888
rect 419592 990876 419598 990888
rect 438670 990876 438676 990888
rect 419592 990848 438676 990876
rect 419592 990836 419598 990848
rect 438670 990836 438676 990848
rect 438728 990836 438734 990888
rect 450262 990836 450268 990888
rect 450320 990876 450326 990888
rect 463602 990876 463608 990888
rect 450320 990848 463608 990876
rect 450320 990836 450326 990848
rect 463602 990836 463608 990848
rect 463660 990836 463666 990888
rect 143258 990808 143264 990820
rect 130396 990780 143264 990808
rect 143258 990768 143264 990780
rect 143316 990768 143322 990820
rect 173802 990768 173808 990820
rect 173860 990808 173866 990820
rect 179322 990808 179328 990820
rect 173860 990780 179328 990808
rect 173860 990768 173866 990780
rect 179322 990768 179328 990780
rect 179380 990768 179386 990820
rect 246942 990768 246948 990820
rect 247000 990808 247006 990820
rect 284662 990808 284668 990820
rect 247000 990780 284668 990808
rect 247000 990768 247006 990780
rect 284662 990768 284668 990780
rect 284720 990808 284726 990820
rect 286962 990808 286968 990820
rect 284720 990780 286968 990808
rect 284720 990768 284726 990780
rect 286962 990768 286968 990780
rect 287020 990768 287026 990820
rect 391756 990768 391808 990820
rect 476120 990768 476172 990820
rect 527548 990768 527600 990820
rect 629300 990768 629352 990820
rect 187602 990700 187608 990752
rect 187660 990740 187666 990752
rect 187694 990740 187700 990752
rect 187660 990712 187700 990740
rect 187660 990700 187666 990712
rect 187694 990700 187700 990712
rect 187752 990700 187758 990752
rect 202874 990700 202880 990752
rect 202932 990740 202938 990752
rect 233050 990740 233056 990752
rect 202932 990712 233056 990740
rect 202932 990700 202938 990712
rect 233050 990700 233056 990712
rect 233108 990700 233114 990752
rect 244188 990700 244240 990752
rect 295800 990700 295852 990752
rect 386328 990700 386380 990752
rect 482922 990700 482928 990752
rect 482980 990740 482986 990752
rect 526898 990740 526904 990752
rect 482980 990712 526904 990740
rect 482980 990700 482986 990712
rect 526898 990700 526904 990712
rect 526956 990740 526962 990752
rect 628650 990740 628656 990752
rect 526956 990712 628656 990740
rect 526956 990700 526962 990712
rect 628650 990700 628656 990712
rect 628708 990700 628714 990752
rect 79508 990632 79560 990684
rect 79968 990632 80020 990684
rect 130936 990632 130988 990684
rect 182364 990632 182416 990684
rect 233700 990632 233752 990684
rect 285312 990632 285364 990684
rect 333520 990632 333572 990684
rect 387156 990632 387208 990684
rect 391756 990632 391808 990684
rect 391860 990644 405596 990672
rect 89996 990564 90048 990616
rect 110506 990564 110512 990616
rect 110564 990604 110570 990616
rect 130102 990604 130108 990616
rect 110564 990576 130108 990604
rect 110564 990564 110570 990576
rect 130102 990564 130108 990576
rect 130160 990564 130166 990616
rect 179322 990564 179328 990616
rect 179380 990604 179386 990616
rect 181714 990604 181720 990616
rect 179380 990576 181720 990604
rect 179380 990564 179386 990576
rect 181714 990564 181720 990576
rect 181772 990564 181778 990616
rect 186688 990564 186740 990616
rect 194692 990564 194744 990616
rect 386506 990604 386512 990616
rect 386419 990576 386512 990604
rect 386506 990564 386512 990576
rect 386564 990604 386570 990616
rect 391860 990604 391888 990644
rect 386564 990576 391888 990604
rect 386564 990564 386570 990576
rect 164148 990496 164200 990548
rect 192852 990496 192904 990548
rect 193220 990496 193272 990548
rect 212448 990496 212500 990548
rect 231860 990496 231912 990548
rect 286962 990496 286968 990548
rect 287020 990536 287026 990548
rect 386524 990536 386552 990564
rect 287020 990508 386552 990536
rect 405568 990536 405596 990644
rect 596088 990632 596140 990684
rect 419534 990604 419540 990616
rect 405752 990576 419540 990604
rect 405752 990536 405780 990576
rect 419534 990564 419540 990576
rect 419592 990564 419598 990616
rect 438762 990564 438768 990616
rect 438820 990604 438826 990616
rect 450262 990604 450268 990616
rect 438820 990576 450268 990604
rect 438820 990564 438826 990576
rect 450262 990564 450268 990576
rect 450320 990564 450326 990616
rect 469312 990564 469364 990616
rect 405568 990508 405780 990536
rect 287020 990496 287026 990508
rect 141332 990428 141384 990480
rect 143258 990428 143264 990480
rect 143316 990468 143322 990480
rect 160094 990468 160100 990480
rect 143316 990440 160100 990468
rect 143316 990428 143322 990440
rect 160094 990428 160100 990440
rect 160152 990428 160158 990480
rect 181714 990428 181720 990480
rect 181772 990468 181778 990480
rect 187602 990468 187608 990480
rect 181772 990440 187608 990468
rect 181772 990428 181778 990440
rect 187602 990428 187608 990440
rect 187660 990428 187666 990480
rect 187694 990428 187700 990480
rect 187752 990468 187758 990480
rect 202874 990468 202880 990480
rect 187752 990440 202880 990468
rect 187752 990428 187758 990440
rect 202874 990428 202880 990440
rect 202932 990428 202938 990480
rect 233050 990428 233056 990480
rect 233108 990468 233114 990480
rect 246942 990468 246948 990480
rect 233108 990440 246948 990468
rect 233108 990428 233114 990440
rect 246942 990428 246948 990440
rect 247000 990428 247006 990480
rect 469036 990496 469088 990548
rect 483020 990496 483072 990548
rect 560208 990496 560260 990548
rect 576860 990564 576912 990616
rect 623688 990564 623740 990616
rect 623872 990496 623924 990548
rect 639788 990496 639840 990548
rect 154396 990360 154448 990412
rect 154580 990360 154632 990412
rect 386328 990360 386380 990412
rect 397644 990360 397696 990412
rect 424968 990360 425020 990412
rect 540980 990428 541032 990480
rect 483020 990360 483072 990412
rect 486608 990360 486660 990412
rect 507768 990292 507820 990344
rect 507860 990292 507912 990344
rect 521660 990360 521712 990412
rect 540888 990360 540940 990412
rect 154580 990224 154632 990276
rect 164148 990224 164200 990276
rect 397644 990224 397696 990276
rect 405740 990224 405792 990276
rect 521660 990224 521712 990276
rect 537852 990224 537904 990276
rect 540888 990224 540940 990276
rect 42248 990156 42300 990208
rect 79968 990156 80020 990208
rect 639788 990156 639840 990208
rect 673644 990156 673696 990208
rect 42426 990088 42432 990140
rect 42484 990128 42490 990140
rect 79042 990128 79048 990140
rect 42484 990100 79048 990128
rect 42484 990088 42490 990100
rect 79042 990088 79048 990100
rect 79100 990088 79106 990140
rect 89996 990088 90048 990140
rect 405740 990088 405792 990140
rect 424968 990088 425020 990140
rect 628650 990088 628656 990140
rect 628708 990088 628714 990140
rect 629300 990088 629352 990140
rect 673552 990088 673604 990140
rect 42524 990020 42576 990072
rect 628668 990060 628696 990088
rect 673454 990060 673460 990072
rect 628668 990032 673460 990060
rect 673454 990020 673460 990032
rect 673512 990020 673518 990072
rect 41788 969348 41840 969400
rect 42340 969348 42392 969400
rect 41788 968464 41840 968516
rect 42524 968464 42576 968516
rect 673454 965268 673460 965320
rect 673512 965308 673518 965320
rect 675386 965308 675392 965320
rect 673512 965280 675392 965308
rect 673512 965268 673518 965280
rect 675386 965268 675392 965280
rect 675444 965268 675450 965320
rect 673552 964724 673604 964776
rect 675392 964724 675444 964776
rect 41788 962412 41840 962464
rect 42340 962412 42392 962464
rect 41782 956428 41788 956480
rect 41840 956468 41846 956480
rect 42426 956468 42432 956480
rect 41840 956440 42432 956468
rect 41840 956428 41846 956440
rect 42426 956428 42432 956440
rect 42484 956428 42490 956480
rect 673644 953300 673696 953352
rect 675392 953300 675444 953352
rect 44272 930112 44324 930164
rect 45468 930112 45520 930164
rect 39672 922904 39724 922956
rect 44272 922904 44324 922956
rect 39856 914676 39908 914728
rect 41420 914676 41472 914728
rect 42248 914676 42300 914728
rect 673552 910732 673604 910784
rect 677784 910732 677836 910784
rect 673178 908012 673184 908064
rect 673236 908052 673242 908064
rect 673454 908052 673460 908064
rect 673236 908024 673460 908052
rect 673236 908012 673242 908024
rect 673454 908012 673460 908024
rect 673512 908012 673518 908064
rect 673178 888768 673184 888820
rect 673236 888808 673242 888820
rect 673454 888808 673460 888820
rect 673236 888780 673460 888808
rect 673236 888768 673242 888780
rect 673454 888768 673460 888780
rect 673512 888768 673518 888820
rect 39856 879792 39908 879844
rect 40132 879792 40184 879844
rect 44180 879792 44232 879844
rect 45836 879792 45888 879844
rect 41420 875576 41472 875628
rect 42248 875576 42300 875628
rect 673552 875508 673604 875560
rect 675392 875508 675444 875560
rect 673644 875032 673696 875084
rect 673644 874896 673696 874948
rect 673730 869388 673736 869440
rect 673788 869428 673794 869440
rect 675202 869428 675208 869440
rect 673788 869400 675208 869428
rect 673788 869388 673794 869400
rect 675202 869388 675208 869400
rect 675260 869388 675266 869440
rect 673644 864968 673696 865020
rect 673828 864968 673880 865020
rect 675392 864968 675444 865020
rect 673546 836272 673552 836324
rect 673604 836312 673610 836324
rect 673604 836284 673684 836312
rect 673604 836272 673610 836284
rect 673656 836256 673684 836284
rect 673638 836204 673644 836256
rect 673696 836204 673702 836256
rect 673546 830764 673552 830816
rect 673604 830804 673610 830816
rect 673638 830804 673644 830816
rect 673604 830776 673644 830804
rect 673604 830764 673610 830776
rect 673638 830764 673644 830776
rect 673696 830764 673702 830816
rect 673546 821040 673552 821092
rect 673604 821080 673610 821092
rect 674098 821080 674104 821092
rect 673604 821052 674104 821080
rect 673604 821040 673610 821052
rect 674098 821040 674104 821052
rect 674156 821040 674162 821092
rect 42248 807304 42300 807356
rect 42708 807304 42760 807356
rect 44548 805944 44600 805996
rect 44732 805944 44784 805996
rect 41788 798328 41840 798380
rect 42524 798328 42576 798380
rect 674098 797580 674104 797632
rect 674156 797620 674162 797632
rect 675294 797620 675300 797632
rect 674156 797592 675300 797620
rect 674156 797580 674162 797592
rect 675294 797580 675300 797592
rect 675352 797580 675358 797632
rect 41788 787856 41840 787908
rect 42432 787856 42484 787908
rect 42708 787856 42760 787908
rect 42242 787176 42248 787228
rect 42300 787216 42306 787228
rect 42610 787216 42616 787228
rect 42300 787188 42616 787216
rect 42300 787176 42306 787188
rect 42610 787176 42616 787188
rect 42668 787176 42674 787228
rect 674006 786428 674012 786480
rect 674064 786468 674070 786480
rect 675294 786468 675300 786480
rect 674064 786440 675300 786468
rect 674064 786428 674070 786440
rect 675294 786428 675300 786440
rect 675352 786428 675358 786480
rect 673644 785272 673696 785324
rect 675392 785272 675444 785324
rect 673000 778336 673052 778388
rect 673092 778200 673144 778252
rect 673460 774868 673512 774920
rect 673828 774868 673880 774920
rect 675392 774868 675444 774920
rect 672816 772760 672868 772812
rect 673092 772760 673144 772812
rect 42524 768612 42576 768664
rect 42708 768612 42760 768664
rect 673546 768612 673552 768664
rect 673604 768652 673610 768664
rect 674006 768652 674012 768664
rect 673604 768624 674012 768652
rect 673604 768612 673610 768624
rect 674006 768612 674012 768624
rect 674064 768612 674070 768664
rect 41788 754468 41840 754520
rect 42524 754468 42576 754520
rect 42708 754468 42760 754520
rect 41782 744404 41788 744456
rect 41840 744444 41846 744456
rect 42610 744444 42616 744456
rect 41840 744416 42616 744444
rect 41840 744404 41846 744416
rect 42610 744404 42616 744416
rect 42668 744404 42674 744456
rect 673546 741888 673552 741940
rect 673604 741928 673610 741940
rect 674190 741928 674196 741940
rect 673604 741900 674196 741928
rect 673604 741888 673610 741900
rect 674190 741888 674196 741900
rect 674248 741928 674254 741940
rect 675386 741928 675392 741940
rect 674248 741900 675392 741928
rect 674248 741888 674254 741900
rect 675386 741888 675392 741900
rect 675444 741888 675450 741940
rect 673644 741344 673696 741396
rect 675392 741344 675444 741396
rect 673000 739712 673052 739764
rect 673184 739576 673236 739628
rect 673460 730124 673512 730176
rect 675392 730124 675444 730176
rect 673828 729988 673880 730040
rect 675116 729988 675168 730040
rect 674006 720400 674012 720452
rect 674064 720440 674070 720452
rect 674190 720440 674196 720452
rect 674064 720412 674196 720440
rect 674064 720400 674070 720412
rect 674190 720400 674196 720412
rect 674248 720400 674254 720452
rect 41788 711288 41840 711340
rect 42524 711288 42576 711340
rect 674006 710676 674012 710728
rect 674064 710716 674070 710728
rect 675294 710716 675300 710728
rect 674064 710688 675300 710716
rect 674064 710676 674070 710688
rect 675294 710676 675300 710688
rect 675352 710676 675358 710728
rect 42248 700952 42300 701004
rect 42524 700952 42576 701004
rect 41782 700816 41788 700868
rect 41840 700856 41846 700868
rect 42610 700856 42616 700868
rect 41840 700828 42616 700856
rect 41840 700816 41846 700828
rect 42610 700816 42616 700828
rect 42668 700816 42674 700868
rect 673638 695920 673644 695972
rect 673696 695960 673702 695972
rect 675386 695960 675392 695972
rect 673696 695932 675392 695960
rect 673696 695920 673702 695932
rect 675386 695920 675392 695932
rect 675444 695920 675450 695972
rect 673092 695512 673144 695564
rect 673184 695512 673236 695564
rect 44640 695444 44692 695496
rect 44916 695444 44968 695496
rect 673552 695308 673604 695360
rect 673828 695308 673880 695360
rect 675392 695308 675444 695360
rect 44732 676200 44784 676252
rect 44916 676200 44968 676252
rect 42340 669128 42392 669180
rect 41788 669060 41840 669112
rect 673184 662464 673236 662516
rect 44548 662396 44600 662448
rect 44732 662396 44784 662448
rect 673184 662328 673236 662380
rect 41788 657636 41840 657688
rect 42524 657636 42576 657688
rect 41782 657092 41788 657144
rect 41840 657132 41846 657144
rect 42334 657132 42340 657144
rect 41840 657104 42340 657132
rect 41840 657092 41846 657104
rect 42334 657092 42340 657104
rect 42392 657132 42398 657144
rect 42610 657132 42616 657144
rect 42392 657104 42616 657132
rect 42392 657092 42398 657104
rect 42610 657092 42616 657104
rect 42668 657092 42674 657144
rect 44640 656820 44692 656872
rect 44824 656820 44876 656872
rect 673638 651720 673644 651772
rect 673696 651760 673702 651772
rect 675386 651760 675392 651772
rect 673696 651732 675392 651760
rect 673696 651720 673702 651732
rect 675386 651720 675392 651732
rect 675444 651720 675450 651772
rect 673552 651108 673604 651160
rect 675392 651108 675444 651160
rect 673460 639684 673512 639736
rect 675392 639684 675444 639736
rect 672816 637508 672868 637560
rect 673092 637508 673144 637560
rect 42524 633496 42576 633548
rect 42524 633292 42576 633344
rect 42334 633224 42340 633276
rect 42392 633264 42398 633276
rect 42610 633264 42616 633276
rect 42392 633236 42616 633264
rect 42392 633224 42398 633236
rect 42610 633224 42616 633236
rect 42668 633224 42674 633276
rect 41788 625880 41840 625932
rect 42432 625880 42484 625932
rect 672816 618264 672868 618316
rect 673000 618264 673052 618316
rect 41874 614456 41880 614508
rect 41932 614496 41938 614508
rect 42242 614496 42248 614508
rect 41932 614468 42248 614496
rect 41932 614456 41938 614468
rect 42242 614456 42248 614468
rect 42300 614496 42306 614508
rect 42610 614496 42616 614508
rect 42300 614468 42616 614496
rect 42300 614456 42306 614468
rect 42610 614456 42616 614468
rect 42668 614456 42674 614508
rect 41788 614388 41840 614440
rect 42524 614388 42576 614440
rect 673638 606704 673644 606756
rect 673696 606744 673702 606756
rect 675386 606744 675392 606756
rect 673696 606716 675392 606744
rect 673696 606704 673702 606716
rect 675386 606704 675392 606716
rect 675444 606704 675450 606756
rect 673552 605616 673604 605668
rect 675300 605616 675352 605668
rect 44640 604528 44692 604580
rect 44640 604392 44692 604444
rect 673552 604392 673604 604444
rect 673828 604392 673880 604444
rect 672816 598952 672868 599004
rect 673092 598952 673144 599004
rect 673460 594872 673512 594924
rect 675392 594872 675444 594924
rect 673092 585148 673144 585200
rect 673000 585080 673052 585132
rect 42242 584196 42248 584248
rect 42300 584236 42306 584248
rect 42610 584236 42616 584248
rect 42300 584208 42616 584236
rect 42300 584196 42306 584208
rect 42610 584196 42616 584208
rect 42668 584196 42674 584248
rect 41788 581680 41840 581732
rect 42432 581680 42484 581732
rect 41788 572228 41840 572280
rect 42248 572228 42300 572280
rect 42524 572228 42576 572280
rect 41782 571616 41788 571668
rect 41840 571656 41846 571668
rect 42610 571656 42616 571668
rect 41840 571628 42616 571656
rect 41840 571616 41846 571628
rect 42610 571616 42616 571628
rect 42668 571616 42674 571668
rect 672816 569916 672868 569968
rect 673000 569916 673052 569968
rect 673552 565836 673604 565888
rect 673920 565836 673972 565888
rect 673638 561484 673644 561536
rect 673696 561524 673702 561536
rect 675386 561524 675392 561536
rect 673696 561496 675392 561524
rect 673696 561484 673702 561496
rect 675386 561484 675392 561496
rect 675444 561484 675450 561536
rect 672816 560260 672868 560312
rect 673000 560260 673052 560312
rect 673552 559920 673604 559972
rect 673920 559920 673972 559972
rect 675392 559920 675444 559972
rect 673460 550468 673512 550520
rect 675392 550468 675444 550520
rect 673000 546524 673052 546576
rect 673092 546320 673144 546372
rect 44732 540948 44784 541000
rect 44916 540948 44968 541000
rect 41788 538500 41840 538552
rect 42432 538500 42484 538552
rect 41782 528436 41788 528488
rect 41840 528476 41846 528488
rect 42426 528476 42432 528488
rect 41840 528448 42432 528476
rect 41840 528436 41846 528448
rect 42426 528436 42432 528448
rect 42484 528476 42490 528488
rect 42610 528476 42616 528488
rect 42484 528448 42616 528476
rect 42484 528436 42490 528448
rect 42610 528436 42616 528448
rect 42668 528436 42674 528488
rect 673092 527144 673144 527196
rect 673184 527008 673236 527060
rect 673736 522928 673788 522980
rect 673920 522928 673972 522980
rect 673184 521568 673236 521620
rect 676128 521568 676180 521620
rect 44548 496816 44600 496868
rect 44732 496816 44784 496868
rect 673736 463632 673788 463684
rect 677692 463632 677744 463684
rect 39396 458192 39448 458244
rect 44272 458192 44324 458244
rect 673000 449896 673052 449948
rect 673368 449896 673420 449948
rect 39856 448264 39908 448316
rect 42248 448264 42300 448316
rect 676220 440172 676272 440224
rect 677692 440172 677744 440224
rect 42248 413380 42300 413432
rect 42616 413380 42668 413432
rect 672816 412496 672868 412548
rect 676220 412496 676272 412548
rect 41788 410932 41840 410984
rect 42524 410932 42576 410984
rect 672540 405628 672592 405680
rect 672724 405628 672776 405680
rect 673460 401548 673512 401600
rect 675300 401548 675352 401600
rect 41788 401480 41840 401532
rect 42248 401480 42300 401532
rect 42616 401480 42668 401532
rect 41966 400120 41972 400172
rect 42024 400160 42030 400172
rect 42426 400160 42432 400172
rect 42024 400132 42432 400160
rect 42024 400120 42030 400132
rect 42426 400120 42432 400132
rect 42484 400120 42490 400172
rect 672540 386384 672592 386436
rect 672816 386384 672868 386436
rect 673546 384004 673552 384056
rect 673604 384044 673610 384056
rect 675386 384044 675392 384056
rect 673604 384016 675392 384044
rect 673604 384004 673610 384016
rect 675386 384004 675392 384016
rect 675444 384004 675450 384056
rect 673644 382712 673696 382764
rect 675392 382712 675444 382764
rect 42340 380876 42392 380928
rect 42616 380876 42668 380928
rect 673828 372308 673880 372360
rect 675392 372308 675444 372360
rect 41788 368636 41840 368688
rect 42524 368636 42576 368688
rect 42524 367004 42576 367056
rect 42800 366936 42852 366988
rect 41788 357484 41840 357536
rect 42340 357484 42392 357536
rect 42616 357484 42668 357536
rect 41782 356668 41788 356720
rect 41840 356708 41846 356720
rect 42426 356708 42432 356720
rect 41840 356680 42432 356708
rect 41840 356668 41846 356680
rect 42426 356668 42432 356680
rect 42484 356668 42490 356720
rect 672632 353336 672684 353388
rect 672540 353200 672592 353252
rect 42708 347692 42760 347744
rect 42892 347692 42944 347744
rect 672540 347692 672592 347744
rect 672724 347692 672776 347744
rect 673644 338512 673696 338564
rect 675392 338512 675444 338564
rect 42340 334636 42392 334688
rect 42616 334636 42668 334688
rect 42616 328448 42668 328500
rect 42892 328448 42944 328500
rect 672448 328448 672500 328500
rect 672724 328448 672776 328500
rect 673828 327088 673880 327140
rect 675392 327088 675444 327140
rect 41788 324504 41840 324556
rect 42524 324436 42576 324488
rect 42340 314576 42392 314628
rect 42616 314508 42668 314560
rect 41788 314440 41840 314492
rect 42524 314440 42576 314492
rect 42800 314440 42852 314492
rect 41782 313760 41788 313812
rect 41840 313800 41846 313812
rect 42426 313800 42432 313812
rect 41840 313772 42432 313800
rect 41840 313760 41846 313772
rect 42426 313760 42432 313772
rect 42484 313760 42490 313812
rect 672540 309068 672592 309120
rect 672816 309068 672868 309120
rect 42426 307912 42432 307964
rect 42484 307952 42490 307964
rect 42702 307952 42708 307964
rect 42484 307924 42708 307952
rect 42484 307912 42490 307924
rect 42702 307912 42708 307924
rect 42760 307912 42766 307964
rect 673460 304920 673512 304972
rect 673828 304920 673880 304972
rect 42616 295332 42668 295384
rect 42800 295332 42852 295384
rect 673644 293496 673696 293548
rect 675024 293496 675076 293548
rect 673822 293156 673828 293208
rect 673880 293196 673886 293208
rect 675386 293196 675392 293208
rect 673880 293168 675392 293196
rect 673880 293156 673886 293168
rect 675386 293156 675392 293168
rect 675444 293156 675450 293208
rect 672632 289824 672684 289876
rect 672816 289824 672868 289876
rect 673460 283024 673512 283076
rect 674932 283024 674984 283076
rect 675392 283024 675444 283076
rect 41788 282276 41840 282328
rect 42432 282276 42484 282328
rect 42616 282276 42668 282328
rect 42702 282208 42708 282260
rect 42760 282208 42766 282260
rect 42720 282056 42748 282208
rect 42702 282004 42708 282056
rect 42760 282004 42766 282056
rect 673920 276020 673972 276072
rect 675208 276020 675260 276072
rect 42524 275952 42576 276004
rect 42800 275952 42852 276004
rect 41788 270784 41840 270836
rect 42524 270784 42576 270836
rect 41782 270240 41788 270292
rect 41840 270280 41846 270292
rect 42334 270280 42340 270292
rect 41840 270252 42340 270280
rect 41840 270240 41846 270252
rect 42334 270240 42340 270252
rect 42392 270280 42398 270292
rect 42702 270280 42708 270292
rect 42392 270252 42708 270280
rect 42392 270240 42398 270252
rect 42702 270240 42708 270252
rect 42760 270240 42766 270292
rect 673736 266296 673788 266348
rect 674932 266296 674984 266348
rect 673822 248140 673828 248192
rect 673880 248180 673886 248192
rect 675386 248180 675392 248192
rect 673880 248152 675392 248180
rect 673880 248140 673886 248152
rect 675386 248140 675392 248152
rect 675444 248140 675450 248192
rect 673644 247460 673696 247512
rect 673920 247460 673972 247512
rect 675392 247460 675444 247512
rect 42334 246984 42340 247036
rect 42392 247024 42398 247036
rect 42702 247024 42708 247036
rect 42392 246996 42708 247024
rect 42392 246984 42398 246996
rect 42702 246984 42708 246996
rect 42760 246984 42766 247036
rect 41788 239028 41840 239080
rect 42432 239028 42484 239080
rect 42616 239028 42668 239080
rect 673736 237668 673788 237720
rect 675392 237668 675444 237720
rect 41788 228624 41840 228676
rect 42524 228624 42576 228676
rect 41782 228012 41788 228064
rect 41840 228052 41846 228064
rect 42426 228052 42432 228064
rect 41840 228024 42432 228052
rect 41840 228012 41846 228024
rect 42426 228012 42432 228024
rect 42484 228052 42490 228064
rect 42702 228052 42708 228064
rect 42484 228024 42708 228052
rect 42484 228012 42490 228024
rect 42702 228012 42708 228024
rect 42760 228012 42766 228064
rect 42248 227876 42300 227928
rect 42524 227876 42576 227928
rect 672724 212508 672776 212560
rect 672908 212508 672960 212560
rect 673546 203872 673552 203924
rect 673604 203912 673610 203924
rect 673822 203912 673828 203924
rect 673604 203884 673828 203912
rect 673604 203872 673610 203884
rect 673822 203872 673828 203884
rect 673880 203912 673886 203924
rect 675386 203912 675392 203924
rect 673880 203884 675392 203912
rect 673880 203872 673886 203884
rect 675386 203872 675392 203884
rect 675444 203872 675450 203924
rect 673460 203328 673512 203380
rect 673644 203328 673696 203380
rect 675392 203328 675444 203380
rect 672540 198704 672592 198756
rect 672724 198704 672776 198756
rect 41788 196732 41840 196784
rect 42340 196732 42392 196784
rect 41788 195848 41840 195900
rect 42616 195848 42668 195900
rect 44640 195848 44692 195900
rect 673736 191972 673788 192024
rect 674012 191972 674064 192024
rect 41788 189796 41840 189848
rect 42340 189796 42392 189848
rect 42242 184220 42248 184272
rect 42300 184260 42306 184272
rect 42426 184260 42432 184272
rect 42300 184232 42432 184260
rect 42300 184220 42306 184232
rect 42426 184220 42432 184232
rect 42484 184220 42490 184272
rect 44456 173884 44508 173936
rect 44732 173884 44784 173936
rect 672724 173884 672776 173936
rect 672908 173884 672960 173936
rect 673828 173884 673880 173936
rect 674012 173884 674064 173936
rect 44732 160148 44784 160200
rect 672540 160080 672592 160132
rect 672724 160080 672776 160132
rect 673644 160080 673696 160132
rect 673828 160080 673880 160132
rect 44640 160012 44692 160064
rect 673546 158312 673552 158364
rect 673604 158352 673610 158364
rect 675386 158352 675392 158364
rect 673604 158324 675392 158352
rect 673604 158312 673610 158324
rect 675386 158312 675392 158324
rect 675444 158312 675450 158364
rect 673460 157292 673512 157344
rect 675392 157292 675444 157344
rect 44640 154504 44692 154556
rect 44732 154504 44784 154556
rect 673644 147840 673696 147892
rect 674012 147840 674064 147892
rect 675392 147840 675444 147892
rect 44732 140768 44784 140820
rect 44640 140700 44692 140752
rect 44732 121524 44784 121576
rect 44640 121388 44692 121440
rect 672724 115880 672776 115932
rect 672816 115880 672868 115932
rect 673546 112752 673552 112804
rect 673604 112792 673610 112804
rect 675386 112792 675392 112804
rect 673604 112764 675392 112792
rect 673604 112752 673610 112764
rect 675386 112752 675392 112764
rect 675444 112752 675450 112804
rect 673460 112072 673512 112124
rect 675392 112072 675444 112124
rect 672816 102144 672868 102196
rect 673644 102144 673696 102196
rect 673828 102144 673880 102196
rect 672724 102076 672776 102128
rect 673644 102008 673696 102060
rect 675392 102008 675444 102060
rect 44272 96568 44324 96620
rect 44548 96568 44600 96620
rect 672816 82900 672868 82952
rect 672816 82696 672868 82748
rect 44272 77256 44324 77308
rect 44364 77256 44416 77308
rect 39672 75216 39724 75268
rect 39672 74944 39724 74996
rect 39580 67940 39632 67992
rect 41420 67940 41472 67992
rect 41420 64608 41472 64660
rect 42708 64608 42760 64660
rect 39672 52368 39724 52420
rect 39856 52368 39908 52420
rect 45468 47880 45520 47932
rect 179420 47880 179472 47932
rect 518808 47880 518860 47932
rect 673644 47880 673696 47932
rect 39856 47812 39908 47864
rect 189172 47812 189224 47864
rect 527450 47812 527456 47864
rect 527508 47852 527514 47864
rect 673546 47852 673552 47864
rect 527508 47824 673552 47852
rect 527508 47812 527514 47824
rect 673546 47812 673552 47824
rect 673604 47812 673610 47864
rect 45560 47744 45612 47796
rect 149060 47744 149112 47796
rect 528652 47744 528704 47796
rect 672816 47744 672868 47796
rect 39764 47676 39816 47728
rect 86316 47676 86368 47728
rect 179420 47472 179472 47524
rect 195980 47540 196032 47592
rect 198648 47540 198700 47592
rect 198740 47540 198792 47592
rect 212540 47608 212592 47660
rect 270500 47608 270552 47660
rect 303620 47540 303672 47592
rect 304540 47540 304592 47592
rect 359372 47540 359424 47592
rect 361488 47540 361540 47592
rect 231768 47472 231820 47524
rect 251180 47472 251232 47524
rect 270408 47472 270460 47524
rect 289728 47404 289780 47456
rect 86316 47336 86368 47388
rect 199016 47336 199068 47388
rect 201408 47336 201460 47388
rect 251180 47336 251232 47388
rect 270408 47336 270460 47388
rect 364156 47404 364208 47456
rect 416780 47472 416832 47524
rect 303620 47336 303672 47388
rect 361488 47336 361540 47388
rect 414204 47336 414256 47388
rect 417976 47336 418028 47388
rect 418068 47336 418120 47388
rect 471980 47336 472032 47388
rect 526812 47336 526864 47388
rect 199654 47268 199660 47320
rect 199712 47308 199718 47320
rect 199712 47280 276060 47308
rect 199712 47268 199718 47280
rect 217968 47200 218020 47252
rect 240140 47200 240192 47252
rect 276032 47240 276060 47280
rect 285588 47268 285640 47320
rect 307576 47268 307628 47320
rect 362408 47268 362460 47320
rect 364156 47268 364208 47320
rect 406752 47268 406804 47320
rect 461492 47268 461544 47320
rect 516324 47268 516376 47320
rect 518808 47268 518860 47320
rect 276032 47212 285720 47240
rect 200856 47132 200908 47184
rect 242900 47132 242952 47184
rect 149060 47064 149112 47116
rect 154580 47064 154632 47116
rect 173808 46996 173860 47048
rect 188528 47064 188580 47116
rect 192852 47064 192904 47116
rect 186688 46928 186740 46980
rect 194692 46928 194744 46980
rect 201408 47064 201460 47116
rect 247408 47064 247460 47116
rect 285588 47064 285640 47116
rect 285692 47104 285720 47212
rect 309416 47200 309468 47252
rect 352564 47200 352616 47252
rect 364248 47200 364300 47252
rect 407396 47200 407448 47252
rect 416780 47200 416832 47252
rect 417240 47200 417292 47252
rect 418068 47200 418120 47252
rect 419080 47200 419132 47252
rect 462136 47200 462188 47252
rect 473820 47200 473872 47252
rect 516968 47200 517020 47252
rect 299480 47132 299532 47184
rect 305736 47132 305788 47184
rect 351920 47132 351972 47184
rect 360568 47132 360620 47184
rect 406752 47132 406804 47184
rect 468294 47172 468300 47184
rect 417896 47144 468300 47172
rect 417896 47116 417924 47144
rect 468294 47132 468300 47144
rect 468352 47172 468358 47184
rect 527450 47172 527456 47184
rect 468352 47144 527456 47172
rect 468352 47132 468358 47144
rect 527450 47132 527456 47144
rect 527508 47132 527514 47184
rect 303890 47104 303896 47116
rect 285692 47076 303896 47104
rect 303890 47064 303896 47076
rect 303948 47104 303954 47116
rect 308214 47104 308220 47116
rect 303948 47076 308220 47104
rect 303948 47064 303954 47076
rect 308214 47064 308220 47076
rect 308272 47104 308278 47116
rect 358722 47104 358728 47116
rect 308272 47076 358728 47104
rect 308272 47064 308278 47076
rect 358722 47064 358728 47076
rect 358780 47104 358786 47116
rect 363046 47104 363052 47116
rect 358780 47076 363052 47104
rect 358780 47064 358786 47076
rect 363046 47064 363052 47076
rect 363104 47104 363110 47116
rect 413554 47104 413560 47116
rect 363104 47076 413560 47104
rect 363104 47064 363110 47076
rect 413554 47064 413560 47076
rect 413612 47104 413618 47116
rect 417878 47104 417884 47116
rect 413612 47076 417884 47104
rect 413612 47064 413618 47076
rect 417878 47064 417884 47076
rect 417936 47064 417942 47116
rect 417976 47064 418028 47116
rect 468944 47064 468996 47116
rect 523776 47064 523828 47116
rect 569132 47064 569184 47116
rect 201592 46996 201644 47048
rect 217968 46996 218020 47048
rect 514484 46928 514536 46980
rect 522488 46928 522540 46980
rect 526812 46928 526864 46980
rect 634820 46928 634872 46980
rect 42242 45636 42248 45688
rect 42300 45676 42306 45688
rect 145098 45676 145104 45688
rect 42300 45648 145104 45676
rect 42300 45636 42306 45648
rect 145098 45636 145104 45648
rect 145156 45636 145162 45688
rect 42708 45568 42760 45620
rect 140964 45568 141016 45620
rect 242900 45500 242952 45552
rect 297732 45500 297784 45552
rect 579160 45500 579212 45552
rect 673460 45500 673512 45552
rect 145098 44208 145104 44260
rect 145156 44248 145162 44260
rect 195330 44248 195336 44260
rect 145156 44220 195336 44248
rect 145156 44208 145162 44220
rect 195330 44208 195336 44220
rect 195388 44208 195394 44260
rect 140964 44140 141016 44192
rect 254032 44140 254084 44192
rect 569224 44140 569276 44192
rect 299480 41964 299532 42016
rect 302240 41964 302292 42016
rect 305000 41964 305052 42016
rect 411536 41964 411588 42016
rect 414572 41964 414624 42016
rect 415860 41964 415912 42016
rect 418252 41964 418304 42016
rect 466368 41964 466420 42016
rect 469404 41964 469456 42016
rect 470692 41964 470744 42016
rect 473084 41964 473136 42016
rect 189264 41828 189316 41880
rect 191104 41828 191156 41880
rect 192300 41828 192352 41880
rect 195422 41828 195428 41880
rect 195480 41868 195486 41880
rect 199562 41868 199568 41880
rect 195480 41840 199568 41868
rect 195480 41828 195486 41840
rect 199562 41828 199568 41840
rect 199620 41828 199626 41880
rect 193588 41760 193640 41812
rect 196440 41760 196492 41812
rect 198464 41760 198516 41812
rect 200120 41760 200172 41812
rect 253940 41556 253992 41608
rect 296904 41896 296956 41948
rect 352656 41896 352708 41948
rect 355508 41896 355560 41948
rect 356980 41896 357032 41948
rect 359832 41896 359884 41948
rect 361120 41896 361172 41948
rect 407488 41896 407540 41948
rect 410248 41896 410300 41948
rect 411162 41896 411168 41948
rect 411220 41936 411226 41948
rect 411220 41908 415624 41936
rect 411220 41896 411226 41908
rect 297916 41828 297968 41880
rect 300676 41828 300728 41880
rect 352012 41828 352064 41880
rect 354312 41828 354364 41880
rect 360476 41828 360528 41880
rect 295432 41760 295484 41812
rect 303160 41760 303212 41812
rect 305276 41760 305328 41812
rect 306564 41760 306616 41812
rect 308680 41760 308732 41812
rect 350172 41760 350224 41812
rect 357992 41760 358044 41812
rect 409322 41828 409328 41880
rect 409380 41868 409386 41880
rect 412358 41868 412364 41880
rect 409380 41840 412364 41868
rect 409380 41828 409386 41840
rect 412358 41828 412364 41840
rect 412416 41868 412422 41880
rect 415486 41868 415492 41880
rect 412416 41840 415492 41868
rect 412416 41828 412422 41840
rect 415486 41828 415492 41840
rect 415544 41828 415550 41880
rect 415596 41868 415624 41908
rect 462320 41896 462372 41948
rect 465080 41896 465132 41948
rect 465994 41896 466000 41948
rect 466052 41936 466058 41948
rect 474366 41936 474372 41948
rect 466052 41908 474372 41936
rect 466052 41896 466058 41908
rect 474366 41896 474372 41908
rect 474424 41896 474430 41948
rect 523218 41896 523224 41948
rect 523276 41936 523282 41948
rect 527358 41936 527364 41948
rect 523276 41908 527364 41936
rect 523276 41896 523282 41908
rect 527358 41896 527364 41908
rect 527416 41896 527422 41948
rect 419534 41868 419540 41880
rect 415596 41840 419540 41868
rect 419534 41828 419540 41840
rect 419592 41828 419598 41880
rect 459836 41828 459888 41880
rect 467564 41828 467616 41880
rect 468478 41828 468484 41880
rect 468536 41868 468542 41880
rect 472526 41868 472532 41880
rect 468536 41840 472532 41868
rect 468536 41828 468542 41840
rect 472526 41828 472532 41840
rect 472584 41828 472590 41880
rect 518894 41828 518900 41880
rect 518952 41868 518958 41880
rect 524874 41868 524880 41880
rect 518952 41840 524880 41868
rect 518952 41828 518958 41840
rect 524874 41828 524880 41840
rect 524932 41828 524938 41880
rect 363512 41760 363564 41812
rect 405004 41760 405056 41812
rect 412732 41760 412784 41812
rect 464154 41760 464160 41812
rect 464212 41800 464218 41812
rect 467190 41800 467196 41812
rect 464212 41772 467196 41800
rect 464212 41760 464218 41772
rect 467190 41760 467196 41772
rect 467248 41800 467254 41812
rect 470042 41800 470048 41812
rect 467248 41772 470048 41800
rect 467248 41760 467254 41772
rect 470042 41760 470048 41772
rect 470100 41760 470106 41812
rect 517060 41760 517112 41812
rect 520096 41760 520148 41812
rect 521384 41760 521436 41812
rect 524420 41760 524472 41812
rect 525708 41760 525760 41812
rect 527916 41760 527968 41812
rect 133098 40196 133150 40248
rect 143816 40196 143868 40248
rect 140996 40060 141048 40112
rect 143072 40060 143124 40112
rect 143356 40060 143408 40112
rect 252100 39652 252152 39704
rect 254032 39652 254084 39704
<< via1 >>
rect 463792 992264 463844 992316
rect 475476 992264 475528 992316
rect 482928 992264 482980 992316
rect 130292 990836 130344 990888
rect 79048 990768 79100 990820
rect 110420 990768 110472 990820
rect 130108 990768 130160 990820
rect 419540 990836 419592 990888
rect 438676 990836 438728 990888
rect 450268 990836 450320 990888
rect 463608 990836 463660 990888
rect 143264 990768 143316 990820
rect 173808 990768 173860 990820
rect 179328 990768 179380 990820
rect 246948 990768 247000 990820
rect 284668 990768 284720 990820
rect 286968 990768 287020 990820
rect 187608 990700 187660 990752
rect 187700 990700 187752 990752
rect 202880 990700 202932 990752
rect 233056 990700 233108 990752
rect 482928 990700 482980 990752
rect 526904 990700 526956 990752
rect 628656 990700 628708 990752
rect 110512 990564 110564 990616
rect 130108 990564 130160 990616
rect 179328 990564 179380 990616
rect 181720 990564 181772 990616
rect 386512 990564 386564 990616
rect 286968 990496 287020 990548
rect 419540 990564 419592 990616
rect 438768 990564 438820 990616
rect 450268 990564 450320 990616
rect 143264 990428 143316 990480
rect 160100 990428 160152 990480
rect 181720 990428 181772 990480
rect 187608 990428 187660 990480
rect 187700 990428 187752 990480
rect 202880 990428 202932 990480
rect 233056 990428 233108 990480
rect 246948 990428 247000 990480
rect 42432 990088 42484 990140
rect 79048 990088 79100 990140
rect 628656 990088 628708 990140
rect 673460 990020 673512 990072
rect 673460 965268 673512 965320
rect 675392 965268 675444 965320
rect 41788 956428 41840 956480
rect 42432 956428 42484 956480
rect 673184 908012 673236 908064
rect 673460 908012 673512 908064
rect 673184 888768 673236 888820
rect 673460 888768 673512 888820
rect 673736 869388 673788 869440
rect 675208 869388 675260 869440
rect 673552 836272 673604 836324
rect 673644 836204 673696 836256
rect 673552 830764 673604 830816
rect 673644 830764 673696 830816
rect 673552 821040 673604 821092
rect 674104 821040 674156 821092
rect 674104 797580 674156 797632
rect 675300 797580 675352 797632
rect 42248 787176 42300 787228
rect 42616 787176 42668 787228
rect 674012 786428 674064 786480
rect 675300 786428 675352 786480
rect 673552 768612 673604 768664
rect 674012 768612 674064 768664
rect 41788 744404 41840 744456
rect 42616 744404 42668 744456
rect 673552 741888 673604 741940
rect 674196 741888 674248 741940
rect 675392 741888 675444 741940
rect 674012 720400 674064 720452
rect 674196 720400 674248 720452
rect 674012 710676 674064 710728
rect 675300 710676 675352 710728
rect 41788 700816 41840 700868
rect 42616 700816 42668 700868
rect 673644 695920 673696 695972
rect 675392 695920 675444 695972
rect 41788 657092 41840 657144
rect 42340 657092 42392 657144
rect 42616 657092 42668 657144
rect 673644 651720 673696 651772
rect 675392 651720 675444 651772
rect 42340 633224 42392 633276
rect 42616 633224 42668 633276
rect 41880 614456 41932 614508
rect 42248 614456 42300 614508
rect 42616 614456 42668 614508
rect 673644 606704 673696 606756
rect 675392 606704 675444 606756
rect 42248 584196 42300 584248
rect 42616 584196 42668 584248
rect 41788 571616 41840 571668
rect 42616 571616 42668 571668
rect 673644 561484 673696 561536
rect 675392 561484 675444 561536
rect 41788 528436 41840 528488
rect 42432 528436 42484 528488
rect 42616 528436 42668 528488
rect 41972 400120 42024 400172
rect 42432 400120 42484 400172
rect 673552 384004 673604 384056
rect 675392 384004 675444 384056
rect 41788 356668 41840 356720
rect 42432 356668 42484 356720
rect 41788 313760 41840 313812
rect 42432 313760 42484 313812
rect 42432 307912 42484 307964
rect 42708 307912 42760 307964
rect 673828 293156 673880 293208
rect 675392 293156 675444 293208
rect 42708 282208 42760 282260
rect 42708 282004 42760 282056
rect 41788 270240 41840 270292
rect 42340 270240 42392 270292
rect 42708 270240 42760 270292
rect 673828 248140 673880 248192
rect 675392 248140 675444 248192
rect 42340 246984 42392 247036
rect 42708 246984 42760 247036
rect 41788 228012 41840 228064
rect 42432 228012 42484 228064
rect 42708 228012 42760 228064
rect 673552 203872 673604 203924
rect 673828 203872 673880 203924
rect 675392 203872 675444 203924
rect 42248 184220 42300 184272
rect 42432 184220 42484 184272
rect 673552 158312 673604 158364
rect 675392 158312 675444 158364
rect 673552 112752 673604 112804
rect 675392 112752 675444 112804
rect 527456 47812 527508 47864
rect 673552 47812 673604 47864
rect 199660 47268 199712 47320
rect 468300 47132 468352 47184
rect 527456 47132 527508 47184
rect 303896 47064 303948 47116
rect 308220 47064 308272 47116
rect 358728 47064 358780 47116
rect 363052 47064 363104 47116
rect 413560 47064 413612 47116
rect 417884 47064 417936 47116
rect 42248 45636 42300 45688
rect 145104 45636 145156 45688
rect 145104 44208 145156 44260
rect 195336 44208 195388 44260
rect 195428 41828 195480 41880
rect 199568 41828 199620 41880
rect 411168 41896 411220 41948
rect 409328 41828 409380 41880
rect 412364 41828 412416 41880
rect 415492 41828 415544 41880
rect 466000 41896 466052 41948
rect 474372 41896 474424 41948
rect 523224 41896 523276 41948
rect 527364 41896 527416 41948
rect 419540 41828 419592 41880
rect 468484 41828 468536 41880
rect 472532 41828 472584 41880
rect 518900 41828 518952 41880
rect 524880 41828 524932 41880
rect 464160 41760 464212 41812
rect 467196 41760 467248 41812
rect 470048 41760 470100 41812
<< obsm1 >>
rect 76171 996231 92229 1037600
rect 127571 996231 143629 1037600
rect 178971 996231 195029 1037600
rect 230371 996231 246429 1037600
rect 281971 996231 298029 1037600
rect 333437 998007 348124 1037545
rect 383771 996231 399829 1037600
rect 472771 996231 488829 1037600
rect 524171 996231 540229 1037600
rect 575637 998007 590324 1037545
rect 625971 996231 642029 1037600
rect 84010 995596 84016 995648
rect 84068 995636 84074 995648
rect 91738 995636 91744 995648
rect 84068 995608 91744 995636
rect 84068 995596 84074 995608
rect 91738 995596 91744 995608
rect 91796 995596 91802 995648
rect 238202 995596 238208 995648
rect 238260 995636 238266 995648
rect 245930 995636 245936 995648
rect 238260 995608 245936 995636
rect 238260 995596 238266 995608
rect 245930 995596 245936 995608
rect 245988 995596 245994 995648
rect 531958 995596 531964 995648
rect 532016 995636 532022 995648
rect 539686 995636 539692 995648
rect 532016 995608 539692 995636
rect 532016 995596 532022 995608
rect 539686 995596 539692 995608
rect 539744 995596 539750 995648
rect 135346 995460 135352 995512
rect 135404 995500 135410 995512
rect 143166 995500 143172 995512
rect 135404 995472 143172 995500
rect 135404 995460 135410 995472
rect 143166 995460 143172 995472
rect 143224 995460 143230 995512
rect 633802 995460 633808 995512
rect 633860 995500 633866 995512
rect 641530 995500 641536 995512
rect 633860 995472 641536 995500
rect 633860 995460 633866 995472
rect 641530 995460 641536 995472
rect 641588 995460 641594 995512
rect 289630 995256 289636 995308
rect 289688 995296 289694 995308
rect 297634 995296 297640 995308
rect 289688 995268 297640 995296
rect 289688 995256 289694 995268
rect 297634 995256 297640 995268
rect 297692 995256 297698 995308
rect 391474 995256 391480 995308
rect 391532 995296 391538 995308
rect 399478 995296 399484 995308
rect 391532 995268 399484 995296
rect 391532 995256 391538 995268
rect 399478 995256 399484 995268
rect 399536 995256 399542 995308
rect 480438 995256 480444 995308
rect 480496 995296 480502 995308
rect 488442 995296 488448 995308
rect 480496 995268 488448 995296
rect 480496 995256 480502 995268
rect 488442 995256 488448 995268
rect 488500 995256 488506 995308
rect 231854 995052 231860 995104
rect 231912 995092 231918 995104
rect 244182 995092 244188 995104
rect 231912 995064 244188 995092
rect 231912 995052 231918 995064
rect 244182 995052 244188 995064
rect 244240 995052 244246 995104
rect 141418 992060 141424 992112
rect 141476 992100 141482 992112
rect 154390 992100 154396 992112
rect 141476 992072 154396 992100
rect 141476 992060 141482 992072
rect 154390 992060 154396 992072
rect 154448 992060 154454 992112
rect 391750 990768 391756 990820
rect 391808 990808 391814 990820
rect 476114 990808 476120 990820
rect 391808 990780 476120 990808
rect 391808 990768 391814 990780
rect 476114 990768 476120 990780
rect 476172 990808 476178 990820
rect 527542 990808 527548 990820
rect 476172 990780 527548 990808
rect 476172 990768 476178 990780
rect 527542 990768 527548 990780
rect 527600 990808 527606 990820
rect 629294 990808 629300 990820
rect 527600 990780 629300 990808
rect 527600 990768 527606 990780
rect 629294 990768 629300 990780
rect 629352 990768 629358 990820
rect 244182 990700 244188 990752
rect 244240 990740 244246 990752
rect 295794 990740 295800 990752
rect 244240 990712 295800 990740
rect 244240 990700 244246 990712
rect 295794 990700 295800 990712
rect 295852 990740 295858 990752
rect 386322 990740 386328 990752
rect 295852 990712 386328 990740
rect 295852 990700 295858 990712
rect 386322 990700 386328 990712
rect 386380 990700 386386 990752
rect 79502 990632 79508 990684
rect 79560 990672 79566 990684
rect 79962 990672 79968 990684
rect 79560 990644 79968 990672
rect 79560 990632 79566 990644
rect 79962 990632 79968 990644
rect 80020 990672 80026 990684
rect 130930 990672 130936 990684
rect 80020 990644 130936 990672
rect 80020 990632 80026 990644
rect 130930 990632 130936 990644
rect 130988 990672 130994 990684
rect 182358 990672 182364 990684
rect 130988 990644 182364 990672
rect 130988 990632 130994 990644
rect 182358 990632 182364 990644
rect 182416 990672 182422 990684
rect 233694 990672 233700 990684
rect 182416 990644 233700 990672
rect 182416 990632 182422 990644
rect 233694 990632 233700 990644
rect 233752 990672 233758 990684
rect 285306 990672 285312 990684
rect 233752 990644 285312 990672
rect 233752 990632 233758 990644
rect 285306 990632 285312 990644
rect 285364 990672 285370 990684
rect 333514 990672 333520 990684
rect 285364 990644 333520 990672
rect 285364 990632 285370 990644
rect 333514 990632 333520 990644
rect 333572 990672 333578 990684
rect 387150 990672 387156 990684
rect 333572 990644 387156 990672
rect 333572 990632 333578 990644
rect 387150 990632 387156 990644
rect 387208 990672 387214 990684
rect 391750 990672 391756 990684
rect 387208 990644 391756 990672
rect 387208 990632 387214 990644
rect 391750 990632 391756 990644
rect 391808 990632 391814 990684
rect 89990 990564 89996 990616
rect 90048 990604 90054 990616
rect 90048 990576 91140 990604
rect 90048 990564 90054 990576
rect 91112 990536 91140 990576
rect 186682 990564 186688 990616
rect 186740 990604 186746 990616
rect 194686 990604 194692 990616
rect 186740 990576 194692 990604
rect 186740 990564 186746 990576
rect 194686 990564 194692 990576
rect 194744 990564 194750 990616
rect 91112 990508 110368 990536
rect 110340 990468 110368 990508
rect 164142 990496 164148 990548
rect 164200 990536 164206 990548
rect 192846 990536 192852 990548
rect 164200 990508 192852 990536
rect 164200 990496 164206 990508
rect 192846 990496 192852 990508
rect 192904 990536 192910 990548
rect 193214 990536 193220 990548
rect 192904 990508 193220 990536
rect 192904 990496 192910 990508
rect 193214 990496 193220 990508
rect 193272 990496 193278 990548
rect 212442 990496 212448 990548
rect 212500 990536 212506 990548
rect 231854 990536 231860 990548
rect 212500 990508 231860 990536
rect 212500 990496 212506 990508
rect 231854 990496 231860 990508
rect 231912 990496 231918 990548
rect 596082 990632 596088 990684
rect 596140 990672 596146 990684
rect 596140 990644 598980 990672
rect 596140 990632 596146 990644
rect 469306 990564 469312 990616
rect 469364 990604 469370 990616
rect 576854 990604 576860 990616
rect 469364 990576 483060 990604
rect 469364 990564 469370 990576
rect 483032 990548 483060 990576
rect 565740 990576 576860 990604
rect 469030 990536 469036 990548
rect 449820 990508 469036 990536
rect 141326 990468 141332 990480
rect 110340 990440 141332 990468
rect 141326 990428 141332 990440
rect 141384 990428 141390 990480
rect 449820 990468 449848 990508
rect 469030 990496 469036 990508
rect 469088 990496 469094 990548
rect 483014 990496 483020 990548
rect 483072 990496 483078 990548
rect 560202 990496 560208 990548
rect 560260 990536 560266 990548
rect 565740 990536 565768 990576
rect 576854 990564 576860 990576
rect 576912 990564 576918 990616
rect 560260 990508 565768 990536
rect 598952 990536 598980 990644
rect 623682 990604 623688 990616
rect 604564 990576 623688 990604
rect 604564 990536 604592 990576
rect 623682 990564 623688 990576
rect 623740 990564 623746 990616
rect 598952 990508 604592 990536
rect 560260 990496 560266 990508
rect 623866 990496 623872 990548
rect 623924 990536 623930 990548
rect 639782 990536 639788 990548
rect 623924 990508 639788 990536
rect 623924 990496 623930 990508
rect 639782 990496 639788 990508
rect 639840 990496 639846 990548
rect 540974 990468 540980 990480
rect 430592 990440 449848 990468
rect 540900 990440 540980 990468
rect 154390 990360 154396 990412
rect 154448 990400 154454 990412
rect 154574 990400 154580 990412
rect 154448 990372 154580 990400
rect 154448 990360 154454 990372
rect 154574 990360 154580 990372
rect 154632 990360 154638 990412
rect 386322 990360 386328 990412
rect 386380 990400 386386 990412
rect 397638 990400 397644 990412
rect 386380 990372 397644 990400
rect 386380 990360 386386 990372
rect 397638 990360 397644 990372
rect 397696 990360 397702 990412
rect 424962 990360 424968 990412
rect 425020 990400 425026 990412
rect 430592 990400 430620 990440
rect 540900 990412 540928 990440
rect 540974 990428 540980 990440
rect 541032 990428 541038 990480
rect 425020 990372 430620 990400
rect 425020 990360 425026 990372
rect 483014 990360 483020 990412
rect 483072 990400 483078 990412
rect 486602 990400 486608 990412
rect 483072 990372 486608 990400
rect 483072 990360 483078 990372
rect 486602 990360 486608 990372
rect 486660 990400 486666 990412
rect 521654 990400 521660 990412
rect 486660 990372 502288 990400
rect 486660 990360 486666 990372
rect 502260 990332 502288 990372
rect 511920 990372 521660 990400
rect 507762 990332 507768 990344
rect 502260 990304 507768 990332
rect 507762 990292 507768 990304
rect 507820 990292 507826 990344
rect 507854 990292 507860 990344
rect 507912 990332 507918 990344
rect 511920 990332 511948 990372
rect 521654 990360 521660 990372
rect 521712 990360 521718 990412
rect 540882 990360 540888 990412
rect 540940 990360 540946 990412
rect 507912 990304 511948 990332
rect 507912 990292 507918 990304
rect 154574 990224 154580 990276
rect 154632 990264 154638 990276
rect 164142 990264 164148 990276
rect 154632 990236 164148 990264
rect 154632 990224 154638 990236
rect 164142 990224 164148 990236
rect 164200 990224 164206 990276
rect 397638 990224 397644 990276
rect 397696 990264 397702 990276
rect 405734 990264 405740 990276
rect 397696 990236 405740 990264
rect 397696 990224 397702 990236
rect 405734 990224 405740 990236
rect 405792 990224 405798 990276
rect 521654 990224 521660 990276
rect 521712 990264 521718 990276
rect 537846 990264 537852 990276
rect 521712 990236 537852 990264
rect 521712 990224 521718 990236
rect 537846 990224 537852 990236
rect 537904 990264 537910 990276
rect 540882 990264 540888 990276
rect 537904 990236 540888 990264
rect 537904 990224 537910 990236
rect 540882 990224 540888 990236
rect 540940 990224 540946 990276
rect 42242 990156 42248 990208
rect 42300 990196 42306 990208
rect 79962 990196 79968 990208
rect 42300 990168 79968 990196
rect 42300 990156 42306 990168
rect 79962 990156 79968 990168
rect 80020 990156 80026 990208
rect 639782 990156 639788 990208
rect 639840 990196 639846 990208
rect 673638 990196 673644 990208
rect 639840 990168 673644 990196
rect 639840 990156 639846 990168
rect 673638 990156 673644 990168
rect 673696 990156 673702 990208
rect 89990 990088 89996 990140
rect 90048 990088 90054 990140
rect 405734 990088 405740 990140
rect 405792 990128 405798 990140
rect 424962 990128 424968 990140
rect 405792 990100 424968 990128
rect 405792 990088 405798 990100
rect 424962 990088 424968 990100
rect 425020 990088 425026 990140
rect 629294 990088 629300 990140
rect 629352 990128 629358 990140
rect 673546 990128 673552 990140
rect 629352 990100 673552 990128
rect 629352 990088 629358 990100
rect 673546 990088 673552 990100
rect 673604 990088 673610 990140
rect 42518 990020 42524 990072
rect 42576 990060 42582 990072
rect 90008 990060 90036 990088
rect 42576 990032 90036 990060
rect 42576 990020 42582 990032
rect 0 954171 41369 970229
rect 41782 969348 41788 969400
rect 41840 969388 41846 969400
rect 42334 969388 42340 969400
rect 41840 969360 42340 969388
rect 41840 969348 41846 969360
rect 42334 969348 42340 969360
rect 42392 969348 42398 969400
rect 41782 968464 41788 968516
rect 41840 968504 41846 968516
rect 42518 968504 42524 968516
rect 41840 968476 42524 968504
rect 41840 968464 41846 968476
rect 42518 968464 42524 968476
rect 42576 968464 42582 968516
rect 673546 964724 673552 964776
rect 673604 964764 673610 964776
rect 675386 964764 675392 964776
rect 673604 964736 675392 964764
rect 673604 964724 673610 964736
rect 675386 964724 675392 964736
rect 675444 964724 675450 964776
rect 41782 962412 41788 962464
rect 41840 962452 41846 962464
rect 42334 962452 42340 962464
rect 41840 962424 42340 962452
rect 41840 962412 41846 962424
rect 42334 962412 42340 962424
rect 42392 962412 42398 962464
rect 673638 953300 673644 953352
rect 673696 953340 673702 953352
rect 675386 953340 675392 953352
rect 673696 953312 675392 953340
rect 673696 953300 673702 953312
rect 675386 953300 675392 953312
rect 675444 953300 675450 953352
rect 676231 951571 717600 967629
rect 44266 930112 44272 930164
rect 44324 930152 44330 930164
rect 45462 930152 45468 930164
rect 44324 930124 45468 930152
rect 44324 930112 44330 930124
rect 45462 930112 45468 930124
rect 45520 930112 45526 930164
rect 32 912024 39593 926957
rect 39666 922904 39672 922956
rect 39724 922944 39730 922956
rect 44266 922944 44272 922956
rect 39724 922916 44272 922944
rect 39724 922904 39730 922916
rect 44266 922904 44272 922916
rect 44324 922904 44330 922956
rect 39850 914676 39856 914728
rect 39908 914716 39914 914728
rect 41414 914716 41420 914728
rect 39908 914688 41420 914716
rect 39908 914676 39914 914688
rect 41414 914676 41420 914688
rect 41472 914716 41478 914728
rect 42242 914716 42248 914728
rect 41472 914688 42248 914716
rect 41472 914676 41478 914688
rect 42242 914676 42248 914688
rect 42300 914676 42306 914728
rect 673546 910732 673552 910784
rect 673604 910772 673610 910784
rect 677778 910772 677784 910784
rect 673604 910744 677784 910772
rect 673604 910732 673610 910744
rect 677778 910732 677784 910744
rect 677836 910732 677842 910784
rect 678007 907643 717568 922576
rect 55 869837 39593 884383
rect 39850 879792 39856 879844
rect 39908 879832 39914 879844
rect 40126 879832 40132 879844
rect 39908 879804 40132 879832
rect 39908 879792 39914 879804
rect 40126 879792 40132 879804
rect 40184 879832 40190 879844
rect 44174 879832 44180 879844
rect 40184 879804 44180 879832
rect 40184 879792 40190 879804
rect 44174 879792 44180 879804
rect 44232 879832 44238 879844
rect 45830 879832 45836 879844
rect 44232 879804 45836 879832
rect 44232 879792 44238 879804
rect 45830 879792 45836 879804
rect 45888 879792 45894 879844
rect 41414 875576 41420 875628
rect 41472 875616 41478 875628
rect 42242 875616 42248 875628
rect 41472 875588 42248 875616
rect 41472 875576 41478 875588
rect 42242 875576 42248 875588
rect 42300 875576 42306 875628
rect 673546 875508 673552 875560
rect 673604 875548 673610 875560
rect 675386 875548 675392 875560
rect 673604 875520 675392 875548
rect 673604 875508 673610 875520
rect 675386 875508 675392 875520
rect 675444 875508 675450 875560
rect 673638 875032 673644 875084
rect 673696 875032 673702 875084
rect 673656 874948 673684 875032
rect 673638 874896 673644 874948
rect 673696 874896 673702 874948
rect 673638 864968 673644 865020
rect 673696 865008 673702 865020
rect 673822 865008 673828 865020
rect 673696 864980 673828 865008
rect 673696 864968 673702 864980
rect 673822 864968 673828 864980
rect 673880 865008 673886 865020
rect 675386 865008 675392 865020
rect 673880 864980 675392 865008
rect 673880 864968 673886 864980
rect 675386 864968 675392 864980
rect 675444 864968 675450 865020
rect 676231 862371 717600 878429
rect 55 827637 39593 842324
rect 678007 818817 717545 833363
rect 42242 807304 42248 807356
rect 42300 807344 42306 807356
rect 42702 807344 42708 807356
rect 42300 807316 42708 807344
rect 42300 807304 42306 807316
rect 42702 807304 42708 807316
rect 42760 807304 42766 807356
rect 44542 805944 44548 805996
rect 44600 805984 44606 805996
rect 44726 805984 44732 805996
rect 44600 805956 44732 805984
rect 44600 805944 44606 805956
rect 44726 805944 44732 805956
rect 44784 805944 44790 805996
rect 0 784371 41369 800429
rect 41782 798328 41788 798380
rect 41840 798368 41846 798380
rect 42518 798368 42524 798380
rect 41840 798340 42524 798368
rect 41840 798328 41846 798340
rect 42518 798328 42524 798340
rect 42576 798328 42582 798380
rect 41782 787856 41788 787908
rect 41840 787896 41846 787908
rect 42426 787896 42432 787908
rect 41840 787868 42432 787896
rect 41840 787856 41846 787868
rect 42426 787856 42432 787868
rect 42484 787896 42490 787908
rect 42702 787896 42708 787908
rect 42484 787868 42708 787896
rect 42484 787856 42490 787868
rect 42702 787856 42708 787868
rect 42760 787856 42766 787908
rect 673638 785272 673644 785324
rect 673696 785312 673702 785324
rect 675386 785312 675392 785324
rect 673696 785284 675392 785312
rect 673696 785272 673702 785284
rect 675386 785272 675392 785284
rect 675444 785272 675450 785324
rect 672994 778336 673000 778388
rect 673052 778336 673058 778388
rect 673012 778240 673040 778336
rect 673086 778240 673092 778252
rect 673012 778212 673092 778240
rect 673086 778200 673092 778212
rect 673144 778200 673150 778252
rect 673454 774868 673460 774920
rect 673512 774908 673518 774920
rect 673822 774908 673828 774920
rect 673512 774880 673828 774908
rect 673512 774868 673518 774880
rect 673822 774868 673828 774880
rect 673880 774908 673886 774920
rect 675386 774908 675392 774920
rect 673880 774880 675392 774908
rect 673880 774868 673886 774880
rect 675386 774868 675392 774880
rect 675444 774868 675450 774920
rect 676231 773171 717600 789229
rect 672810 772760 672816 772812
rect 672868 772800 672874 772812
rect 673086 772800 673092 772812
rect 672868 772772 673092 772800
rect 672868 772760 672874 772772
rect 673086 772760 673092 772772
rect 673144 772760 673150 772812
rect 42518 768612 42524 768664
rect 42576 768652 42582 768664
rect 42702 768652 42708 768664
rect 42576 768624 42708 768652
rect 42576 768612 42582 768624
rect 42702 768612 42708 768624
rect 42760 768612 42766 768664
rect 0 741171 41369 757229
rect 41782 754468 41788 754520
rect 41840 754508 41846 754520
rect 42518 754508 42524 754520
rect 41840 754480 42524 754508
rect 41840 754468 41846 754480
rect 42518 754468 42524 754480
rect 42576 754508 42582 754520
rect 42702 754508 42708 754520
rect 42576 754480 42708 754508
rect 42576 754468 42582 754480
rect 42702 754468 42708 754480
rect 42760 754468 42766 754520
rect 673638 741344 673644 741396
rect 673696 741384 673702 741396
rect 675386 741384 675392 741396
rect 673696 741356 675392 741384
rect 673696 741344 673702 741356
rect 675386 741344 675392 741356
rect 675444 741344 675450 741396
rect 672994 739712 673000 739764
rect 673052 739712 673058 739764
rect 673012 739616 673040 739712
rect 673178 739616 673184 739628
rect 673012 739588 673184 739616
rect 673178 739576 673184 739588
rect 673236 739576 673242 739628
rect 673454 730124 673460 730176
rect 673512 730164 673518 730176
rect 675386 730164 675392 730176
rect 673512 730136 675392 730164
rect 673512 730124 673518 730136
rect 675386 730124 675392 730136
rect 675444 730124 675450 730176
rect 673822 729988 673828 730040
rect 673880 730028 673886 730040
rect 675110 730028 675116 730040
rect 673880 730000 675116 730028
rect 673880 729988 673886 730000
rect 675110 729988 675116 730000
rect 675168 729988 675174 730040
rect 676231 728171 717600 744229
rect 0 697971 41369 714029
rect 41782 711288 41788 711340
rect 41840 711328 41846 711340
rect 42518 711328 42524 711340
rect 41840 711300 42524 711328
rect 41840 711288 41846 711300
rect 42518 711288 42524 711300
rect 42576 711288 42582 711340
rect 42242 700952 42248 701004
rect 42300 700992 42306 701004
rect 42518 700992 42524 701004
rect 42300 700964 42524 700992
rect 42300 700952 42306 700964
rect 42518 700952 42524 700964
rect 42576 700952 42582 701004
rect 673086 695512 673092 695564
rect 673144 695552 673150 695564
rect 673178 695552 673184 695564
rect 673144 695524 673184 695552
rect 673144 695512 673150 695524
rect 673178 695512 673184 695524
rect 673236 695512 673242 695564
rect 44634 695444 44640 695496
rect 44692 695484 44698 695496
rect 44910 695484 44916 695496
rect 44692 695456 44916 695484
rect 44692 695444 44698 695456
rect 44910 695444 44916 695456
rect 44968 695444 44974 695496
rect 673546 695308 673552 695360
rect 673604 695348 673610 695360
rect 673822 695348 673828 695360
rect 673604 695320 673828 695348
rect 673604 695308 673610 695320
rect 673822 695308 673828 695320
rect 673880 695348 673886 695360
rect 675386 695348 675392 695360
rect 673880 695320 675392 695348
rect 673880 695308 673886 695320
rect 675386 695308 675392 695320
rect 675444 695308 675450 695360
rect 676231 683171 717600 699229
rect 44726 676200 44732 676252
rect 44784 676240 44790 676252
rect 44910 676240 44916 676252
rect 44784 676212 44916 676240
rect 44784 676200 44790 676212
rect 44910 676200 44916 676212
rect 44968 676200 44974 676252
rect 0 654771 41369 670829
rect 42334 669168 42340 669180
rect 41800 669140 42340 669168
rect 41800 669112 41828 669140
rect 42334 669128 42340 669140
rect 42392 669128 42398 669180
rect 41782 669060 41788 669112
rect 41840 669060 41846 669112
rect 673178 662464 673184 662516
rect 673236 662464 673242 662516
rect 44542 662396 44548 662448
rect 44600 662436 44606 662448
rect 44726 662436 44732 662448
rect 44600 662408 44732 662436
rect 44600 662396 44606 662408
rect 44726 662396 44732 662408
rect 44784 662396 44790 662448
rect 673196 662380 673224 662464
rect 673178 662328 673184 662380
rect 673236 662328 673242 662380
rect 41782 657636 41788 657688
rect 41840 657676 41846 657688
rect 42518 657676 42524 657688
rect 41840 657648 42524 657676
rect 41840 657636 41846 657648
rect 42518 657636 42524 657648
rect 42576 657636 42582 657688
rect 44634 656820 44640 656872
rect 44692 656860 44698 656872
rect 44818 656860 44824 656872
rect 44692 656832 44824 656860
rect 44692 656820 44698 656832
rect 44818 656820 44824 656832
rect 44876 656820 44882 656872
rect 673546 651108 673552 651160
rect 673604 651148 673610 651160
rect 675386 651148 675392 651160
rect 673604 651120 675392 651148
rect 673604 651108 673610 651120
rect 675386 651108 675392 651120
rect 675444 651108 675450 651160
rect 673454 639684 673460 639736
rect 673512 639724 673518 639736
rect 675386 639724 675392 639736
rect 673512 639696 675392 639724
rect 673512 639684 673518 639696
rect 675386 639684 675392 639696
rect 675444 639684 675450 639736
rect 676231 637971 717600 654029
rect 672810 637508 672816 637560
rect 672868 637548 672874 637560
rect 673086 637548 673092 637560
rect 672868 637520 673092 637548
rect 672868 637508 672874 637520
rect 673086 637508 673092 637520
rect 673144 637508 673150 637560
rect 42518 633496 42524 633548
rect 42576 633496 42582 633548
rect 42536 633344 42564 633496
rect 42518 633292 42524 633344
rect 42576 633292 42582 633344
rect 0 611571 41369 627629
rect 41782 625880 41788 625932
rect 41840 625920 41846 625932
rect 42426 625920 42432 625932
rect 41840 625892 42432 625920
rect 41840 625880 41846 625892
rect 42426 625880 42432 625892
rect 42484 625880 42490 625932
rect 672810 618264 672816 618316
rect 672868 618304 672874 618316
rect 672994 618304 673000 618316
rect 672868 618276 673000 618304
rect 672868 618264 672874 618276
rect 672994 618264 673000 618276
rect 673052 618264 673058 618316
rect 41782 614388 41788 614440
rect 41840 614428 41846 614440
rect 42518 614428 42524 614440
rect 41840 614400 42524 614428
rect 41840 614388 41846 614400
rect 42518 614388 42524 614400
rect 42576 614388 42582 614440
rect 673546 605616 673552 605668
rect 673604 605656 673610 605668
rect 675294 605656 675300 605668
rect 673604 605628 675300 605656
rect 673604 605616 673610 605628
rect 675294 605616 675300 605628
rect 675352 605616 675358 605668
rect 44634 604528 44640 604580
rect 44692 604528 44698 604580
rect 44652 604444 44680 604528
rect 44634 604392 44640 604444
rect 44692 604392 44698 604444
rect 673546 604392 673552 604444
rect 673604 604432 673610 604444
rect 673822 604432 673828 604444
rect 673604 604404 673828 604432
rect 673604 604392 673610 604404
rect 673822 604392 673828 604404
rect 673880 604392 673886 604444
rect 672810 598952 672816 599004
rect 672868 598992 672874 599004
rect 673086 598992 673092 599004
rect 672868 598964 673092 598992
rect 672868 598952 672874 598964
rect 673086 598952 673092 598964
rect 673144 598952 673150 599004
rect 673454 594872 673460 594924
rect 673512 594912 673518 594924
rect 675386 594912 675392 594924
rect 673512 594884 675392 594912
rect 673512 594872 673518 594884
rect 675386 594872 675392 594884
rect 675444 594872 675450 594924
rect 676231 592971 717600 609029
rect 673086 585188 673092 585200
rect 673012 585160 673092 585188
rect 673012 585132 673040 585160
rect 673086 585148 673092 585160
rect 673144 585148 673150 585200
rect 672994 585080 673000 585132
rect 673052 585080 673058 585132
rect 0 568371 41369 584429
rect 41782 581680 41788 581732
rect 41840 581720 41846 581732
rect 42426 581720 42432 581732
rect 41840 581692 42432 581720
rect 41840 581680 41846 581692
rect 42426 581680 42432 581692
rect 42484 581680 42490 581732
rect 41782 572228 41788 572280
rect 41840 572268 41846 572280
rect 42242 572268 42248 572280
rect 41840 572240 42248 572268
rect 41840 572228 41846 572240
rect 42242 572228 42248 572240
rect 42300 572268 42306 572280
rect 42518 572268 42524 572280
rect 42300 572240 42524 572268
rect 42300 572228 42306 572240
rect 42518 572228 42524 572240
rect 42576 572228 42582 572280
rect 672810 569916 672816 569968
rect 672868 569956 672874 569968
rect 672994 569956 673000 569968
rect 672868 569928 673000 569956
rect 672868 569916 672874 569928
rect 672994 569916 673000 569928
rect 673052 569916 673058 569968
rect 673546 565836 673552 565888
rect 673604 565876 673610 565888
rect 673914 565876 673920 565888
rect 673604 565848 673920 565876
rect 673604 565836 673610 565848
rect 673914 565836 673920 565848
rect 673972 565836 673978 565888
rect 672810 560260 672816 560312
rect 672868 560300 672874 560312
rect 672994 560300 673000 560312
rect 672868 560272 673000 560300
rect 672868 560260 672874 560272
rect 672994 560260 673000 560272
rect 673052 560260 673058 560312
rect 673546 559920 673552 559972
rect 673604 559960 673610 559972
rect 673914 559960 673920 559972
rect 673604 559932 673920 559960
rect 673604 559920 673610 559932
rect 673914 559920 673920 559932
rect 673972 559960 673978 559972
rect 675386 559960 675392 559972
rect 673972 559932 675392 559960
rect 673972 559920 673978 559932
rect 675386 559920 675392 559932
rect 675444 559920 675450 559972
rect 673454 550468 673460 550520
rect 673512 550508 673518 550520
rect 675386 550508 675392 550520
rect 673512 550480 675392 550508
rect 673512 550468 673518 550480
rect 675386 550468 675392 550480
rect 675444 550468 675450 550520
rect 676231 547771 717600 563829
rect 672994 546524 673000 546576
rect 673052 546564 673058 546576
rect 673052 546536 673132 546564
rect 673052 546524 673058 546536
rect 673104 546372 673132 546536
rect 673086 546320 673092 546372
rect 673144 546320 673150 546372
rect 0 525171 41369 541229
rect 44726 540948 44732 541000
rect 44784 540988 44790 541000
rect 44910 540988 44916 541000
rect 44784 540960 44916 540988
rect 44784 540948 44790 540960
rect 44910 540948 44916 540960
rect 44968 540948 44974 541000
rect 41782 538500 41788 538552
rect 41840 538540 41846 538552
rect 42426 538540 42432 538552
rect 41840 538512 42432 538540
rect 41840 538500 41846 538512
rect 42426 538500 42432 538512
rect 42484 538500 42490 538552
rect 673086 527144 673092 527196
rect 673144 527144 673150 527196
rect 673104 527048 673132 527144
rect 673178 527048 673184 527060
rect 673104 527020 673184 527048
rect 673178 527008 673184 527020
rect 673236 527008 673242 527060
rect 673730 522928 673736 522980
rect 673788 522968 673794 522980
rect 673914 522968 673920 522980
rect 673788 522940 673920 522968
rect 673788 522928 673794 522940
rect 673914 522928 673920 522940
rect 673972 522928 673978 522980
rect 673178 521568 673184 521620
rect 673236 521608 673242 521620
rect 676122 521608 676128 521620
rect 673236 521580 676128 521608
rect 673236 521568 673242 521580
rect 676122 521568 676128 521580
rect 676180 521568 676186 521620
rect 678007 504217 717545 518763
rect 55 483037 39593 497583
rect 44542 496816 44548 496868
rect 44600 496856 44606 496868
rect 44726 496856 44732 496868
rect 44600 496828 44732 496856
rect 44600 496816 44606 496828
rect 44726 496816 44732 496828
rect 44784 496816 44790 496868
rect 673730 463632 673736 463684
rect 673788 463672 673794 463684
rect 677686 463672 677692 463684
rect 673788 463644 677692 463672
rect 673788 463632 673794 463644
rect 677686 463632 677692 463644
rect 677744 463632 677750 463684
rect 678007 459843 717568 474776
rect 39390 458192 39396 458244
rect 39448 458232 39454 458244
rect 44266 458232 44272 458244
rect 39448 458204 44272 458232
rect 39448 458192 39454 458204
rect 44266 458192 44272 458204
rect 44324 458192 44330 458244
rect 32 440824 39593 455757
rect 672994 449896 673000 449948
rect 673052 449936 673058 449948
rect 673362 449936 673368 449948
rect 673052 449908 673368 449936
rect 673052 449896 673058 449908
rect 673362 449896 673368 449908
rect 673420 449896 673426 449948
rect 39850 448264 39856 448316
rect 39908 448304 39914 448316
rect 42242 448304 42248 448316
rect 39908 448276 42248 448304
rect 39908 448264 39914 448276
rect 42242 448264 42248 448276
rect 42300 448264 42306 448316
rect 676214 440172 676220 440224
rect 676272 440212 676278 440224
rect 677686 440212 677692 440224
rect 676272 440184 677692 440212
rect 676272 440172 676278 440184
rect 677686 440172 677692 440184
rect 677744 440172 677750 440224
rect 678007 415876 717545 430563
rect 0 397571 41369 413629
rect 42242 413380 42248 413432
rect 42300 413420 42306 413432
rect 42610 413420 42616 413432
rect 42300 413392 42616 413420
rect 42300 413380 42306 413392
rect 42610 413380 42616 413392
rect 42668 413380 42674 413432
rect 672810 412496 672816 412548
rect 672868 412536 672874 412548
rect 676214 412536 676220 412548
rect 672868 412508 676220 412536
rect 672868 412496 672874 412508
rect 676214 412496 676220 412508
rect 676272 412496 676278 412548
rect 41782 410932 41788 410984
rect 41840 410972 41846 410984
rect 42518 410972 42524 410984
rect 41840 410944 42524 410972
rect 41840 410932 41846 410944
rect 42518 410932 42524 410944
rect 42576 410932 42582 410984
rect 672534 405628 672540 405680
rect 672592 405668 672598 405680
rect 672718 405668 672724 405680
rect 672592 405640 672724 405668
rect 672592 405628 672598 405640
rect 672718 405628 672724 405640
rect 672776 405628 672782 405680
rect 673454 401548 673460 401600
rect 673512 401588 673518 401600
rect 675294 401588 675300 401600
rect 673512 401560 675300 401588
rect 673512 401548 673518 401560
rect 675294 401548 675300 401560
rect 675352 401548 675358 401600
rect 41782 401480 41788 401532
rect 41840 401520 41846 401532
rect 42242 401520 42248 401532
rect 41840 401492 42248 401520
rect 41840 401480 41846 401492
rect 42242 401480 42248 401492
rect 42300 401520 42306 401532
rect 42610 401520 42616 401532
rect 42300 401492 42616 401520
rect 42300 401480 42306 401492
rect 42610 401480 42616 401492
rect 42668 401480 42674 401532
rect 672534 386384 672540 386436
rect 672592 386424 672598 386436
rect 672810 386424 672816 386436
rect 672592 386396 672816 386424
rect 672592 386384 672598 386396
rect 672810 386384 672816 386396
rect 672868 386384 672874 386436
rect 673638 382712 673644 382764
rect 673696 382752 673702 382764
rect 675386 382752 675392 382764
rect 673696 382724 675392 382752
rect 673696 382712 673702 382724
rect 675386 382712 675392 382724
rect 675444 382712 675450 382764
rect 42334 380876 42340 380928
rect 42392 380916 42398 380928
rect 42610 380916 42616 380928
rect 42392 380888 42616 380916
rect 42392 380876 42398 380888
rect 42610 380876 42616 380888
rect 42668 380876 42674 380928
rect 673822 372308 673828 372360
rect 673880 372348 673886 372360
rect 675386 372348 675392 372360
rect 673880 372320 675392 372348
rect 673880 372308 673886 372320
rect 675386 372308 675392 372320
rect 675444 372308 675450 372360
rect 676231 370571 717600 386629
rect 0 354371 41369 370429
rect 41782 368636 41788 368688
rect 41840 368676 41846 368688
rect 42518 368676 42524 368688
rect 41840 368648 42524 368676
rect 41840 368636 41846 368648
rect 42518 368636 42524 368648
rect 42576 368636 42582 368688
rect 42518 367004 42524 367056
rect 42576 367004 42582 367056
rect 42536 366976 42564 367004
rect 42794 366976 42800 366988
rect 42536 366948 42800 366976
rect 42794 366936 42800 366948
rect 42852 366936 42858 366988
rect 41782 357484 41788 357536
rect 41840 357524 41846 357536
rect 42334 357524 42340 357536
rect 41840 357496 42340 357524
rect 41840 357484 41846 357496
rect 42334 357484 42340 357496
rect 42392 357524 42398 357536
rect 42610 357524 42616 357536
rect 42392 357496 42616 357524
rect 42392 357484 42398 357496
rect 42610 357484 42616 357496
rect 42668 357484 42674 357536
rect 672626 353376 672632 353388
rect 672552 353348 672632 353376
rect 672552 353252 672580 353348
rect 672626 353336 672632 353348
rect 672684 353336 672690 353388
rect 672534 353200 672540 353252
rect 672592 353200 672598 353252
rect 42702 347692 42708 347744
rect 42760 347732 42766 347744
rect 42886 347732 42892 347744
rect 42760 347704 42892 347732
rect 42760 347692 42766 347704
rect 42886 347692 42892 347704
rect 42944 347692 42950 347744
rect 672534 347692 672540 347744
rect 672592 347732 672598 347744
rect 672718 347732 672724 347744
rect 672592 347704 672724 347732
rect 672592 347692 672598 347704
rect 672718 347692 672724 347704
rect 672776 347692 672782 347744
rect 673638 338512 673644 338564
rect 673696 338552 673702 338564
rect 675386 338552 675392 338564
rect 673696 338524 675392 338552
rect 673696 338512 673702 338524
rect 675386 338512 675392 338524
rect 675444 338512 675450 338564
rect 42334 334636 42340 334688
rect 42392 334676 42398 334688
rect 42610 334676 42616 334688
rect 42392 334648 42616 334676
rect 42392 334636 42398 334648
rect 42610 334636 42616 334648
rect 42668 334636 42674 334688
rect 42610 328448 42616 328500
rect 42668 328488 42674 328500
rect 42886 328488 42892 328500
rect 42668 328460 42892 328488
rect 42668 328448 42674 328460
rect 42886 328448 42892 328460
rect 42944 328448 42950 328500
rect 672442 328448 672448 328500
rect 672500 328488 672506 328500
rect 672718 328488 672724 328500
rect 672500 328460 672724 328488
rect 672500 328448 672506 328460
rect 672718 328448 672724 328460
rect 672776 328448 672782 328500
rect 0 311171 41369 327229
rect 673822 327088 673828 327140
rect 673880 327128 673886 327140
rect 675386 327128 675392 327140
rect 673880 327100 675392 327128
rect 673880 327088 673886 327100
rect 675386 327088 675392 327100
rect 675444 327088 675450 327140
rect 676231 325371 717600 341429
rect 41782 324504 41788 324556
rect 41840 324544 41846 324556
rect 41840 324516 42564 324544
rect 41840 324504 41846 324516
rect 42536 324488 42564 324516
rect 42518 324436 42524 324488
rect 42576 324436 42582 324488
rect 42334 314576 42340 314628
rect 42392 314576 42398 314628
rect 42352 314548 42380 314576
rect 42610 314548 42616 314560
rect 41800 314520 42616 314548
rect 41800 314492 41828 314520
rect 42610 314508 42616 314520
rect 42668 314508 42674 314560
rect 41782 314440 41788 314492
rect 41840 314440 41846 314492
rect 42518 314440 42524 314492
rect 42576 314480 42582 314492
rect 42794 314480 42800 314492
rect 42576 314452 42800 314480
rect 42576 314440 42582 314452
rect 42794 314440 42800 314452
rect 42852 314440 42858 314492
rect 672534 309068 672540 309120
rect 672592 309108 672598 309120
rect 672810 309108 672816 309120
rect 672592 309080 672816 309108
rect 672592 309068 672598 309080
rect 672810 309068 672816 309080
rect 672868 309068 672874 309120
rect 673454 304920 673460 304972
rect 673512 304960 673518 304972
rect 673822 304960 673828 304972
rect 673512 304932 673828 304960
rect 673512 304920 673518 304932
rect 673822 304920 673828 304932
rect 673880 304920 673886 304972
rect 42610 295332 42616 295384
rect 42668 295372 42674 295384
rect 42794 295372 42800 295384
rect 42668 295344 42800 295372
rect 42668 295332 42674 295344
rect 42794 295332 42800 295344
rect 42852 295332 42858 295384
rect 673638 293496 673644 293548
rect 673696 293536 673702 293548
rect 675018 293536 675024 293548
rect 673696 293508 675024 293536
rect 673696 293496 673702 293508
rect 675018 293496 675024 293508
rect 675076 293496 675082 293548
rect 672626 289824 672632 289876
rect 672684 289864 672690 289876
rect 672810 289864 672816 289876
rect 672684 289836 672816 289864
rect 672684 289824 672690 289836
rect 672810 289824 672816 289836
rect 672868 289824 672874 289876
rect 0 267971 41369 284029
rect 673454 283024 673460 283076
rect 673512 283064 673518 283076
rect 674926 283064 674932 283076
rect 673512 283036 674932 283064
rect 673512 283024 673518 283036
rect 674926 283024 674932 283036
rect 674984 283064 674990 283076
rect 675386 283064 675392 283076
rect 674984 283036 675392 283064
rect 674984 283024 674990 283036
rect 675386 283024 675392 283036
rect 675444 283024 675450 283076
rect 41782 282276 41788 282328
rect 41840 282316 41846 282328
rect 42426 282316 42432 282328
rect 41840 282288 42432 282316
rect 41840 282276 41846 282288
rect 42426 282276 42432 282288
rect 42484 282316 42490 282328
rect 42610 282316 42616 282328
rect 42484 282288 42616 282316
rect 42484 282276 42490 282288
rect 42610 282276 42616 282288
rect 42668 282276 42674 282328
rect 676231 280371 717600 296429
rect 673914 276020 673920 276072
rect 673972 276060 673978 276072
rect 675202 276060 675208 276072
rect 673972 276032 675208 276060
rect 673972 276020 673978 276032
rect 675202 276020 675208 276032
rect 675260 276020 675266 276072
rect 42518 275952 42524 276004
rect 42576 275992 42582 276004
rect 42794 275992 42800 276004
rect 42576 275964 42800 275992
rect 42576 275952 42582 275964
rect 42794 275952 42800 275964
rect 42852 275952 42858 276004
rect 41782 270784 41788 270836
rect 41840 270824 41846 270836
rect 42518 270824 42524 270836
rect 41840 270796 42524 270824
rect 41840 270784 41846 270796
rect 42518 270784 42524 270796
rect 42576 270784 42582 270836
rect 673730 266296 673736 266348
rect 673788 266336 673794 266348
rect 674926 266336 674932 266348
rect 673788 266308 674932 266336
rect 673788 266296 673794 266308
rect 674926 266296 674932 266308
rect 674984 266296 674990 266348
rect 673638 247460 673644 247512
rect 673696 247500 673702 247512
rect 673914 247500 673920 247512
rect 673696 247472 673920 247500
rect 673696 247460 673702 247472
rect 673914 247460 673920 247472
rect 673972 247500 673978 247512
rect 675386 247500 675392 247512
rect 673972 247472 675392 247500
rect 673972 247460 673978 247472
rect 675386 247460 675392 247472
rect 675444 247460 675450 247512
rect 0 224771 41369 240829
rect 41782 239028 41788 239080
rect 41840 239068 41846 239080
rect 42426 239068 42432 239080
rect 41840 239040 42432 239068
rect 41840 239028 41846 239040
rect 42426 239028 42432 239040
rect 42484 239068 42490 239080
rect 42610 239068 42616 239080
rect 42484 239040 42616 239068
rect 42484 239028 42490 239040
rect 42610 239028 42616 239040
rect 42668 239028 42674 239080
rect 673730 237668 673736 237720
rect 673788 237708 673794 237720
rect 675386 237708 675392 237720
rect 673788 237680 675392 237708
rect 673788 237668 673794 237680
rect 675386 237668 675392 237680
rect 675444 237668 675450 237720
rect 676231 235371 717600 251429
rect 41782 228624 41788 228676
rect 41840 228664 41846 228676
rect 42518 228664 42524 228676
rect 41840 228636 42524 228664
rect 41840 228624 41846 228636
rect 42518 228624 42524 228636
rect 42576 228624 42582 228676
rect 42242 227876 42248 227928
rect 42300 227916 42306 227928
rect 42518 227916 42524 227928
rect 42300 227888 42524 227916
rect 42300 227876 42306 227888
rect 42518 227876 42524 227888
rect 42576 227876 42582 227928
rect 672718 212508 672724 212560
rect 672776 212548 672782 212560
rect 672902 212548 672908 212560
rect 672776 212520 672908 212548
rect 672776 212508 672782 212520
rect 672902 212508 672908 212520
rect 672960 212508 672966 212560
rect 673454 203328 673460 203380
rect 673512 203368 673518 203380
rect 673638 203368 673644 203380
rect 673512 203340 673644 203368
rect 673512 203328 673518 203340
rect 673638 203328 673644 203340
rect 673696 203368 673702 203380
rect 675386 203368 675392 203380
rect 673696 203340 675392 203368
rect 673696 203328 673702 203340
rect 675386 203328 675392 203340
rect 675444 203328 675450 203380
rect 672534 198704 672540 198756
rect 672592 198744 672598 198756
rect 672718 198744 672724 198756
rect 672592 198716 672724 198744
rect 672592 198704 672598 198716
rect 672718 198704 672724 198716
rect 672776 198704 672782 198756
rect 0 181571 41369 197629
rect 41782 196732 41788 196784
rect 41840 196772 41846 196784
rect 42334 196772 42340 196784
rect 41840 196744 42340 196772
rect 41840 196732 41846 196744
rect 42334 196732 42340 196744
rect 42392 196732 42398 196784
rect 41782 195848 41788 195900
rect 41840 195888 41846 195900
rect 42610 195888 42616 195900
rect 41840 195860 42616 195888
rect 41840 195848 41846 195860
rect 42610 195848 42616 195860
rect 42668 195888 42674 195900
rect 44634 195888 44640 195900
rect 42668 195860 44640 195888
rect 42668 195848 42674 195860
rect 44634 195848 44640 195860
rect 44692 195848 44698 195900
rect 673730 191972 673736 192024
rect 673788 192012 673794 192024
rect 674006 192012 674012 192024
rect 673788 191984 674012 192012
rect 673788 191972 673794 191984
rect 674006 191972 674012 191984
rect 674064 191972 674070 192024
rect 676231 190171 717600 206229
rect 41782 189796 41788 189848
rect 41840 189836 41846 189848
rect 42334 189836 42340 189848
rect 41840 189808 42340 189836
rect 41840 189796 41846 189808
rect 42334 189796 42340 189808
rect 42392 189796 42398 189848
rect 44450 173884 44456 173936
rect 44508 173924 44514 173936
rect 44726 173924 44732 173936
rect 44508 173896 44732 173924
rect 44508 173884 44514 173896
rect 44726 173884 44732 173896
rect 44784 173884 44790 173936
rect 672718 173884 672724 173936
rect 672776 173924 672782 173936
rect 672902 173924 672908 173936
rect 672776 173896 672908 173924
rect 672776 173884 672782 173896
rect 672902 173884 672908 173896
rect 672960 173884 672966 173936
rect 673822 173884 673828 173936
rect 673880 173924 673886 173936
rect 674006 173924 674012 173936
rect 673880 173896 674012 173924
rect 673880 173884 673886 173896
rect 674006 173884 674012 173896
rect 674064 173884 674070 173936
rect 44726 160188 44732 160200
rect 44652 160160 44732 160188
rect 44652 160064 44680 160160
rect 44726 160148 44732 160160
rect 44784 160148 44790 160200
rect 672534 160080 672540 160132
rect 672592 160120 672598 160132
rect 672718 160120 672724 160132
rect 672592 160092 672724 160120
rect 672592 160080 672598 160092
rect 672718 160080 672724 160092
rect 672776 160080 672782 160132
rect 673638 160080 673644 160132
rect 673696 160120 673702 160132
rect 673822 160120 673828 160132
rect 673696 160092 673828 160120
rect 673696 160080 673702 160092
rect 673822 160080 673828 160092
rect 673880 160080 673886 160132
rect 44634 160012 44640 160064
rect 44692 160012 44698 160064
rect 673454 157292 673460 157344
rect 673512 157332 673518 157344
rect 675386 157332 675392 157344
rect 673512 157304 675392 157332
rect 673512 157292 673518 157304
rect 675386 157292 675392 157304
rect 675444 157292 675450 157344
rect 44634 154504 44640 154556
rect 44692 154544 44698 154556
rect 44726 154544 44732 154556
rect 44692 154516 44732 154544
rect 44692 154504 44698 154516
rect 44726 154504 44732 154516
rect 44784 154504 44790 154556
rect 673638 147840 673644 147892
rect 673696 147880 673702 147892
rect 674006 147880 674012 147892
rect 673696 147852 674012 147880
rect 673696 147840 673702 147852
rect 674006 147840 674012 147852
rect 674064 147880 674070 147892
rect 675386 147880 675392 147892
rect 674064 147852 675392 147880
rect 674064 147840 674070 147852
rect 675386 147840 675392 147852
rect 675444 147840 675450 147892
rect 676231 145171 717600 161229
rect 44726 140808 44732 140820
rect 44652 140780 44732 140808
rect 44652 140752 44680 140780
rect 44726 140768 44732 140780
rect 44784 140768 44790 140820
rect 44634 140700 44640 140752
rect 44692 140700 44698 140752
rect 55 110237 39593 124783
rect 44726 121564 44732 121576
rect 44652 121536 44732 121564
rect 44652 121440 44680 121536
rect 44726 121524 44732 121536
rect 44784 121524 44790 121576
rect 44634 121388 44640 121440
rect 44692 121388 44698 121440
rect 672718 115880 672724 115932
rect 672776 115920 672782 115932
rect 672810 115920 672816 115932
rect 672776 115892 672816 115920
rect 672776 115880 672782 115892
rect 672810 115880 672816 115892
rect 672868 115880 672874 115932
rect 673454 112072 673460 112124
rect 673512 112112 673518 112124
rect 675386 112112 675392 112124
rect 673512 112084 675392 112112
rect 673512 112072 673518 112084
rect 675386 112072 675392 112084
rect 675444 112072 675450 112124
rect 672810 102184 672816 102196
rect 672736 102156 672816 102184
rect 672736 102128 672764 102156
rect 672810 102144 672816 102156
rect 672868 102144 672874 102196
rect 673638 102144 673644 102196
rect 673696 102184 673702 102196
rect 673822 102184 673828 102196
rect 673696 102156 673828 102184
rect 673696 102144 673702 102156
rect 673822 102144 673828 102156
rect 673880 102144 673886 102196
rect 672718 102076 672724 102128
rect 672776 102076 672782 102128
rect 673638 102008 673644 102060
rect 673696 102048 673702 102060
rect 675386 102048 675392 102060
rect 673696 102020 675392 102048
rect 673696 102008 673702 102020
rect 675386 102008 675392 102020
rect 675444 102008 675450 102060
rect 676231 99971 717600 116029
rect 44266 96568 44272 96620
rect 44324 96608 44330 96620
rect 44542 96608 44548 96620
rect 44324 96580 44548 96608
rect 44324 96568 44330 96580
rect 44542 96568 44548 96580
rect 44600 96568 44606 96620
rect 32 68024 39593 82957
rect 672810 82900 672816 82952
rect 672868 82900 672874 82952
rect 672828 82748 672856 82900
rect 672810 82696 672816 82748
rect 672868 82696 672874 82748
rect 44266 77256 44272 77308
rect 44324 77296 44330 77308
rect 44358 77296 44364 77308
rect 44324 77268 44364 77296
rect 44324 77256 44330 77268
rect 44358 77256 44364 77268
rect 44416 77256 44422 77308
rect 39666 75216 39672 75268
rect 39724 75216 39730 75268
rect 39684 74996 39712 75216
rect 39666 74944 39672 74996
rect 39724 74944 39730 74996
rect 39574 67940 39580 67992
rect 39632 67980 39638 67992
rect 41414 67980 41420 67992
rect 39632 67952 41420 67980
rect 39632 67940 39638 67952
rect 41414 67940 41420 67952
rect 41472 67940 41478 67992
rect 41414 64608 41420 64660
rect 41472 64648 41478 64660
rect 42702 64648 42708 64660
rect 41472 64620 42708 64648
rect 41472 64608 41478 64620
rect 42702 64608 42708 64620
rect 42760 64608 42766 64660
rect 39666 52368 39672 52420
rect 39724 52408 39730 52420
rect 39850 52408 39856 52420
rect 39724 52380 39856 52408
rect 39724 52368 39730 52380
rect 39850 52368 39856 52380
rect 39908 52368 39914 52420
rect 45462 47880 45468 47932
rect 45520 47920 45526 47932
rect 179414 47920 179420 47932
rect 45520 47892 179420 47920
rect 45520 47880 45526 47892
rect 179414 47880 179420 47892
rect 179472 47880 179478 47932
rect 518802 47880 518808 47932
rect 518860 47920 518866 47932
rect 673638 47920 673644 47932
rect 518860 47892 673644 47920
rect 518860 47880 518866 47892
rect 673638 47880 673644 47892
rect 673696 47880 673702 47932
rect 39850 47812 39856 47864
rect 39908 47852 39914 47864
rect 189166 47852 189172 47864
rect 39908 47824 189172 47852
rect 39908 47812 39914 47824
rect 189166 47812 189172 47824
rect 189224 47812 189230 47864
rect 45554 47744 45560 47796
rect 45612 47784 45618 47796
rect 149054 47784 149060 47796
rect 45612 47756 149060 47784
rect 45612 47744 45618 47756
rect 149054 47744 149060 47756
rect 149112 47744 149118 47796
rect 528646 47744 528652 47796
rect 528704 47784 528710 47796
rect 672810 47784 672816 47796
rect 528704 47756 672816 47784
rect 528704 47744 528710 47756
rect 672810 47744 672816 47756
rect 672868 47744 672874 47796
rect 39758 47676 39764 47728
rect 39816 47716 39822 47728
rect 86310 47716 86316 47728
rect 39816 47688 86316 47716
rect 39816 47676 39822 47688
rect 86310 47676 86316 47688
rect 86368 47676 86374 47728
rect 212534 47648 212540 47660
rect 198936 47620 212540 47648
rect 195974 47580 195980 47592
rect 193232 47552 195980 47580
rect 179414 47472 179420 47524
rect 179472 47512 179478 47524
rect 193232 47512 193260 47552
rect 195974 47540 195980 47552
rect 196032 47580 196038 47592
rect 198642 47580 198648 47592
rect 196032 47552 198648 47580
rect 196032 47540 196038 47552
rect 198642 47540 198648 47552
rect 198700 47540 198706 47592
rect 198734 47540 198740 47592
rect 198792 47580 198798 47592
rect 198936 47580 198964 47620
rect 212534 47608 212540 47620
rect 212592 47608 212598 47660
rect 270494 47608 270500 47660
rect 270552 47608 270558 47660
rect 270512 47580 270540 47608
rect 198792 47552 198964 47580
rect 270420 47552 270540 47580
rect 198792 47540 198798 47552
rect 270420 47524 270448 47552
rect 303614 47540 303620 47592
rect 303672 47580 303678 47592
rect 304534 47580 304540 47592
rect 303672 47552 304540 47580
rect 303672 47540 303678 47552
rect 304534 47540 304540 47552
rect 304592 47580 304598 47592
rect 359366 47580 359372 47592
rect 304592 47552 359372 47580
rect 304592 47540 304598 47552
rect 359366 47540 359372 47552
rect 359424 47580 359430 47592
rect 361482 47580 361488 47592
rect 359424 47552 361488 47580
rect 359424 47540 359430 47552
rect 361482 47540 361488 47552
rect 361540 47540 361546 47592
rect 179472 47484 193260 47512
rect 179472 47472 179478 47484
rect 231762 47472 231768 47524
rect 231820 47512 231826 47524
rect 251174 47512 251180 47524
rect 231820 47484 231992 47512
rect 231820 47472 231826 47484
rect 231964 47444 231992 47484
rect 237392 47484 251180 47512
rect 237392 47444 237420 47484
rect 251174 47472 251180 47484
rect 251232 47472 251238 47524
rect 270402 47472 270408 47524
rect 270460 47472 270466 47524
rect 416774 47512 416780 47524
rect 400232 47484 416780 47512
rect 231964 47416 237420 47444
rect 289722 47404 289728 47456
rect 289780 47444 289786 47456
rect 289780 47416 295288 47444
rect 289780 47404 289786 47416
rect 86310 47336 86316 47388
rect 86368 47376 86374 47388
rect 199010 47376 199016 47388
rect 86368 47348 199016 47376
rect 86368 47336 86374 47348
rect 199010 47336 199016 47348
rect 199068 47376 199074 47388
rect 201402 47376 201408 47388
rect 199068 47348 201408 47376
rect 199068 47336 199074 47348
rect 201402 47336 201408 47348
rect 201460 47336 201466 47388
rect 251174 47336 251180 47388
rect 251232 47376 251238 47388
rect 270402 47376 270408 47388
rect 251232 47348 270408 47376
rect 251232 47336 251238 47348
rect 270402 47336 270408 47348
rect 270460 47336 270466 47388
rect 295260 47376 295288 47416
rect 364150 47404 364156 47456
rect 364208 47444 364214 47456
rect 400232 47444 400260 47484
rect 416774 47472 416780 47484
rect 416832 47472 416838 47524
rect 364208 47416 400260 47444
rect 364208 47404 364214 47416
rect 303614 47376 303620 47388
rect 295260 47348 303620 47376
rect 303614 47336 303620 47348
rect 303672 47336 303678 47388
rect 361482 47336 361488 47388
rect 361540 47376 361546 47388
rect 414198 47376 414204 47388
rect 361540 47348 414204 47376
rect 361540 47336 361546 47348
rect 414198 47336 414204 47348
rect 414256 47376 414262 47388
rect 417970 47376 417976 47388
rect 414256 47348 417976 47376
rect 414256 47336 414262 47348
rect 417970 47336 417976 47348
rect 418028 47336 418034 47388
rect 418062 47336 418068 47388
rect 418120 47376 418126 47388
rect 471974 47376 471980 47388
rect 418120 47348 471980 47376
rect 418120 47336 418126 47348
rect 471974 47336 471980 47348
rect 472032 47376 472038 47388
rect 526806 47376 526812 47388
rect 472032 47348 526812 47376
rect 472032 47336 472038 47348
rect 526806 47336 526812 47348
rect 526864 47336 526870 47388
rect 217962 47200 217968 47252
rect 218020 47240 218026 47252
rect 240134 47240 240140 47252
rect 218020 47212 240140 47240
rect 218020 47200 218026 47212
rect 240134 47200 240140 47212
rect 240192 47200 240198 47252
rect 285582 47268 285588 47320
rect 285640 47308 285646 47320
rect 307570 47308 307576 47320
rect 285640 47280 307576 47308
rect 285640 47268 285646 47280
rect 307570 47268 307576 47280
rect 307628 47308 307634 47320
rect 362402 47308 362408 47320
rect 307628 47280 362408 47308
rect 307628 47268 307634 47280
rect 362402 47268 362408 47280
rect 362460 47308 362466 47320
rect 364150 47308 364156 47320
rect 362460 47280 364156 47308
rect 362460 47268 362466 47280
rect 364150 47268 364156 47280
rect 364208 47268 364214 47320
rect 406746 47268 406752 47320
rect 406804 47308 406810 47320
rect 461486 47308 461492 47320
rect 406804 47280 461492 47308
rect 406804 47268 406810 47280
rect 461486 47268 461492 47280
rect 461544 47308 461550 47320
rect 516318 47308 516324 47320
rect 461544 47280 516324 47308
rect 461544 47268 461550 47280
rect 516318 47268 516324 47280
rect 516376 47308 516382 47320
rect 518802 47308 518808 47320
rect 516376 47280 518808 47308
rect 516376 47268 516382 47280
rect 518802 47268 518808 47280
rect 518860 47268 518866 47320
rect 200850 47132 200856 47184
rect 200908 47172 200914 47184
rect 242894 47172 242900 47184
rect 200908 47144 242900 47172
rect 200908 47132 200914 47144
rect 242894 47132 242900 47144
rect 242952 47132 242958 47184
rect 149054 47064 149060 47116
rect 149112 47104 149118 47116
rect 154574 47104 154580 47116
rect 149112 47076 154580 47104
rect 149112 47064 149118 47076
rect 154574 47064 154580 47076
rect 154632 47064 154638 47116
rect 188522 47104 188528 47116
rect 186608 47076 188528 47104
rect 173802 46996 173808 47048
rect 173860 47036 173866 47048
rect 173860 47008 179368 47036
rect 173860 46996 173866 47008
rect 179340 46968 179368 47008
rect 186608 46968 186636 47076
rect 188522 47064 188528 47076
rect 188580 47104 188586 47116
rect 192846 47104 192852 47116
rect 188580 47076 192852 47104
rect 188580 47064 188586 47076
rect 192846 47064 192852 47076
rect 192904 47104 192910 47116
rect 192904 47076 198688 47104
rect 192904 47064 192910 47076
rect 179340 46940 186636 46968
rect 186682 46928 186688 46980
rect 186740 46968 186746 46980
rect 194686 46968 194692 46980
rect 186740 46940 194692 46968
rect 186740 46928 186746 46940
rect 194686 46928 194692 46940
rect 194744 46928 194750 46980
rect 198660 46968 198688 47076
rect 201402 47064 201408 47116
rect 201460 47104 201466 47116
rect 247402 47104 247408 47116
rect 201460 47076 247408 47104
rect 201460 47064 201466 47076
rect 247402 47064 247408 47076
rect 247460 47104 247466 47116
rect 285582 47104 285588 47116
rect 247460 47076 285588 47104
rect 247460 47064 247466 47076
rect 285582 47064 285588 47076
rect 285640 47064 285646 47116
rect 309410 47200 309416 47252
rect 309468 47240 309474 47252
rect 352558 47240 352564 47252
rect 309468 47212 352564 47240
rect 309468 47200 309474 47212
rect 352558 47200 352564 47212
rect 352616 47200 352622 47252
rect 364242 47200 364248 47252
rect 364300 47240 364306 47252
rect 407390 47240 407396 47252
rect 364300 47212 407396 47240
rect 364300 47200 364306 47212
rect 407390 47200 407396 47212
rect 407448 47200 407454 47252
rect 416774 47200 416780 47252
rect 416832 47240 416838 47252
rect 417234 47240 417240 47252
rect 416832 47212 417240 47240
rect 416832 47200 416838 47212
rect 417234 47200 417240 47212
rect 417292 47240 417298 47252
rect 418062 47240 418068 47252
rect 417292 47212 418068 47240
rect 417292 47200 417298 47212
rect 418062 47200 418068 47212
rect 418120 47200 418126 47252
rect 419074 47200 419080 47252
rect 419132 47240 419138 47252
rect 462130 47240 462136 47252
rect 419132 47212 462136 47240
rect 419132 47200 419138 47212
rect 462130 47200 462136 47212
rect 462188 47200 462194 47252
rect 473814 47200 473820 47252
rect 473872 47240 473878 47252
rect 516962 47240 516968 47252
rect 473872 47212 516968 47240
rect 473872 47200 473878 47212
rect 516962 47200 516968 47212
rect 517020 47200 517026 47252
rect 299474 47132 299480 47184
rect 299532 47172 299538 47184
rect 305730 47172 305736 47184
rect 299532 47144 305736 47172
rect 299532 47132 299538 47144
rect 305730 47132 305736 47144
rect 305788 47172 305794 47184
rect 351914 47172 351920 47184
rect 305788 47144 351920 47172
rect 305788 47132 305794 47144
rect 351914 47132 351920 47144
rect 351972 47132 351978 47184
rect 360562 47132 360568 47184
rect 360620 47172 360626 47184
rect 406746 47172 406752 47184
rect 360620 47144 406752 47172
rect 360620 47132 360626 47144
rect 406746 47132 406752 47144
rect 406804 47132 406810 47184
rect 417970 47064 417976 47116
rect 418028 47104 418034 47116
rect 468938 47104 468944 47116
rect 418028 47076 468944 47104
rect 418028 47064 418034 47076
rect 468938 47064 468944 47076
rect 468996 47104 469002 47116
rect 523770 47104 523776 47116
rect 468996 47076 523776 47104
rect 468996 47064 469002 47076
rect 523770 47064 523776 47076
rect 523828 47104 523834 47116
rect 569126 47104 569132 47116
rect 523828 47076 569132 47104
rect 523828 47064 523834 47076
rect 569126 47064 569132 47076
rect 569184 47064 569190 47116
rect 201586 47036 201592 47048
rect 198752 47008 201592 47036
rect 198752 46968 198780 47008
rect 201586 46996 201592 47008
rect 201644 47036 201650 47048
rect 217962 47036 217968 47048
rect 201644 47008 217968 47036
rect 201644 46996 201650 47008
rect 217962 46996 217968 47008
rect 218020 46996 218026 47048
rect 198660 46940 198780 46968
rect 514478 46928 514484 46980
rect 514536 46968 514542 46980
rect 522482 46968 522488 46980
rect 514536 46940 522488 46968
rect 514536 46928 514542 46940
rect 522482 46928 522488 46940
rect 522540 46928 522546 46980
rect 526806 46928 526812 46980
rect 526864 46968 526870 46980
rect 634814 46968 634820 46980
rect 526864 46940 634820 46968
rect 526864 46928 526870 46940
rect 634814 46928 634820 46940
rect 634872 46928 634878 46980
rect 42702 45568 42708 45620
rect 42760 45608 42766 45620
rect 140958 45608 140964 45620
rect 42760 45580 140964 45608
rect 42760 45568 42766 45580
rect 140958 45568 140964 45580
rect 141016 45568 141022 45620
rect 242894 45500 242900 45552
rect 242952 45540 242958 45552
rect 297726 45540 297732 45552
rect 242952 45512 297732 45540
rect 242952 45500 242958 45512
rect 297726 45500 297732 45512
rect 297784 45500 297790 45552
rect 579154 45500 579160 45552
rect 579212 45540 579218 45552
rect 673454 45540 673460 45552
rect 579212 45512 673460 45540
rect 579212 45500 579218 45512
rect 673454 45500 673460 45512
rect 673512 45500 673518 45552
rect 140958 44140 140964 44192
rect 141016 44180 141022 44192
rect 254026 44180 254032 44192
rect 141016 44152 254032 44180
rect 141016 44140 141022 44152
rect 254026 44140 254032 44152
rect 254084 44180 254090 44192
rect 569218 44180 569224 44192
rect 254084 44152 569224 44180
rect 254084 44140 254090 44152
rect 569218 44140 569224 44152
rect 569276 44140 569282 44192
rect 299474 42004 299480 42016
rect 296916 41976 299480 42004
rect 296916 41948 296944 41976
rect 299474 41964 299480 41976
rect 299532 41964 299538 42016
rect 302234 41964 302240 42016
rect 302292 42004 302298 42016
rect 304994 42004 305000 42016
rect 302292 41976 305000 42004
rect 302292 41964 302298 41976
rect 304994 41964 305000 41976
rect 305052 41964 305058 42016
rect 411530 42004 411536 42016
rect 410260 41976 411536 42004
rect 410260 41948 410288 41976
rect 411530 41964 411536 41976
rect 411588 42004 411594 42016
rect 414566 42004 414572 42016
rect 411588 41976 414572 42004
rect 411588 41964 411594 41976
rect 414566 41964 414572 41976
rect 414624 42004 414630 42016
rect 415854 42004 415860 42016
rect 414624 41976 415860 42004
rect 414624 41964 414630 41976
rect 415854 41964 415860 41976
rect 415912 42004 415918 42016
rect 418246 42004 418252 42016
rect 415912 41976 418252 42004
rect 415912 41964 415918 41976
rect 418246 41964 418252 41976
rect 418304 41964 418310 42016
rect 466362 42004 466368 42016
rect 465092 41976 466368 42004
rect 465092 41948 465120 41976
rect 466362 41964 466368 41976
rect 466420 42004 466426 42016
rect 469398 42004 469404 42016
rect 466420 41976 469404 42004
rect 466420 41964 466426 41976
rect 469398 41964 469404 41976
rect 469456 42004 469462 42016
rect 470686 42004 470692 42016
rect 469456 41976 470692 42004
rect 469456 41964 469462 41976
rect 470686 41964 470692 41976
rect 470744 42004 470750 42016
rect 473078 42004 473084 42016
rect 470744 41976 473084 42004
rect 470744 41964 470750 41976
rect 473078 41964 473084 41976
rect 473136 41964 473142 42016
rect 296898 41936 296904 41948
rect 295352 41908 296904 41936
rect 189258 41828 189264 41880
rect 189316 41868 189322 41880
rect 191098 41868 191104 41880
rect 189316 41840 191104 41868
rect 189316 41828 189322 41840
rect 191098 41828 191104 41840
rect 191156 41868 191162 41880
rect 192294 41868 192300 41880
rect 191156 41840 192300 41868
rect 191156 41828 191162 41840
rect 192294 41828 192300 41840
rect 192352 41868 192358 41880
rect 192352 41840 193628 41868
rect 192352 41828 192358 41840
rect 193600 41812 193628 41840
rect 193582 41760 193588 41812
rect 193640 41800 193646 41812
rect 196434 41800 196440 41812
rect 193640 41772 196440 41800
rect 193640 41760 193646 41772
rect 196434 41760 196440 41772
rect 196492 41760 196498 41812
rect 198458 41760 198464 41812
rect 198516 41800 198522 41812
rect 200114 41800 200120 41812
rect 198516 41772 200120 41800
rect 198516 41760 198522 41772
rect 200114 41760 200120 41772
rect 200172 41760 200178 41812
rect 253934 41556 253940 41608
rect 253992 41596 253998 41608
rect 253992 41568 256740 41596
rect 253992 41556 253998 41568
rect 256712 41528 256740 41568
rect 256712 41500 275968 41528
rect 275940 41460 275968 41500
rect 295352 41460 295380 41908
rect 296898 41896 296904 41908
rect 296956 41896 296962 41948
rect 352650 41896 352656 41948
rect 352708 41936 352714 41948
rect 355502 41936 355508 41948
rect 352708 41908 355508 41936
rect 352708 41896 352714 41908
rect 355502 41896 355508 41908
rect 355560 41896 355566 41948
rect 356974 41896 356980 41948
rect 357032 41936 357038 41948
rect 359826 41936 359832 41948
rect 357032 41908 359832 41936
rect 357032 41896 357038 41908
rect 359826 41896 359832 41908
rect 359884 41936 359890 41948
rect 361114 41936 361120 41948
rect 359884 41908 361120 41936
rect 359884 41896 359890 41908
rect 361114 41896 361120 41908
rect 361172 41896 361178 41948
rect 407482 41896 407488 41948
rect 407540 41936 407546 41948
rect 410242 41936 410248 41948
rect 407540 41908 410248 41936
rect 407540 41896 407546 41908
rect 410242 41896 410248 41908
rect 410300 41896 410306 41948
rect 297910 41828 297916 41880
rect 297968 41868 297974 41880
rect 300670 41868 300676 41880
rect 297968 41840 300676 41868
rect 297968 41828 297974 41840
rect 300670 41828 300676 41840
rect 300728 41828 300734 41880
rect 352006 41828 352012 41880
rect 352064 41868 352070 41880
rect 354306 41868 354312 41880
rect 352064 41840 354312 41868
rect 352064 41828 352070 41840
rect 354306 41828 354312 41840
rect 354364 41868 354370 41880
rect 360470 41868 360476 41880
rect 354364 41840 360476 41868
rect 354364 41828 354370 41840
rect 360470 41828 360476 41840
rect 360528 41828 360534 41880
rect 295426 41760 295432 41812
rect 295484 41800 295490 41812
rect 303154 41800 303160 41812
rect 295484 41772 303160 41800
rect 295484 41760 295490 41772
rect 303154 41760 303160 41772
rect 303212 41760 303218 41812
rect 305270 41760 305276 41812
rect 305328 41800 305334 41812
rect 306558 41800 306564 41812
rect 305328 41772 306564 41800
rect 305328 41760 305334 41772
rect 306558 41760 306564 41772
rect 306616 41800 306622 41812
rect 308674 41800 308680 41812
rect 306616 41772 308680 41800
rect 306616 41760 306622 41772
rect 308674 41760 308680 41772
rect 308732 41760 308738 41812
rect 350166 41760 350172 41812
rect 350224 41800 350230 41812
rect 357986 41800 357992 41812
rect 350224 41772 357992 41800
rect 350224 41760 350230 41772
rect 357986 41760 357992 41772
rect 358044 41760 358050 41812
rect 361132 41800 361160 41896
rect 462314 41896 462320 41948
rect 462372 41936 462378 41948
rect 465074 41936 465080 41948
rect 462372 41908 465080 41936
rect 462372 41896 462378 41908
rect 465074 41896 465080 41908
rect 465132 41896 465138 41948
rect 459830 41828 459836 41880
rect 459888 41868 459894 41880
rect 467558 41868 467564 41880
rect 459888 41840 467564 41868
rect 459888 41828 459894 41840
rect 467558 41828 467564 41840
rect 467616 41828 467622 41880
rect 363506 41800 363512 41812
rect 361132 41772 363512 41800
rect 363506 41760 363512 41772
rect 363564 41760 363570 41812
rect 404998 41760 405004 41812
rect 405056 41800 405062 41812
rect 412726 41800 412732 41812
rect 405056 41772 412732 41800
rect 405056 41760 405062 41772
rect 412726 41760 412732 41772
rect 412784 41760 412790 41812
rect 517054 41760 517060 41812
rect 517112 41800 517118 41812
rect 520090 41800 520096 41812
rect 517112 41772 520096 41800
rect 517112 41760 517118 41772
rect 520090 41760 520096 41772
rect 520148 41800 520154 41812
rect 521378 41800 521384 41812
rect 520148 41772 521384 41800
rect 520148 41760 520154 41772
rect 521378 41760 521384 41772
rect 521436 41800 521442 41812
rect 524414 41800 524420 41812
rect 521436 41772 524420 41800
rect 521436 41760 521442 41772
rect 524414 41760 524420 41772
rect 524472 41800 524478 41812
rect 525702 41800 525708 41812
rect 524472 41772 525708 41800
rect 524472 41760 524478 41772
rect 525702 41760 525708 41772
rect 525760 41800 525766 41812
rect 527910 41800 527916 41812
rect 525760 41772 527916 41800
rect 525760 41760 525766 41772
rect 527910 41760 527916 41772
rect 527968 41760 527974 41812
rect 275940 41432 295380 41460
rect 133092 40196 133098 40248
rect 133150 40236 133156 40248
rect 143810 40236 143816 40248
rect 133150 40208 143816 40236
rect 133150 40196 133156 40208
rect 143810 40196 143816 40208
rect 143868 40196 143874 40248
rect 140990 40060 140996 40112
rect 141048 40100 141054 40112
rect 143066 40100 143072 40112
rect 141048 40072 143072 40100
rect 141048 40060 141054 40072
rect 142586 40000 142614 40072
rect 143066 40060 143072 40072
rect 143124 40100 143130 40112
rect 143350 40100 143356 40112
rect 143124 40072 143356 40100
rect 143124 40060 143130 40072
rect 143350 40060 143356 40072
rect 143408 40100 143414 40112
rect 143408 40072 144684 40100
rect 143408 40060 143414 40072
rect 144656 40000 144684 40072
rect 79076 55 93763 39593
rect 132600 37949 142517 40000
rect 142573 38005 142619 40000
rect 142675 37949 147600 40000
rect 132600 158 147600 37949
rect 186371 0 202429 41369
rect 252094 39652 252100 39704
rect 252152 39692 252158 39704
rect 254026 39692 254032 39704
rect 252152 39664 254032 39692
rect 252152 39652 252158 39664
rect 254026 39652 254032 39664
rect 254084 39652 254090 39704
rect 241243 32 256176 39593
rect 294971 0 311029 41369
rect 349771 0 365829 41369
rect 404571 0 420629 41369
rect 459371 0 475429 41369
rect 514171 0 530229 41369
rect 569276 55 583963 39593
rect 623217 55 637763 39593
<< metal2 >>
rect 45926 996512 45982 996568
rect 41713 969217 42193 969273
rect 41713 967377 42193 967433
rect 41713 965537 42193 965593
rect 41713 964341 42193 964397
rect 41713 963697 42193 963753
rect 41713 963053 42193 963109
rect 41713 962501 42193 962557
rect 41713 961213 42193 961269
rect 41713 960569 42193 960625
rect 41713 960017 42193 960073
rect 41713 959373 42193 959429
rect 41713 958729 42193 958785
rect 41713 958177 42193 958233
rect 42432 990140 42484 990146
rect 45466 990120 45522 990176
rect 42432 990082 42484 990088
rect 41713 956889 42193 956945
rect 41800 956486 41828 956889
rect 41788 956480 41840 956486
rect 41788 956422 41840 956428
rect 41713 956337 42193 956393
rect 41713 955693 42193 955749
rect 41713 955049 42193 955105
rect 42444 956486 42472 990082
rect 42432 956480 42484 956486
rect 42432 956422 42484 956428
rect 39670 908112 39726 908168
rect 40406 907976 40462 908032
rect 40406 888936 40462 888992
rect 40130 879960 40186 880016
rect 41418 875064 41474 875120
rect 39854 837528 39910 837584
rect 39854 832632 39910 832688
rect 39670 827464 39726 827520
rect 41713 799417 42193 799473
rect 41713 797577 42193 797633
rect 41713 795737 42193 795793
rect 41713 794541 42193 794597
rect 41713 793897 42193 793953
rect 41713 793253 42193 793309
rect 41713 792701 42193 792757
rect 41713 791413 42193 791469
rect 41713 790769 42193 790825
rect 41713 790217 42193 790273
rect 41713 789573 42193 789629
rect 41713 788929 42193 788985
rect 41713 788377 42193 788433
rect 42444 788066 42472 956422
rect 42260 788038 42472 788066
rect 42260 787250 42288 788038
rect 41800 787234 42288 787250
rect 41800 787228 42300 787234
rect 41800 787222 42248 787228
rect 41800 787145 41828 787222
rect 42248 787170 42300 787176
rect 41713 787089 42193 787145
rect 42260 787139 42288 787170
rect 41722 787086 41828 787089
rect 41713 786537 42193 786593
rect 41713 785893 42193 785949
rect 41713 785249 42193 785305
rect 42616 787228 42668 787234
rect 42616 787170 42668 787176
rect 41713 756217 42193 756273
rect 41713 754377 42193 754433
rect 41713 752537 42193 752593
rect 41713 751341 42193 751397
rect 41713 750697 42193 750753
rect 41713 750053 42193 750109
rect 41713 749501 42193 749557
rect 41713 748213 42193 748269
rect 41713 747569 42193 747625
rect 41713 747017 42193 747073
rect 41713 746373 42193 746429
rect 41713 745729 42193 745785
rect 41713 745177 42193 745233
rect 41788 744456 41840 744462
rect 41788 744398 41840 744404
rect 41800 743945 41828 744398
rect 41713 743889 42193 743945
rect 41713 743337 42193 743393
rect 41713 742693 42193 742749
rect 41713 742049 42193 742105
rect 42628 744462 42656 787170
rect 42616 744456 42668 744462
rect 42616 744398 42668 744404
rect 41713 713017 42193 713073
rect 41713 711177 42193 711233
rect 41713 709337 42193 709393
rect 41713 708141 42193 708197
rect 41713 707497 42193 707553
rect 41713 706853 42193 706909
rect 41713 706301 42193 706357
rect 41713 705013 42193 705069
rect 41713 704369 42193 704425
rect 41713 703817 42193 703873
rect 41713 703173 42193 703229
rect 41713 702529 42193 702585
rect 41713 701977 42193 702033
rect 41788 700868 41840 700874
rect 41788 700810 41840 700816
rect 41800 700754 41828 700810
rect 41722 700745 41828 700754
rect 41713 700689 42193 700745
rect 41713 700137 42193 700193
rect 41713 699493 42193 699549
rect 41713 698849 42193 698905
rect 41713 669817 42193 669873
rect 41713 667977 42193 668033
rect 41713 666137 42193 666193
rect 41713 664941 42193 664997
rect 41713 664297 42193 664353
rect 41713 663653 42193 663709
rect 41713 663101 42193 663157
rect 41713 661813 42193 661869
rect 41713 661169 42193 661225
rect 41713 660617 42193 660673
rect 41713 659973 42193 660029
rect 41713 659329 42193 659385
rect 41713 658777 42193 658833
rect 41713 657489 42193 657545
rect 41722 657478 41828 657489
rect 41800 657150 41828 657478
rect 41788 657144 41840 657150
rect 41788 657086 41840 657092
rect 42340 657144 42392 657150
rect 42340 657086 42392 657092
rect 41713 656937 42193 656993
rect 41713 656293 42193 656349
rect 41713 655649 42193 655705
rect 42352 633282 42380 657086
rect 42340 633276 42392 633282
rect 42340 633218 42392 633224
rect 41713 626617 42193 626673
rect 41713 624777 42193 624833
rect 41713 622937 42193 622993
rect 41713 621741 42193 621797
rect 41713 621097 42193 621153
rect 41713 620453 42193 620509
rect 41713 619901 42193 619957
rect 42628 700874 42656 744398
rect 42616 700868 42668 700874
rect 42616 700810 42668 700816
rect 42628 657150 42656 700810
rect 42616 657144 42668 657150
rect 42616 657086 42668 657092
rect 41713 618613 42193 618669
rect 41713 617969 42193 618025
rect 41713 617417 42193 617473
rect 41713 616773 42193 616829
rect 41713 616129 42193 616185
rect 41713 615577 42193 615633
rect 41880 614508 41932 614514
rect 41880 614450 41932 614456
rect 42248 614508 42300 614514
rect 42248 614450 42300 614456
rect 41892 614345 41920 614450
rect 41713 614289 42193 614345
rect 41713 613737 42193 613793
rect 41713 613093 42193 613149
rect 41713 612449 42193 612505
rect 42260 584254 42288 614450
rect 42248 584248 42300 584254
rect 42248 584190 42300 584196
rect 41713 583417 42193 583473
rect 41713 581577 42193 581633
rect 41713 579737 42193 579793
rect 41713 578541 42193 578597
rect 41713 577897 42193 577953
rect 41713 577253 42193 577309
rect 41713 576701 42193 576757
rect 42616 633276 42668 633282
rect 42616 633218 42668 633224
rect 42628 614514 42656 633218
rect 42616 614508 42668 614514
rect 42616 614450 42668 614456
rect 41713 575413 42193 575469
rect 41713 574769 42193 574825
rect 41713 574217 42193 574273
rect 41713 573573 42193 573629
rect 41713 572929 42193 572985
rect 41713 572377 42193 572433
rect 41788 571668 41840 571674
rect 41788 571610 41840 571616
rect 41800 571146 41828 571610
rect 41722 571145 41828 571146
rect 41713 571089 42193 571145
rect 41713 570537 42193 570593
rect 41713 569893 42193 569949
rect 41713 569249 42193 569305
rect 41713 540217 42193 540273
rect 41713 538377 42193 538433
rect 41713 536537 42193 536593
rect 41713 535341 42193 535397
rect 41713 534697 42193 534753
rect 41713 534053 42193 534109
rect 41713 533501 42193 533557
rect 41713 532213 42193 532269
rect 41713 531569 42193 531625
rect 41713 531017 42193 531073
rect 41713 530373 42193 530429
rect 41713 529729 42193 529785
rect 41713 529177 42193 529233
rect 42616 584248 42668 584254
rect 42616 584190 42668 584196
rect 42628 571674 42656 584190
rect 42616 571668 42668 571674
rect 42616 571610 42668 571616
rect 41788 528488 41840 528494
rect 41788 528430 41840 528436
rect 41800 527945 41828 528430
rect 41713 527889 42193 527945
rect 41713 527337 42193 527393
rect 41713 526693 42193 526749
rect 41713 526049 42193 526105
rect 39762 492904 39818 492960
rect 39946 455368 40002 455424
rect 39670 451832 39726 451888
rect 39670 440952 39726 441008
rect 42432 528488 42484 528494
rect 42432 528430 42484 528436
rect 41713 412617 42193 412673
rect 41713 410777 42193 410833
rect 41713 408937 42193 408993
rect 41713 407741 42193 407797
rect 41713 407097 42193 407153
rect 41713 406453 42193 406509
rect 41713 405901 42193 405957
rect 41713 404613 42193 404669
rect 41713 403969 42193 404025
rect 41713 403417 42193 403473
rect 41713 402773 42193 402829
rect 41713 402129 42193 402185
rect 41713 401577 42193 401633
rect 41713 400289 42193 400345
rect 41984 400178 42012 400289
rect 41972 400172 42024 400178
rect 42246 400152 42302 400208
rect 42444 400178 42472 528430
rect 42628 528494 42656 571610
rect 42616 528488 42668 528494
rect 42616 528430 42668 528436
rect 42432 400172 42484 400178
rect 41972 400114 42024 400120
rect 42432 400114 42484 400120
rect 41713 399737 42193 399793
rect 41713 399093 42193 399149
rect 41713 398449 42193 398505
rect 41713 369417 42193 369473
rect 41713 367577 42193 367633
rect 41713 365737 42193 365793
rect 41713 364541 42193 364597
rect 41713 363897 42193 363953
rect 41713 363253 42193 363309
rect 41713 362701 42193 362757
rect 41713 361413 42193 361469
rect 41713 360769 42193 360825
rect 41713 360217 42193 360273
rect 41713 359573 42193 359629
rect 41713 358929 42193 358985
rect 41713 358377 42193 358433
rect 41713 357089 42193 357145
rect 41800 356726 41828 357089
rect 42444 356726 42472 400114
rect 42614 400152 42670 400208
rect 41788 356720 41840 356726
rect 41788 356662 41840 356668
rect 42432 356720 42484 356726
rect 42432 356662 42484 356668
rect 41713 356537 42193 356593
rect 41713 355893 42193 355949
rect 41713 355249 42193 355305
rect 41713 326217 42193 326273
rect 41713 324377 42193 324433
rect 41713 322537 42193 322593
rect 41713 321341 42193 321397
rect 41713 320697 42193 320753
rect 41713 320053 42193 320109
rect 41713 319501 42193 319557
rect 41713 318213 42193 318269
rect 41713 317569 42193 317625
rect 41713 317017 42193 317073
rect 41713 316373 42193 316429
rect 41713 315729 42193 315785
rect 41713 315177 42193 315233
rect 41713 313889 42193 313945
rect 41800 313818 41828 313889
rect 42444 313818 42472 356662
rect 41788 313812 41840 313818
rect 41788 313754 41840 313760
rect 42432 313812 42484 313818
rect 42432 313754 42484 313760
rect 41713 313337 42193 313393
rect 41713 312693 42193 312749
rect 41713 312049 42193 312105
rect 42444 307970 42472 313754
rect 42432 307964 42484 307970
rect 42432 307906 42484 307912
rect 42708 307964 42760 307970
rect 42708 307906 42760 307912
rect 41713 283017 42193 283073
rect 41713 281177 42193 281233
rect 41713 279337 42193 279393
rect 41713 278141 42193 278197
rect 41713 277497 42193 277553
rect 41713 276853 42193 276909
rect 41713 276301 42193 276357
rect 41713 275013 42193 275069
rect 41713 274369 42193 274425
rect 41713 273817 42193 273873
rect 41713 273173 42193 273229
rect 41713 272529 42193 272585
rect 41713 271977 42193 272033
rect 41713 270689 42193 270745
rect 41800 270298 41828 270689
rect 41788 270292 41840 270298
rect 41788 270234 41840 270240
rect 42340 270292 42392 270298
rect 42340 270234 42392 270240
rect 41713 270137 42193 270193
rect 41713 269493 42193 269549
rect 41713 268849 42193 268905
rect 42352 247042 42380 270234
rect 42340 247036 42392 247042
rect 42340 246978 42392 246984
rect 41713 239817 42193 239873
rect 41713 237977 42193 238033
rect 41713 236137 42193 236193
rect 41713 234941 42193 234997
rect 41713 234297 42193 234353
rect 41713 233653 42193 233709
rect 41713 233101 42193 233157
rect 42720 282266 42748 307906
rect 42708 282260 42760 282266
rect 42708 282202 42760 282208
rect 42708 282056 42760 282062
rect 42708 281998 42760 282004
rect 41713 231813 42193 231869
rect 41713 231169 42193 231225
rect 41713 230617 42193 230673
rect 41713 229973 42193 230029
rect 41713 229329 42193 229385
rect 41713 228777 42193 228833
rect 42720 270298 42748 281998
rect 42708 270292 42760 270298
rect 42708 270234 42760 270240
rect 42708 247036 42760 247042
rect 42708 246978 42760 246984
rect 41788 228064 41840 228070
rect 41788 228006 41840 228012
rect 42432 228064 42484 228070
rect 42432 228006 42484 228012
rect 41800 227545 41828 228006
rect 41713 227489 42193 227545
rect 41713 226937 42193 226993
rect 41713 226293 42193 226349
rect 41713 225649 42193 225705
rect 41713 196617 42193 196673
rect 41713 194777 42193 194833
rect 41713 192937 42193 192993
rect 41713 191741 42193 191797
rect 41713 191097 42193 191153
rect 41713 190453 42193 190509
rect 41713 189901 42193 189957
rect 41713 188613 42193 188669
rect 41713 187969 42193 188025
rect 41713 187417 42193 187473
rect 41713 186773 42193 186829
rect 41713 186129 42193 186185
rect 41713 185577 42193 185633
rect 41713 184289 42193 184345
rect 41892 184226 41920 184289
rect 42260 184278 42288 184309
rect 42248 184272 42300 184278
rect 41892 184220 42248 184226
rect 41892 184214 42300 184220
rect 41892 184198 42288 184214
rect 41713 183737 42193 183793
rect 41713 183093 42193 183149
rect 41713 182449 42193 182505
rect 39762 120128 39818 120184
rect 41418 115912 41474 115968
rect 39394 84224 39450 84280
rect 42260 45694 42288 184198
rect 42444 184278 42472 228006
rect 42720 228070 42748 246978
rect 42708 228064 42760 228070
rect 42708 228006 42760 228012
rect 42432 184272 42484 184278
rect 42432 184214 42484 184220
rect 44362 917224 44418 917280
rect 333518 997600 333574 997656
rect 77049 995407 77105 995887
rect 77693 995407 77749 995887
rect 78337 995407 78393 995887
rect 78889 995452 78945 995887
rect 78876 995407 78945 995452
rect 80177 995407 80233 995887
rect 80729 995407 80785 995887
rect 81373 995407 81429 995887
rect 82017 995407 82073 995887
rect 82569 995407 82625 995887
rect 83213 995407 83269 995887
rect 84501 995407 84557 995887
rect 85053 995407 85109 995887
rect 85697 995407 85753 995887
rect 86341 995407 86397 995887
rect 87537 995407 87593 995887
rect 89377 995407 89433 995887
rect 91217 995407 91273 995887
rect 128449 995407 128505 995887
rect 129093 995407 129149 995887
rect 129737 995407 129793 995887
rect 130289 995407 130345 995887
rect 131577 995407 131633 995887
rect 132129 995407 132185 995887
rect 132773 995407 132829 995887
rect 133417 995407 133473 995887
rect 133969 995407 134025 995887
rect 134613 995407 134669 995887
rect 135901 995407 135957 995887
rect 136453 995407 136509 995887
rect 137097 995407 137153 995887
rect 137741 995407 137797 995887
rect 138937 995407 138993 995887
rect 140777 995407 140833 995887
rect 142617 995407 142673 995887
rect 179849 995407 179905 995887
rect 180493 995407 180549 995887
rect 181137 995407 181193 995887
rect 181689 995466 181745 995887
rect 181689 995407 181760 995466
rect 182977 995407 183033 995887
rect 183529 995407 183585 995887
rect 184173 995407 184229 995887
rect 184817 995407 184873 995887
rect 185369 995407 185425 995887
rect 186013 995407 186069 995887
rect 187301 995407 187357 995887
rect 187853 995407 187909 995887
rect 188497 995407 188553 995887
rect 189141 995407 189197 995887
rect 190337 995407 190393 995887
rect 192177 995407 192233 995887
rect 194017 995407 194073 995887
rect 231249 995407 231305 995887
rect 231893 995407 231949 995887
rect 232537 995407 232593 995887
rect 233089 995466 233145 995887
rect 233068 995407 233145 995466
rect 234377 995407 234433 995887
rect 234929 995407 234985 995887
rect 235573 995407 235629 995887
rect 236217 995407 236273 995887
rect 236769 995407 236825 995887
rect 237413 995407 237469 995887
rect 238701 995407 238757 995887
rect 239253 995407 239309 995887
rect 239897 995407 239953 995887
rect 240541 995407 240597 995887
rect 241737 995407 241793 995887
rect 243577 995407 243633 995887
rect 245417 995407 245473 995887
rect 282849 995407 282905 995887
rect 283493 995407 283549 995887
rect 284137 995407 284193 995887
rect 284689 995452 284745 995887
rect 284680 995407 284745 995452
rect 285977 995407 286033 995887
rect 286529 995407 286585 995887
rect 287173 995407 287229 995887
rect 287817 995407 287873 995887
rect 288369 995407 288425 995887
rect 289013 995407 289069 995887
rect 290301 995407 290357 995887
rect 290853 995407 290909 995887
rect 291497 995407 291553 995887
rect 292141 995407 292197 995887
rect 293337 995407 293393 995887
rect 295177 995407 295233 995887
rect 297017 995407 297073 995887
rect 78876 992202 78904 995407
rect 78876 992174 79088 992202
rect 79060 990826 79088 992174
rect 79048 990820 79100 990826
rect 79048 990762 79100 990768
rect 79060 990146 79088 990762
rect 130304 990894 130332 995407
rect 130292 990888 130344 990894
rect 130292 990830 130344 990836
rect 110420 990820 110472 990826
rect 110420 990762 110472 990768
rect 130108 990820 130160 990826
rect 130108 990762 130160 990768
rect 110432 990706 110460 990762
rect 110432 990678 110552 990706
rect 110524 990622 110552 990678
rect 130120 990622 130148 990762
rect 110512 990616 110564 990622
rect 110512 990558 110564 990564
rect 130108 990616 130160 990622
rect 130108 990558 130160 990564
rect 143264 990820 143316 990826
rect 143264 990762 143316 990768
rect 143276 990486 143304 990762
rect 143264 990480 143316 990486
rect 143264 990422 143316 990428
rect 173808 990820 173860 990826
rect 173808 990762 173860 990768
rect 179328 990820 179380 990826
rect 179328 990762 179380 990768
rect 173820 990729 173848 990762
rect 160098 990720 160154 990729
rect 160098 990655 160154 990664
rect 173806 990720 173862 990729
rect 173806 990655 173862 990664
rect 160112 990486 160140 990655
rect 179340 990622 179368 990762
rect 181732 990622 181760 995407
rect 187608 990752 187660 990758
rect 187608 990694 187660 990700
rect 187700 990752 187752 990758
rect 187700 990694 187752 990700
rect 179328 990616 179380 990622
rect 179328 990558 179380 990564
rect 181720 990616 181772 990622
rect 181720 990558 181772 990564
rect 160100 990480 160152 990486
rect 160100 990422 160152 990428
rect 181732 990486 181760 990558
rect 187620 990486 187648 990694
rect 187712 990486 187740 990694
rect 202880 990752 202932 990758
rect 202880 990694 202932 990700
rect 193218 990548 193274 990584
rect 193218 990528 193220 990548
rect 193272 990528 193274 990548
rect 202892 990486 202920 990694
rect 212446 990548 212502 990584
rect 233068 990758 233096 995407
rect 233056 990752 233108 990758
rect 233056 990694 233108 990700
rect 212446 990528 212448 990548
rect 212500 990528 212502 990548
rect 233068 990486 233096 990694
rect 284680 990826 284708 995407
rect 246948 990820 247000 990826
rect 246948 990762 247000 990768
rect 284668 990820 284720 990826
rect 284668 990762 284720 990768
rect 246960 990486 246988 990762
rect 286968 990820 287020 990826
rect 286968 990762 287020 990768
rect 286980 990554 287008 990762
rect 585690 996376 585746 996432
rect 672630 996512 672686 996568
rect 672446 996376 672502 996432
rect 384649 995407 384705 995887
rect 385293 995407 385349 995887
rect 385937 995407 385993 995887
rect 386489 995452 386545 995887
rect 386489 995407 386552 995452
rect 387777 995407 387833 995887
rect 388329 995407 388385 995887
rect 388973 995407 389029 995887
rect 389617 995407 389673 995887
rect 390169 995407 390225 995887
rect 390813 995407 390869 995887
rect 392101 995407 392157 995887
rect 392653 995407 392709 995887
rect 393297 995407 393353 995887
rect 393941 995407 393997 995887
rect 395137 995407 395193 995887
rect 396977 995407 397033 995887
rect 398817 995407 398873 995887
rect 473649 995407 473705 995887
rect 474293 995407 474349 995887
rect 474937 995407 474993 995887
rect 475489 995452 475545 995887
rect 475488 995407 475545 995452
rect 476777 995407 476833 995887
rect 477329 995407 477385 995887
rect 477973 995407 478029 995887
rect 478617 995407 478673 995887
rect 479169 995407 479225 995887
rect 479813 995407 479869 995887
rect 481101 995407 481157 995887
rect 481653 995407 481709 995887
rect 482297 995407 482353 995887
rect 482941 995407 482997 995887
rect 484137 995407 484193 995887
rect 485977 995407 486033 995887
rect 487817 995407 487873 995887
rect 525049 995407 525105 995887
rect 525693 995407 525749 995887
rect 526337 995407 526393 995887
rect 526889 995407 526945 995887
rect 528177 995407 528233 995887
rect 528729 995407 528785 995887
rect 529373 995407 529429 995887
rect 530017 995407 530073 995887
rect 530569 995407 530625 995887
rect 531213 995407 531269 995887
rect 532501 995407 532557 995887
rect 533053 995407 533109 995887
rect 533697 995407 533753 995887
rect 534341 995407 534397 995887
rect 535537 995407 535593 995887
rect 537377 995407 537433 995887
rect 537850 995424 537906 995480
rect 538034 995424 538090 995480
rect 286968 990548 287020 990554
rect 286968 990490 287020 990496
rect 181720 990480 181772 990486
rect 181720 990422 181772 990428
rect 187608 990480 187660 990486
rect 187608 990422 187660 990428
rect 187700 990480 187752 990486
rect 187700 990422 187752 990428
rect 202880 990480 202932 990486
rect 202880 990422 202932 990428
rect 233056 990480 233108 990486
rect 233056 990422 233108 990428
rect 246948 990480 247000 990486
rect 246948 990422 247000 990428
rect 386524 990622 386552 995407
rect 386512 990616 386564 990622
rect 386512 990558 386564 990564
rect 475488 992322 475516 995407
rect 463792 992316 463844 992322
rect 463792 992258 463844 992264
rect 475476 992316 475528 992322
rect 475476 992258 475528 992264
rect 419540 990888 419592 990894
rect 419540 990830 419592 990836
rect 438676 990888 438728 990894
rect 438676 990830 438728 990836
rect 450268 990888 450320 990894
rect 450268 990830 450320 990836
rect 463608 990888 463660 990894
rect 463804 990842 463832 992258
rect 463660 990836 463832 990842
rect 463608 990830 463832 990836
rect 419552 990622 419580 990830
rect 419540 990616 419592 990622
rect 419540 990558 419592 990564
rect 438688 990570 438716 990830
rect 450280 990622 450308 990830
rect 463620 990814 463832 990830
rect 482928 992316 482980 992322
rect 482928 992258 482980 992264
rect 482940 990758 482968 992258
rect 482928 990752 482980 990758
rect 482928 990694 482980 990700
rect 438768 990616 438820 990622
rect 438688 990564 438768 990570
rect 438688 990558 438820 990564
rect 450268 990616 450320 990622
rect 450268 990558 450320 990564
rect 438688 990542 438808 990558
rect 526916 990758 526944 995407
rect 526904 990752 526956 990758
rect 526904 990694 526956 990700
rect 539217 995407 539273 995887
rect 626849 995407 626905 995887
rect 627493 995407 627549 995887
rect 628137 995407 628193 995887
rect 628689 995466 628745 995887
rect 628668 995407 628745 995466
rect 629977 995407 630033 995887
rect 630529 995407 630585 995887
rect 631173 995407 631229 995887
rect 631817 995407 631873 995887
rect 632369 995407 632425 995887
rect 633013 995407 633069 995887
rect 634301 995407 634357 995887
rect 634853 995407 634909 995887
rect 635497 995407 635553 995887
rect 636141 995407 636197 995887
rect 637337 995407 637393 995887
rect 639177 995407 639233 995887
rect 641017 995407 641073 995887
rect 628668 990758 628696 995407
rect 628656 990752 628708 990758
rect 628656 990694 628708 990700
rect 576858 990564 576860 990584
rect 576912 990564 576914 990584
rect 576858 990528 576914 990564
rect 596086 990528 596142 990584
rect 540978 990428 540980 990448
rect 541032 990428 541034 990448
rect 540978 990392 541034 990428
rect 560206 990392 560262 990448
rect 628668 990146 628696 990694
rect 79048 990140 79100 990146
rect 79048 990082 79100 990088
rect 628656 990140 628708 990146
rect 628656 990082 628708 990088
rect 44454 835216 44510 835272
rect 672538 828688 672594 828744
rect 44730 828008 44786 828064
rect 673460 990072 673512 990078
rect 673460 990014 673512 990020
rect 673472 965326 673500 990014
rect 673460 965320 673512 965326
rect 673460 965262 673512 965268
rect 673366 908112 673422 908168
rect 673184 908064 673236 908070
rect 673184 908006 673236 908012
rect 673196 888826 673224 908006
rect 673184 888820 673236 888826
rect 673184 888762 673236 888768
rect 672630 826104 672686 826160
rect 673274 826104 673330 826160
rect 673182 823656 673238 823712
rect 672998 792104 673054 792160
rect 673182 792104 673238 792160
rect 672814 753480 672870 753536
rect 672998 753480 673054 753536
rect 672998 618160 673054 618216
rect 672814 618024 672870 618080
rect 44546 560224 44602 560280
rect 44914 560224 44970 560280
rect 673090 511400 673146 511456
rect 673274 511400 673330 511456
rect 672998 509088 673054 509144
rect 44454 493176 44510 493232
rect 44546 488552 44602 488608
rect 44362 448568 44418 448624
rect 673274 502288 673330 502344
rect 673472 908070 673500 965262
rect 675407 966695 675887 966751
rect 675407 966051 675887 966107
rect 675407 965407 675887 965463
rect 675392 965320 675444 965326
rect 675392 965262 675444 965268
rect 675404 964911 675432 965262
rect 675404 964883 675887 964911
rect 675407 964855 675887 964883
rect 675407 963567 675887 963623
rect 675407 963015 675887 963071
rect 675407 962371 675887 962427
rect 675407 961727 675887 961783
rect 675407 961175 675887 961231
rect 675407 960531 675887 960587
rect 673460 908064 673512 908070
rect 673460 908006 673512 908012
rect 673460 888820 673512 888826
rect 673460 888762 673512 888768
rect 673472 888729 673500 888762
rect 673458 888720 673514 888729
rect 673458 888655 673514 888664
rect 675407 959243 675887 959299
rect 675407 958691 675887 958747
rect 675407 958047 675887 958103
rect 675407 957403 675887 957459
rect 675407 956207 675887 956263
rect 675407 954367 675887 954423
rect 675407 952527 675887 952583
rect 677874 918584 677930 918640
rect 677598 915320 677654 915376
rect 677598 912736 677654 912792
rect 677874 912736 677930 912792
rect 677874 908112 677930 908168
rect 677782 907704 677838 907760
rect 675298 888720 675354 888729
rect 675298 888655 675354 888664
rect 675312 875697 675340 888655
rect 675407 877495 675887 877551
rect 675407 876851 675887 876907
rect 675407 876207 675887 876263
rect 675407 875697 675887 875711
rect 675220 875669 675887 875697
rect 675220 869446 675248 875669
rect 675407 875655 675887 875669
rect 675407 874367 675887 874423
rect 675407 873815 675887 873871
rect 675407 873171 675887 873227
rect 675407 872527 675887 872583
rect 675407 871975 675887 872031
rect 675407 871331 675887 871387
rect 673736 869440 673788 869446
rect 673736 869382 673788 869388
rect 675208 869440 675260 869446
rect 675208 869382 675260 869388
rect 673748 855522 673776 869382
rect 673656 855494 673776 855522
rect 673656 850082 673684 855494
rect 673564 850054 673684 850082
rect 673564 836330 673592 850054
rect 673552 836324 673604 836330
rect 673552 836266 673604 836272
rect 673644 836256 673696 836262
rect 673644 836198 673696 836204
rect 673656 830822 673684 836198
rect 673552 830816 673604 830822
rect 673552 830758 673604 830764
rect 673644 830816 673696 830822
rect 673644 830758 673696 830764
rect 673564 821098 673592 830758
rect 673552 821092 673604 821098
rect 673552 821034 673604 821040
rect 673552 768664 673604 768670
rect 673552 768606 673604 768612
rect 673564 741946 673592 768606
rect 673552 741940 673604 741946
rect 673552 741882 673604 741888
rect 675407 870043 675887 870099
rect 675407 869491 675887 869547
rect 675407 868847 675887 868903
rect 675407 868203 675887 868259
rect 675407 867007 675887 867063
rect 675407 865167 675887 865223
rect 675407 863327 675887 863383
rect 676126 828688 676182 828744
rect 676126 823656 676182 823712
rect 674104 821092 674156 821098
rect 674104 821034 674156 821040
rect 674116 797638 674144 821034
rect 674104 797632 674156 797638
rect 674104 797574 674156 797580
rect 675300 797632 675352 797638
rect 675300 797574 675352 797580
rect 675312 786497 675340 797574
rect 675407 788295 675887 788351
rect 675407 787651 675887 787707
rect 675407 787007 675887 787063
rect 675407 786497 675887 786511
rect 675312 786486 675887 786497
rect 674012 786480 674064 786486
rect 674012 786422 674064 786428
rect 675300 786480 675887 786486
rect 675352 786469 675887 786480
rect 675407 786455 675887 786469
rect 675300 786422 675352 786428
rect 674024 768670 674052 786422
rect 675312 786386 675340 786422
rect 675407 785167 675887 785223
rect 675407 784615 675887 784671
rect 675407 783971 675887 784027
rect 675407 783327 675887 783383
rect 675407 782775 675887 782831
rect 675407 782131 675887 782187
rect 675407 780843 675887 780899
rect 675407 780291 675887 780347
rect 675407 779647 675887 779703
rect 675407 779003 675887 779059
rect 675407 777807 675887 777863
rect 675407 775967 675887 776023
rect 675407 774127 675887 774183
rect 674012 768664 674064 768670
rect 674012 768606 674064 768612
rect 675407 743295 675887 743351
rect 675407 742651 675887 742707
rect 675407 742007 675887 742063
rect 674196 741940 674248 741946
rect 674196 741882 674248 741888
rect 675392 741940 675444 741946
rect 675392 741882 675444 741888
rect 673644 695972 673696 695978
rect 673644 695914 673696 695920
rect 673458 685344 673514 685400
rect 673656 651778 673684 695914
rect 674208 720458 674236 741882
rect 675404 741511 675432 741882
rect 675404 741483 675887 741511
rect 675407 741455 675887 741483
rect 675407 740167 675887 740223
rect 675407 739615 675887 739671
rect 675407 738971 675887 739027
rect 675407 738327 675887 738383
rect 675407 737775 675887 737831
rect 675407 737131 675887 737187
rect 675407 735843 675887 735899
rect 675407 735291 675887 735347
rect 675407 734647 675887 734703
rect 675407 734003 675887 734059
rect 675407 732807 675887 732863
rect 675407 730967 675887 731023
rect 675407 729127 675887 729183
rect 674012 720452 674064 720458
rect 674012 720394 674064 720400
rect 674196 720452 674248 720458
rect 674196 720394 674248 720400
rect 674024 710734 674052 720394
rect 674012 710728 674064 710734
rect 674012 710670 674064 710676
rect 675300 710728 675352 710734
rect 675300 710670 675352 710676
rect 675312 696497 675340 710670
rect 675407 698295 675887 698351
rect 675407 697651 675887 697707
rect 675407 697007 675887 697063
rect 675407 696497 675887 696511
rect 675312 696469 675887 696497
rect 675404 696455 675887 696469
rect 675404 695978 675432 696455
rect 675392 695972 675444 695978
rect 675392 695914 675444 695920
rect 675407 695167 675887 695223
rect 675407 694615 675887 694671
rect 675407 693971 675887 694027
rect 675407 693327 675887 693383
rect 675407 692775 675887 692831
rect 675407 692131 675887 692187
rect 675407 690843 675887 690899
rect 675407 690291 675887 690347
rect 675407 689647 675887 689703
rect 675407 689003 675887 689059
rect 675407 687807 675887 687863
rect 675407 685967 675887 686023
rect 675390 685344 675446 685400
rect 675407 684127 675887 684183
rect 675407 653095 675887 653151
rect 675407 652451 675887 652507
rect 675407 651807 675887 651863
rect 673644 651772 673696 651778
rect 673644 651714 673696 651720
rect 675392 651772 675444 651778
rect 675392 651714 675444 651720
rect 673656 606762 673684 651714
rect 675404 651311 675432 651714
rect 675404 651283 675887 651311
rect 675407 651255 675887 651283
rect 675407 649967 675887 650023
rect 675407 649415 675887 649471
rect 675407 648771 675887 648827
rect 675407 648127 675887 648183
rect 675407 647575 675887 647631
rect 675407 646931 675887 646987
rect 675407 645643 675887 645699
rect 675407 645091 675887 645147
rect 675407 644447 675887 644503
rect 675407 643803 675887 643859
rect 675407 642607 675887 642663
rect 675407 640767 675887 640823
rect 675407 638927 675887 638983
rect 675407 608095 675887 608151
rect 675407 607451 675887 607507
rect 675407 606807 675887 606863
rect 673644 606756 673696 606762
rect 673644 606698 673696 606704
rect 675392 606756 675444 606762
rect 675392 606698 675444 606704
rect 673656 561542 673684 606698
rect 675404 606311 675432 606698
rect 675404 606283 675887 606311
rect 675407 606255 675887 606283
rect 675407 604967 675887 605023
rect 675407 604415 675887 604471
rect 675407 603771 675887 603827
rect 675407 603127 675887 603183
rect 675407 602575 675887 602631
rect 675407 601931 675887 601987
rect 675407 600643 675887 600699
rect 675407 600091 675887 600147
rect 675407 599447 675887 599503
rect 675407 598803 675887 598859
rect 675407 597607 675887 597663
rect 675407 595767 675887 595823
rect 675407 593927 675887 593983
rect 675407 562895 675887 562951
rect 675407 562251 675887 562307
rect 675407 561607 675887 561663
rect 673644 561536 673696 561542
rect 673644 561478 673696 561484
rect 675392 561536 675444 561542
rect 675392 561478 675444 561484
rect 675404 561111 675432 561478
rect 675404 561068 675887 561111
rect 675407 561055 675887 561068
rect 675407 559767 675887 559823
rect 675407 559215 675887 559271
rect 675407 558571 675887 558627
rect 675407 557927 675887 557983
rect 675407 557375 675887 557431
rect 675407 556731 675887 556787
rect 675407 555443 675887 555499
rect 675407 554891 675887 554947
rect 675407 554247 675887 554303
rect 675407 553603 675887 553659
rect 675407 552407 675887 552463
rect 675407 550567 675887 550623
rect 675407 548727 675887 548783
rect 676126 514120 676182 514176
rect 676126 509088 676182 509144
rect 673642 502288 673698 502344
rect 673366 483112 673422 483168
rect 673366 482976 673422 483032
rect 678058 477536 678114 477592
rect 677874 469920 677930 469976
rect 673366 467472 673422 467528
rect 673274 463664 673330 463720
rect 673458 463664 673514 463720
rect 673458 463528 673514 463584
rect 673734 463528 673790 463584
rect 673090 427896 673146 427952
rect 673550 444352 673606 444408
rect 673734 444352 673790 444408
rect 673366 420824 673422 420880
rect 677414 427896 677470 427952
rect 677598 425720 677654 425776
rect 673552 384056 673604 384062
rect 673552 383998 673604 384004
rect 673564 338745 673592 383998
rect 675407 385695 675887 385751
rect 675407 385051 675887 385107
rect 675407 384407 675887 384463
rect 675392 384056 675444 384062
rect 675392 383998 675444 384004
rect 675404 383911 675432 383998
rect 675404 383860 675887 383911
rect 675407 383855 675887 383860
rect 673550 338736 673606 338745
rect 673550 338671 673606 338680
rect 672538 314744 672594 314800
rect 672538 314472 672594 314528
rect 673564 293298 673592 338671
rect 675407 382567 675887 382623
rect 675407 382015 675887 382071
rect 675407 381371 675887 381427
rect 675407 380727 675887 380783
rect 675407 380175 675887 380231
rect 675407 379531 675887 379587
rect 675407 378243 675887 378299
rect 675407 377691 675887 377747
rect 675407 377047 675887 377103
rect 675407 376403 675887 376459
rect 675407 375207 675887 375263
rect 675407 373367 675887 373423
rect 675407 371527 675887 371583
rect 675407 340495 675887 340551
rect 675407 339851 675887 339907
rect 675407 339207 675887 339263
rect 675390 338736 675446 338745
rect 675446 338680 675887 338711
rect 675390 338671 675887 338680
rect 675407 338655 675887 338671
rect 675407 337367 675887 337423
rect 675407 336815 675887 336871
rect 675407 336171 675887 336227
rect 675407 335527 675887 335583
rect 675407 334975 675887 335031
rect 675407 334331 675887 334387
rect 675407 333043 675887 333099
rect 675407 332491 675887 332547
rect 675407 331847 675887 331903
rect 675407 331203 675887 331259
rect 675407 330007 675887 330063
rect 675407 328167 675887 328223
rect 675407 326327 675887 326383
rect 675407 295495 675887 295551
rect 675407 294851 675887 294907
rect 675407 294207 675887 294263
rect 675407 293692 675887 293711
rect 675404 293655 675887 293692
rect 673564 293270 673868 293298
rect 673840 293214 673868 293270
rect 673828 293208 673880 293214
rect 673828 293150 673880 293156
rect 672538 231784 672594 231840
rect 672906 231784 672962 231840
rect 673552 203924 673604 203930
rect 673552 203866 673604 203872
rect 44454 193160 44510 193216
rect 44638 193160 44694 193216
rect 672538 193160 672594 193216
rect 672906 193160 672962 193216
rect 673564 158370 673592 203866
rect 673840 248198 673868 293150
rect 675404 293214 675432 293655
rect 675392 293208 675444 293214
rect 675392 293150 675444 293156
rect 675022 292984 675078 293040
rect 675206 292984 675262 293040
rect 675390 292984 675446 293040
rect 673828 248192 673880 248198
rect 673828 248134 673880 248140
rect 673840 203930 673868 248134
rect 675407 292367 675887 292423
rect 675407 291815 675887 291871
rect 675407 291171 675887 291227
rect 675407 290527 675887 290583
rect 675407 289975 675887 290031
rect 675407 289331 675887 289387
rect 675407 288043 675887 288099
rect 675407 287491 675887 287547
rect 675407 286847 675887 286903
rect 675407 286203 675887 286259
rect 675407 285007 675887 285063
rect 675407 283167 675887 283223
rect 675407 281327 675887 281383
rect 675407 250495 675887 250551
rect 675407 249851 675887 249907
rect 675407 249207 675887 249263
rect 675407 248676 675887 248711
rect 675404 248655 675887 248676
rect 675404 248198 675432 248655
rect 675392 248192 675444 248198
rect 675392 248134 675444 248140
rect 675407 247367 675887 247423
rect 675407 246815 675887 246871
rect 675407 246171 675887 246227
rect 675407 245527 675887 245583
rect 675407 244975 675887 245031
rect 675407 244331 675887 244387
rect 675407 243043 675887 243099
rect 675407 242491 675887 242547
rect 675407 241847 675887 241903
rect 675407 241203 675887 241259
rect 675407 240007 675887 240063
rect 675407 238167 675887 238223
rect 675407 236327 675887 236383
rect 675407 205295 675887 205351
rect 675407 204651 675887 204707
rect 675407 204007 675887 204063
rect 673828 203924 673880 203930
rect 673828 203866 673880 203872
rect 675392 203924 675444 203930
rect 675392 203866 675444 203872
rect 675404 203511 675432 203866
rect 675404 203483 675887 203511
rect 675407 203455 675887 203483
rect 675407 202167 675887 202223
rect 675407 201615 675887 201671
rect 675407 200971 675887 201027
rect 675407 200327 675887 200383
rect 675407 199775 675887 199831
rect 675407 199131 675887 199187
rect 673734 192344 673790 192400
rect 675407 197843 675887 197899
rect 675407 197291 675887 197347
rect 675407 196647 675887 196703
rect 675407 196003 675887 196059
rect 675407 194807 675887 194863
rect 675407 192967 675887 193023
rect 675390 192344 675446 192400
rect 675407 191127 675887 191183
rect 675407 160295 675887 160351
rect 673552 158364 673604 158370
rect 673552 158306 673604 158312
rect 44178 120128 44234 120184
rect 42338 115912 42394 115968
rect 44178 110472 44234 110528
rect 45466 110472 45522 110528
rect 44270 75792 44326 75848
rect 44270 73208 44326 73264
rect 44270 68176 44326 68232
rect 42248 45688 42300 45694
rect 42248 45630 42300 45636
rect 673564 112810 673592 158306
rect 675407 159651 675887 159707
rect 675407 159007 675887 159063
rect 675407 158508 675887 158511
rect 675404 158455 675887 158508
rect 675404 158370 675432 158455
rect 675392 158364 675444 158370
rect 675392 158306 675444 158312
rect 675407 157167 675887 157223
rect 675407 156615 675887 156671
rect 675407 155971 675887 156027
rect 675407 155327 675887 155383
rect 675407 154775 675887 154831
rect 675407 154131 675887 154187
rect 675407 152843 675887 152899
rect 675407 152291 675887 152347
rect 675407 151647 675887 151703
rect 675407 151003 675887 151059
rect 675407 149807 675887 149863
rect 675407 147967 675887 148023
rect 675407 146127 675887 146183
rect 673552 112804 673604 112810
rect 673552 112746 673604 112752
rect 45558 68176 45614 68232
rect 154578 47116 154634 47152
rect 154578 47096 154580 47116
rect 154632 47096 154634 47116
rect 173806 47096 173862 47152
rect 145104 45688 145156 45694
rect 145104 45630 145156 45636
rect 145116 44266 145144 45630
rect 145104 44260 145156 44266
rect 145104 44202 145156 44208
rect 86314 40160 86370 40216
rect 145116 40202 145144 44202
rect 212538 47660 212594 47696
rect 212538 47640 212540 47660
rect 212592 47640 212594 47660
rect 231582 47640 231638 47696
rect 270498 47660 270554 47696
rect 270498 47640 270500 47660
rect 270552 47640 270554 47660
rect 195336 44260 195388 44266
rect 195336 44202 195388 44208
rect 195348 42193 195376 44202
rect 289634 47640 289690 47696
rect 199660 47320 199712 47326
rect 199660 47262 199712 47268
rect 199672 42193 199700 47262
rect 187327 41713 187383 42193
rect 194043 41713 194099 42193
rect 195331 41834 195387 42193
rect 195428 41880 195480 41886
rect 195331 41828 195428 41834
rect 195331 41822 195480 41828
rect 195331 41806 195468 41822
rect 195331 41713 195387 41806
rect 199568 41880 199620 41886
rect 199655 41834 199711 42193
rect 199620 41828 199711 41834
rect 199568 41822 199711 41828
rect 199580 41806 199711 41822
rect 199655 41713 199711 41806
rect 149058 40296 149114 40352
rect 145103 40174 145144 40202
rect 145103 40000 145131 40174
rect 145091 39706 145143 40000
rect 240138 39888 240194 39944
rect 241242 39752 241298 39808
rect 242898 39752 242954 39808
rect 253938 39888 253994 39944
rect 303896 47116 303948 47122
rect 303896 47058 303948 47064
rect 303908 42193 303936 47058
rect 308220 47116 308272 47122
rect 308220 47058 308272 47064
rect 308232 42193 308260 47058
rect 358728 47116 358780 47122
rect 358728 47058 358780 47064
rect 358740 42193 358768 47058
rect 363052 47116 363104 47122
rect 363052 47058 363104 47064
rect 363064 42193 363092 47058
rect 413560 47116 413612 47122
rect 413560 47058 413612 47064
rect 413572 42193 413600 47058
rect 417884 47116 417936 47122
rect 417884 47058 417936 47064
rect 417896 42193 417924 47058
rect 468300 47184 468352 47190
rect 468300 47126 468352 47132
rect 468312 42193 468340 47126
rect 527456 47864 527508 47870
rect 527456 47806 527508 47812
rect 527468 47190 527496 47806
rect 527456 47184 527508 47190
rect 527456 47126 527508 47132
rect 527468 42193 527496 47126
rect 302643 41713 302699 42193
rect 303908 41806 303987 42193
rect 303931 41713 303987 41806
rect 306967 41713 307023 42193
rect 308232 41806 308311 42193
rect 308255 41713 308311 41806
rect 310095 41713 310151 42193
rect 357443 41713 357499 42193
rect 358731 41713 358787 42193
rect 361767 41713 361823 42193
rect 363055 41713 363111 42193
rect 364895 41713 364951 42193
rect 405527 41713 405583 42193
rect 409207 41834 409263 42193
rect 409328 41880 409380 41886
rect 409207 41828 409328 41834
rect 409207 41822 409380 41828
rect 409207 41806 409368 41822
rect 409207 41713 409263 41806
rect 411047 41834 411103 42193
rect 411168 41948 411220 41954
rect 411168 41890 411220 41896
rect 411180 41834 411208 41890
rect 411047 41806 411208 41834
rect 412243 41834 412299 42193
rect 412364 41880 412416 41886
rect 412243 41828 412364 41834
rect 412243 41822 412416 41828
rect 411047 41713 411103 41806
rect 412243 41806 412404 41822
rect 412243 41713 412299 41806
rect 413531 41820 413600 42193
rect 413531 41713 413587 41820
rect 415371 41834 415427 42193
rect 415492 41880 415544 41886
rect 415371 41828 415492 41834
rect 415371 41822 415544 41828
rect 415371 41806 415532 41822
rect 415371 41713 415427 41806
rect 416567 41713 416623 42193
rect 417855 41820 417924 42193
rect 419540 41880 419592 41886
rect 419695 41834 419751 42193
rect 419592 41828 419751 41834
rect 419540 41822 419751 41828
rect 417855 41713 417911 41820
rect 419552 41806 419751 41822
rect 419695 41713 419751 41806
rect 460327 41713 460383 42193
rect 464007 41834 464063 42193
rect 464007 41818 464200 41834
rect 464007 41812 464212 41818
rect 464007 41806 464160 41812
rect 464007 41713 464063 41806
rect 464160 41754 464212 41760
rect 465847 41834 465903 42193
rect 466000 41948 466052 41954
rect 466000 41890 466052 41896
rect 466012 41834 466040 41890
rect 465847 41806 466040 41834
rect 465847 41713 465903 41806
rect 467043 41834 467099 42193
rect 467043 41818 467236 41834
rect 467043 41812 467248 41818
rect 467043 41806 467196 41812
rect 467043 41713 467099 41806
rect 468312 41834 468387 42193
rect 468484 41880 468536 41886
rect 468312 41828 468484 41834
rect 468312 41822 468536 41828
rect 468312 41806 468524 41822
rect 470171 41834 470227 42193
rect 470060 41818 470227 41834
rect 467196 41754 467248 41760
rect 468331 41713 468387 41806
rect 470048 41812 470227 41818
rect 470100 41806 470227 41812
rect 470048 41754 470100 41760
rect 470171 41713 470227 41806
rect 471367 41713 471423 42193
rect 472532 41880 472584 41886
rect 472655 41834 472711 42193
rect 472584 41828 472711 41834
rect 472532 41822 472711 41828
rect 472544 41806 472711 41822
rect 474372 41948 474424 41954
rect 474372 41890 474424 41896
rect 474384 41834 474412 41890
rect 474495 41834 474551 42193
rect 474384 41806 474551 41834
rect 472655 41713 472711 41806
rect 474495 41713 474551 41806
rect 515127 41713 515183 42193
rect 518807 41834 518863 42193
rect 518900 41880 518952 41886
rect 518807 41828 518900 41834
rect 518807 41822 518952 41828
rect 518807 41806 518940 41822
rect 518807 41713 518863 41806
rect 520647 41713 520703 42193
rect 521843 41713 521899 42193
rect 523131 41834 523187 42193
rect 523224 41948 523276 41954
rect 523224 41890 523276 41896
rect 523236 41834 523264 41890
rect 523131 41806 523264 41834
rect 523131 41713 523187 41806
rect 524880 41880 524932 41886
rect 524971 41834 525027 42193
rect 524932 41828 525027 41834
rect 524880 41822 525027 41828
rect 524892 41806 525027 41822
rect 524971 41713 525027 41806
rect 526167 41713 526223 42193
rect 527455 41970 527511 42193
rect 527376 41954 527511 41970
rect 527364 41948 527511 41954
rect 527416 41942 527511 41948
rect 527364 41890 527416 41896
rect 527455 41713 527511 41942
rect 529295 41713 529351 42193
rect 622950 40432 623006 40488
rect 569222 40160 569278 40216
rect 579158 40160 579214 40216
rect 673564 47870 673592 112746
rect 675407 115095 675887 115151
rect 675407 114451 675887 114507
rect 675407 113807 675887 113863
rect 675407 113283 675887 113311
rect 675404 113255 675887 113283
rect 675404 112810 675432 113255
rect 675392 112804 675444 112810
rect 675392 112746 675444 112752
rect 675407 111967 675887 112023
rect 675407 111415 675887 111471
rect 675407 110771 675887 110827
rect 675407 110127 675887 110183
rect 675407 109575 675887 109631
rect 675407 108931 675887 108987
rect 675407 107643 675887 107699
rect 675407 107091 675887 107147
rect 675407 106447 675887 106503
rect 675407 105803 675887 105859
rect 675407 104607 675887 104663
rect 675407 102767 675887 102823
rect 675407 100927 675887 100983
rect 673552 47864 673604 47870
rect 673552 47806 673604 47812
rect 632978 40160 633034 40216
rect 634818 40160 634874 40216
rect 622950 39616 623006 39672
<< via2 >>
rect 160098 990664 160154 990720
rect 173806 990664 173862 990720
rect 193220 990528 193272 990548
rect 212448 990528 212500 990548
rect 576860 990564 576912 990584
rect 540980 990428 541032 990448
rect 673458 888664 673514 888720
rect 675298 888664 675354 888720
rect 673550 338680 673606 338736
rect 675390 338680 675446 338736
rect 154580 47096 154632 47116
rect 212540 47640 212592 47660
rect 270500 47640 270552 47660
<< obsm2 >>
rect 45926 996568 45982 996577
rect 45926 996503 45982 996512
rect 42248 990208 42300 990214
rect 42248 990150 42300 990156
rect 45466 990176 45522 990185
rect 0 969973 41713 970183
rect 0 969805 41657 969973
rect 41713 969861 42193 969917
rect 0 969329 41713 969805
rect 41800 969406 41828 969861
rect 41788 969400 41840 969406
rect 41788 969342 41840 969348
rect 0 969161 41657 969329
rect 0 968685 41713 969161
rect 0 968517 41657 968685
rect 41713 968573 42193 968629
rect 0 968133 41713 968517
rect 41788 968516 41840 968522
rect 41788 968458 41840 968464
rect 0 967965 41657 968133
rect 41800 968077 41828 968458
rect 41713 968021 42193 968077
rect 0 967489 41713 967965
rect 0 967321 41657 967489
rect 0 966845 41713 967321
rect 0 966677 41657 966845
rect 41713 966733 42193 966789
rect 0 966293 41713 966677
rect 0 966125 41657 966293
rect 41713 966181 42193 966237
rect 0 965649 41713 966125
rect 0 965481 41657 965649
rect 0 965005 41713 965481
rect 0 964837 41657 965005
rect 41713 964893 42193 964949
rect 0 964453 41713 964837
rect 0 964285 41657 964453
rect 0 963809 41713 964285
rect 0 963641 41657 963809
rect 0 963165 41713 963641
rect 0 962997 41657 963165
rect 0 962613 41713 962997
rect 0 962445 41657 962613
rect 41788 962464 41840 962470
rect 0 961969 41713 962445
rect 41788 962406 41840 962412
rect 0 961801 41657 961969
rect 41800 961913 41828 962406
rect 41713 961857 42193 961913
rect 41722 961846 41828 961857
rect 0 961325 41713 961801
rect 0 961157 41657 961325
rect 0 960681 41713 961157
rect 0 960513 41657 960681
rect 0 960129 41713 960513
rect 0 959961 41657 960129
rect 0 959485 41713 959961
rect 0 959317 41657 959485
rect 0 958841 41713 959317
rect 0 958673 41657 958841
rect 0 958289 41713 958673
rect 0 958121 41657 958289
rect 0 957645 41713 958121
rect 0 957477 41657 957645
rect 41713 957533 42193 957589
rect 0 957001 41713 957477
rect 41892 957386 41920 957533
rect 42260 957386 42288 990150
rect 45466 990111 45522 990120
rect 42340 969400 42392 969406
rect 42340 969342 42392 969348
rect 42352 962470 42380 969342
rect 42340 962464 42392 962470
rect 42340 962406 42392 962412
rect 41892 957358 42288 957386
rect 0 956833 41657 957001
rect 0 956449 41713 956833
rect 0 956281 41657 956449
rect 0 955805 41713 956281
rect 0 955637 41657 955805
rect 0 955161 41713 955637
rect 0 954993 41657 955161
rect 0 954609 41713 954993
rect 0 954441 41657 954609
rect 41713 954497 42193 954553
rect 0 954242 41713 954441
rect 714 922887 38812 926940
rect 38868 922978 39600 926940
rect 38868 922962 39712 922978
rect 38868 922956 39724 922962
rect 38868 922950 39672 922956
rect 38868 922943 39600 922950
rect 39672 922898 39724 922904
rect 714 920944 39593 922887
rect 714 918832 39479 920944
rect 39535 919034 39600 920888
rect 39535 919006 39896 919034
rect 39535 918888 39600 919006
rect 714 916155 39593 918832
rect 714 912098 39247 916155
rect 39303 912234 39600 916099
rect 39868 914734 39896 919006
rect 42260 914734 42288 957358
rect 42524 990072 42576 990078
rect 42524 990014 42576 990020
rect 42536 968522 42564 990014
rect 42524 968516 42576 968522
rect 42524 968458 42576 968464
rect 39856 914728 39908 914734
rect 39856 914670 39908 914676
rect 41420 914728 41472 914734
rect 41420 914670 41472 914676
rect 42248 914728 42300 914734
rect 42248 914670 42300 914676
rect 39303 912206 39712 912234
rect 39303 912100 39600 912206
rect 39684 908177 39712 912206
rect 39670 908168 39726 908177
rect 39670 908103 39726 908112
rect 40406 908032 40462 908041
rect 40406 907967 40462 907976
rect 40420 889001 40448 907967
rect 40406 888992 40462 889001
rect 40406 888927 40462 888936
rect 985 879822 34812 884658
rect 34868 879878 40000 884658
rect 40130 880016 40186 880025
rect 40130 879951 40186 879960
rect 39868 879850 39896 879878
rect 40144 879850 40172 879951
rect 39856 879844 39908 879850
rect 985 874735 39593 879822
rect 39856 879786 39908 879792
rect 40132 879844 40184 879850
rect 40132 879786 40184 879792
rect 41432 875634 41460 914670
rect 41420 875628 41472 875634
rect 41420 875570 41472 875576
rect 42248 875628 42300 875634
rect 42248 875570 42300 875576
rect 41432 875129 41460 875570
rect 41418 875120 41474 875129
rect 41418 875055 41474 875064
rect 985 869853 39533 874735
rect 39589 869899 40000 874679
rect 985 837622 34812 842458
rect 34868 837678 40000 842458
rect 985 832535 39593 837622
rect 39854 837584 39910 837593
rect 39854 837519 39910 837528
rect 39868 832697 39896 837519
rect 39854 832688 39910 832697
rect 39854 832623 39910 832632
rect 985 827653 39533 832535
rect 39589 827699 40000 832479
rect 39684 827529 39712 827699
rect 39670 827520 39726 827529
rect 39670 827455 39726 827464
rect 42260 807362 42288 875570
rect 42248 807356 42300 807362
rect 42248 807298 42300 807304
rect 0 800173 41713 800383
rect 0 800005 41657 800173
rect 41713 800061 42193 800117
rect 0 799529 41713 800005
rect 41800 799898 41828 800061
rect 41800 799870 42288 799898
rect 0 799361 41657 799529
rect 0 798885 41713 799361
rect 0 798717 41657 798885
rect 41713 798773 42193 798829
rect 0 798333 41713 798717
rect 41788 798380 41840 798386
rect 0 798165 41657 798333
rect 41788 798322 41840 798328
rect 41800 798277 41828 798322
rect 41713 798221 42193 798277
rect 0 797689 41713 798165
rect 0 797521 41657 797689
rect 0 797045 41713 797521
rect 0 796877 41657 797045
rect 41713 796933 42193 796989
rect 0 796493 41713 796877
rect 0 796325 41657 796493
rect 41713 796381 42193 796437
rect 0 795849 41713 796325
rect 0 795681 41657 795849
rect 0 795205 41713 795681
rect 0 795037 41657 795205
rect 41713 795093 42193 795149
rect 0 794653 41713 795037
rect 0 794485 41657 794653
rect 0 794009 41713 794485
rect 0 793841 41657 794009
rect 0 793365 41713 793841
rect 0 793197 41657 793365
rect 0 792813 41713 793197
rect 0 792645 41657 792813
rect 0 792169 41713 792645
rect 42260 792282 42288 799870
rect 41800 792254 42288 792282
rect 0 792001 41657 792169
rect 41800 792113 41828 792254
rect 41713 792057 42193 792113
rect 0 791525 41713 792001
rect 0 791357 41657 791525
rect 0 790881 41713 791357
rect 0 790713 41657 790881
rect 0 790329 41713 790713
rect 0 790161 41657 790329
rect 0 789685 41713 790161
rect 0 789517 41657 789685
rect 0 789041 41713 789517
rect 0 788873 41657 789041
rect 0 788489 41713 788873
rect 0 788321 41657 788489
rect 0 787845 41713 788321
rect 42536 798386 42564 968458
rect 45480 930170 45508 990111
rect 44272 930164 44324 930170
rect 44272 930106 44324 930112
rect 45468 930164 45520 930170
rect 45468 930106 45520 930112
rect 44284 922962 44312 930106
rect 44272 922956 44324 922962
rect 44272 922898 44324 922904
rect 44180 879844 44232 879850
rect 44180 879786 44232 879792
rect 42708 807356 42760 807362
rect 42708 807298 42760 807304
rect 42524 798380 42576 798386
rect 42524 798322 42576 798328
rect 41788 787908 41840 787914
rect 41788 787850 41840 787856
rect 0 787677 41657 787845
rect 41800 787794 41828 787850
rect 41722 787789 41828 787794
rect 41713 787733 42193 787789
rect 0 787201 41713 787677
rect 42432 787908 42484 787914
rect 42432 787850 42484 787856
rect 0 787033 41657 787201
rect 0 786649 41713 787033
rect 42444 786978 42472 787850
rect 42260 786950 42472 786978
rect 0 786481 41657 786649
rect 0 786005 41713 786481
rect 0 785837 41657 786005
rect 0 785361 41713 785837
rect 0 785193 41657 785361
rect 0 784809 41713 785193
rect 0 784641 41657 784809
rect 41713 784697 42193 784753
rect 0 784442 41713 784641
rect 0 756973 41713 757183
rect 42260 757058 42288 786950
rect 42536 768670 42564 798322
rect 42720 787914 42748 807298
rect 42708 787908 42760 787914
rect 42708 787850 42760 787856
rect 42524 768664 42576 768670
rect 42524 768606 42576 768612
rect 42260 757030 42380 757058
rect 0 756805 41657 756973
rect 41722 756917 42288 756922
rect 41713 756894 42288 756917
rect 41713 756861 42193 756894
rect 0 756329 41713 756805
rect 0 756161 41657 756329
rect 0 755685 41713 756161
rect 0 755517 41657 755685
rect 41713 755573 42193 755629
rect 0 755133 41713 755517
rect 0 754965 41657 755133
rect 41713 755021 42193 755077
rect 0 754489 41713 754965
rect 41800 754526 41828 755021
rect 41788 754520 41840 754526
rect 0 754321 41657 754489
rect 41788 754462 41840 754468
rect 0 753845 41713 754321
rect 0 753677 41657 753845
rect 41713 753733 42193 753789
rect 0 753293 41713 753677
rect 0 753125 41657 753293
rect 41713 753181 42193 753237
rect 0 752649 41713 753125
rect 0 752481 41657 752649
rect 0 752005 41713 752481
rect 0 751837 41657 752005
rect 41713 751893 42193 751949
rect 0 751453 41713 751837
rect 0 751285 41657 751453
rect 0 750809 41713 751285
rect 0 750641 41657 750809
rect 0 750165 41713 750641
rect 0 749997 41657 750165
rect 0 749613 41713 749997
rect 0 749445 41657 749613
rect 0 748969 41713 749445
rect 42260 749034 42288 756894
rect 41800 749006 42288 749034
rect 0 748801 41657 748969
rect 41800 748913 41828 749006
rect 41713 748857 42193 748913
rect 0 748325 41713 748801
rect 0 748157 41657 748325
rect 0 747681 41713 748157
rect 0 747513 41657 747681
rect 0 747129 41713 747513
rect 0 746961 41657 747129
rect 0 746485 41713 746961
rect 0 746317 41657 746485
rect 0 745841 41713 746317
rect 0 745673 41657 745841
rect 0 745289 41713 745673
rect 0 745121 41657 745289
rect 0 744645 41713 745121
rect 42352 744682 42380 757030
rect 42524 754520 42576 754526
rect 42524 754462 42576 754468
rect 41800 744654 42380 744682
rect 0 744477 41657 744645
rect 41800 744589 41828 744654
rect 41713 744533 42193 744589
rect 0 744001 41713 744477
rect 0 743833 41657 744001
rect 0 743449 41713 743833
rect 0 743281 41657 743449
rect 0 742805 41713 743281
rect 0 742637 41657 742805
rect 0 742161 41713 742637
rect 0 741993 41657 742161
rect 0 741609 41713 741993
rect 0 741441 41657 741609
rect 41713 741497 42193 741553
rect 0 741242 41713 741441
rect 0 713773 41713 713983
rect 42260 713810 42288 744654
rect 42536 744546 42564 754462
rect 42352 744518 42564 744546
rect 42352 713946 42380 744518
rect 42708 768664 42760 768670
rect 42708 768606 42760 768612
rect 42720 754526 42748 768606
rect 42708 754520 42760 754526
rect 42708 754462 42760 754468
rect 42352 713918 42564 713946
rect 42260 713782 42380 713810
rect 0 713605 41657 713773
rect 41713 713703 42193 713717
rect 41713 713675 42288 713703
rect 41713 713661 42193 713675
rect 0 713129 41713 713605
rect 0 712961 41657 713129
rect 0 712485 41713 712961
rect 0 712317 41657 712485
rect 41713 712373 42193 712429
rect 0 711933 41713 712317
rect 0 711765 41657 711933
rect 41713 711821 42193 711877
rect 0 711289 41713 711765
rect 41800 711346 41828 711821
rect 41788 711340 41840 711346
rect 0 711121 41657 711289
rect 41788 711282 41840 711288
rect 0 710645 41713 711121
rect 0 710477 41657 710645
rect 41713 710533 42193 710589
rect 0 710093 41713 710477
rect 0 709925 41657 710093
rect 41713 709981 42193 710037
rect 0 709449 41713 709925
rect 0 709281 41657 709449
rect 0 708805 41713 709281
rect 0 708637 41657 708805
rect 41713 708693 42193 708749
rect 0 708253 41713 708637
rect 0 708085 41657 708253
rect 0 707609 41713 708085
rect 0 707441 41657 707609
rect 0 706965 41713 707441
rect 0 706797 41657 706965
rect 0 706413 41713 706797
rect 0 706245 41657 706413
rect 0 705769 41713 706245
rect 42260 705786 42288 713675
rect 0 705601 41657 705769
rect 41800 705758 42288 705786
rect 41800 705713 41828 705758
rect 41713 705657 42193 705713
rect 42352 705699 42380 713782
rect 42536 711346 42564 713918
rect 42524 711340 42576 711346
rect 42524 711282 42576 711288
rect 42260 705671 42380 705699
rect 0 705125 41713 705601
rect 0 704957 41657 705125
rect 0 704481 41713 704957
rect 0 704313 41657 704481
rect 0 703929 41713 704313
rect 0 703761 41657 703929
rect 0 703285 41713 703761
rect 0 703117 41657 703285
rect 0 702641 41713 703117
rect 0 702473 41657 702641
rect 0 702089 41713 702473
rect 0 701921 41657 702089
rect 0 701445 41713 701921
rect 0 701277 41657 701445
rect 41713 701375 42193 701389
rect 42260 701375 42288 705671
rect 42536 705514 42564 711282
rect 41713 701347 42288 701375
rect 41713 701333 42193 701347
rect 0 700801 41713 701277
rect 42260 701010 42288 701347
rect 42352 705486 42564 705514
rect 42248 701004 42300 701010
rect 42248 700946 42300 700952
rect 0 700633 41657 700801
rect 0 700249 41713 700633
rect 0 700081 41657 700249
rect 0 699605 41713 700081
rect 0 699437 41657 699605
rect 0 698961 41713 699437
rect 0 698793 41657 698961
rect 0 698409 41713 698793
rect 0 698241 41657 698409
rect 41713 698297 42193 698353
rect 0 698042 41713 698241
rect 0 670573 41713 670783
rect 0 670405 41657 670573
rect 41713 670503 42193 670517
rect 41713 670475 42288 670503
rect 41713 670461 42193 670475
rect 0 669929 41713 670405
rect 0 669761 41657 669929
rect 0 669285 41713 669761
rect 0 669117 41657 669285
rect 41713 669173 42193 669229
rect 0 668733 41713 669117
rect 41788 669112 41840 669118
rect 41788 669054 41840 669060
rect 0 668565 41657 668733
rect 41800 668677 41828 669054
rect 41713 668621 42193 668677
rect 0 668089 41713 668565
rect 0 667921 41657 668089
rect 0 667445 41713 667921
rect 0 667277 41657 667445
rect 41713 667333 42193 667389
rect 0 666893 41713 667277
rect 0 666725 41657 666893
rect 41713 666781 42193 666837
rect 0 666249 41713 666725
rect 0 666081 41657 666249
rect 0 665605 41713 666081
rect 0 665437 41657 665605
rect 41713 665493 42193 665549
rect 0 665053 41713 665437
rect 0 664885 41657 665053
rect 0 664409 41713 664885
rect 0 664241 41657 664409
rect 0 663765 41713 664241
rect 0 663597 41657 663765
rect 0 663213 41713 663597
rect 0 663045 41657 663213
rect 0 662569 41713 663045
rect 0 662401 41657 662569
rect 42260 662538 42288 670475
rect 42352 669186 42380 705486
rect 42524 701004 42576 701010
rect 42524 700946 42576 700952
rect 42340 669180 42392 669186
rect 42340 669122 42392 669128
rect 41708 662510 42288 662538
rect 41708 662485 42193 662510
rect 41713 662457 42193 662485
rect 42352 662499 42380 669122
rect 42352 662471 42472 662499
rect 0 661925 41713 662401
rect 0 661757 41657 661925
rect 0 661281 41713 661757
rect 0 661113 41657 661281
rect 0 660729 41713 661113
rect 0 660561 41657 660729
rect 0 660085 41713 660561
rect 0 659917 41657 660085
rect 0 659441 41713 659917
rect 0 659273 41657 659441
rect 0 658889 41713 659273
rect 0 658721 41657 658889
rect 0 658245 41713 658721
rect 0 658077 41657 658245
rect 41713 658133 42193 658189
rect 0 657601 41713 658077
rect 41800 657694 41828 658133
rect 41788 657688 41840 657694
rect 41788 657630 41840 657636
rect 0 657433 41657 657601
rect 0 657049 41713 657433
rect 0 656881 41657 657049
rect 0 656405 41713 656881
rect 0 656237 41657 656405
rect 0 655761 41713 656237
rect 0 655593 41657 655761
rect 0 655209 41713 655593
rect 0 655041 41657 655209
rect 41713 655097 42193 655153
rect 0 654842 41713 655041
rect 0 627373 41713 627583
rect 0 627205 41657 627373
rect 41713 627314 42193 627317
rect 41713 627286 42288 627314
rect 41713 627261 42193 627286
rect 0 626729 41713 627205
rect 0 626561 41657 626729
rect 0 626085 41713 626561
rect 0 625917 41657 626085
rect 41713 625973 42193 626029
rect 41788 625932 41840 625938
rect 0 625533 41713 625917
rect 41788 625874 41840 625880
rect 0 625365 41657 625533
rect 41800 625477 41828 625874
rect 41713 625421 42193 625477
rect 0 624889 41713 625365
rect 0 624721 41657 624889
rect 0 624245 41713 624721
rect 0 624077 41657 624245
rect 41713 624133 42193 624189
rect 0 623693 41713 624077
rect 0 623525 41657 623693
rect 41713 623581 42193 623637
rect 0 623049 41713 623525
rect 0 622881 41657 623049
rect 0 622405 41713 622881
rect 0 622237 41657 622405
rect 41713 622293 42193 622349
rect 0 621853 41713 622237
rect 0 621685 41657 621853
rect 0 621209 41713 621685
rect 0 621041 41657 621209
rect 0 620565 41713 621041
rect 0 620397 41657 620565
rect 0 620013 41713 620397
rect 0 619845 41657 620013
rect 0 619369 41713 619845
rect 42260 619426 42288 627286
rect 42444 625938 42472 662471
rect 42536 657694 42564 700946
rect 42524 657688 42576 657694
rect 42524 657630 42576 657636
rect 42536 633554 42564 657630
rect 42524 633548 42576 633554
rect 42524 633490 42576 633496
rect 42524 633344 42576 633350
rect 42524 633286 42576 633292
rect 42432 625932 42484 625938
rect 42432 625874 42484 625880
rect 41800 619398 42288 619426
rect 0 619201 41657 619369
rect 41800 619313 41828 619398
rect 41713 619257 42193 619313
rect 0 618725 41713 619201
rect 0 618557 41657 618725
rect 0 618081 41713 618557
rect 0 617913 41657 618081
rect 0 617529 41713 617913
rect 0 617361 41657 617529
rect 0 616885 41713 617361
rect 0 616717 41657 616885
rect 0 616241 41713 616717
rect 0 616073 41657 616241
rect 0 615689 41713 616073
rect 0 615521 41657 615689
rect 0 615045 41713 615521
rect 0 614877 41657 615045
rect 41713 614933 42193 614989
rect 0 614401 41713 614877
rect 41800 614446 41828 614933
rect 41788 614440 41840 614446
rect 0 614233 41657 614401
rect 41788 614382 41840 614388
rect 0 613849 41713 614233
rect 0 613681 41657 613849
rect 0 613205 41713 613681
rect 0 613037 41657 613205
rect 0 612561 41713 613037
rect 0 612393 41657 612561
rect 0 612009 41713 612393
rect 0 611841 41657 612009
rect 41713 611897 42193 611953
rect 0 611642 41713 611841
rect 0 584173 41713 584383
rect 0 584005 41657 584173
rect 41713 584103 42193 584117
rect 41713 584075 42288 584103
rect 41713 584061 42193 584075
rect 0 583529 41713 584005
rect 0 583361 41657 583529
rect 0 582885 41713 583361
rect 0 582717 41657 582885
rect 41713 582773 42193 582829
rect 0 582333 41713 582717
rect 0 582165 41657 582333
rect 41713 582221 42193 582277
rect 0 581689 41713 582165
rect 41800 581738 41828 582221
rect 41788 581732 41840 581738
rect 0 581521 41657 581689
rect 41788 581674 41840 581680
rect 0 581045 41713 581521
rect 0 580877 41657 581045
rect 41713 580933 42193 580989
rect 0 580493 41713 580877
rect 0 580325 41657 580493
rect 41713 580381 42193 580437
rect 0 579849 41713 580325
rect 0 579681 41657 579849
rect 0 579205 41713 579681
rect 0 579037 41657 579205
rect 41713 579093 42193 579149
rect 0 578653 41713 579037
rect 0 578485 41657 578653
rect 0 578009 41713 578485
rect 0 577841 41657 578009
rect 0 577365 41713 577841
rect 0 577197 41657 577365
rect 0 576813 41713 577197
rect 0 576645 41657 576813
rect 0 576169 41713 576645
rect 42260 576178 42288 584075
rect 42444 581738 42472 625874
rect 42536 614446 42564 633286
rect 42524 614440 42576 614446
rect 42524 614382 42576 614388
rect 42432 581732 42484 581738
rect 42432 581674 42484 581680
rect 0 576001 41657 576169
rect 41892 576150 42288 576178
rect 41892 576113 41920 576150
rect 41713 576057 42193 576113
rect 0 575525 41713 576001
rect 0 575357 41657 575525
rect 0 574881 41713 575357
rect 0 574713 41657 574881
rect 0 574329 41713 574713
rect 0 574161 41657 574329
rect 0 573685 41713 574161
rect 0 573517 41657 573685
rect 0 573041 41713 573517
rect 0 572873 41657 573041
rect 0 572489 41713 572873
rect 0 572321 41657 572489
rect 0 571845 41713 572321
rect 41788 572280 41840 572286
rect 41788 572222 41840 572228
rect 42248 572280 42300 572286
rect 42248 572222 42300 572228
rect 0 571677 41657 571845
rect 41800 571789 41828 572222
rect 41713 571733 42193 571789
rect 0 571201 41713 571677
rect 0 571033 41657 571201
rect 0 570649 41713 571033
rect 0 570481 41657 570649
rect 0 570005 41713 570481
rect 0 569837 41657 570005
rect 0 569361 41713 569837
rect 0 569193 41657 569361
rect 0 568809 41713 569193
rect 0 568641 41657 568809
rect 41713 568697 42193 568753
rect 0 568442 41713 568641
rect 0 540973 41713 541183
rect 42260 541090 42288 572222
rect 42260 541062 42380 541090
rect 0 540805 41657 540973
rect 41713 540903 42193 540917
rect 41713 540875 42288 540903
rect 41713 540861 42193 540875
rect 0 540329 41713 540805
rect 0 540161 41657 540329
rect 0 539685 41713 540161
rect 0 539517 41657 539685
rect 41713 539573 42193 539629
rect 0 539133 41713 539517
rect 0 538965 41657 539133
rect 41713 539021 42193 539077
rect 0 538489 41713 538965
rect 41800 538558 41828 539021
rect 41788 538552 41840 538558
rect 41788 538494 41840 538500
rect 0 538321 41657 538489
rect 0 537845 41713 538321
rect 0 537677 41657 537845
rect 41713 537733 42193 537789
rect 0 537293 41713 537677
rect 0 537125 41657 537293
rect 41713 537181 42193 537237
rect 0 536649 41713 537125
rect 0 536481 41657 536649
rect 0 536005 41713 536481
rect 0 535837 41657 536005
rect 41713 535893 42193 535949
rect 0 535453 41713 535837
rect 0 535285 41657 535453
rect 0 534809 41713 535285
rect 0 534641 41657 534809
rect 0 534165 41713 534641
rect 0 533997 41657 534165
rect 0 533613 41713 533997
rect 0 533445 41657 533613
rect 0 532969 41713 533445
rect 0 532801 41657 532969
rect 42260 532930 42288 540875
rect 41708 532902 42288 532930
rect 41708 532885 42193 532902
rect 41713 532857 42193 532885
rect 0 532325 41713 532801
rect 0 532157 41657 532325
rect 0 531681 41713 532157
rect 0 531513 41657 531681
rect 0 531129 41713 531513
rect 0 530961 41657 531129
rect 0 530485 41713 530961
rect 0 530317 41657 530485
rect 0 529841 41713 530317
rect 0 529673 41657 529841
rect 0 529289 41713 529673
rect 0 529121 41657 529289
rect 0 528645 41713 529121
rect 42352 528850 42380 541062
rect 42444 538558 42472 581674
rect 42536 572286 42564 614382
rect 42524 572280 42576 572286
rect 42524 572222 42576 572228
rect 42432 538552 42484 538558
rect 42484 538500 42564 538506
rect 42432 538494 42564 538500
rect 42444 538478 42564 538494
rect 41892 528822 42380 528850
rect 0 528477 41657 528645
rect 41892 528589 41920 528822
rect 41713 528533 42193 528589
rect 0 528001 41713 528477
rect 0 527833 41657 528001
rect 0 527449 41713 527833
rect 0 527281 41657 527449
rect 0 526805 41713 527281
rect 0 526637 41657 526805
rect 0 526161 41713 526637
rect 0 525993 41657 526161
rect 0 525609 41713 525993
rect 0 525441 41657 525609
rect 41713 525497 42193 525553
rect 0 525242 41713 525441
rect 985 493022 34812 497858
rect 34868 493078 40000 497858
rect 985 487935 39593 493022
rect 39776 492969 39804 493078
rect 39762 492960 39818 492969
rect 39762 492895 39818 492904
rect 985 483053 39533 487935
rect 39589 483099 40000 487879
rect 39396 458244 39448 458250
rect 39396 458186 39448 458192
rect 39408 455740 39436 458186
rect 714 451687 38812 455740
rect 38868 451874 39600 455740
rect 39946 455424 40002 455433
rect 39946 455359 40002 455368
rect 39670 451888 39726 451897
rect 38868 451846 39670 451874
rect 38868 451743 39600 451846
rect 39670 451823 39726 451832
rect 714 449744 39593 451687
rect 714 447632 39479 449744
rect 39535 447794 39600 449688
rect 39856 448316 39908 448322
rect 39856 448258 39908 448264
rect 39868 447794 39896 448258
rect 39535 447766 39896 447794
rect 39535 447688 39600 447766
rect 714 444955 39593 447632
rect 714 440900 39247 444955
rect 39303 440994 39600 444899
rect 39670 441008 39726 441017
rect 39303 440966 39670 440994
rect 39303 440900 39600 440966
rect 39960 440994 39988 455359
rect 42260 448322 42288 528822
rect 42248 448316 42300 448322
rect 42248 448258 42300 448264
rect 39726 440966 39988 440994
rect 39670 440943 39726 440952
rect 0 413373 41713 413583
rect 42260 413438 42288 448258
rect 42248 413432 42300 413438
rect 42248 413374 42300 413380
rect 0 413205 41657 413373
rect 41713 413303 42193 413317
rect 41713 413275 42288 413303
rect 41713 413261 42193 413275
rect 0 412729 41713 413205
rect 0 412561 41657 412729
rect 0 412085 41713 412561
rect 0 411917 41657 412085
rect 41713 411973 42193 412029
rect 0 411533 41713 411917
rect 0 411365 41657 411533
rect 41722 411477 41828 411482
rect 41713 411421 42193 411477
rect 0 410889 41713 411365
rect 41800 410990 41828 411421
rect 41788 410984 41840 410990
rect 41788 410926 41840 410932
rect 0 410721 41657 410889
rect 0 410245 41713 410721
rect 0 410077 41657 410245
rect 41713 410133 42193 410189
rect 0 409693 41713 410077
rect 0 409525 41657 409693
rect 41713 409581 42193 409637
rect 0 409049 41713 409525
rect 0 408881 41657 409049
rect 0 408405 41713 408881
rect 0 408237 41657 408405
rect 41713 408293 42193 408349
rect 0 407853 41713 408237
rect 0 407685 41657 407853
rect 0 407209 41713 407685
rect 0 407041 41657 407209
rect 0 406565 41713 407041
rect 0 406397 41657 406565
rect 0 406013 41713 406397
rect 0 405845 41657 406013
rect 0 405369 41713 405845
rect 0 405201 41657 405369
rect 41713 405299 42193 405313
rect 42260 405299 42288 413275
rect 41713 405271 42288 405299
rect 41713 405257 42193 405271
rect 0 404725 41713 405201
rect 0 404557 41657 404725
rect 0 404081 41713 404557
rect 0 403913 41657 404081
rect 0 403529 41713 403913
rect 0 403361 41657 403529
rect 0 402885 41713 403361
rect 0 402717 41657 402885
rect 0 402241 41713 402717
rect 0 402073 41657 402241
rect 0 401689 41713 402073
rect 0 401521 41657 401689
rect 41788 401532 41840 401538
rect 0 401045 41713 401521
rect 41788 401474 41840 401480
rect 42248 401532 42300 401538
rect 42248 401474 42300 401480
rect 0 400877 41657 401045
rect 41800 400989 41828 401474
rect 41713 400933 42193 400989
rect 0 400401 41713 400877
rect 0 400233 41657 400401
rect 0 399849 41713 400233
rect 42260 400217 42288 401474
rect 42246 400208 42302 400217
rect 42536 410990 42564 538478
rect 42616 413432 42668 413438
rect 42616 413374 42668 413380
rect 42524 410984 42576 410990
rect 42524 410926 42576 410932
rect 42246 400143 42302 400152
rect 0 399681 41657 399849
rect 0 399205 41713 399681
rect 0 399037 41657 399205
rect 0 398561 41713 399037
rect 0 398393 41657 398561
rect 0 398009 41713 398393
rect 0 397841 41657 398009
rect 41713 397897 42193 397953
rect 0 397642 41713 397841
rect 42340 380928 42392 380934
rect 42340 380870 42392 380876
rect 0 370173 41713 370383
rect 0 370005 41657 370173
rect 41713 370103 42193 370117
rect 41713 370075 42288 370103
rect 41713 370061 42193 370075
rect 0 369529 41713 370005
rect 0 369361 41657 369529
rect 0 368885 41713 369361
rect 0 368717 41657 368885
rect 41713 368773 42193 368829
rect 0 368333 41713 368717
rect 41788 368688 41840 368694
rect 41788 368630 41840 368636
rect 0 368165 41657 368333
rect 41800 368277 41828 368630
rect 41713 368221 42193 368277
rect 0 367689 41713 368165
rect 0 367521 41657 367689
rect 0 367045 41713 367521
rect 0 366877 41657 367045
rect 41713 366933 42193 366989
rect 0 366493 41713 366877
rect 0 366325 41657 366493
rect 41713 366381 42193 366437
rect 0 365849 41713 366325
rect 0 365681 41657 365849
rect 0 365205 41713 365681
rect 0 365037 41657 365205
rect 41713 365093 42193 365149
rect 0 364653 41713 365037
rect 0 364485 41657 364653
rect 0 364009 41713 364485
rect 0 363841 41657 364009
rect 0 363365 41713 363841
rect 0 363197 41657 363365
rect 0 362813 41713 363197
rect 0 362645 41657 362813
rect 0 362169 41713 362645
rect 42260 362250 42288 370075
rect 41892 362222 42288 362250
rect 0 362001 41657 362169
rect 41892 362114 41920 362222
rect 41722 362113 41920 362114
rect 41713 362057 42193 362113
rect 0 361525 41713 362001
rect 0 361357 41657 361525
rect 0 360881 41713 361357
rect 0 360713 41657 360881
rect 0 360329 41713 360713
rect 0 360161 41657 360329
rect 0 359685 41713 360161
rect 0 359517 41657 359685
rect 0 359041 41713 359517
rect 0 358873 41657 359041
rect 0 358489 41713 358873
rect 0 358321 41657 358489
rect 0 357845 41713 358321
rect 0 357677 41657 357845
rect 41713 357733 42193 357789
rect 0 357201 41713 357677
rect 41800 357542 41828 357733
rect 42352 357542 42380 380870
rect 41788 357536 41840 357542
rect 41788 357478 41840 357484
rect 42340 357536 42392 357542
rect 42340 357478 42392 357484
rect 0 357033 41657 357201
rect 0 356649 41713 357033
rect 42536 368694 42564 410926
rect 42628 401538 42656 413374
rect 42616 401532 42668 401538
rect 42616 401474 42668 401480
rect 42614 400208 42670 400217
rect 42614 400143 42670 400152
rect 42628 380934 42656 400143
rect 42616 380928 42668 380934
rect 42616 380870 42668 380876
rect 42524 368688 42576 368694
rect 42524 368630 42576 368636
rect 42536 367062 42564 368630
rect 42524 367056 42576 367062
rect 42524 366998 42576 367004
rect 42800 366988 42852 366994
rect 42800 366930 42852 366936
rect 42616 357536 42668 357542
rect 42616 357478 42668 357484
rect 0 356481 41657 356649
rect 0 356005 41713 356481
rect 0 355837 41657 356005
rect 0 355361 41713 355837
rect 0 355193 41657 355361
rect 0 354809 41713 355193
rect 0 354641 41657 354809
rect 41713 354697 42193 354753
rect 0 354442 41713 354641
rect 42340 334688 42392 334694
rect 42340 334630 42392 334636
rect 0 326973 41713 327183
rect 0 326805 41657 326973
rect 41713 326890 42193 326917
rect 41713 326862 42288 326890
rect 41713 326861 42193 326862
rect 0 326329 41713 326805
rect 0 326161 41657 326329
rect 0 325685 41713 326161
rect 0 325517 41657 325685
rect 41713 325573 42193 325629
rect 0 325133 41713 325517
rect 0 324965 41657 325133
rect 41713 325021 42193 325077
rect 0 324489 41713 324965
rect 41800 324562 41828 325021
rect 41788 324556 41840 324562
rect 41788 324498 41840 324504
rect 0 324321 41657 324489
rect 0 323845 41713 324321
rect 0 323677 41657 323845
rect 41713 323733 42193 323789
rect 0 323293 41713 323677
rect 0 323125 41657 323293
rect 41713 323181 42193 323237
rect 0 322649 41713 323125
rect 0 322481 41657 322649
rect 0 322005 41713 322481
rect 0 321837 41657 322005
rect 41713 321893 42193 321949
rect 0 321453 41713 321837
rect 0 321285 41657 321453
rect 0 320809 41713 321285
rect 0 320641 41657 320809
rect 0 320165 41713 320641
rect 0 319997 41657 320165
rect 0 319613 41713 319997
rect 0 319445 41657 319613
rect 0 318969 41713 319445
rect 0 318801 41657 318969
rect 41713 318899 42193 318913
rect 42260 318899 42288 326862
rect 41713 318871 42288 318899
rect 41713 318857 42193 318871
rect 0 318325 41713 318801
rect 0 318157 41657 318325
rect 0 317681 41713 318157
rect 0 317513 41657 317681
rect 0 317129 41713 317513
rect 0 316961 41657 317129
rect 0 316485 41713 316961
rect 0 316317 41657 316485
rect 0 315841 41713 316317
rect 0 315673 41657 315841
rect 0 315289 41713 315673
rect 0 315121 41657 315289
rect 0 314645 41713 315121
rect 0 314477 41657 314645
rect 42352 314634 42380 334630
rect 42340 314628 42392 314634
rect 41713 314533 42193 314589
rect 42340 314570 42392 314576
rect 41800 314498 41828 314533
rect 41788 314492 41840 314498
rect 0 314001 41713 314477
rect 41788 314434 41840 314440
rect 0 313833 41657 314001
rect 0 313449 41713 313833
rect 42628 334694 42656 357478
rect 42812 347834 42840 366930
rect 42720 347806 42840 347834
rect 42720 347750 42748 347806
rect 42708 347744 42760 347750
rect 42708 347686 42760 347692
rect 42892 347744 42944 347750
rect 42892 347686 42944 347692
rect 42616 334688 42668 334694
rect 42616 334630 42668 334636
rect 42904 328506 42932 347686
rect 42616 328500 42668 328506
rect 42616 328442 42668 328448
rect 42892 328500 42944 328506
rect 42892 328442 42944 328448
rect 42524 324488 42576 324494
rect 42628 324442 42656 328442
rect 42576 324436 42656 324442
rect 42524 324430 42656 324436
rect 42536 324414 42656 324430
rect 42536 314498 42564 324414
rect 42616 314560 42668 314566
rect 42616 314502 42668 314508
rect 42524 314492 42576 314498
rect 42524 314434 42576 314440
rect 0 313281 41657 313449
rect 0 312805 41713 313281
rect 0 312637 41657 312805
rect 0 312161 41713 312637
rect 0 311993 41657 312161
rect 0 311609 41713 311993
rect 0 311441 41657 311609
rect 41713 311497 42193 311553
rect 0 311242 41713 311441
rect 42628 295474 42656 314502
rect 42800 314492 42852 314498
rect 42800 314434 42852 314440
rect 42536 295446 42656 295474
rect 0 283773 41713 283983
rect 0 283605 41657 283773
rect 41713 283661 42193 283717
rect 0 283129 41713 283605
rect 41892 283234 41920 283661
rect 41892 283206 42288 283234
rect 0 282961 41657 283129
rect 0 282485 41713 282961
rect 0 282317 41657 282485
rect 41713 282373 42193 282429
rect 41788 282328 41840 282334
rect 0 281933 41713 282317
rect 41788 282270 41840 282276
rect 0 281765 41657 281933
rect 41800 281877 41828 282270
rect 41713 281821 42193 281877
rect 0 281289 41713 281765
rect 0 281121 41657 281289
rect 0 280645 41713 281121
rect 0 280477 41657 280645
rect 41713 280533 42193 280589
rect 0 280093 41713 280477
rect 0 279925 41657 280093
rect 41713 279981 42193 280037
rect 0 279449 41713 279925
rect 0 279281 41657 279449
rect 0 278805 41713 279281
rect 0 278637 41657 278805
rect 41713 278693 42193 278749
rect 0 278253 41713 278637
rect 0 278085 41657 278253
rect 0 277609 41713 278085
rect 0 277441 41657 277609
rect 0 276965 41713 277441
rect 0 276797 41657 276965
rect 0 276413 41713 276797
rect 0 276245 41657 276413
rect 0 275769 41713 276245
rect 0 275601 41657 275769
rect 41713 275657 42193 275713
rect 41800 275618 41828 275657
rect 42260 275618 42288 283206
rect 42432 282328 42484 282334
rect 42432 282270 42484 282276
rect 0 275125 41713 275601
rect 41800 275590 42288 275618
rect 0 274957 41657 275125
rect 0 274481 41713 274957
rect 0 274313 41657 274481
rect 0 273929 41713 274313
rect 0 273761 41657 273929
rect 0 273285 41713 273761
rect 0 273117 41657 273285
rect 0 272641 41713 273117
rect 0 272473 41657 272641
rect 0 272089 41713 272473
rect 0 271921 41657 272089
rect 0 271445 41713 271921
rect 0 271277 41657 271445
rect 41722 271389 41828 271402
rect 41713 271333 42193 271389
rect 0 270801 41713 271277
rect 41800 270842 41828 271333
rect 41788 270836 41840 270842
rect 0 270633 41657 270801
rect 41788 270778 41840 270784
rect 0 270249 41713 270633
rect 0 270081 41657 270249
rect 0 269605 41713 270081
rect 0 269437 41657 269605
rect 0 268961 41713 269437
rect 0 268793 41657 268961
rect 0 268409 41713 268793
rect 0 268241 41657 268409
rect 41713 268297 42193 268353
rect 0 268042 41713 268241
rect 0 240573 41713 240783
rect 0 240405 41657 240573
rect 41722 240517 42288 240530
rect 41713 240502 42288 240517
rect 41713 240461 42193 240502
rect 0 239929 41713 240405
rect 0 239761 41657 239929
rect 0 239285 41713 239761
rect 0 239117 41657 239285
rect 41713 239173 42193 239229
rect 0 238733 41713 239117
rect 41788 239080 41840 239086
rect 41788 239022 41840 239028
rect 0 238565 41657 238733
rect 41800 238677 41828 239022
rect 41713 238621 42193 238677
rect 0 238089 41713 238565
rect 0 237921 41657 238089
rect 0 237445 41713 237921
rect 0 237277 41657 237445
rect 41713 237333 42193 237389
rect 0 236893 41713 237277
rect 0 236725 41657 236893
rect 41713 236781 42193 236837
rect 0 236249 41713 236725
rect 0 236081 41657 236249
rect 0 235605 41713 236081
rect 0 235437 41657 235605
rect 41713 235493 42193 235549
rect 0 235053 41713 235437
rect 0 234885 41657 235053
rect 0 234409 41713 234885
rect 0 234241 41657 234409
rect 0 233765 41713 234241
rect 0 233597 41657 233765
rect 0 233213 41713 233597
rect 0 233045 41657 233213
rect 0 232569 41713 233045
rect 42260 232642 42288 240502
rect 42444 239086 42472 282270
rect 42536 282146 42564 295446
rect 42616 295384 42668 295390
rect 42616 295326 42668 295332
rect 42628 282334 42656 295326
rect 42616 282328 42668 282334
rect 42616 282270 42668 282276
rect 42812 295390 42840 314434
rect 42800 295384 42852 295390
rect 42800 295326 42852 295332
rect 42536 282118 42840 282146
rect 42524 276004 42576 276010
rect 42524 275946 42576 275952
rect 42536 270842 42564 275946
rect 42524 270836 42576 270842
rect 42524 270778 42576 270784
rect 42432 239080 42484 239086
rect 42432 239022 42484 239028
rect 41892 232614 42288 232642
rect 0 232401 41657 232569
rect 41892 232513 41920 232614
rect 41713 232457 42193 232513
rect 0 231925 41713 232401
rect 0 231757 41657 231925
rect 0 231281 41713 231757
rect 0 231113 41657 231281
rect 0 230729 41713 231113
rect 0 230561 41657 230729
rect 0 230085 41713 230561
rect 0 229917 41657 230085
rect 0 229441 41713 229917
rect 0 229273 41657 229441
rect 0 228889 41713 229273
rect 0 228721 41657 228889
rect 0 228245 41713 228721
rect 42536 228682 42564 270778
rect 42812 276010 42840 282118
rect 42800 276004 42852 276010
rect 42800 275946 42852 275952
rect 42616 239080 42668 239086
rect 42616 239022 42668 239028
rect 41788 228676 41840 228682
rect 41788 228618 41840 228624
rect 42524 228676 42576 228682
rect 42524 228618 42576 228624
rect 0 228077 41657 228245
rect 41800 228189 41828 228618
rect 41713 228133 42193 228189
rect 41722 228126 41828 228133
rect 0 227601 41713 228077
rect 0 227433 41657 227601
rect 42248 227928 42300 227934
rect 42248 227870 42300 227876
rect 0 227049 41713 227433
rect 0 226881 41657 227049
rect 0 226405 41713 226881
rect 0 226237 41657 226405
rect 0 225761 41713 226237
rect 0 225593 41657 225761
rect 0 225209 41713 225593
rect 0 225041 41657 225209
rect 41713 225097 42193 225153
rect 0 224842 41713 225041
rect 0 197373 41713 197583
rect 0 197205 41657 197373
rect 41713 197261 42193 197317
rect 41722 197254 41828 197261
rect 0 196729 41713 197205
rect 41800 196790 41828 197254
rect 41788 196784 41840 196790
rect 0 196561 41657 196729
rect 41788 196726 41840 196732
rect 0 196085 41713 196561
rect 0 195917 41657 196085
rect 41713 195973 42193 196029
rect 0 195533 41713 195917
rect 41788 195900 41840 195906
rect 41788 195842 41840 195848
rect 0 195365 41657 195533
rect 41800 195477 41828 195842
rect 41713 195421 42193 195477
rect 0 194889 41713 195365
rect 0 194721 41657 194889
rect 0 194245 41713 194721
rect 0 194077 41657 194245
rect 41713 194133 42193 194189
rect 0 193693 41713 194077
rect 0 193525 41657 193693
rect 41713 193581 42193 193637
rect 0 193049 41713 193525
rect 0 192881 41657 193049
rect 0 192405 41713 192881
rect 0 192237 41657 192405
rect 41713 192293 42193 192349
rect 0 191853 41713 192237
rect 0 191685 41657 191853
rect 0 191209 41713 191685
rect 0 191041 41657 191209
rect 0 190565 41713 191041
rect 0 190397 41657 190565
rect 0 190013 41713 190397
rect 0 189845 41657 190013
rect 41788 189848 41840 189854
rect 0 189369 41713 189845
rect 41788 189790 41840 189796
rect 0 189201 41657 189369
rect 41800 189313 41828 189790
rect 41713 189257 42193 189313
rect 0 188725 41713 189201
rect 0 188557 41657 188725
rect 0 188081 41713 188557
rect 0 187913 41657 188081
rect 0 187529 41713 187913
rect 0 187361 41657 187529
rect 0 186885 41713 187361
rect 0 186717 41657 186885
rect 0 186241 41713 186717
rect 0 186073 41657 186241
rect 0 185689 41713 186073
rect 0 185521 41657 185689
rect 0 185045 41713 185521
rect 0 184877 41657 185045
rect 41713 184933 42193 184989
rect 0 184401 41713 184877
rect 41800 184498 41828 184933
rect 42260 184498 42288 227870
rect 42340 196784 42392 196790
rect 42340 196726 42392 196732
rect 42352 189854 42380 196726
rect 42340 189848 42392 189854
rect 42340 189790 42392 189796
rect 41800 184470 42380 184498
rect 0 184233 41657 184401
rect 0 183849 41713 184233
rect 0 183681 41657 183849
rect 0 183205 41713 183681
rect 0 183037 41657 183205
rect 0 182561 41713 183037
rect 0 182393 41657 182561
rect 0 182009 41713 182393
rect 0 181841 41657 182009
rect 41713 181897 42193 181953
rect 0 181642 41713 181841
rect 985 120222 34812 125058
rect 34868 120278 40000 125058
rect 985 115135 39593 120222
rect 39776 120193 39804 120278
rect 39762 120184 39818 120193
rect 39762 120119 39818 120128
rect 41418 115968 41474 115977
rect 41418 115903 41474 115912
rect 985 110253 39533 115135
rect 39589 110299 40000 115079
rect 39394 84280 39450 84289
rect 39394 84215 39450 84224
rect 39408 82940 39436 84215
rect 714 78887 38812 82940
rect 38868 78962 39600 82940
rect 38868 78943 39712 78962
rect 39500 78934 39712 78943
rect 714 76944 39593 78887
rect 714 74832 39479 76944
rect 39535 75154 39600 76888
rect 39684 75274 39712 78934
rect 39672 75268 39724 75274
rect 39672 75210 39724 75216
rect 39535 75126 39804 75154
rect 39535 74990 39620 75126
rect 39672 74996 39724 75002
rect 39535 74888 39600 74990
rect 39672 74938 39724 74944
rect 714 72155 39593 74832
rect 714 68098 39247 72155
rect 39303 68218 39600 72099
rect 39303 68100 39620 68218
rect 39592 67998 39620 68100
rect 39580 67992 39632 67998
rect 39580 67934 39632 67940
rect 39684 52426 39712 74938
rect 39672 52420 39724 52426
rect 39672 52362 39724 52368
rect 39776 47734 39804 75126
rect 41432 67998 41460 115903
rect 41420 67992 41472 67998
rect 41420 67934 41472 67940
rect 41432 64666 41460 67934
rect 41420 64660 41472 64666
rect 41420 64602 41472 64608
rect 39856 52420 39908 52426
rect 39856 52362 39908 52368
rect 39868 47870 39896 52362
rect 39856 47864 39908 47870
rect 39856 47806 39908 47812
rect 39764 47728 39816 47734
rect 39764 47670 39816 47676
rect 42352 115977 42380 184470
rect 42536 227934 42564 228618
rect 42524 227928 42576 227934
rect 42524 227870 42576 227876
rect 42628 195906 42656 239022
rect 42616 195900 42668 195906
rect 42616 195842 42668 195848
rect 44192 120193 44220 879786
rect 44284 458250 44312 922898
rect 44362 917280 44418 917289
rect 44362 917215 44418 917224
rect 44272 458244 44324 458250
rect 44272 458186 44324 458192
rect 44376 448633 44404 917215
rect 45940 879866 45968 996503
rect 76242 995943 92183 1037600
rect 76242 995887 76441 995943
rect 76609 995887 76993 995943
rect 77161 995887 77637 995943
rect 77805 995887 78281 995943
rect 78449 995887 78833 995943
rect 79001 995887 79477 995943
rect 79645 995887 80121 995943
rect 80289 995887 80673 995943
rect 80841 995887 81317 995943
rect 81485 995887 81961 995943
rect 82129 995887 82513 995943
rect 82681 995887 83157 995943
rect 83325 995887 83801 995943
rect 83969 995887 84445 995943
rect 84613 995887 84997 995943
rect 85165 995887 85641 995943
rect 85809 995887 86285 995943
rect 86453 995887 86837 995943
rect 87005 995887 87481 995943
rect 87649 995887 88125 995943
rect 88293 995887 88677 995943
rect 88845 995887 89321 995943
rect 89489 995887 89965 995943
rect 90133 995887 90517 995943
rect 90685 995887 91161 995943
rect 91329 995887 91805 995943
rect 91973 995887 92183 995943
rect 127642 995943 143583 1037600
rect 127642 995887 127841 995943
rect 128009 995887 128393 995943
rect 128561 995887 129037 995943
rect 129205 995887 129681 995943
rect 129849 995887 130233 995943
rect 130401 995887 130877 995943
rect 131045 995887 131521 995943
rect 131689 995887 132073 995943
rect 132241 995887 132717 995943
rect 132885 995887 133361 995943
rect 133529 995887 133913 995943
rect 134081 995887 134557 995943
rect 134725 995887 135201 995943
rect 135369 995887 135845 995943
rect 136013 995887 136397 995943
rect 136565 995887 137041 995943
rect 137209 995887 137685 995943
rect 137853 995887 138237 995943
rect 138405 995887 138881 995943
rect 139049 995887 139525 995943
rect 139693 995887 140077 995943
rect 140245 995887 140721 995943
rect 140889 995887 141365 995943
rect 141533 995887 141917 995943
rect 142085 995887 142561 995943
rect 142729 995887 143205 995943
rect 143373 995887 143583 995943
rect 179042 995943 194983 1037600
rect 179042 995887 179241 995943
rect 179409 995887 179793 995943
rect 179961 995887 180437 995943
rect 180605 995887 181081 995943
rect 181249 995887 181633 995943
rect 181801 995887 182277 995943
rect 182445 995887 182921 995943
rect 183089 995887 183473 995943
rect 183641 995887 184117 995943
rect 184285 995887 184761 995943
rect 184929 995887 185313 995943
rect 185481 995887 185957 995943
rect 186125 995887 186601 995943
rect 186769 995887 187245 995943
rect 187413 995887 187797 995943
rect 187965 995887 188441 995943
rect 188609 995887 189085 995943
rect 189253 995887 189637 995943
rect 189805 995887 190281 995943
rect 190449 995887 190925 995943
rect 191093 995887 191477 995943
rect 191645 995887 192121 995943
rect 192289 995887 192765 995943
rect 192933 995887 193317 995943
rect 193485 995887 193961 995943
rect 194129 995887 194605 995943
rect 194773 995887 194983 995943
rect 230442 995943 246383 1037600
rect 230442 995887 230641 995943
rect 230809 995887 231193 995943
rect 231361 995887 231837 995943
rect 232005 995887 232481 995943
rect 232649 995887 233033 995943
rect 233201 995887 233677 995943
rect 233845 995887 234321 995943
rect 234489 995887 234873 995943
rect 235041 995887 235517 995943
rect 235685 995887 236161 995943
rect 236329 995887 236713 995943
rect 236881 995887 237357 995943
rect 237525 995887 238001 995943
rect 238169 995887 238645 995943
rect 238813 995887 239197 995943
rect 239365 995887 239841 995943
rect 240009 995887 240485 995943
rect 240653 995887 241037 995943
rect 241205 995887 241681 995943
rect 241849 995887 242325 995943
rect 242493 995887 242877 995943
rect 243045 995887 243521 995943
rect 243689 995887 244165 995943
rect 244333 995887 244717 995943
rect 244885 995887 245361 995943
rect 245529 995887 246005 995943
rect 246173 995887 246383 995943
rect 282042 995943 297983 1037600
rect 333453 1002788 348258 1036615
rect 333453 998067 343422 1002788
rect 333499 997656 338279 998011
rect 338335 998007 343422 998067
rect 333499 997600 333518 997656
rect 333574 997600 338279 997656
rect 343478 997600 348258 1002732
rect 333518 997591 333574 997600
rect 282042 995887 282241 995943
rect 282409 995887 282793 995943
rect 282961 995887 283437 995943
rect 283605 995887 284081 995943
rect 284249 995887 284633 995943
rect 284801 995887 285277 995943
rect 285445 995887 285921 995943
rect 286089 995887 286473 995943
rect 286641 995887 287117 995943
rect 287285 995887 287761 995943
rect 287929 995887 288313 995943
rect 288481 995887 288957 995943
rect 289125 995887 289601 995943
rect 289769 995887 290245 995943
rect 290413 995887 290797 995943
rect 290965 995887 291441 995943
rect 291609 995887 292085 995943
rect 292253 995887 292637 995943
rect 292805 995887 293281 995943
rect 293449 995887 293925 995943
rect 294093 995887 294477 995943
rect 294645 995887 295121 995943
rect 295289 995887 295765 995943
rect 295933 995887 296317 995943
rect 296485 995887 296961 995943
rect 297129 995887 297605 995943
rect 297773 995887 297983 995943
rect 76497 995407 76553 995887
rect 79533 995452 79589 995887
rect 79520 995407 79589 995452
rect 83857 995661 83913 995887
rect 83857 995654 84056 995661
rect 83857 995648 84068 995654
rect 83857 995633 84016 995648
rect 83857 995407 83913 995633
rect 84016 995590 84068 995596
rect 86893 995407 86949 995887
rect 88181 995407 88237 995887
rect 88733 995407 88789 995887
rect 90021 995452 90077 995887
rect 90008 995407 90077 995452
rect 90573 995407 90629 995887
rect 91744 995648 91796 995654
rect 91744 995590 91796 995596
rect 91756 995466 91784 995590
rect 91861 995466 91917 995887
rect 91756 995438 91917 995466
rect 91861 995407 91917 995438
rect 127897 995407 127953 995887
rect 130933 995407 130989 995887
rect 135257 995466 135313 995887
rect 135352 995512 135404 995518
rect 135257 995460 135352 995466
rect 135257 995454 135404 995460
rect 135257 995438 135392 995454
rect 135257 995407 135313 995438
rect 138293 995407 138349 995887
rect 139581 995407 139637 995887
rect 140133 995407 140189 995887
rect 141421 995407 141477 995887
rect 141973 995407 142029 995887
rect 143172 995512 143224 995518
rect 143261 995466 143317 995887
rect 143224 995460 143317 995466
rect 143172 995454 143317 995460
rect 143184 995438 143317 995454
rect 143261 995407 143317 995438
rect 179297 995407 179353 995887
rect 182333 995466 182389 995887
rect 182333 995407 182404 995466
rect 186657 995466 186713 995887
rect 186657 995407 186728 995466
rect 189693 995407 189749 995887
rect 190981 995407 191037 995887
rect 191533 995407 191589 995887
rect 192821 995466 192877 995887
rect 192821 995407 192892 995466
rect 193373 995407 193429 995887
rect 194661 995466 194717 995887
rect 194661 995407 194732 995466
rect 230697 995407 230753 995887
rect 233733 995466 233789 995887
rect 233712 995407 233789 995466
rect 238057 995466 238113 995887
rect 238208 995648 238260 995654
rect 238208 995590 238260 995596
rect 238220 995466 238248 995590
rect 238057 995438 238248 995466
rect 238057 995407 238113 995438
rect 241093 995407 241149 995887
rect 242381 995407 242437 995887
rect 242933 995407 242989 995887
rect 244221 995466 244277 995887
rect 244200 995407 244277 995466
rect 244773 995407 244829 995887
rect 245936 995648 245988 995654
rect 245936 995590 245988 995596
rect 245948 995466 245976 995590
rect 246061 995466 246117 995887
rect 245948 995438 246117 995466
rect 246061 995407 246117 995438
rect 282297 995407 282353 995887
rect 285333 995452 285389 995887
rect 285324 995407 285389 995452
rect 289657 995452 289713 995887
rect 289648 995407 289713 995452
rect 292693 995407 292749 995887
rect 293981 995407 294037 995887
rect 294533 995407 294589 995887
rect 295821 995452 295877 995887
rect 295812 995407 295877 995452
rect 296373 995407 296429 995887
rect 297661 995452 297717 995887
rect 297652 995407 297717 995452
rect 79520 990690 79548 995407
rect 79508 990684 79560 990690
rect 79508 990626 79560 990632
rect 79968 990684 80020 990690
rect 79968 990626 80020 990632
rect 79980 990214 80008 990626
rect 90008 990622 90036 995407
rect 130948 990690 130976 995407
rect 141436 992118 141464 995407
rect 141424 992112 141476 992118
rect 141424 992054 141476 992060
rect 154396 992112 154448 992118
rect 154396 992054 154448 992060
rect 141436 990978 141464 992054
rect 141344 990950 141464 990978
rect 130936 990684 130988 990690
rect 130936 990626 130988 990632
rect 89996 990616 90048 990622
rect 89996 990558 90048 990564
rect 79968 990208 80020 990214
rect 79968 990150 80020 990156
rect 90008 990146 90036 990558
rect 141344 990486 141372 990950
rect 141332 990480 141384 990486
rect 141332 990422 141384 990428
rect 154408 990418 154436 992054
rect 182376 990690 182404 995407
rect 182364 990684 182416 990690
rect 182364 990626 182416 990632
rect 186700 990622 186728 995407
rect 186688 990616 186740 990622
rect 186688 990558 186740 990564
rect 164148 990548 164200 990554
rect 164148 990490 164200 990496
rect 154396 990412 154448 990418
rect 154396 990354 154448 990360
rect 154580 990412 154632 990418
rect 154580 990354 154632 990360
rect 154592 990282 154620 990354
rect 164160 990282 164188 990490
rect 192864 990554 192892 995407
rect 194704 990622 194732 995407
rect 231860 995104 231912 995110
rect 231860 995046 231912 995052
rect 194692 990616 194744 990622
rect 193218 990584 193274 990593
rect 192852 990548 192904 990554
rect 194692 990558 194744 990564
rect 193218 990519 193220 990528
rect 192852 990490 192904 990496
rect 193272 990519 193274 990528
rect 193220 990490 193272 990496
rect 212446 990584 212502 990593
rect 231872 990554 231900 995046
rect 212446 990519 212448 990528
rect 212500 990519 212502 990528
rect 231860 990548 231912 990554
rect 212448 990490 212500 990496
rect 231860 990490 231912 990496
rect 233712 990690 233740 995407
rect 244200 995110 244228 995407
rect 244188 995104 244240 995110
rect 244188 995046 244240 995052
rect 244200 990758 244228 995046
rect 244188 990752 244240 990758
rect 244188 990694 244240 990700
rect 233700 990684 233752 990690
rect 233700 990626 233752 990632
rect 285324 990690 285352 995407
rect 289648 995314 289676 995407
rect 289636 995308 289688 995314
rect 289636 995250 289688 995256
rect 285312 990684 285364 990690
rect 285312 990626 285364 990632
rect 295812 990758 295840 995407
rect 297652 995314 297680 995407
rect 297640 995308 297692 995314
rect 297640 995250 297692 995256
rect 295800 990752 295852 990758
rect 295800 990694 295852 990700
rect 333532 990690 333560 997591
rect 383842 995943 399783 1037600
rect 383842 995887 384041 995943
rect 384209 995887 384593 995943
rect 384761 995887 385237 995943
rect 385405 995887 385881 995943
rect 386049 995887 386433 995943
rect 386601 995887 387077 995943
rect 387245 995887 387721 995943
rect 387889 995887 388273 995943
rect 388441 995887 388917 995943
rect 389085 995887 389561 995943
rect 389729 995887 390113 995943
rect 390281 995887 390757 995943
rect 390925 995887 391401 995943
rect 391569 995887 392045 995943
rect 392213 995887 392597 995943
rect 392765 995887 393241 995943
rect 393409 995887 393885 995943
rect 394053 995887 394437 995943
rect 394605 995887 395081 995943
rect 395249 995887 395725 995943
rect 395893 995887 396277 995943
rect 396445 995887 396921 995943
rect 397089 995887 397565 995943
rect 397733 995887 398117 995943
rect 398285 995887 398761 995943
rect 398929 995887 399405 995943
rect 399573 995887 399783 995943
rect 472842 995943 488783 1037600
rect 472842 995887 473041 995943
rect 473209 995887 473593 995943
rect 473761 995887 474237 995943
rect 474405 995887 474881 995943
rect 475049 995887 475433 995943
rect 475601 995887 476077 995943
rect 476245 995887 476721 995943
rect 476889 995887 477273 995943
rect 477441 995887 477917 995943
rect 478085 995887 478561 995943
rect 478729 995887 479113 995943
rect 479281 995887 479757 995943
rect 479925 995887 480401 995943
rect 480569 995887 481045 995943
rect 481213 995887 481597 995943
rect 481765 995887 482241 995943
rect 482409 995887 482885 995943
rect 483053 995887 483437 995943
rect 483605 995887 484081 995943
rect 484249 995887 484725 995943
rect 484893 995887 485277 995943
rect 485445 995887 485921 995943
rect 486089 995887 486565 995943
rect 486733 995887 487117 995943
rect 487285 995887 487761 995943
rect 487929 995887 488405 995943
rect 488573 995887 488783 995943
rect 524242 995943 540183 1037600
rect 575653 1002788 590458 1036615
rect 575653 998067 585622 1002788
rect 575699 997600 580479 998011
rect 580535 998007 585622 998067
rect 585678 997600 590458 1002732
rect 585704 996441 585732 997600
rect 585690 996432 585746 996441
rect 585690 996367 585746 996376
rect 524242 995887 524441 995943
rect 524609 995887 524993 995943
rect 525161 995887 525637 995943
rect 525805 995887 526281 995943
rect 526449 995887 526833 995943
rect 527001 995887 527477 995943
rect 527645 995887 528121 995943
rect 528289 995887 528673 995943
rect 528841 995887 529317 995943
rect 529485 995887 529961 995943
rect 530129 995887 530513 995943
rect 530681 995887 531157 995943
rect 531325 995887 531801 995943
rect 531969 995887 532445 995943
rect 532613 995887 532997 995943
rect 533165 995887 533641 995943
rect 533809 995887 534285 995943
rect 534453 995887 534837 995943
rect 535005 995887 535481 995943
rect 535649 995887 536125 995943
rect 536293 995887 536677 995943
rect 536845 995887 537321 995943
rect 537489 995887 537965 995943
rect 538133 995887 538517 995943
rect 538685 995887 539161 995943
rect 539329 995887 539805 995943
rect 539973 995887 540183 995943
rect 626042 995943 641983 1037600
rect 672630 996568 672686 996577
rect 672630 996503 672686 996512
rect 672446 996432 672502 996441
rect 672446 996367 672502 996376
rect 626042 995887 626241 995943
rect 626409 995887 626793 995943
rect 626961 995887 627437 995943
rect 627605 995887 628081 995943
rect 628249 995887 628633 995943
rect 628801 995887 629277 995943
rect 629445 995887 629921 995943
rect 630089 995887 630473 995943
rect 630641 995887 631117 995943
rect 631285 995887 631761 995943
rect 631929 995887 632313 995943
rect 632481 995887 632957 995943
rect 633125 995887 633601 995943
rect 633769 995887 634245 995943
rect 634413 995887 634797 995943
rect 634965 995887 635441 995943
rect 635609 995887 636085 995943
rect 636253 995887 636637 995943
rect 636805 995887 637281 995943
rect 637449 995887 637925 995943
rect 638093 995887 638477 995943
rect 638645 995887 639121 995943
rect 639289 995887 639765 995943
rect 639933 995887 640317 995943
rect 640485 995887 640961 995943
rect 641129 995887 641605 995943
rect 641773 995887 641983 995943
rect 384097 995407 384153 995887
rect 387133 995452 387189 995887
rect 387133 995407 387196 995452
rect 391457 995452 391513 995887
rect 391457 995407 391520 995452
rect 394493 995407 394549 995887
rect 395781 995407 395837 995887
rect 396333 995407 396389 995887
rect 397621 995452 397677 995887
rect 397621 995407 397684 995452
rect 398173 995407 398229 995887
rect 399461 995452 399517 995887
rect 399461 995407 399524 995452
rect 473097 995407 473153 995887
rect 476133 995452 476189 995887
rect 476132 995407 476189 995452
rect 480457 995452 480513 995887
rect 480456 995407 480513 995452
rect 483493 995407 483549 995887
rect 484781 995407 484837 995887
rect 485333 995407 485389 995887
rect 486621 995452 486677 995887
rect 486620 995407 486677 995452
rect 487173 995407 487229 995887
rect 488461 995452 488517 995887
rect 488460 995407 488517 995452
rect 524497 995407 524553 995887
rect 527533 995407 527589 995887
rect 531857 995466 531913 995887
rect 531964 995648 532016 995654
rect 531964 995590 532016 995596
rect 531976 995466 532004 995590
rect 531857 995438 532004 995466
rect 531857 995407 531913 995438
rect 534893 995407 534949 995887
rect 536181 995407 536237 995887
rect 536733 995407 536789 995887
rect 538021 995489 538077 995887
rect 537850 995480 537906 995489
rect 537850 995415 537906 995424
rect 538021 995480 538090 995489
rect 538021 995424 538034 995480
rect 538021 995415 538090 995424
rect 386328 990752 386380 990758
rect 386328 990694 386380 990700
rect 333520 990684 333572 990690
rect 333520 990626 333572 990632
rect 386340 990418 386368 990694
rect 387168 990690 387196 995407
rect 391492 995314 391520 995407
rect 391480 995308 391532 995314
rect 391480 995250 391532 995256
rect 391756 990820 391808 990826
rect 391756 990762 391808 990768
rect 391768 990690 391796 990762
rect 387156 990684 387208 990690
rect 387156 990626 387208 990632
rect 391756 990684 391808 990690
rect 391756 990626 391808 990632
rect 397656 990418 397684 995407
rect 399496 995314 399524 995407
rect 399484 995308 399536 995314
rect 399484 995250 399536 995256
rect 476132 990826 476160 995407
rect 480456 995314 480484 995407
rect 480444 995308 480496 995314
rect 480444 995250 480496 995256
rect 476120 990820 476172 990826
rect 476120 990762 476172 990768
rect 469312 990616 469364 990622
rect 469048 990564 469312 990570
rect 469048 990558 469364 990564
rect 469048 990554 469352 990558
rect 469036 990548 469352 990554
rect 469088 990542 469352 990548
rect 483020 990548 483072 990554
rect 469036 990490 469088 990496
rect 483020 990490 483072 990496
rect 483032 990418 483060 990490
rect 486620 990418 486648 995407
rect 488460 995314 488488 995407
rect 488448 995308 488500 995314
rect 488448 995250 488500 995256
rect 527560 990826 527588 995407
rect 527548 990820 527600 990826
rect 527548 990762 527600 990768
rect 386328 990412 386380 990418
rect 386328 990354 386380 990360
rect 397644 990412 397696 990418
rect 397644 990354 397696 990360
rect 424968 990412 425020 990418
rect 424968 990354 425020 990360
rect 483020 990412 483072 990418
rect 483020 990354 483072 990360
rect 486608 990412 486660 990418
rect 486608 990354 486660 990360
rect 521660 990412 521712 990418
rect 521660 990354 521712 990360
rect 397656 990282 397684 990354
rect 154580 990276 154632 990282
rect 154580 990218 154632 990224
rect 164148 990276 164200 990282
rect 164148 990218 164200 990224
rect 397644 990276 397696 990282
rect 397644 990218 397696 990224
rect 405740 990276 405792 990282
rect 405740 990218 405792 990224
rect 405752 990146 405780 990218
rect 424980 990146 425008 990354
rect 507768 990344 507820 990350
rect 507860 990344 507912 990350
rect 507820 990292 507860 990298
rect 507768 990286 507912 990292
rect 507780 990270 507900 990286
rect 521672 990282 521700 990354
rect 537864 990282 537892 995415
rect 538021 995407 538077 995415
rect 538573 995407 538629 995887
rect 539692 995648 539744 995654
rect 539692 995590 539744 995596
rect 539704 995466 539732 995590
rect 539861 995466 539917 995887
rect 539704 995438 539917 995466
rect 539861 995407 539917 995438
rect 626297 995407 626353 995887
rect 629333 995466 629389 995887
rect 629312 995407 629389 995466
rect 633657 995466 633713 995887
rect 633808 995512 633860 995518
rect 633657 995460 633808 995466
rect 633657 995454 633860 995460
rect 633657 995438 633848 995454
rect 633657 995407 633713 995438
rect 636693 995407 636749 995887
rect 637981 995407 638037 995887
rect 638533 995407 638589 995887
rect 639821 995466 639877 995887
rect 639800 995407 639877 995466
rect 640373 995407 640429 995887
rect 641536 995512 641588 995518
rect 641661 995466 641717 995887
rect 641588 995460 641717 995466
rect 641536 995454 641717 995460
rect 641548 995438 641717 995454
rect 641661 995407 641717 995438
rect 629312 990826 629340 995407
rect 629300 990820 629352 990826
rect 629300 990762 629352 990768
rect 596088 990684 596140 990690
rect 596088 990626 596140 990632
rect 576860 990616 576912 990622
rect 576858 990584 576860 990593
rect 596100 990593 596128 990626
rect 623688 990616 623740 990622
rect 576912 990584 576914 990593
rect 560208 990548 560260 990554
rect 576858 990519 576914 990528
rect 596086 990584 596142 990593
rect 623740 990564 623912 990570
rect 623688 990558 623912 990564
rect 623700 990554 623912 990558
rect 623700 990548 623924 990554
rect 623700 990542 623872 990548
rect 596086 990519 596142 990528
rect 560208 990490 560260 990496
rect 623872 990490 623924 990496
rect 540980 990480 541032 990486
rect 540978 990448 540980 990457
rect 560220 990457 560248 990490
rect 541032 990448 541034 990457
rect 540888 990412 540940 990418
rect 540978 990383 541034 990392
rect 560206 990448 560262 990457
rect 560206 990383 560262 990392
rect 540888 990354 540940 990360
rect 540900 990282 540928 990354
rect 521660 990276 521712 990282
rect 521660 990218 521712 990224
rect 537852 990276 537904 990282
rect 537852 990218 537904 990224
rect 540888 990276 540940 990282
rect 540888 990218 540940 990224
rect 629312 990146 629340 990762
rect 639800 990554 639828 995407
rect 639788 990548 639840 990554
rect 639788 990490 639840 990496
rect 639800 990214 639828 990490
rect 639788 990208 639840 990214
rect 639788 990150 639840 990156
rect 89996 990140 90048 990146
rect 89996 990082 90048 990088
rect 405740 990140 405792 990146
rect 405740 990082 405792 990088
rect 424968 990140 425020 990146
rect 424968 990082 425020 990088
rect 629300 990140 629352 990146
rect 629300 990082 629352 990088
rect 45848 879850 45968 879866
rect 45836 879844 45968 879850
rect 45888 879838 45968 879844
rect 45836 879786 45888 879792
rect 44454 835272 44510 835281
rect 44454 835207 44510 835216
rect 44468 493241 44496 835207
rect 672460 828730 672488 996367
rect 672538 828744 672594 828753
rect 672460 828702 672538 828730
rect 672538 828679 672594 828688
rect 44730 828064 44786 828073
rect 44730 827999 44786 828008
rect 44744 806002 44772 827999
rect 672644 826169 672672 996503
rect 673644 990208 673696 990214
rect 673644 990150 673696 990156
rect 673552 990140 673604 990146
rect 673552 990082 673604 990088
rect 673366 908168 673422 908177
rect 673366 908103 673422 908112
rect 672630 826160 672686 826169
rect 672630 826095 672686 826104
rect 673274 826160 673330 826169
rect 673274 826095 673330 826104
rect 673182 823712 673238 823721
rect 673182 823647 673238 823656
rect 44548 805996 44600 806002
rect 44548 805938 44600 805944
rect 44732 805996 44784 806002
rect 44732 805938 44784 805944
rect 44560 786570 44588 805938
rect 673196 792169 673224 823647
rect 672998 792160 673054 792169
rect 672998 792095 673054 792104
rect 673182 792160 673238 792169
rect 673182 792095 673238 792104
rect 44560 786542 44772 786570
rect 44744 778274 44772 786542
rect 673012 778394 673040 792095
rect 673000 778388 673052 778394
rect 673000 778330 673052 778336
rect 44652 778246 44772 778274
rect 673092 778252 673144 778258
rect 44652 759098 44680 778246
rect 673092 778194 673144 778200
rect 673104 772818 673132 778194
rect 672816 772812 672868 772818
rect 672816 772754 672868 772760
rect 673092 772812 673144 772818
rect 673092 772754 673144 772760
rect 44560 759070 44680 759098
rect 44560 701026 44588 759070
rect 672828 753545 672856 772754
rect 672814 753536 672870 753545
rect 672814 753471 672870 753480
rect 672998 753536 673054 753545
rect 672998 753471 673054 753480
rect 673012 739770 673040 753471
rect 673000 739764 673052 739770
rect 673000 739706 673052 739712
rect 673184 739628 673236 739634
rect 673184 739570 673236 739576
rect 673196 714762 673224 739570
rect 673104 714734 673224 714762
rect 44560 700998 44680 701026
rect 44652 695502 44680 700998
rect 673104 695570 673132 714734
rect 673092 695564 673144 695570
rect 673092 695506 673144 695512
rect 673184 695564 673236 695570
rect 673184 695506 673236 695512
rect 44640 695496 44692 695502
rect 44640 695438 44692 695444
rect 44916 695496 44968 695502
rect 44916 695438 44968 695444
rect 44928 676258 44956 695438
rect 44732 676252 44784 676258
rect 44732 676194 44784 676200
rect 44916 676252 44968 676258
rect 44916 676194 44968 676200
rect 44560 662454 44588 662485
rect 44744 662454 44772 676194
rect 673196 662522 673224 695506
rect 673184 662516 673236 662522
rect 673184 662458 673236 662464
rect 44548 662448 44600 662454
rect 44732 662448 44784 662454
rect 44600 662396 44680 662402
rect 44548 662390 44680 662396
rect 44732 662390 44784 662396
rect 44560 662374 44680 662390
rect 44652 656878 44680 662374
rect 673184 662380 673236 662386
rect 673184 662322 673236 662328
rect 44640 656872 44692 656878
rect 44640 656814 44692 656820
rect 44824 656872 44876 656878
rect 44824 656814 44876 656820
rect 44836 642818 44864 656814
rect 673196 643090 673224 662322
rect 44652 642790 44864 642818
rect 673104 643062 673224 643090
rect 44652 604586 44680 642790
rect 673104 637566 673132 643062
rect 672816 637560 672868 637566
rect 672816 637502 672868 637508
rect 673092 637560 673144 637566
rect 673092 637502 673144 637508
rect 672828 618322 672856 637502
rect 672816 618316 672868 618322
rect 672816 618258 672868 618264
rect 673000 618316 673052 618322
rect 673000 618258 673052 618264
rect 673012 618225 673040 618258
rect 672998 618216 673054 618225
rect 672998 618151 673054 618160
rect 672814 618080 672870 618089
rect 672814 618015 672870 618024
rect 44640 604580 44692 604586
rect 44640 604522 44692 604528
rect 44640 604444 44692 604450
rect 44640 604386 44692 604392
rect 44652 585154 44680 604386
rect 672828 599010 672856 618015
rect 672816 599004 672868 599010
rect 672816 598946 672868 598952
rect 673092 599004 673144 599010
rect 673092 598946 673144 598952
rect 673104 585206 673132 598946
rect 44560 585126 44680 585154
rect 673092 585200 673144 585206
rect 673092 585142 673144 585148
rect 673000 585132 673052 585138
rect 44560 560289 44588 585126
rect 673000 585074 673052 585080
rect 673012 569974 673040 585074
rect 672816 569968 672868 569974
rect 672816 569910 672868 569916
rect 673000 569968 673052 569974
rect 673000 569910 673052 569916
rect 672828 560318 672856 569910
rect 672816 560312 672868 560318
rect 44546 560280 44602 560289
rect 44546 560215 44602 560224
rect 44914 560280 44970 560289
rect 672816 560254 672868 560260
rect 673000 560312 673052 560318
rect 673000 560254 673052 560260
rect 44914 560215 44970 560224
rect 44928 541006 44956 560215
rect 673012 546582 673040 560254
rect 673000 546576 673052 546582
rect 673000 546518 673052 546524
rect 673092 546372 673144 546378
rect 673092 546314 673144 546320
rect 44732 541000 44784 541006
rect 44732 540942 44784 540948
rect 44916 541000 44968 541006
rect 44916 540942 44968 540948
rect 44744 496874 44772 540942
rect 673104 527202 673132 546314
rect 673092 527196 673144 527202
rect 673092 527138 673144 527144
rect 673184 527060 673236 527066
rect 673184 527002 673236 527008
rect 673196 521626 673224 527002
rect 673184 521620 673236 521626
rect 673184 521562 673236 521568
rect 673288 511465 673316 826095
rect 673090 511456 673146 511465
rect 673090 511391 673146 511400
rect 673274 511456 673330 511465
rect 673274 511391 673330 511400
rect 672998 509144 673054 509153
rect 672998 509079 673054 509088
rect 44548 496868 44600 496874
rect 44548 496810 44600 496816
rect 44732 496868 44784 496874
rect 44732 496810 44784 496816
rect 44454 493232 44510 493241
rect 44454 493167 44510 493176
rect 44560 488617 44588 496810
rect 44546 488608 44602 488617
rect 44546 488543 44602 488552
rect 673012 449954 673040 509079
rect 673000 449948 673052 449954
rect 673000 449890 673052 449896
rect 44362 448624 44418 448633
rect 44362 448559 44418 448568
rect 673104 427961 673132 511391
rect 673274 502344 673330 502353
rect 673274 502279 673330 502288
rect 673288 463729 673316 502279
rect 673380 483177 673408 908103
rect 673564 964782 673592 990082
rect 673552 964776 673604 964782
rect 673552 964718 673604 964724
rect 673564 910790 673592 964718
rect 673656 953358 673684 990150
rect 675887 967359 717600 967558
rect 675407 967247 675887 967303
rect 675943 967191 717600 967359
rect 675887 966807 717600 967191
rect 675943 966639 717600 966807
rect 675887 966163 717600 966639
rect 675943 965995 717600 966163
rect 675887 965519 717600 965995
rect 675943 965351 717600 965519
rect 675887 964967 717600 965351
rect 675943 964799 717600 964967
rect 675392 964776 675444 964782
rect 675392 964718 675444 964724
rect 675404 964267 675432 964718
rect 675887 964323 717600 964799
rect 675404 964239 675887 964267
rect 675407 964211 675887 964239
rect 675943 964155 717600 964323
rect 675887 963679 717600 964155
rect 675943 963511 717600 963679
rect 675887 963127 717600 963511
rect 675943 962959 717600 963127
rect 675887 962483 717600 962959
rect 675943 962315 717600 962483
rect 675887 961839 717600 962315
rect 675943 961671 717600 961839
rect 675887 961287 717600 961671
rect 675943 961119 717600 961287
rect 675887 960643 717600 961119
rect 675943 960475 717600 960643
rect 675887 959999 717600 960475
rect 675407 959929 675887 959943
rect 675312 959901 675887 959929
rect 673644 953352 673696 953358
rect 673644 953294 673696 953300
rect 673552 910784 673604 910790
rect 673552 910726 673604 910732
rect 673564 875566 673592 910726
rect 673552 875560 673604 875566
rect 673552 875502 673604 875508
rect 673656 875090 673684 953294
rect 675312 951810 675340 959901
rect 675407 959887 675887 959901
rect 675943 959831 717600 959999
rect 675887 959355 717600 959831
rect 675943 959187 717600 959355
rect 675887 958803 717600 959187
rect 675943 958635 717600 958803
rect 675887 958159 717600 958635
rect 675943 957991 717600 958159
rect 675887 957515 717600 957991
rect 675943 957347 717600 957515
rect 675887 956963 717600 957347
rect 675407 956851 675887 956907
rect 675943 956795 717600 956963
rect 675887 956319 717600 956795
rect 675943 956151 717600 956319
rect 675887 955675 717600 956151
rect 675407 955563 675887 955619
rect 675943 955507 717600 955675
rect 675887 955123 717600 955507
rect 675407 955011 675887 955067
rect 675943 954955 717600 955123
rect 675887 954479 717600 954955
rect 675943 954311 717600 954479
rect 675887 953835 717600 954311
rect 675407 953751 675887 953779
rect 675404 953723 675887 953751
rect 675404 953358 675432 953723
rect 675943 953667 717600 953835
rect 675392 953352 675444 953358
rect 675392 953294 675444 953300
rect 675887 953283 717600 953667
rect 675407 953171 675887 953227
rect 675943 953115 717600 953283
rect 675887 952639 717600 953115
rect 675943 952471 717600 952639
rect 675887 951995 717600 952471
rect 675407 951932 675887 951939
rect 675404 951883 675887 951932
rect 675404 951810 675432 951883
rect 675943 951827 717600 951995
rect 675312 951782 675432 951810
rect 675887 951617 717600 951827
rect 677874 918640 677930 918649
rect 678000 918626 678297 922500
rect 677930 918598 678297 918626
rect 677874 918575 677930 918584
rect 678000 918501 678297 918598
rect 678353 918445 716886 922502
rect 678007 915768 716886 918445
rect 677598 915376 677654 915385
rect 677598 915311 677654 915320
rect 677612 912801 677640 915311
rect 678000 914002 678065 915712
rect 677796 913974 678065 914002
rect 677598 912792 677654 912801
rect 677598 912727 677654 912736
rect 677796 910790 677824 913974
rect 678000 913712 678065 913974
rect 678121 913656 716886 915768
rect 677874 912792 677930 912801
rect 677874 912727 677930 912736
rect 677784 910784 677836 910790
rect 677784 910726 677836 910732
rect 677888 908177 677916 912727
rect 678007 911713 716886 913656
rect 677874 908168 677930 908177
rect 677874 908103 677930 908112
rect 677782 907760 677838 907769
rect 678000 907746 678732 911657
rect 677838 907718 678732 907746
rect 677782 907695 677838 907704
rect 678000 907660 678732 907718
rect 678788 907660 716886 911713
rect 675887 878159 717600 878358
rect 675407 878047 675887 878103
rect 675943 877991 717600 878159
rect 675887 877607 717600 877991
rect 675943 877439 717600 877607
rect 675887 876963 717600 877439
rect 675943 876795 717600 876963
rect 675887 876319 717600 876795
rect 675943 876151 717600 876319
rect 675887 875767 717600 876151
rect 673644 875084 673696 875090
rect 673644 875026 673696 875032
rect 673644 874948 673696 874954
rect 673644 874890 673696 874896
rect 673656 865026 673684 874890
rect 675943 875599 717600 875767
rect 675392 875560 675444 875566
rect 675392 875502 675444 875508
rect 675404 875067 675432 875502
rect 675887 875123 717600 875599
rect 675404 875039 675887 875067
rect 675407 875011 675887 875039
rect 675943 874955 717600 875123
rect 675887 874479 717600 874955
rect 675943 874311 717600 874479
rect 675887 873927 717600 874311
rect 675943 873759 717600 873927
rect 675887 873283 717600 873759
rect 675943 873115 717600 873283
rect 675887 872639 717600 873115
rect 675943 872471 717600 872639
rect 675887 872087 717600 872471
rect 675943 871919 717600 872087
rect 675887 871443 717600 871919
rect 675943 871275 717600 871443
rect 675887 870799 717600 871275
rect 675407 870740 675887 870743
rect 675404 870687 675887 870740
rect 675404 870210 675432 870687
rect 675943 870631 717600 870799
rect 675312 870182 675432 870210
rect 673644 865020 673696 865026
rect 673644 864962 673696 864968
rect 673828 865020 673880 865026
rect 673828 864962 673880 864968
rect 673644 785324 673696 785330
rect 673644 785266 673696 785272
rect 673460 774920 673512 774926
rect 673460 774862 673512 774868
rect 673472 730182 673500 774862
rect 673656 741402 673684 785266
rect 673840 774926 673868 864962
rect 675312 862730 675340 870182
rect 675887 870155 717600 870631
rect 675943 869987 717600 870155
rect 675887 869603 717600 869987
rect 675943 869435 717600 869603
rect 675887 868959 717600 869435
rect 675943 868791 717600 868959
rect 675887 868315 717600 868791
rect 675943 868147 717600 868315
rect 675887 867763 717600 868147
rect 675407 867651 675887 867707
rect 675943 867595 717600 867763
rect 675887 867119 717600 867595
rect 675943 866951 717600 867119
rect 675887 866475 717600 866951
rect 675407 866363 675887 866419
rect 675943 866307 717600 866475
rect 675887 865923 717600 866307
rect 675407 865811 675887 865867
rect 675943 865755 717600 865923
rect 675887 865279 717600 865755
rect 675943 865111 717600 865279
rect 675392 865020 675444 865026
rect 675392 864962 675444 864968
rect 675404 864579 675432 864962
rect 675887 864635 717600 865111
rect 675404 864551 675887 864579
rect 675407 864523 675887 864551
rect 675943 864467 717600 864635
rect 675887 864083 717600 864467
rect 675407 863971 675887 864027
rect 675943 863915 717600 864083
rect 675887 863439 717600 863915
rect 675943 863271 717600 863439
rect 675887 862795 717600 863271
rect 675407 862730 675887 862739
rect 675312 862702 675887 862730
rect 675407 862683 675887 862702
rect 675943 862627 717600 862795
rect 675887 862417 717600 862627
rect 676126 828744 676182 828753
rect 676126 828679 676182 828688
rect 676140 823721 676168 828679
rect 677600 828521 678011 833301
rect 678067 828465 716615 833347
rect 676126 823712 676182 823721
rect 676126 823647 676182 823656
rect 678007 823378 716615 828465
rect 677600 818542 682732 823322
rect 682788 818542 716615 823378
rect 675887 788959 717600 789158
rect 675407 788847 675887 788903
rect 675943 788791 717600 788959
rect 675887 788407 717600 788791
rect 675943 788239 717600 788407
rect 675887 787763 717600 788239
rect 675943 787595 717600 787763
rect 675887 787119 717600 787595
rect 675943 786951 717600 787119
rect 675887 786567 717600 786951
rect 673828 774920 673880 774926
rect 673828 774862 673880 774868
rect 675943 786399 717600 786567
rect 675887 785923 717600 786399
rect 675407 785839 675887 785867
rect 675404 785811 675887 785839
rect 675404 785330 675432 785811
rect 675943 785755 717600 785923
rect 675392 785324 675444 785330
rect 675887 785279 717600 785755
rect 675392 785266 675444 785272
rect 675943 785111 717600 785279
rect 675887 784727 717600 785111
rect 675943 784559 717600 784727
rect 675887 784083 717600 784559
rect 675943 783915 717600 784083
rect 675887 783439 717600 783915
rect 675943 783271 717600 783439
rect 675887 782887 717600 783271
rect 675943 782719 717600 782887
rect 675887 782243 717600 782719
rect 675943 782075 717600 782243
rect 675887 781599 717600 782075
rect 675407 781538 675887 781543
rect 675312 781510 675887 781538
rect 675312 773514 675340 781510
rect 675407 781487 675887 781510
rect 675943 781431 717600 781599
rect 675887 780955 717600 781431
rect 675943 780787 717600 780955
rect 675887 780403 717600 780787
rect 675943 780235 717600 780403
rect 675887 779759 717600 780235
rect 675943 779591 717600 779759
rect 675887 779115 717600 779591
rect 675943 778947 717600 779115
rect 675887 778563 717600 778947
rect 675407 778451 675887 778507
rect 675943 778395 717600 778563
rect 675887 777919 717600 778395
rect 675943 777751 717600 777919
rect 675887 777275 717600 777751
rect 675407 777163 675887 777219
rect 675943 777107 717600 777275
rect 675887 776723 717600 777107
rect 675407 776611 675887 776667
rect 675943 776555 717600 776723
rect 675887 776079 717600 776555
rect 675943 775911 717600 776079
rect 675887 775435 717600 775911
rect 675407 775351 675887 775379
rect 675404 775323 675887 775351
rect 675404 774926 675432 775323
rect 675943 775267 717600 775435
rect 675392 774920 675444 774926
rect 675887 774883 717600 775267
rect 675392 774862 675444 774868
rect 675407 774771 675887 774827
rect 675943 774715 717600 774883
rect 675887 774239 717600 774715
rect 675943 774071 717600 774239
rect 675887 773595 717600 774071
rect 675407 773514 675887 773539
rect 675312 773486 675887 773514
rect 675407 773483 675887 773486
rect 675943 773427 717600 773595
rect 675887 773217 717600 773427
rect 675887 743959 717600 744158
rect 675407 743847 675887 743903
rect 675943 743791 717600 743959
rect 675887 743407 717600 743791
rect 675943 743239 717600 743407
rect 675887 742763 717600 743239
rect 675943 742595 717600 742763
rect 675887 742119 717600 742595
rect 675943 741951 717600 742119
rect 673644 741396 673696 741402
rect 673644 741338 673696 741344
rect 673460 730176 673512 730182
rect 673460 730118 673512 730124
rect 673472 685409 673500 730118
rect 673828 730040 673880 730046
rect 673828 729982 673880 729988
rect 673552 695360 673604 695366
rect 673552 695302 673604 695308
rect 673458 685400 673514 685409
rect 673458 685335 673514 685344
rect 673472 639742 673500 685335
rect 673564 651166 673592 695302
rect 673840 695366 673868 729982
rect 675887 741567 717600 741951
rect 675392 741396 675444 741402
rect 675943 741399 717600 741567
rect 675392 741338 675444 741344
rect 675404 740874 675432 741338
rect 675887 740923 717600 741399
rect 675128 740867 675432 740874
rect 675128 740846 675887 740867
rect 675128 730046 675156 740846
rect 675407 740811 675887 740846
rect 675943 740755 717600 740923
rect 675887 740279 717600 740755
rect 675943 740111 717600 740279
rect 675887 739727 717600 740111
rect 675943 739559 717600 739727
rect 675887 739083 717600 739559
rect 675943 738915 717600 739083
rect 675887 738439 717600 738915
rect 675943 738271 717600 738439
rect 675887 737887 717600 738271
rect 675943 737719 717600 737887
rect 675887 737243 717600 737719
rect 675943 737075 717600 737243
rect 675887 736599 717600 737075
rect 675407 736522 675887 736543
rect 675312 736494 675887 736522
rect 675116 730040 675168 730046
rect 675116 729982 675168 729988
rect 675312 729042 675340 736494
rect 675407 736487 675887 736494
rect 675943 736431 717600 736599
rect 675887 735955 717600 736431
rect 675943 735787 717600 735955
rect 675887 735403 717600 735787
rect 675943 735235 717600 735403
rect 675887 734759 717600 735235
rect 675943 734591 717600 734759
rect 675887 734115 717600 734591
rect 675943 733947 717600 734115
rect 675887 733563 717600 733947
rect 675407 733451 675887 733507
rect 675943 733395 717600 733563
rect 675887 732919 717600 733395
rect 675943 732751 717600 732919
rect 675887 732275 717600 732751
rect 675407 732163 675887 732219
rect 675943 732107 717600 732275
rect 675887 731723 717600 732107
rect 675407 731611 675887 731667
rect 675943 731555 717600 731723
rect 675887 731079 717600 731555
rect 675943 730911 717600 731079
rect 675887 730435 717600 730911
rect 675407 730351 675887 730379
rect 675404 730323 675887 730351
rect 675404 730182 675432 730323
rect 675943 730267 717600 730435
rect 675392 730176 675444 730182
rect 675392 730118 675444 730124
rect 675887 729883 717600 730267
rect 675407 729771 675887 729827
rect 675943 729715 717600 729883
rect 675887 729239 717600 729715
rect 675943 729071 717600 729239
rect 675312 729014 675432 729042
rect 675404 728539 675432 729014
rect 675887 728595 717600 729071
rect 675404 728484 675887 728539
rect 675407 728483 675887 728484
rect 675943 728427 717600 728595
rect 675887 728217 717600 728427
rect 675887 698959 717600 699158
rect 675407 698847 675887 698903
rect 675943 698791 717600 698959
rect 675887 698407 717600 698791
rect 675943 698239 717600 698407
rect 675887 697763 717600 698239
rect 675943 697595 717600 697763
rect 675887 697119 717600 697595
rect 675943 696951 717600 697119
rect 675887 696567 717600 696951
rect 675943 696399 717600 696567
rect 675887 695923 717600 696399
rect 675407 695844 675887 695867
rect 675404 695811 675887 695844
rect 675404 695366 675432 695811
rect 675943 695755 717600 695923
rect 673828 695360 673880 695366
rect 673828 695302 673880 695308
rect 675392 695360 675444 695366
rect 675392 695302 675444 695308
rect 675887 695279 717600 695755
rect 675943 695111 717600 695279
rect 675887 694727 717600 695111
rect 675943 694559 717600 694727
rect 675887 694083 717600 694559
rect 675943 693915 717600 694083
rect 675887 693439 717600 693915
rect 675943 693271 717600 693439
rect 675887 692887 717600 693271
rect 675943 692719 717600 692887
rect 675887 692243 717600 692719
rect 675943 692075 717600 692243
rect 675312 691614 675432 691642
rect 675312 683525 675340 691614
rect 675404 691543 675432 691614
rect 675887 691599 717600 692075
rect 675404 691492 675887 691543
rect 675407 691487 675887 691492
rect 675943 691431 717600 691599
rect 675887 690955 717600 691431
rect 675943 690787 717600 690955
rect 675887 690403 717600 690787
rect 675943 690235 717600 690403
rect 675887 689759 717600 690235
rect 675943 689591 717600 689759
rect 675887 689115 717600 689591
rect 675943 688947 717600 689115
rect 675887 688563 717600 688947
rect 675407 688451 675887 688507
rect 675943 688395 717600 688563
rect 675887 687919 717600 688395
rect 675943 687751 717600 687919
rect 675887 687275 717600 687751
rect 675407 687163 675887 687219
rect 675943 687107 717600 687275
rect 675887 686723 717600 687107
rect 675407 686611 675887 686667
rect 675943 686555 717600 686723
rect 675887 686079 717600 686555
rect 675943 685911 717600 686079
rect 675887 685435 717600 685911
rect 675390 685400 675446 685409
rect 675446 685344 675887 685379
rect 675390 685335 675887 685344
rect 675407 685323 675887 685335
rect 675943 685267 717600 685435
rect 675887 684883 717600 685267
rect 675407 684771 675887 684827
rect 675943 684715 717600 684883
rect 675887 684239 717600 684715
rect 675943 684071 717600 684239
rect 675887 683595 717600 684071
rect 675407 683525 675887 683539
rect 675312 683497 675887 683525
rect 675407 683483 675887 683497
rect 675943 683427 717600 683595
rect 675887 683217 717600 683427
rect 675887 653759 717600 653958
rect 675407 653647 675887 653703
rect 675943 653591 717600 653759
rect 675887 653207 717600 653591
rect 675943 653039 717600 653207
rect 675887 652563 717600 653039
rect 675943 652395 717600 652563
rect 675887 651919 717600 652395
rect 675943 651751 717600 651919
rect 673552 651160 673604 651166
rect 673552 651102 673604 651108
rect 673460 639736 673512 639742
rect 673460 639678 673512 639684
rect 673472 594930 673500 639678
rect 673564 605674 673592 651102
rect 675887 651367 717600 651751
rect 675943 651199 717600 651367
rect 675392 651160 675444 651166
rect 675392 651102 675444 651108
rect 675404 650667 675432 651102
rect 675887 650723 717600 651199
rect 675404 650639 675887 650667
rect 675407 650611 675887 650639
rect 675943 650555 717600 650723
rect 675887 650079 717600 650555
rect 675943 649911 717600 650079
rect 675887 649527 717600 649911
rect 675943 649359 717600 649527
rect 675887 648883 717600 649359
rect 675943 648715 717600 648883
rect 675887 648239 717600 648715
rect 675943 648071 717600 648239
rect 675887 647687 717600 648071
rect 675943 647519 717600 647687
rect 675887 647043 717600 647519
rect 675943 646875 717600 647043
rect 675887 646399 717600 646875
rect 675407 646340 675887 646343
rect 675404 646287 675887 646340
rect 675404 645810 675432 646287
rect 675943 646231 717600 646399
rect 675312 645782 675432 645810
rect 675312 638330 675340 645782
rect 675887 645755 717600 646231
rect 675943 645587 717600 645755
rect 675887 645203 717600 645587
rect 675943 645035 717600 645203
rect 675887 644559 717600 645035
rect 675943 644391 717600 644559
rect 675887 643915 717600 644391
rect 675943 643747 717600 643915
rect 675887 643363 717600 643747
rect 675407 643251 675887 643307
rect 675943 643195 717600 643363
rect 675887 642719 717600 643195
rect 675943 642551 717600 642719
rect 675887 642075 717600 642551
rect 675407 641963 675887 642019
rect 675943 641907 717600 642075
rect 675887 641523 717600 641907
rect 675407 641411 675887 641467
rect 675943 641355 717600 641523
rect 675887 640879 717600 641355
rect 675943 640711 717600 640879
rect 675887 640235 717600 640711
rect 675407 640151 675887 640179
rect 675404 640123 675887 640151
rect 675404 639742 675432 640123
rect 675943 640067 717600 640235
rect 675392 639736 675444 639742
rect 675392 639678 675444 639684
rect 675887 639683 717600 640067
rect 675407 639571 675887 639627
rect 675943 639515 717600 639683
rect 675887 639039 717600 639515
rect 675943 638871 717600 639039
rect 675887 638395 717600 638871
rect 675407 638330 675887 638339
rect 675312 638302 675887 638330
rect 675407 638283 675887 638302
rect 675943 638227 717600 638395
rect 675887 638017 717600 638227
rect 675887 608759 717600 608958
rect 675407 608647 675887 608703
rect 675943 608591 717600 608759
rect 675887 608207 717600 608591
rect 675943 608039 717600 608207
rect 675887 607563 717600 608039
rect 675943 607395 717600 607563
rect 675887 606919 717600 607395
rect 675943 606751 717600 606919
rect 673552 605668 673604 605674
rect 673552 605610 673604 605616
rect 673564 604450 673592 605610
rect 673552 604444 673604 604450
rect 673552 604386 673604 604392
rect 673460 594924 673512 594930
rect 673460 594866 673512 594872
rect 673472 550526 673500 594866
rect 673552 565888 673604 565894
rect 673552 565830 673604 565836
rect 673564 559978 673592 565830
rect 675887 606367 717600 606751
rect 675943 606199 717600 606367
rect 675887 605723 717600 606199
rect 675300 605668 675352 605674
rect 675407 605653 675887 605667
rect 675352 605625 675887 605653
rect 675300 605610 675352 605616
rect 675407 605611 675887 605625
rect 675943 605555 717600 605723
rect 675887 605079 717600 605555
rect 675943 604911 717600 605079
rect 675887 604527 717600 604911
rect 673828 604444 673880 604450
rect 673828 604386 673880 604392
rect 673840 585154 673868 604386
rect 675943 604359 717600 604527
rect 675887 603883 717600 604359
rect 675943 603715 717600 603883
rect 675887 603239 717600 603715
rect 675943 603071 717600 603239
rect 675887 602687 717600 603071
rect 675943 602519 717600 602687
rect 675887 602043 717600 602519
rect 675943 601875 717600 602043
rect 675887 601399 717600 601875
rect 675407 601338 675887 601343
rect 675312 601310 675887 601338
rect 675312 593314 675340 601310
rect 675407 601287 675887 601310
rect 675943 601231 717600 601399
rect 675887 600755 717600 601231
rect 675943 600587 717600 600755
rect 675887 600203 717600 600587
rect 675943 600035 717600 600203
rect 675887 599559 717600 600035
rect 675943 599391 717600 599559
rect 675887 598915 717600 599391
rect 675943 598747 717600 598915
rect 675887 598363 717600 598747
rect 675407 598251 675887 598307
rect 675943 598195 717600 598363
rect 675887 597719 717600 598195
rect 675943 597551 717600 597719
rect 675887 597075 717600 597551
rect 675407 596963 675887 597019
rect 675943 596907 717600 597075
rect 675887 596523 717600 596907
rect 675407 596411 675887 596467
rect 675943 596355 717600 596523
rect 675887 595879 717600 596355
rect 675943 595711 717600 595879
rect 675887 595235 717600 595711
rect 675407 595151 675887 595179
rect 675404 595123 675887 595151
rect 675404 594930 675432 595123
rect 675943 595067 717600 595235
rect 675392 594924 675444 594930
rect 675392 594866 675444 594872
rect 675887 594683 717600 595067
rect 675407 594571 675887 594627
rect 675943 594515 717600 594683
rect 675887 594039 717600 594515
rect 675943 593871 717600 594039
rect 675887 593395 717600 593871
rect 675407 593314 675887 593339
rect 675312 593286 675887 593314
rect 675407 593283 675887 593286
rect 675943 593227 717600 593395
rect 675887 593017 717600 593227
rect 673840 585126 673960 585154
rect 673932 565894 673960 585126
rect 673920 565888 673972 565894
rect 673920 565830 673972 565836
rect 675887 563559 717600 563758
rect 675407 563447 675887 563503
rect 675943 563391 717600 563559
rect 675887 563007 717600 563391
rect 675943 562839 717600 563007
rect 675887 562363 717600 562839
rect 675943 562195 717600 562363
rect 675887 561719 717600 562195
rect 675943 561551 717600 561719
rect 675887 561167 717600 561551
rect 675943 560999 717600 561167
rect 675887 560523 717600 560999
rect 675407 560439 675887 560467
rect 675404 560411 675887 560439
rect 675404 559978 675432 560411
rect 675943 560355 717600 560523
rect 673552 559972 673604 559978
rect 673552 559914 673604 559920
rect 673920 559972 673972 559978
rect 673920 559914 673972 559920
rect 675392 559972 675444 559978
rect 675392 559914 675444 559920
rect 673460 550520 673512 550526
rect 673460 550462 673512 550468
rect 673932 522986 673960 559914
rect 675887 559879 717600 560355
rect 675943 559711 717600 559879
rect 675887 559327 717600 559711
rect 675943 559159 717600 559327
rect 675887 558683 717600 559159
rect 675943 558515 717600 558683
rect 675887 558039 717600 558515
rect 675943 557871 717600 558039
rect 675887 557487 717600 557871
rect 675943 557319 717600 557487
rect 675887 556843 717600 557319
rect 675943 556675 717600 556843
rect 675887 556199 717600 556675
rect 675407 556129 675887 556143
rect 675312 556101 675887 556129
rect 675312 548125 675340 556101
rect 675407 556087 675887 556101
rect 675943 556031 717600 556199
rect 675887 555555 717600 556031
rect 675943 555387 717600 555555
rect 675887 555003 717600 555387
rect 675943 554835 717600 555003
rect 675887 554359 717600 554835
rect 675943 554191 717600 554359
rect 675887 553715 717600 554191
rect 675943 553547 717600 553715
rect 675887 553163 717600 553547
rect 675407 553051 675887 553107
rect 675943 552995 717600 553163
rect 675887 552519 717600 552995
rect 675943 552351 717600 552519
rect 675887 551875 717600 552351
rect 675407 551763 675887 551819
rect 675943 551707 717600 551875
rect 675887 551323 717600 551707
rect 675407 551211 675887 551267
rect 675943 551155 717600 551323
rect 675887 550679 717600 551155
rect 675392 550520 675444 550526
rect 675943 550511 717600 550679
rect 675392 550462 675444 550468
rect 675404 549979 675432 550462
rect 675887 550035 717600 550511
rect 675404 549951 675887 549979
rect 675407 549923 675887 549951
rect 675943 549867 717600 550035
rect 675887 549483 717600 549867
rect 675407 549371 675887 549427
rect 675943 549315 717600 549483
rect 675887 548839 717600 549315
rect 675943 548671 717600 548839
rect 675887 548195 717600 548671
rect 675407 548125 675887 548139
rect 675312 548097 675887 548125
rect 675407 548083 675887 548097
rect 675943 548027 717600 548195
rect 675887 547817 717600 548027
rect 673736 522980 673788 522986
rect 673736 522922 673788 522928
rect 673920 522980 673972 522986
rect 673920 522922 673972 522928
rect 673748 511850 673776 522922
rect 676128 521620 676180 521626
rect 676128 521562 676180 521568
rect 676140 514185 676168 521562
rect 676126 514176 676182 514185
rect 676126 514111 676182 514120
rect 673656 511822 673776 511850
rect 673656 502353 673684 511822
rect 676140 509153 676168 514111
rect 677600 513921 678011 518701
rect 678067 513865 716615 518747
rect 676126 509144 676182 509153
rect 676126 509079 676182 509088
rect 678007 508778 716615 513865
rect 677600 503942 682732 508722
rect 682788 503942 716615 508778
rect 673642 502344 673698 502353
rect 673642 502279 673698 502288
rect 673366 483168 673422 483177
rect 673366 483103 673422 483112
rect 673366 483032 673422 483041
rect 673366 482967 673422 482976
rect 673380 467537 673408 482967
rect 678058 477592 678114 477601
rect 678058 477527 678114 477536
rect 678072 474700 678100 477527
rect 678000 470778 678297 474700
rect 677888 470750 678297 470778
rect 677888 469985 677916 470750
rect 678000 470701 678297 470750
rect 678353 470645 716886 474700
rect 677874 469976 677930 469985
rect 677874 469911 677930 469920
rect 678007 467968 716886 470645
rect 673366 467528 673422 467537
rect 673366 467463 673422 467472
rect 678000 466018 678065 467912
rect 677704 465990 678065 466018
rect 673274 463720 673330 463729
rect 673274 463655 673330 463664
rect 673458 463720 673514 463729
rect 677704 463690 677732 465990
rect 678000 465912 678065 465990
rect 678121 465856 716886 467968
rect 678007 463913 716886 465856
rect 673458 463655 673514 463664
rect 673736 463684 673788 463690
rect 673472 463593 673500 463655
rect 673736 463626 673788 463632
rect 677692 463684 677744 463690
rect 677692 463626 677744 463632
rect 673748 463593 673776 463626
rect 673458 463584 673514 463593
rect 673458 463519 673514 463528
rect 673734 463584 673790 463593
rect 673734 463519 673790 463528
rect 673368 449948 673420 449954
rect 673368 449890 673420 449896
rect 673090 427952 673146 427961
rect 673090 427887 673146 427896
rect 673380 420889 673408 449890
rect 673748 444417 673776 463519
rect 678000 459898 678732 463857
rect 677704 459870 678732 459898
rect 673550 444408 673606 444417
rect 673550 444343 673606 444352
rect 673734 444408 673790 444417
rect 673734 444343 673790 444352
rect 673564 430658 673592 444343
rect 677704 440230 677732 459870
rect 678000 459860 678732 459870
rect 678788 459860 716886 463913
rect 676220 440224 676272 440230
rect 676220 440166 676272 440172
rect 677692 440224 677744 440230
rect 677692 440166 677744 440172
rect 673564 430630 673684 430658
rect 673656 430522 673684 430630
rect 673564 430494 673684 430522
rect 673366 420880 673422 420889
rect 673366 420815 673422 420824
rect 672816 412548 672868 412554
rect 672816 412490 672868 412496
rect 672828 411210 672856 412490
rect 673564 411346 673592 430494
rect 676232 412554 676260 440166
rect 677414 427952 677470 427961
rect 677414 427887 677470 427896
rect 677428 425762 677456 427887
rect 677600 425785 678011 430501
rect 677598 425776 678011 425785
rect 677428 425734 677598 425762
rect 677654 425721 678011 425776
rect 677598 425711 677654 425720
rect 678067 425665 716615 430547
rect 678007 420578 716615 425665
rect 677600 415742 682732 420522
rect 682788 415742 716615 420578
rect 676220 412548 676272 412554
rect 676220 412490 676272 412496
rect 672736 411182 672856 411210
rect 673472 411318 673592 411346
rect 672736 405686 672764 411182
rect 672540 405680 672592 405686
rect 672540 405622 672592 405628
rect 672724 405680 672776 405686
rect 672724 405622 672776 405628
rect 672552 386442 672580 405622
rect 673472 401606 673500 411318
rect 673460 401600 673512 401606
rect 673460 401542 673512 401548
rect 675300 401600 675352 401606
rect 675300 401542 675352 401548
rect 672540 386436 672592 386442
rect 672540 386378 672592 386384
rect 672816 386436 672868 386442
rect 672816 386378 672868 386384
rect 672828 372586 672856 386378
rect 672644 372558 672856 372586
rect 672644 353394 672672 372558
rect 672632 353388 672684 353394
rect 672632 353330 672684 353336
rect 672540 353252 672592 353258
rect 672540 353194 672592 353200
rect 672552 347750 672580 353194
rect 672540 347744 672592 347750
rect 672540 347686 672592 347692
rect 672724 347744 672776 347750
rect 672724 347686 672776 347692
rect 672736 328506 672764 347686
rect 675312 383253 675340 401542
rect 675887 386359 717600 386558
rect 675407 386247 675887 386303
rect 675943 386191 717600 386359
rect 675887 385807 717600 386191
rect 675943 385639 717600 385807
rect 675887 385163 717600 385639
rect 675943 384995 717600 385163
rect 675887 384519 717600 384995
rect 675943 384351 717600 384519
rect 675887 383967 717600 384351
rect 675943 383799 717600 383967
rect 675887 383323 717600 383799
rect 675407 383253 675887 383267
rect 675312 383225 675887 383253
rect 675404 383211 675887 383225
rect 675404 382770 675432 383211
rect 675943 383155 717600 383323
rect 673644 382764 673696 382770
rect 673644 382706 673696 382712
rect 675392 382764 675444 382770
rect 675392 382706 675444 382712
rect 672448 328500 672500 328506
rect 672448 328442 672500 328448
rect 672724 328500 672776 328506
rect 672724 328442 672776 328448
rect 672460 314786 672488 328442
rect 672538 314800 672594 314809
rect 672460 314758 672538 314786
rect 672538 314735 672594 314744
rect 672538 314528 672594 314537
rect 672538 314463 672594 314472
rect 672552 309126 672580 314463
rect 672540 309120 672592 309126
rect 672540 309062 672592 309068
rect 672816 309120 672868 309126
rect 672816 309062 672868 309068
rect 672828 289882 672856 309062
rect 673460 304972 673512 304978
rect 673460 304914 673512 304920
rect 672632 289876 672684 289882
rect 672632 289818 672684 289824
rect 672816 289876 672868 289882
rect 672816 289818 672868 289824
rect 672644 276060 672672 289818
rect 673472 283082 673500 304914
rect 673656 338570 673684 382706
rect 675887 382679 717600 383155
rect 675943 382511 717600 382679
rect 675887 382127 717600 382511
rect 675943 381959 717600 382127
rect 675887 381483 717600 381959
rect 675943 381315 717600 381483
rect 675887 380839 717600 381315
rect 675943 380671 717600 380839
rect 675887 380287 717600 380671
rect 675943 380119 717600 380287
rect 675887 379643 717600 380119
rect 675943 379475 717600 379643
rect 675887 378999 717600 379475
rect 675407 378929 675887 378943
rect 675312 378901 675887 378929
rect 673828 372360 673880 372366
rect 673828 372302 673880 372308
rect 673644 338564 673696 338570
rect 673644 338506 673696 338512
rect 673656 293554 673684 338506
rect 673840 327146 673868 372302
rect 675312 370925 675340 378901
rect 675407 378887 675887 378901
rect 675943 378831 717600 378999
rect 675887 378355 717600 378831
rect 675943 378187 717600 378355
rect 675887 377803 717600 378187
rect 675943 377635 717600 377803
rect 675887 377159 717600 377635
rect 675943 376991 717600 377159
rect 675887 376515 717600 376991
rect 675943 376347 717600 376515
rect 675887 375963 717600 376347
rect 675407 375851 675887 375907
rect 675943 375795 717600 375963
rect 675887 375319 717600 375795
rect 675943 375151 717600 375319
rect 675887 374675 717600 375151
rect 675407 374563 675887 374619
rect 675943 374507 717600 374675
rect 675887 374123 717600 374507
rect 675407 374011 675887 374067
rect 675943 373955 717600 374123
rect 675887 373479 717600 373955
rect 675943 373311 717600 373479
rect 675887 372835 717600 373311
rect 675407 372751 675887 372779
rect 675404 372723 675887 372751
rect 675404 372366 675432 372723
rect 675943 372667 717600 372835
rect 675392 372360 675444 372366
rect 675392 372302 675444 372308
rect 675887 372283 717600 372667
rect 675407 372171 675887 372227
rect 675943 372115 717600 372283
rect 675887 371639 717600 372115
rect 675943 371471 717600 371639
rect 675887 370995 717600 371471
rect 675407 370925 675887 370939
rect 675312 370897 675887 370925
rect 675407 370883 675887 370897
rect 675943 370827 717600 370995
rect 675887 370617 717600 370827
rect 675887 341159 717600 341358
rect 675407 341047 675887 341103
rect 675943 340991 717600 341159
rect 675887 340607 717600 340991
rect 675943 340439 717600 340607
rect 675887 339963 717600 340439
rect 675943 339795 717600 339963
rect 675887 339319 717600 339795
rect 675943 339151 717600 339319
rect 675887 338767 717600 339151
rect 675943 338599 717600 338767
rect 675392 338564 675444 338570
rect 675392 338506 675444 338512
rect 675404 338067 675432 338506
rect 675887 338123 717600 338599
rect 675404 338028 675887 338067
rect 675407 338011 675887 338028
rect 675943 337955 717600 338123
rect 675887 337479 717600 337955
rect 675943 337311 717600 337479
rect 675887 336927 717600 337311
rect 675943 336759 717600 336927
rect 675887 336283 717600 336759
rect 675943 336115 717600 336283
rect 675887 335639 717600 336115
rect 675943 335471 717600 335639
rect 675887 335087 717600 335471
rect 675943 334919 717600 335087
rect 675887 334443 717600 334919
rect 675943 334275 717600 334443
rect 675887 333799 717600 334275
rect 675407 333729 675887 333743
rect 675312 333701 675887 333729
rect 673828 327140 673880 327146
rect 673828 327082 673880 327088
rect 673840 304978 673868 327082
rect 675312 325725 675340 333701
rect 675407 333687 675887 333701
rect 675943 333631 717600 333799
rect 675887 333155 717600 333631
rect 675943 332987 717600 333155
rect 675887 332603 717600 332987
rect 675943 332435 717600 332603
rect 675887 331959 717600 332435
rect 675943 331791 717600 331959
rect 675887 331315 717600 331791
rect 675943 331147 717600 331315
rect 675887 330763 717600 331147
rect 675407 330651 675887 330707
rect 675943 330595 717600 330763
rect 675887 330119 717600 330595
rect 675943 329951 717600 330119
rect 675887 329475 717600 329951
rect 675407 329363 675887 329419
rect 675943 329307 717600 329475
rect 675887 328923 717600 329307
rect 675407 328811 675887 328867
rect 675943 328755 717600 328923
rect 675887 328279 717600 328755
rect 675943 328111 717600 328279
rect 675887 327635 717600 328111
rect 675407 327556 675887 327579
rect 675404 327523 675887 327556
rect 675404 327146 675432 327523
rect 675943 327467 717600 327635
rect 675392 327140 675444 327146
rect 675392 327082 675444 327088
rect 675887 327083 717600 327467
rect 675407 326971 675887 327027
rect 675943 326915 717600 327083
rect 675887 326439 717600 326915
rect 675943 326271 717600 326439
rect 675887 325795 717600 326271
rect 675407 325725 675887 325739
rect 675312 325697 675887 325725
rect 675407 325683 675887 325697
rect 675943 325627 717600 325795
rect 675887 325417 717600 325627
rect 673828 304972 673880 304978
rect 673828 304914 673880 304920
rect 675887 296159 717600 296358
rect 675407 296047 675887 296103
rect 675943 295991 717600 296159
rect 675887 295607 717600 295991
rect 675943 295439 717600 295607
rect 675887 294963 717600 295439
rect 675943 294795 717600 294963
rect 675887 294319 717600 294795
rect 675943 294151 717600 294319
rect 675887 293767 717600 294151
rect 673644 293548 673696 293554
rect 673644 293490 673696 293496
rect 675024 293548 675076 293554
rect 675024 293490 675076 293496
rect 673460 283076 673512 283082
rect 673460 283018 673512 283024
rect 672644 276032 672764 276060
rect 672736 256714 672764 276032
rect 673736 266348 673788 266354
rect 673736 266290 673788 266296
rect 672552 256686 672764 256714
rect 672552 231849 672580 256686
rect 673644 247512 673696 247518
rect 673644 247454 673696 247460
rect 672538 231840 672594 231849
rect 672538 231775 672594 231784
rect 672906 231840 672962 231849
rect 672906 231775 672962 231784
rect 672920 212566 672948 231775
rect 672724 212560 672776 212566
rect 672724 212502 672776 212508
rect 672908 212560 672960 212566
rect 672908 212502 672960 212508
rect 672736 198762 672764 212502
rect 673460 203380 673512 203386
rect 673460 203322 673512 203328
rect 672540 198756 672592 198762
rect 672540 198698 672592 198704
rect 672724 198756 672776 198762
rect 672724 198698 672776 198704
rect 44640 195900 44692 195906
rect 44640 195842 44692 195848
rect 44652 193225 44680 195842
rect 672552 193225 672580 198698
rect 44454 193216 44510 193225
rect 44454 193151 44510 193160
rect 44638 193216 44694 193225
rect 44638 193151 44694 193160
rect 672538 193216 672594 193225
rect 672538 193151 672594 193160
rect 672906 193216 672962 193225
rect 672906 193151 672962 193160
rect 44468 173942 44496 193151
rect 672920 173942 672948 193151
rect 44456 173936 44508 173942
rect 44456 173878 44508 173884
rect 44732 173936 44784 173942
rect 44732 173878 44784 173884
rect 672724 173936 672776 173942
rect 672724 173878 672776 173884
rect 672908 173936 672960 173942
rect 672908 173878 672960 173884
rect 44744 160206 44772 173878
rect 44732 160200 44784 160206
rect 44732 160142 44784 160148
rect 672736 160138 672764 173878
rect 672540 160132 672592 160138
rect 672540 160074 672592 160080
rect 672724 160132 672776 160138
rect 672724 160074 672776 160080
rect 44640 160064 44692 160070
rect 44640 160006 44692 160012
rect 44652 154562 44680 160006
rect 44640 154556 44692 154562
rect 44640 154498 44692 154504
rect 44732 154556 44784 154562
rect 44732 154498 44784 154504
rect 44744 140826 44772 154498
rect 44732 140820 44784 140826
rect 44732 140762 44784 140768
rect 44640 140752 44692 140758
rect 44640 140694 44692 140700
rect 672552 140706 672580 160074
rect 673472 157350 673500 203322
rect 673656 203386 673684 247454
rect 673748 237726 673776 266290
rect 675036 293049 675064 293490
rect 675943 293599 717600 293767
rect 675887 293123 717600 293599
rect 675407 293049 675887 293067
rect 675022 293040 675078 293049
rect 675022 292975 675078 292984
rect 675206 293040 675262 293049
rect 675206 292975 675262 292984
rect 675390 293040 675887 293049
rect 675446 293011 675887 293040
rect 675390 292975 675446 292984
rect 674932 283076 674984 283082
rect 674932 283018 674984 283024
rect 673920 276072 673972 276078
rect 673920 276014 673972 276020
rect 673736 237720 673788 237726
rect 673736 237662 673788 237668
rect 673644 203380 673696 203386
rect 673644 203322 673696 203328
rect 673748 192409 673776 237662
rect 673932 247518 673960 276014
rect 674944 266354 674972 283018
rect 675220 276078 675248 292975
rect 675943 292955 717600 293123
rect 675887 292479 717600 292955
rect 675943 292311 717600 292479
rect 675887 291927 717600 292311
rect 675943 291759 717600 291927
rect 675887 291283 717600 291759
rect 675943 291115 717600 291283
rect 675887 290639 717600 291115
rect 675943 290471 717600 290639
rect 675887 290087 717600 290471
rect 675943 289919 717600 290087
rect 675887 289443 717600 289919
rect 675943 289275 717600 289443
rect 675887 288799 717600 289275
rect 675407 288729 675887 288743
rect 675312 288701 675887 288729
rect 675312 280725 675340 288701
rect 675407 288687 675887 288701
rect 675943 288631 717600 288799
rect 675887 288155 717600 288631
rect 675943 287987 717600 288155
rect 675887 287603 717600 287987
rect 675943 287435 717600 287603
rect 675887 286959 717600 287435
rect 675943 286791 717600 286959
rect 675887 286315 717600 286791
rect 675943 286147 717600 286315
rect 675887 285763 717600 286147
rect 675407 285651 675887 285707
rect 675943 285595 717600 285763
rect 675887 285119 717600 285595
rect 675943 284951 717600 285119
rect 675887 284475 717600 284951
rect 675407 284363 675887 284419
rect 675943 284307 717600 284475
rect 675887 283923 717600 284307
rect 675407 283811 675887 283867
rect 675943 283755 717600 283923
rect 675887 283279 717600 283755
rect 675943 283111 717600 283279
rect 675392 283076 675444 283082
rect 675392 283018 675444 283024
rect 675404 282579 675432 283018
rect 675887 282635 717600 283111
rect 675404 282540 675887 282579
rect 675407 282523 675887 282540
rect 675943 282467 717600 282635
rect 675887 282083 717600 282467
rect 675407 281971 675887 282027
rect 675943 281915 717600 282083
rect 675887 281439 717600 281915
rect 675943 281271 717600 281439
rect 675887 280795 717600 281271
rect 675407 280725 675887 280739
rect 675312 280697 675887 280725
rect 675407 280683 675887 280697
rect 675943 280627 717600 280795
rect 675887 280417 717600 280627
rect 675208 276072 675260 276078
rect 675208 276014 675260 276020
rect 674932 266348 674984 266354
rect 674932 266290 674984 266296
rect 675887 251159 717600 251358
rect 675407 251047 675887 251103
rect 675943 250991 717600 251159
rect 675887 250607 717600 250991
rect 675943 250439 717600 250607
rect 675887 249963 717600 250439
rect 675943 249795 717600 249963
rect 675887 249319 717600 249795
rect 675943 249151 717600 249319
rect 675887 248767 717600 249151
rect 675943 248599 717600 248767
rect 675887 248123 717600 248599
rect 675407 248039 675887 248067
rect 675404 248011 675887 248039
rect 675404 247518 675432 248011
rect 675943 247955 717600 248123
rect 673920 247512 673972 247518
rect 673920 247454 673972 247460
rect 675392 247512 675444 247518
rect 675887 247479 717600 247955
rect 675392 247454 675444 247460
rect 675943 247311 717600 247479
rect 675887 246927 717600 247311
rect 675943 246759 717600 246927
rect 675887 246283 717600 246759
rect 675943 246115 717600 246283
rect 675887 245639 717600 246115
rect 675943 245471 717600 245639
rect 675887 245087 717600 245471
rect 675943 244919 717600 245087
rect 675887 244443 717600 244919
rect 675943 244275 717600 244443
rect 675887 243799 717600 244275
rect 675407 243729 675887 243743
rect 675312 243701 675887 243729
rect 675312 235725 675340 243701
rect 675407 243687 675887 243701
rect 675943 243631 717600 243799
rect 675887 243155 717600 243631
rect 675943 242987 717600 243155
rect 675887 242603 717600 242987
rect 675943 242435 717600 242603
rect 675887 241959 717600 242435
rect 675943 241791 717600 241959
rect 675887 241315 717600 241791
rect 675943 241147 717600 241315
rect 675887 240763 717600 241147
rect 675407 240651 675887 240707
rect 675943 240595 717600 240763
rect 675887 240119 717600 240595
rect 675943 239951 717600 240119
rect 675887 239475 717600 239951
rect 675407 239363 675887 239419
rect 675943 239307 717600 239475
rect 675887 238923 717600 239307
rect 675407 238811 675887 238867
rect 675943 238755 717600 238923
rect 675887 238279 717600 238755
rect 675943 238111 717600 238279
rect 675392 237720 675444 237726
rect 675392 237662 675444 237668
rect 675404 237579 675432 237662
rect 675887 237635 717600 238111
rect 675404 237524 675887 237579
rect 675407 237523 675887 237524
rect 675943 237467 717600 237635
rect 675887 237083 717600 237467
rect 675407 236971 675887 237027
rect 675943 236915 717600 237083
rect 675887 236439 717600 236915
rect 675943 236271 717600 236439
rect 675887 235795 717600 236271
rect 675407 235725 675887 235739
rect 675312 235697 675887 235725
rect 675407 235683 675887 235697
rect 675943 235627 717600 235795
rect 675887 235417 717600 235627
rect 675887 205959 717600 206158
rect 675407 205847 675887 205903
rect 675943 205791 717600 205959
rect 675887 205407 717600 205791
rect 675943 205239 717600 205407
rect 675887 204763 717600 205239
rect 675943 204595 717600 204763
rect 675887 204119 717600 204595
rect 675943 203951 717600 204119
rect 675887 203567 717600 203951
rect 675943 203399 717600 203567
rect 675392 203380 675444 203386
rect 675392 203322 675444 203328
rect 675404 202867 675432 203322
rect 675887 202923 717600 203399
rect 675404 202844 675887 202867
rect 675407 202811 675887 202844
rect 675943 202755 717600 202923
rect 675887 202279 717600 202755
rect 675943 202111 717600 202279
rect 675887 201727 717600 202111
rect 675943 201559 717600 201727
rect 675887 201083 717600 201559
rect 675943 200915 717600 201083
rect 675887 200439 717600 200915
rect 675943 200271 717600 200439
rect 675887 199887 717600 200271
rect 675943 199719 717600 199887
rect 675887 199243 717600 199719
rect 675943 199075 717600 199243
rect 675312 198614 675432 198642
rect 673734 192400 673790 192409
rect 673734 192335 673790 192344
rect 673748 192030 673776 192335
rect 673736 192024 673788 192030
rect 673736 191966 673788 191972
rect 674012 192024 674064 192030
rect 674012 191966 674064 191972
rect 674024 173942 674052 191966
rect 675312 190525 675340 198614
rect 675404 198543 675432 198614
rect 675887 198599 717600 199075
rect 675404 198492 675887 198543
rect 675407 198487 675887 198492
rect 675943 198431 717600 198599
rect 675887 197955 717600 198431
rect 675943 197787 717600 197955
rect 675887 197403 717600 197787
rect 675943 197235 717600 197403
rect 675887 196759 717600 197235
rect 675943 196591 717600 196759
rect 675887 196115 717600 196591
rect 675943 195947 717600 196115
rect 675887 195563 717600 195947
rect 675407 195451 675887 195507
rect 675943 195395 717600 195563
rect 675887 194919 717600 195395
rect 675943 194751 717600 194919
rect 675887 194275 717600 194751
rect 675407 194163 675887 194219
rect 675943 194107 717600 194275
rect 675887 193723 717600 194107
rect 675407 193611 675887 193667
rect 675943 193555 717600 193723
rect 675887 193079 717600 193555
rect 675943 192911 717600 193079
rect 675887 192435 717600 192911
rect 675390 192400 675446 192409
rect 675446 192344 675887 192379
rect 675390 192335 675887 192344
rect 675407 192323 675887 192335
rect 675943 192267 717600 192435
rect 675887 191883 717600 192267
rect 675407 191771 675887 191827
rect 675943 191715 717600 191883
rect 675887 191239 717600 191715
rect 675943 191071 717600 191239
rect 675887 190595 717600 191071
rect 675407 190525 675887 190539
rect 675312 190497 675887 190525
rect 675407 190483 675887 190497
rect 675943 190427 717600 190595
rect 675887 190217 717600 190427
rect 673828 173936 673880 173942
rect 673828 173878 673880 173884
rect 674012 173936 674064 173942
rect 674012 173878 674064 173884
rect 673840 160138 673868 173878
rect 675887 160959 717600 161158
rect 675407 160847 675887 160903
rect 675943 160791 717600 160959
rect 675887 160407 717600 160791
rect 675943 160239 717600 160407
rect 673644 160132 673696 160138
rect 673644 160074 673696 160080
rect 673828 160132 673880 160138
rect 673828 160074 673880 160080
rect 673460 157344 673512 157350
rect 673460 157286 673512 157292
rect 44652 135266 44680 140694
rect 672552 140678 672672 140706
rect 44652 135238 44772 135266
rect 44744 121582 44772 135238
rect 44732 121576 44784 121582
rect 44732 121518 44784 121524
rect 44640 121440 44692 121446
rect 44640 121382 44692 121388
rect 672644 121394 672672 140678
rect 44178 120184 44234 120193
rect 44178 120119 44234 120128
rect 42338 115968 42394 115977
rect 42338 115903 42394 115912
rect 44192 110537 44220 120119
rect 44178 110528 44234 110537
rect 44178 110463 44234 110472
rect 44652 102082 44680 121382
rect 672644 121366 672764 121394
rect 672736 115938 672764 121366
rect 672724 115932 672776 115938
rect 672724 115874 672776 115880
rect 672816 115932 672868 115938
rect 672816 115874 672868 115880
rect 45466 110528 45522 110537
rect 45466 110463 45522 110472
rect 44560 102054 44680 102082
rect 44560 96626 44588 102054
rect 44272 96620 44324 96626
rect 44272 96562 44324 96568
rect 44548 96620 44600 96626
rect 44548 96562 44600 96568
rect 44284 77314 44312 96562
rect 44272 77308 44324 77314
rect 44272 77250 44324 77256
rect 44364 77308 44416 77314
rect 44364 77250 44416 77256
rect 44270 75848 44326 75857
rect 44376 75834 44404 77250
rect 44326 75806 44404 75834
rect 44270 75783 44326 75792
rect 44284 73273 44312 75783
rect 44270 73264 44326 73273
rect 44270 73199 44326 73208
rect 44284 68241 44312 73199
rect 44270 68232 44326 68241
rect 44270 68167 44326 68176
rect 42708 64660 42760 64666
rect 42708 64602 42760 64608
rect 42720 45626 42748 64602
rect 45480 47938 45508 110463
rect 672828 102202 672856 115874
rect 673472 112130 673500 157286
rect 673656 147898 673684 160074
rect 675887 159763 717600 160239
rect 675943 159595 717600 159763
rect 675887 159119 717600 159595
rect 675943 158951 717600 159119
rect 675887 158567 717600 158951
rect 675943 158399 717600 158567
rect 675887 157923 717600 158399
rect 675407 157828 675887 157867
rect 675404 157811 675887 157828
rect 675404 157350 675432 157811
rect 675943 157755 717600 157923
rect 675392 157344 675444 157350
rect 675392 157286 675444 157292
rect 675887 157279 717600 157755
rect 675943 157111 717600 157279
rect 675887 156727 717600 157111
rect 675943 156559 717600 156727
rect 675887 156083 717600 156559
rect 675943 155915 717600 156083
rect 675887 155439 717600 155915
rect 675943 155271 717600 155439
rect 675887 154887 717600 155271
rect 675943 154719 717600 154887
rect 675887 154243 717600 154719
rect 675943 154075 717600 154243
rect 675887 153599 717600 154075
rect 675407 153529 675887 153543
rect 675312 153501 675887 153529
rect 673644 147892 673696 147898
rect 673644 147834 673696 147840
rect 674012 147892 674064 147898
rect 674012 147834 674064 147840
rect 674024 140706 674052 147834
rect 675312 145525 675340 153501
rect 675407 153487 675887 153501
rect 675943 153431 717600 153599
rect 675887 152955 717600 153431
rect 675943 152787 717600 152955
rect 675887 152403 717600 152787
rect 675943 152235 717600 152403
rect 675887 151759 717600 152235
rect 675943 151591 717600 151759
rect 675887 151115 717600 151591
rect 675943 150947 717600 151115
rect 675887 150563 717600 150947
rect 675407 150451 675887 150507
rect 675943 150395 717600 150563
rect 675887 149919 717600 150395
rect 675943 149751 717600 149919
rect 675887 149275 717600 149751
rect 675407 149163 675887 149219
rect 675943 149107 717600 149275
rect 675887 148723 717600 149107
rect 675407 148611 675887 148667
rect 675943 148555 717600 148723
rect 675887 148079 717600 148555
rect 675943 147911 717600 148079
rect 675392 147892 675444 147898
rect 675392 147834 675444 147840
rect 675404 147379 675432 147834
rect 675887 147435 717600 147911
rect 675404 147356 675887 147379
rect 675407 147323 675887 147356
rect 675943 147267 717600 147435
rect 675887 146883 717600 147267
rect 675407 146771 675887 146827
rect 675943 146715 717600 146883
rect 675887 146239 717600 146715
rect 675943 146071 717600 146239
rect 675887 145595 717600 146071
rect 675407 145525 675887 145539
rect 675312 145497 675887 145525
rect 675407 145483 675887 145497
rect 675943 145427 717600 145595
rect 675887 145217 717600 145427
rect 673932 140678 674052 140706
rect 673932 121530 673960 140678
rect 673840 121502 673960 121530
rect 673460 112124 673512 112130
rect 673460 112066 673512 112072
rect 672816 102196 672868 102202
rect 672816 102138 672868 102144
rect 672724 102128 672776 102134
rect 672724 102070 672776 102076
rect 672736 96642 672764 102070
rect 672736 96614 672856 96642
rect 672828 82958 672856 96614
rect 672816 82952 672868 82958
rect 672816 82894 672868 82900
rect 672816 82748 672868 82754
rect 672816 82690 672868 82696
rect 45558 68232 45614 68241
rect 45558 68167 45614 68176
rect 45468 47932 45520 47938
rect 45468 47874 45520 47880
rect 45572 47802 45600 68167
rect 179420 47932 179472 47938
rect 179420 47874 179472 47880
rect 518808 47932 518860 47938
rect 518808 47874 518860 47880
rect 45560 47796 45612 47802
rect 45560 47738 45612 47744
rect 149060 47796 149112 47802
rect 149060 47738 149112 47744
rect 86316 47728 86368 47734
rect 86316 47670 86368 47676
rect 86328 47394 86356 47670
rect 86316 47388 86368 47394
rect 86316 47330 86368 47336
rect 42708 45620 42760 45626
rect 42708 45562 42760 45568
rect 86328 40225 86356 47330
rect 149072 47122 149100 47738
rect 179432 47530 179460 47874
rect 189172 47864 189224 47870
rect 189172 47806 189224 47812
rect 179420 47524 179472 47530
rect 179420 47466 179472 47472
rect 154578 47152 154634 47161
rect 149060 47116 149112 47122
rect 154578 47087 154580 47096
rect 149060 47058 149112 47064
rect 154632 47087 154634 47096
rect 173806 47152 173862 47161
rect 173806 47087 173862 47096
rect 188528 47116 188580 47122
rect 154580 47058 154632 47064
rect 140964 45620 141016 45626
rect 140964 45562 141016 45568
rect 140976 44198 141004 45562
rect 140964 44192 141016 44198
rect 140964 44134 141016 44140
rect 133098 40248 133150 40254
rect 86314 40216 86370 40225
rect 133098 40190 133150 40196
rect 140976 40202 141004 44134
rect 143816 40248 143868 40254
rect 86314 40151 86370 40160
rect 133110 40000 133138 40190
rect 140976 40174 141036 40202
rect 149072 40361 149100 47058
rect 173820 47054 173848 47087
rect 188528 47058 188580 47064
rect 173808 47048 173860 47054
rect 173808 46990 173860 46996
rect 186688 46980 186740 46986
rect 186688 46922 186740 46928
rect 186700 42193 186728 46922
rect 188540 42193 188568 47058
rect 189184 42193 189212 47806
rect 212538 47696 212594 47705
rect 212538 47631 212540 47640
rect 212592 47631 212594 47640
rect 231582 47696 231638 47705
rect 231582 47631 231638 47640
rect 270498 47696 270554 47705
rect 270498 47631 270500 47640
rect 212540 47602 212592 47608
rect 195980 47592 196032 47598
rect 195980 47534 196032 47540
rect 198648 47592 198700 47598
rect 198740 47592 198792 47598
rect 198700 47540 198740 47546
rect 198648 47534 198792 47540
rect 192852 47116 192904 47122
rect 192852 47058 192904 47064
rect 192864 42193 192892 47058
rect 194692 46980 194744 46986
rect 194692 46922 194744 46928
rect 194704 42193 194732 46922
rect 195992 42193 196020 47534
rect 198660 47518 198780 47534
rect 231596 47410 231624 47631
rect 270552 47631 270554 47640
rect 289634 47696 289690 47705
rect 289634 47631 289690 47640
rect 270500 47602 270552 47608
rect 231768 47524 231820 47530
rect 231768 47466 231820 47472
rect 251180 47524 251232 47530
rect 251180 47466 251232 47472
rect 270408 47524 270460 47530
rect 270408 47466 270460 47472
rect 231780 47410 231808 47466
rect 199016 47388 199068 47394
rect 199016 47330 199068 47336
rect 201408 47388 201460 47394
rect 231596 47382 231808 47410
rect 251192 47394 251220 47466
rect 270420 47394 270448 47466
rect 289648 47410 289676 47631
rect 303620 47592 303672 47598
rect 303620 47534 303672 47540
rect 304540 47592 304592 47598
rect 304540 47534 304592 47540
rect 359372 47592 359424 47598
rect 359372 47534 359424 47540
rect 361488 47592 361540 47598
rect 361488 47534 361540 47540
rect 289728 47456 289780 47462
rect 289648 47404 289728 47410
rect 289648 47398 289780 47404
rect 251180 47388 251232 47394
rect 201408 47330 201460 47336
rect 251180 47330 251232 47336
rect 270408 47388 270460 47394
rect 289648 47382 289768 47398
rect 303632 47394 303660 47534
rect 303620 47388 303672 47394
rect 270408 47330 270460 47336
rect 303620 47330 303672 47336
rect 199028 42193 199056 47330
rect 200856 47184 200908 47190
rect 200856 47126 200908 47132
rect 200868 42193 200896 47126
rect 201420 47122 201448 47330
rect 285588 47320 285640 47326
rect 285588 47262 285640 47268
rect 217968 47252 218020 47258
rect 217968 47194 218020 47200
rect 240140 47252 240192 47258
rect 240140 47194 240192 47200
rect 201408 47116 201460 47122
rect 201408 47058 201460 47064
rect 217980 47054 218008 47194
rect 201592 47048 201644 47054
rect 201592 46990 201644 46996
rect 217968 47048 218020 47054
rect 217968 46990 218020 46996
rect 186683 41713 186739 42193
rect 187971 41713 188027 42193
rect 188523 41713 188579 42193
rect 189167 41834 189223 42193
rect 189264 41880 189316 41886
rect 189167 41828 189264 41834
rect 189167 41822 189316 41828
rect 189167 41806 189304 41822
rect 189167 41713 189223 41806
rect 189811 41713 189867 42193
rect 190363 41713 190419 42193
rect 191007 41834 191063 42193
rect 191104 41880 191156 41886
rect 191007 41828 191104 41834
rect 191007 41822 191156 41828
rect 191007 41806 191144 41822
rect 191007 41713 191063 41806
rect 191651 41713 191707 42193
rect 192203 41834 192259 42193
rect 192300 41880 192352 41886
rect 192203 41828 192300 41834
rect 192203 41822 192352 41828
rect 192203 41806 192340 41822
rect 192203 41713 192259 41806
rect 192847 41713 192903 42193
rect 193491 41834 193547 42193
rect 193491 41818 193628 41834
rect 193491 41812 193640 41818
rect 193491 41806 193588 41812
rect 193491 41713 193547 41806
rect 193588 41754 193640 41760
rect 194687 41713 194743 42193
rect 195975 41713 196031 42193
rect 196527 41834 196583 42193
rect 197171 41834 197227 42193
rect 197815 41834 197871 42193
rect 198367 41834 198423 42193
rect 196452 41818 198504 41834
rect 196440 41812 198516 41818
rect 196492 41806 198464 41812
rect 196440 41754 196492 41760
rect 196527 41713 196583 41806
rect 197171 41713 197227 41806
rect 197815 41713 197871 41806
rect 198367 41713 198423 41806
rect 198464 41754 198516 41760
rect 199011 41713 199067 42193
rect 200207 41834 200263 42193
rect 200851 41834 200907 42193
rect 200132 41818 200907 41834
rect 200120 41812 200907 41818
rect 200172 41806 200907 41812
rect 200120 41754 200172 41760
rect 200207 41713 200263 41806
rect 200851 41713 200907 41806
rect 201495 41834 201551 42193
rect 201604 41834 201632 46990
rect 201495 41806 201632 41834
rect 201495 41713 201551 41806
rect 202047 41713 202103 42193
rect 186417 41657 186627 41713
rect 186795 41657 187271 41713
rect 187439 41657 187915 41713
rect 188083 41657 188467 41713
rect 188635 41657 189111 41713
rect 189279 41657 189755 41713
rect 189923 41657 190307 41713
rect 190475 41657 190951 41713
rect 191119 41657 191595 41713
rect 191763 41657 192147 41713
rect 192315 41657 192791 41713
rect 192959 41657 193435 41713
rect 193603 41657 193987 41713
rect 194155 41657 194631 41713
rect 194799 41657 195275 41713
rect 195443 41657 195919 41713
rect 196087 41657 196471 41713
rect 196639 41657 197115 41713
rect 197283 41657 197759 41713
rect 197927 41657 198311 41713
rect 198479 41657 198955 41713
rect 199123 41657 199599 41713
rect 199767 41657 200151 41713
rect 200319 41657 200795 41713
rect 200963 41657 201439 41713
rect 201607 41657 201991 41713
rect 202159 41657 202358 41713
rect 149058 40352 149114 40361
rect 149058 40287 149114 40296
rect 143816 40190 143868 40196
rect 141008 40118 141036 40174
rect 140996 40112 141048 40118
rect 140996 40054 141048 40060
rect 143072 40112 143124 40118
rect 143072 40054 143124 40060
rect 143356 40112 143408 40118
rect 143356 40054 143408 40060
rect 141008 40000 141036 40054
rect 143084 40000 143112 40054
rect 143368 40000 143396 40054
rect 143828 40000 143856 40190
rect 78942 34868 83722 40000
rect 83778 39533 88865 39593
rect 88921 39589 93701 40000
rect 132617 39816 140940 40000
rect 140996 39872 141048 40000
rect 141104 39878 141313 40000
rect 141369 39934 141499 40000
rect 141555 39878 141898 40000
rect 141954 39934 142084 40000
rect 142140 39878 143012 40000
rect 141104 39816 143012 39878
rect 83778 34812 93747 39533
rect 78942 985 93747 34812
rect 132617 39204 143012 39816
rect 132617 39147 142955 39204
rect 143068 39151 143128 40000
rect 143184 39747 144517 40000
rect 144573 39803 144689 40000
rect 144745 39747 145035 40000
rect 143184 39650 145035 39747
rect 145199 39650 147532 40000
rect 143184 39369 147532 39650
rect 143184 39297 144495 39369
rect 145520 39341 147532 39369
rect 143184 39243 144441 39297
rect 144551 39285 145464 39313
rect 144551 39271 145530 39285
rect 145586 39275 147532 39341
rect 144551 39261 145436 39271
rect 143184 39207 144367 39243
rect 144551 39241 144623 39261
rect 144625 39241 144645 39261
rect 145414 39247 145461 39261
rect 145464 39247 145530 39271
rect 143244 39169 144367 39207
rect 144497 39233 144551 39241
rect 144571 39233 144625 39241
rect 144497 39205 144625 39233
rect 145414 39219 145530 39247
rect 145414 39214 145461 39219
rect 144497 39187 144551 39205
rect 144571 39187 144625 39205
rect 143068 39148 143188 39151
rect 132617 39076 141720 39147
rect 143011 39091 143188 39148
rect 143244 39147 144345 39169
rect 144423 39113 144571 39187
rect 144701 39185 145358 39205
rect 144681 39158 145358 39185
rect 145461 39191 145525 39214
rect 145530 39191 145599 39219
rect 145655 39206 147532 39275
rect 145461 39163 145599 39191
rect 144681 39131 145405 39158
rect 145461 39150 145525 39163
rect 145530 39150 145599 39163
rect 144401 39091 144497 39113
rect 132617 39010 141654 39076
rect 141776 39063 144497 39091
rect 141776 39049 141847 39063
rect 143068 39049 143128 39063
rect 144423 39049 144497 39063
rect 144627 39094 145405 39131
rect 145525 39135 145591 39150
rect 145599 39135 145653 39150
rect 144627 39057 145469 39094
rect 145525 39085 145653 39135
rect 145525 39084 145591 39085
rect 141776 39039 144497 39049
rect 141776 39020 141847 39039
rect 141850 39020 141869 39039
rect 144553 39028 145469 39057
rect 141710 39011 141776 39020
rect 141784 39011 141850 39020
rect 132617 37861 141628 39010
rect 141710 38969 141850 39011
rect 144553 38983 145545 39028
rect 141710 38954 141776 38969
rect 141784 38954 141850 38969
rect 141925 38964 145545 38983
rect 141684 38928 141710 38954
rect 141736 38928 141784 38954
rect 141684 38906 141784 38928
rect 132617 37823 141590 37861
rect 132617 36927 141538 37823
rect 141684 37805 141736 38906
rect 141906 38898 145545 38964
rect 141840 38850 145545 38898
rect 141646 37783 141736 37805
rect 141646 37767 141684 37783
rect 141720 37767 141736 37783
rect 141792 38284 145545 38850
rect 141792 38216 145477 38284
rect 145601 38228 145653 39085
rect 141792 38176 145437 38216
rect 145533 38178 145653 38228
rect 141792 38110 145371 38176
rect 145533 38160 145601 38178
rect 145607 38160 145653 38178
rect 145493 38150 145533 38160
rect 145567 38150 145607 38160
rect 145493 38136 145607 38150
rect 145493 38120 145533 38136
rect 145567 38120 145607 38136
rect 141594 37693 141720 37767
rect 141792 37711 145319 38110
rect 145427 38108 145493 38120
rect 145501 38108 145567 38120
rect 145427 38080 145567 38108
rect 145709 38104 147532 39206
rect 145427 38054 145493 38080
rect 145501 38054 145567 38080
rect 145663 38064 147532 38104
rect 132617 36860 141471 36927
rect 141594 36871 141646 37693
rect 141776 37637 145319 37711
rect 132617 35845 141419 36860
rect 141527 36821 141646 36871
rect 141527 36804 141594 36821
rect 141601 36804 141646 36821
rect 141475 36730 141601 36804
rect 141702 36748 145319 37637
rect 141475 35901 141527 36730
rect 141657 36674 145319 36748
rect 141583 35845 145319 36674
rect 132617 34484 145319 35845
rect 145375 37980 145501 38054
rect 145623 37998 147532 38064
rect 145375 34678 145427 37980
rect 145557 37924 147532 37998
rect 145483 34734 147532 37924
rect 145375 34540 145470 34678
rect 132617 34469 145362 34484
rect 132617 33839 145319 34469
rect 145418 34413 145470 34540
rect 145375 34371 145470 34413
rect 145375 34370 145418 34371
rect 145375 34275 145470 34370
rect 132617 33810 145290 33839
rect 132617 33765 145245 33810
rect 145375 33783 145427 34275
rect 145526 34219 147532 34734
rect 132617 32852 145240 33765
rect 145346 33754 145427 33783
rect 145301 33747 145346 33754
rect 145375 33747 145427 33754
rect 145301 33733 145427 33747
rect 145301 33709 145346 33733
rect 145375 33709 145427 33733
rect 145296 33704 145301 33709
rect 145348 33704 145375 33709
rect 145296 33682 145375 33704
rect 132617 32688 145114 32852
rect 145296 32796 145348 33682
rect 145483 33653 147532 34219
rect 145431 33626 147532 33653
rect 145170 32744 145348 32796
rect 145404 32688 147532 33626
rect 132617 158 147532 32688
rect 186417 0 202358 41657
rect 240152 39953 240180 47194
rect 242900 47184 242952 47190
rect 242900 47126 242952 47132
rect 242912 45558 242940 47126
rect 285600 47122 285628 47262
rect 299480 47184 299532 47190
rect 299480 47126 299532 47132
rect 247408 47116 247460 47122
rect 247408 47058 247460 47064
rect 285588 47116 285640 47122
rect 285588 47058 285640 47064
rect 242900 45552 242952 45558
rect 242900 45494 242952 45500
rect 240138 39944 240194 39953
rect 240138 39879 240194 39888
rect 242912 39817 242940 45494
rect 241242 39808 241298 39817
rect 241242 39743 241298 39752
rect 242898 39808 242954 39817
rect 242898 39743 242954 39752
rect 241256 39600 241284 39743
rect 247420 39600 247448 47058
rect 297732 45552 297784 45558
rect 297732 45494 297784 45500
rect 254032 44192 254084 44198
rect 254032 44134 254084 44140
rect 253940 41608 253992 41614
rect 253940 41550 253992 41556
rect 253952 39953 253980 41550
rect 253938 39944 253994 39953
rect 253938 39879 253994 39888
rect 254044 39710 254072 44134
rect 297744 42193 297772 45494
rect 295283 41834 295339 42193
rect 295283 41818 295472 41834
rect 295283 41812 295484 41818
rect 295283 41806 295432 41812
rect 295283 41713 295339 41806
rect 295432 41754 295484 41760
rect 295927 41713 295983 42193
rect 296571 41713 296627 42193
rect 296904 41948 296956 41954
rect 296904 41890 296956 41896
rect 296916 41834 296944 41890
rect 297123 41834 297179 42193
rect 296916 41806 297179 41834
rect 297744 41834 297823 42193
rect 297916 41880 297968 41886
rect 297744 41828 297916 41834
rect 297744 41822 297968 41828
rect 297744 41806 297956 41822
rect 297123 41713 297179 41806
rect 297767 41713 297823 41806
rect 298411 41713 298467 42193
rect 298963 41713 299019 42193
rect 299492 42022 299520 47126
rect 304552 42193 304580 47534
rect 307576 47320 307628 47326
rect 307576 47262 307628 47268
rect 305736 47184 305788 47190
rect 305736 47126 305788 47132
rect 305748 42193 305776 47126
rect 307588 42193 307616 47262
rect 309416 47252 309468 47258
rect 309416 47194 309468 47200
rect 352564 47252 352616 47258
rect 352564 47194 352616 47200
rect 309428 42193 309456 47194
rect 351920 47184 351972 47190
rect 351920 47126 351972 47132
rect 351932 42193 351960 47126
rect 352576 42193 352604 47194
rect 359384 42193 359412 47534
rect 361500 47394 361528 47534
rect 416780 47524 416832 47530
rect 416780 47466 416832 47472
rect 364156 47456 364208 47462
rect 364156 47398 364208 47404
rect 361488 47388 361540 47394
rect 361488 47330 361540 47336
rect 364168 47326 364196 47398
rect 414204 47388 414256 47394
rect 414204 47330 414256 47336
rect 362408 47320 362460 47326
rect 362408 47262 362460 47268
rect 364156 47320 364208 47326
rect 364156 47262 364208 47268
rect 406752 47320 406804 47326
rect 406752 47262 406804 47268
rect 360568 47184 360620 47190
rect 360568 47126 360620 47132
rect 360580 42193 360608 47126
rect 362420 42193 362448 47262
rect 364248 47252 364300 47258
rect 364248 47194 364300 47200
rect 364260 42193 364288 47194
rect 406764 47190 406792 47262
rect 407396 47252 407448 47258
rect 407396 47194 407448 47200
rect 406752 47184 406804 47190
rect 406752 47126 406804 47132
rect 406764 42193 406792 47126
rect 407408 42193 407436 47194
rect 414216 42193 414244 47330
rect 416792 47258 416820 47466
rect 417976 47388 418028 47394
rect 417976 47330 418028 47336
rect 418068 47388 418120 47394
rect 418068 47330 418120 47336
rect 471980 47388 472032 47394
rect 471980 47330 472032 47336
rect 416780 47252 416832 47258
rect 416780 47194 416832 47200
rect 417240 47252 417292 47258
rect 417240 47194 417292 47200
rect 417252 42193 417280 47194
rect 417988 47122 418016 47330
rect 418080 47258 418108 47330
rect 461492 47320 461544 47326
rect 461492 47262 461544 47268
rect 418068 47252 418120 47258
rect 418068 47194 418120 47200
rect 419080 47252 419132 47258
rect 419080 47194 419132 47200
rect 417976 47116 418028 47122
rect 417976 47058 418028 47064
rect 419092 42193 419120 47194
rect 461504 42193 461532 47262
rect 462136 47252 462188 47258
rect 462136 47194 462188 47200
rect 462148 42193 462176 47194
rect 468944 47116 468996 47122
rect 468944 47058 468996 47064
rect 468956 42193 468984 47058
rect 471992 42193 472020 47330
rect 518820 47326 518848 47874
rect 526812 47388 526864 47394
rect 526812 47330 526864 47336
rect 516324 47320 516376 47326
rect 516324 47262 516376 47268
rect 518808 47320 518860 47326
rect 518808 47262 518860 47268
rect 473820 47252 473872 47258
rect 473820 47194 473872 47200
rect 473832 42193 473860 47194
rect 514484 46980 514536 46986
rect 514484 46922 514536 46928
rect 514496 42193 514524 46922
rect 516336 42193 516364 47262
rect 516968 47252 517020 47258
rect 516968 47194 517020 47200
rect 516980 42193 517008 47194
rect 523776 47116 523828 47122
rect 523776 47058 523828 47064
rect 522488 46980 522540 46986
rect 522488 46922 522540 46928
rect 522500 42193 522528 46922
rect 523788 42193 523816 47058
rect 526824 46986 526852 47330
rect 672828 47802 672856 82690
rect 528652 47796 528704 47802
rect 528652 47738 528704 47744
rect 672816 47796 672868 47802
rect 672816 47738 672868 47744
rect 526812 46980 526864 46986
rect 526812 46922 526864 46928
rect 526824 42193 526852 46922
rect 528664 42193 528692 47738
rect 569132 47116 569184 47122
rect 569132 47058 569184 47064
rect 299480 42016 299532 42022
rect 299480 41958 299532 41964
rect 299492 41834 299520 41958
rect 299607 41834 299663 42193
rect 299492 41806 299663 41834
rect 299607 41713 299663 41806
rect 300251 41713 300307 42193
rect 300676 41880 300728 41886
rect 300803 41834 300859 42193
rect 301447 41834 301503 42193
rect 302091 41834 302147 42193
rect 302240 42016 302292 42022
rect 302240 41958 302292 41964
rect 302252 41834 302280 41958
rect 300728 41828 302280 41834
rect 300676 41822 302280 41828
rect 300688 41806 302280 41822
rect 300803 41713 300859 41806
rect 301447 41713 301503 41806
rect 302091 41713 302147 41806
rect 303287 41834 303343 42193
rect 303172 41818 303343 41834
rect 303160 41812 303343 41818
rect 303212 41806 303343 41812
rect 304552 41806 304631 42193
rect 305000 42016 305052 42022
rect 305000 41958 305052 41964
rect 305012 41834 305040 41958
rect 305127 41834 305183 42193
rect 305012 41818 305316 41834
rect 305012 41812 305328 41818
rect 305012 41806 305276 41812
rect 303160 41754 303212 41760
rect 303287 41713 303343 41806
rect 304575 41713 304631 41806
rect 305127 41713 305183 41806
rect 305748 41806 305827 42193
rect 305276 41754 305328 41760
rect 305771 41713 305827 41806
rect 306415 41834 306471 42193
rect 306415 41818 306604 41834
rect 306415 41812 306616 41818
rect 306415 41806 306564 41812
rect 306415 41713 306471 41806
rect 306564 41754 306616 41760
rect 307588 41806 307667 42193
rect 308807 41834 308863 42193
rect 309428 41834 309507 42193
rect 308692 41818 309507 41834
rect 307611 41713 307667 41806
rect 308680 41812 309507 41818
rect 308732 41806 309507 41812
rect 308680 41754 308732 41760
rect 308807 41713 308863 41806
rect 309451 41713 309507 41806
rect 310647 41713 310703 42193
rect 350083 41834 350139 42193
rect 350083 41818 350212 41834
rect 350083 41812 350224 41818
rect 350083 41806 350172 41812
rect 350083 41713 350139 41806
rect 350172 41754 350224 41760
rect 350727 41713 350783 42193
rect 351371 41713 351427 42193
rect 351923 41834 351979 42193
rect 352567 41970 352623 42193
rect 352567 41954 352696 41970
rect 352567 41948 352708 41954
rect 352567 41942 352656 41948
rect 352012 41880 352064 41886
rect 351923 41828 352012 41834
rect 351923 41822 352064 41828
rect 351923 41806 352052 41822
rect 351923 41713 351979 41806
rect 352567 41713 352623 41942
rect 352656 41890 352708 41896
rect 353211 41713 353267 42193
rect 353763 41713 353819 42193
rect 354312 41880 354364 41886
rect 354407 41834 354463 42193
rect 354364 41828 354463 41834
rect 354312 41822 354463 41828
rect 354324 41806 354463 41822
rect 354407 41713 354463 41806
rect 355051 41713 355107 42193
rect 355508 41948 355560 41954
rect 355508 41890 355560 41896
rect 355520 41834 355548 41890
rect 355603 41834 355659 42193
rect 356247 41834 356303 42193
rect 356891 41834 356947 42193
rect 356980 41948 357032 41954
rect 356980 41890 357032 41896
rect 356992 41834 357020 41890
rect 355520 41806 357020 41834
rect 355603 41713 355659 41806
rect 356247 41713 356303 41806
rect 356891 41713 356947 41806
rect 358087 41834 358143 42193
rect 358004 41818 358143 41834
rect 357992 41812 358143 41818
rect 358044 41806 358143 41812
rect 357992 41754 358044 41760
rect 358087 41713 358143 41806
rect 359375 41713 359431 42193
rect 359832 41948 359884 41954
rect 359832 41890 359884 41896
rect 359844 41834 359872 41890
rect 359927 41834 359983 42193
rect 359844 41806 359983 41834
rect 360476 41880 360528 41886
rect 360571 41834 360627 42193
rect 361120 41948 361172 41954
rect 361120 41890 361172 41896
rect 360528 41828 360627 41834
rect 360476 41822 360627 41828
rect 360488 41806 360627 41822
rect 361132 41834 361160 41890
rect 361215 41834 361271 42193
rect 361132 41806 361271 41834
rect 359927 41713 359983 41806
rect 360571 41713 360627 41806
rect 361215 41713 361271 41806
rect 362411 41713 362467 42193
rect 363607 41834 363663 42193
rect 364251 41834 364307 42193
rect 363524 41818 364307 41834
rect 363512 41812 364307 41818
rect 363564 41806 364307 41812
rect 363512 41754 363564 41760
rect 363607 41713 363663 41806
rect 364251 41713 364307 41806
rect 365447 41713 365503 42193
rect 404883 41834 404939 42193
rect 404883 41818 405044 41834
rect 404883 41812 405056 41818
rect 404883 41806 405004 41812
rect 404883 41713 404939 41806
rect 405004 41754 405056 41760
rect 406171 41713 406227 42193
rect 406723 41820 406792 42193
rect 407367 41970 407436 42193
rect 407367 41954 407528 41970
rect 407367 41948 407540 41954
rect 407367 41942 407488 41948
rect 407367 41820 407436 41942
rect 407488 41890 407540 41896
rect 406723 41713 406779 41820
rect 407367 41713 407423 41820
rect 408011 41713 408067 42193
rect 408563 41713 408619 42193
rect 409851 41713 409907 42193
rect 410248 41948 410300 41954
rect 410248 41890 410300 41896
rect 410260 41834 410288 41890
rect 410403 41834 410459 42193
rect 410260 41806 410459 41834
rect 410403 41713 410459 41806
rect 411536 42016 411588 42022
rect 411691 41970 411747 42193
rect 411588 41964 411760 41970
rect 411536 41958 411760 41964
rect 411548 41942 411760 41958
rect 411691 41820 411760 41942
rect 412887 41834 412943 42193
rect 411691 41713 411747 41820
rect 412744 41818 412943 41834
rect 412732 41812 412943 41818
rect 412784 41806 412943 41812
rect 412732 41754 412784 41760
rect 412887 41713 412943 41806
rect 414175 41820 414244 42193
rect 414572 42016 414624 42022
rect 414572 41958 414624 41964
rect 414584 41834 414612 41958
rect 414727 41834 414783 42193
rect 414175 41713 414231 41820
rect 414584 41806 414783 41834
rect 414727 41713 414783 41806
rect 415860 42016 415912 42022
rect 415860 41958 415912 41964
rect 415872 41834 415900 41958
rect 416015 41834 416071 42193
rect 415872 41806 416071 41834
rect 416015 41713 416071 41806
rect 417211 41820 417280 42193
rect 418252 42016 418304 42022
rect 418252 41958 418304 41964
rect 418264 41834 418292 41958
rect 418407 41834 418463 42193
rect 419051 41834 419120 42193
rect 418264 41820 419120 41834
rect 417211 41713 417267 41820
rect 418264 41806 419107 41820
rect 418407 41713 418463 41806
rect 419051 41713 419107 41806
rect 420247 41713 420303 42193
rect 459683 41834 459739 42193
rect 459836 41880 459888 41886
rect 459683 41828 459836 41834
rect 459683 41822 459888 41828
rect 459683 41806 459876 41822
rect 459683 41713 459739 41806
rect 460971 41713 461027 42193
rect 461504 41806 461579 42193
rect 462148 41834 462223 42193
rect 462320 41948 462372 41954
rect 462320 41890 462372 41896
rect 462332 41834 462360 41890
rect 462148 41806 462360 41834
rect 461523 41713 461579 41806
rect 462167 41713 462223 41806
rect 462811 41713 462867 42193
rect 463363 41713 463419 42193
rect 464651 41713 464707 42193
rect 465080 41948 465132 41954
rect 465080 41890 465132 41896
rect 465092 41834 465120 41890
rect 465203 41834 465259 42193
rect 465092 41806 465259 41834
rect 465203 41713 465259 41806
rect 466368 42016 466420 42022
rect 466368 41958 466420 41964
rect 466380 41834 466408 41958
rect 466491 41834 466547 42193
rect 466380 41806 466547 41834
rect 466491 41713 466547 41806
rect 467564 41880 467616 41886
rect 467687 41834 467743 42193
rect 467616 41828 467743 41834
rect 467564 41822 467743 41828
rect 467576 41806 467743 41822
rect 468956 41806 469031 42193
rect 469404 42016 469456 42022
rect 469404 41958 469456 41964
rect 469416 41834 469444 41958
rect 469527 41834 469583 42193
rect 470692 42016 470744 42022
rect 470692 41958 470744 41964
rect 469416 41806 469583 41834
rect 467687 41713 467743 41806
rect 468975 41713 469031 41806
rect 469527 41713 469583 41806
rect 470704 41834 470732 41958
rect 470815 41834 470871 42193
rect 470704 41806 470871 41834
rect 470815 41713 470871 41806
rect 471992 41806 472067 42193
rect 473084 42016 473136 42022
rect 473084 41958 473136 41964
rect 473096 41834 473124 41958
rect 473207 41834 473263 42193
rect 473832 41834 473907 42193
rect 473096 41806 473907 41834
rect 472011 41713 472067 41806
rect 473207 41713 473263 41806
rect 473851 41713 473907 41806
rect 475047 41713 475103 42193
rect 514483 41713 514539 42193
rect 515771 41713 515827 42193
rect 516323 41713 516379 42193
rect 516967 41834 517023 42193
rect 516967 41818 517100 41834
rect 516967 41812 517112 41818
rect 516967 41806 517060 41812
rect 516967 41713 517023 41806
rect 517060 41754 517112 41760
rect 517611 41713 517667 42193
rect 518163 41713 518219 42193
rect 519451 41713 519507 42193
rect 520003 41834 520059 42193
rect 520003 41818 520136 41834
rect 520003 41812 520148 41818
rect 520003 41806 520096 41812
rect 520003 41713 520059 41806
rect 520096 41754 520148 41760
rect 521291 41834 521347 42193
rect 521291 41818 521424 41834
rect 521291 41812 521436 41818
rect 521291 41806 521384 41812
rect 521291 41713 521347 41806
rect 521384 41754 521436 41760
rect 522487 41713 522543 42193
rect 523775 41713 523831 42193
rect 524327 41834 524383 42193
rect 524327 41818 524460 41834
rect 524327 41812 524472 41818
rect 524327 41806 524420 41812
rect 524327 41713 524383 41806
rect 524420 41754 524472 41760
rect 525615 41834 525671 42193
rect 525615 41818 525748 41834
rect 525615 41812 525760 41818
rect 525615 41806 525708 41812
rect 525615 41713 525671 41806
rect 525708 41754 525760 41760
rect 526811 41713 526867 42193
rect 528007 41834 528063 42193
rect 528651 41834 528707 42193
rect 527928 41818 528707 41834
rect 527916 41812 528707 41818
rect 527968 41806 528707 41812
rect 527916 41754 527968 41760
rect 528007 41713 528063 41806
rect 528651 41713 528707 41806
rect 529847 41713 529903 42193
rect 295017 41657 295227 41713
rect 295395 41657 295871 41713
rect 296039 41657 296515 41713
rect 296683 41657 297067 41713
rect 297235 41657 297711 41713
rect 297879 41657 298355 41713
rect 298523 41657 298907 41713
rect 299075 41657 299551 41713
rect 299719 41657 300195 41713
rect 300363 41657 300747 41713
rect 300915 41657 301391 41713
rect 301559 41657 302035 41713
rect 302203 41657 302587 41713
rect 302755 41657 303231 41713
rect 303399 41657 303875 41713
rect 304043 41657 304519 41713
rect 304687 41657 305071 41713
rect 305239 41657 305715 41713
rect 305883 41657 306359 41713
rect 306527 41657 306911 41713
rect 307079 41657 307555 41713
rect 307723 41657 308199 41713
rect 308367 41657 308751 41713
rect 308919 41657 309395 41713
rect 309563 41657 310039 41713
rect 310207 41657 310591 41713
rect 310759 41657 310958 41713
rect 252100 39704 252152 39710
rect 252100 39646 252152 39652
rect 254032 39704 254084 39710
rect 254032 39646 254084 39652
rect 252112 39600 252140 39646
rect 241256 39372 245257 39600
rect 241260 38868 245257 39372
rect 245313 39479 247256 39593
rect 247312 39535 249312 39600
rect 249368 39479 252045 39593
rect 245313 39247 252045 39479
rect 252101 39303 256100 39600
rect 245313 38812 256100 39247
rect 241260 714 256100 38812
rect 295017 0 310958 41657
rect 349817 41657 350027 41713
rect 350195 41657 350671 41713
rect 350839 41657 351315 41713
rect 351483 41657 351867 41713
rect 352035 41657 352511 41713
rect 352679 41657 353155 41713
rect 353323 41657 353707 41713
rect 353875 41657 354351 41713
rect 354519 41657 354995 41713
rect 355163 41657 355547 41713
rect 355715 41657 356191 41713
rect 356359 41657 356835 41713
rect 357003 41657 357387 41713
rect 357555 41657 358031 41713
rect 358199 41657 358675 41713
rect 358843 41657 359319 41713
rect 359487 41657 359871 41713
rect 360039 41657 360515 41713
rect 360683 41657 361159 41713
rect 361327 41657 361711 41713
rect 361879 41657 362355 41713
rect 362523 41657 362999 41713
rect 363167 41657 363551 41713
rect 363719 41657 364195 41713
rect 364363 41657 364839 41713
rect 365007 41657 365391 41713
rect 365559 41657 365758 41713
rect 349817 0 365758 41657
rect 404617 41657 404827 41713
rect 404995 41657 405471 41713
rect 405639 41657 406115 41713
rect 406283 41657 406667 41713
rect 406835 41657 407311 41713
rect 407479 41657 407955 41713
rect 408123 41657 408507 41713
rect 408675 41657 409151 41713
rect 409319 41657 409795 41713
rect 409963 41657 410347 41713
rect 410515 41657 410991 41713
rect 411159 41657 411635 41713
rect 411803 41657 412187 41713
rect 412355 41657 412831 41713
rect 412999 41657 413475 41713
rect 413643 41657 414119 41713
rect 414287 41657 414671 41713
rect 414839 41657 415315 41713
rect 415483 41657 415959 41713
rect 416127 41657 416511 41713
rect 416679 41657 417155 41713
rect 417323 41657 417799 41713
rect 417967 41657 418351 41713
rect 418519 41657 418995 41713
rect 419163 41657 419639 41713
rect 419807 41657 420191 41713
rect 420359 41657 420558 41713
rect 404617 0 420558 41657
rect 459417 41657 459627 41713
rect 459795 41657 460271 41713
rect 460439 41657 460915 41713
rect 461083 41657 461467 41713
rect 461635 41657 462111 41713
rect 462279 41657 462755 41713
rect 462923 41657 463307 41713
rect 463475 41657 463951 41713
rect 464119 41657 464595 41713
rect 464763 41657 465147 41713
rect 465315 41657 465791 41713
rect 465959 41657 466435 41713
rect 466603 41657 466987 41713
rect 467155 41657 467631 41713
rect 467799 41657 468275 41713
rect 468443 41657 468919 41713
rect 469087 41657 469471 41713
rect 469639 41657 470115 41713
rect 470283 41657 470759 41713
rect 470927 41657 471311 41713
rect 471479 41657 471955 41713
rect 472123 41657 472599 41713
rect 472767 41657 473151 41713
rect 473319 41657 473795 41713
rect 473963 41657 474439 41713
rect 474607 41657 474991 41713
rect 475159 41657 475358 41713
rect 459417 0 475358 41657
rect 514217 41657 514427 41713
rect 514595 41657 515071 41713
rect 515239 41657 515715 41713
rect 515883 41657 516267 41713
rect 516435 41657 516911 41713
rect 517079 41657 517555 41713
rect 517723 41657 518107 41713
rect 518275 41657 518751 41713
rect 518919 41657 519395 41713
rect 519563 41657 519947 41713
rect 520115 41657 520591 41713
rect 520759 41657 521235 41713
rect 521403 41657 521787 41713
rect 521955 41657 522431 41713
rect 522599 41657 523075 41713
rect 523243 41657 523719 41713
rect 523887 41657 524271 41713
rect 524439 41657 524915 41713
rect 525083 41657 525559 41713
rect 525727 41657 526111 41713
rect 526279 41657 526755 41713
rect 526923 41657 527399 41713
rect 527567 41657 527951 41713
rect 528119 41657 528595 41713
rect 528763 41657 529239 41713
rect 529407 41657 529791 41713
rect 529959 41657 530158 41713
rect 514217 0 530158 41657
rect 569144 40000 569172 47058
rect 634820 46980 634872 46986
rect 634820 46922 634872 46928
rect 579160 45552 579212 45558
rect 579160 45494 579212 45500
rect 569224 44192 569276 44198
rect 569224 44134 569276 44140
rect 569236 40225 569264 44134
rect 579172 40225 579200 45494
rect 622950 40488 623006 40497
rect 622950 40423 623006 40432
rect 569222 40216 569278 40225
rect 569222 40151 569278 40160
rect 579158 40216 579214 40225
rect 579158 40151 579214 40160
rect 579172 40000 579200 40151
rect 622964 40000 622992 40423
rect 634832 40225 634860 46922
rect 673472 45558 673500 112066
rect 673840 102202 673868 121502
rect 675887 115759 717600 115958
rect 675407 115647 675887 115703
rect 675943 115591 717600 115759
rect 675887 115207 717600 115591
rect 675943 115039 717600 115207
rect 675887 114563 717600 115039
rect 675943 114395 717600 114563
rect 675887 113919 717600 114395
rect 675943 113751 717600 113919
rect 675887 113367 717600 113751
rect 675943 113199 717600 113367
rect 675887 112723 717600 113199
rect 675407 112639 675887 112667
rect 675404 112611 675887 112639
rect 675404 112130 675432 112611
rect 675943 112555 717600 112723
rect 675392 112124 675444 112130
rect 675887 112079 717600 112555
rect 675392 112066 675444 112072
rect 675943 111911 717600 112079
rect 675887 111527 717600 111911
rect 675943 111359 717600 111527
rect 675887 110883 717600 111359
rect 675943 110715 717600 110883
rect 675887 110239 717600 110715
rect 675943 110071 717600 110239
rect 675887 109687 717600 110071
rect 675943 109519 717600 109687
rect 675887 109043 717600 109519
rect 675943 108875 717600 109043
rect 675887 108399 717600 108875
rect 675407 108338 675887 108343
rect 675312 108310 675887 108338
rect 673644 102196 673696 102202
rect 673644 102138 673696 102144
rect 673828 102196 673880 102202
rect 673828 102138 673880 102144
rect 673656 102066 673684 102138
rect 673644 102060 673696 102066
rect 673644 102002 673696 102008
rect 673656 47938 673684 102002
rect 675312 100314 675340 108310
rect 675407 108287 675887 108310
rect 675943 108231 717600 108399
rect 675887 107755 717600 108231
rect 675943 107587 717600 107755
rect 675887 107203 717600 107587
rect 675943 107035 717600 107203
rect 675887 106559 717600 107035
rect 675943 106391 717600 106559
rect 675887 105915 717600 106391
rect 675943 105747 717600 105915
rect 675887 105363 717600 105747
rect 675407 105251 675887 105307
rect 675943 105195 717600 105363
rect 675887 104719 717600 105195
rect 675943 104551 717600 104719
rect 675887 104075 717600 104551
rect 675407 103963 675887 104019
rect 675943 103907 717600 104075
rect 675887 103523 717600 103907
rect 675407 103411 675887 103467
rect 675943 103355 717600 103523
rect 675887 102879 717600 103355
rect 675943 102711 717600 102879
rect 675887 102235 717600 102711
rect 675407 102151 675887 102179
rect 675404 102123 675887 102151
rect 675404 102066 675432 102123
rect 675943 102067 717600 102235
rect 675392 102060 675444 102066
rect 675392 102002 675444 102008
rect 675887 101683 717600 102067
rect 675407 101571 675887 101627
rect 675943 101515 717600 101683
rect 675887 101039 717600 101515
rect 675943 100871 717600 101039
rect 675887 100395 717600 100871
rect 675407 100314 675887 100339
rect 675312 100286 675887 100314
rect 675407 100283 675887 100286
rect 675943 100227 717600 100395
rect 675887 100017 717600 100227
rect 673644 47932 673696 47938
rect 673644 47874 673696 47880
rect 673460 45552 673512 45558
rect 673460 45494 673512 45500
rect 632978 40216 633034 40225
rect 632978 40151 633034 40160
rect 634818 40216 634874 40225
rect 634818 40151 634874 40160
rect 632992 40000 633020 40151
rect 569142 34868 573922 40000
rect 573978 39533 579065 39593
rect 579121 39589 583901 40000
rect 622942 39672 627722 40000
rect 622942 39616 622950 39672
rect 623006 39616 627722 39672
rect 573978 34812 583947 39533
rect 622942 34868 627722 39616
rect 627778 39533 632865 39593
rect 632921 39589 637701 40000
rect 627778 34812 637747 39533
rect 569142 985 583947 34812
rect 622942 985 637747 34812
<< metal3 >>
rect 160093 990722 160159 990725
rect 173801 990722 173867 990725
rect 160093 990720 173867 990722
rect 160093 990664 160098 990720
rect 160154 990664 173806 990720
rect 173862 990664 173867 990720
rect 160093 990662 173867 990664
rect 160093 990659 160159 990662
rect 173801 990659 173867 990662
rect 676260 990116 676324 990180
rect 677548 918580 677612 918644
rect 40540 908108 40604 908172
rect 40540 907972 40604 908036
rect 676260 907700 676324 907764
rect 40356 888796 40420 888860
rect 673453 888722 673519 888725
rect 675293 888722 675359 888725
rect 673453 888720 675359 888722
rect 673453 888664 673458 888720
rect 673514 888664 675298 888720
rect 675354 888664 675359 888720
rect 673453 888662 675359 888664
rect 673453 888659 673519 888662
rect 675293 888659 675359 888662
rect 39988 855748 40052 855812
rect 39804 855476 39868 855540
rect 39804 837584 39868 837588
rect 39804 837528 39854 837584
rect 39804 837524 39868 837528
rect 39988 832628 40052 832692
rect 40356 797676 40420 797740
rect 40356 797540 40420 797604
rect 40356 792100 40420 792164
rect 40540 792100 40604 792164
rect 40540 778500 40604 778564
rect 40356 778228 40420 778292
rect 40356 763132 40420 763196
rect 40724 763132 40788 763196
rect 40356 753476 40420 753540
rect 40724 753476 40788 753540
rect 40356 750620 40420 750684
rect 40356 750348 40420 750412
rect 40172 731308 40236 731372
rect 40724 731172 40788 731236
rect 40356 712268 40420 712332
rect 40724 712268 40788 712332
rect 40356 702068 40420 702132
rect 40908 702068 40972 702132
rect 40540 695268 40604 695332
rect 40908 695268 40972 695332
rect 40172 673372 40236 673436
rect 40540 673372 40604 673436
rect 40540 654332 40604 654396
rect 40172 654196 40236 654260
rect 40356 634748 40420 634812
rect 40908 634748 40972 634812
rect 40540 598980 40604 599044
rect 40908 598980 40972 599044
rect 40172 565932 40236 565996
rect 40172 565660 40236 565724
rect 40172 550564 40236 550628
rect 40540 550564 40604 550628
rect 40540 540908 40604 540972
rect 40908 540908 40972 540972
rect 40908 521868 40972 521932
rect 40172 521732 40236 521796
rect 40172 507996 40236 508060
rect 39988 507724 40052 507788
rect 677548 477532 677612 477596
rect 40172 455364 40236 455428
rect 40172 451828 40236 451892
rect 673545 338738 673611 338741
rect 675385 338738 675451 338741
rect 673545 338736 675451 338738
rect 673545 338680 673550 338736
rect 673606 338680 675390 338736
rect 675446 338680 675451 338736
rect 673545 338678 675451 338680
rect 673545 338675 673611 338678
rect 675385 338675 675451 338678
rect 40172 84220 40236 84284
rect 47646 35175 51144 35977
rect 47652 32987 51182 33577
rect 51646 35175 55144 35977
rect 51652 32987 55182 33577
rect 55646 35175 59144 35977
rect 55652 32987 59182 33577
rect 59646 35175 63144 35977
rect 59652 32987 63182 33577
rect 63646 35175 67144 35977
rect 63652 32987 67182 33577
rect 67646 35175 71144 35977
rect 67652 32987 71182 33577
rect 101446 35175 104944 35977
rect 101452 32987 104982 33577
rect 105446 35175 108944 35977
rect 105452 32987 108982 33577
rect 109446 35175 112944 35977
rect 109452 32987 112982 33577
rect 113446 35175 116944 35977
rect 113452 32987 116982 33577
rect 117446 35175 120944 35977
rect 117452 32987 120982 33577
rect 121446 35175 124944 35977
rect 121452 32987 124982 33577
rect 141667 38031 141813 40000
rect 141667 37971 141873 38031
rect 141667 37911 141820 37971
rect 141873 37911 141966 37971
rect 141667 37818 141966 37911
rect 141820 37046 141966 37818
rect 155246 35175 158744 35977
rect 155252 32987 158782 33577
rect 159246 35175 162744 35977
rect 159252 32987 162782 33577
rect 163246 35175 166744 35977
rect 163252 32987 166782 33577
rect 167246 35175 170744 35977
rect 167252 32987 170782 33577
rect 171246 35175 174744 35977
rect 171252 32987 174782 33577
rect 175246 35175 178744 35977
rect 175252 32987 178782 33577
rect 210046 35175 213544 35977
rect 210052 32987 213582 33577
rect 214046 35175 217544 35977
rect 214052 32987 217582 33577
rect 218046 35175 221544 35977
rect 218052 32987 221582 33577
rect 222046 35175 225544 35977
rect 222052 32987 225582 33577
rect 226046 35175 229544 35977
rect 226052 32987 229582 33577
rect 230046 35175 233544 35977
rect 230052 32987 233582 33577
rect 263846 35175 267344 35977
rect 263852 32987 267382 33577
rect 267846 35175 271344 35977
rect 267852 32987 271382 33577
rect 271846 35175 275344 35977
rect 271852 32987 275382 33577
rect 275846 35175 279344 35977
rect 275852 32987 279382 33577
rect 279846 35175 283344 35977
rect 279852 32987 283382 33577
rect 283846 35175 287344 35977
rect 283852 32987 287382 33577
rect 318646 35175 322144 35977
rect 318652 32987 322182 33577
rect 322646 35175 326144 35977
rect 322652 32987 326182 33577
rect 326646 35175 330144 35977
rect 326652 32987 330182 33577
rect 330646 35175 334144 35977
rect 330652 32987 334182 33577
rect 334646 35175 338144 35977
rect 334652 32987 338182 33577
rect 338646 35175 342144 35977
rect 338652 32987 342182 33577
rect 373446 35175 376944 35977
rect 373452 32987 376982 33577
rect 377446 35175 380944 35977
rect 377452 32987 380982 33577
rect 381446 35175 384944 35977
rect 381452 32987 384982 33577
rect 385446 35175 388944 35977
rect 385452 32987 388982 33577
rect 389446 35175 392944 35977
rect 389452 32987 392982 33577
rect 393446 35175 396944 35977
rect 393452 32987 396982 33577
rect 428246 35175 431744 35977
rect 428252 32987 431782 33577
rect 432246 35175 435744 35977
rect 432252 32987 435782 33577
rect 436246 35175 439744 35977
rect 436252 32987 439782 33577
rect 440246 35175 443744 35977
rect 440252 32987 443782 33577
rect 444246 35175 447744 35977
rect 444252 32987 447782 33577
rect 448246 35175 451744 35977
rect 448252 32987 451782 33577
rect 483046 35175 486544 35977
rect 483052 32987 486582 33577
rect 487046 35175 490544 35977
rect 487052 32987 490582 33577
rect 491046 35175 494544 35977
rect 491052 32987 494582 33577
rect 495046 35175 498544 35977
rect 495052 32987 498582 33577
rect 499046 35175 502544 35977
rect 499052 32987 502582 33577
rect 503046 35175 506544 35977
rect 503052 32987 506582 33577
rect 537846 35175 541344 35977
rect 537852 32987 541382 33577
rect 541846 35175 545344 35977
rect 541852 32987 545382 33577
rect 545846 35175 549344 35977
rect 545852 32987 549382 33577
rect 549846 35175 553344 35977
rect 549852 32987 553382 33577
rect 553846 35175 557344 35977
rect 553852 32987 557382 33577
rect 557846 35175 561344 35977
rect 591646 35175 595144 35977
rect 557852 32987 561382 33577
rect 591652 32987 595182 33577
rect 595646 35175 599144 35977
rect 595652 32987 599182 33577
rect 599646 35175 603144 35977
rect 599652 32987 603182 33577
rect 603646 35175 607144 35977
rect 603652 32987 607182 33577
rect 607646 35175 611144 35977
rect 607652 32987 611182 33577
rect 611646 35175 615144 35977
rect 611652 32987 615182 33577
rect 645446 35175 648944 35977
rect 645452 32987 648982 33577
rect 649446 35175 652944 35977
rect 649452 32987 652982 33577
rect 653446 35175 656944 35977
rect 653452 32987 656982 33577
rect 657446 35175 660944 35977
rect 657452 32987 660982 33577
rect 661446 35175 664944 35977
rect 661452 32987 664982 33577
rect 665446 35175 668944 35977
rect 665452 32987 668982 33577
<< obsm3 >>
rect 76262 997338 92114 1037600
rect 127662 997338 143514 1037600
rect 179062 997338 194914 1037600
rect 230462 997338 246314 1037600
rect 282062 997338 297914 1037600
rect 333448 1002850 348258 1037600
rect 333499 997656 338279 1002770
rect 338359 1000165 343398 1002850
rect 338359 1000076 338499 1000165
rect 340859 1000156 343398 1000165
rect 333499 997600 333518 997656
rect 333574 997600 338279 997656
rect 338579 997600 340779 1000085
rect 340859 1000076 340898 1000156
rect 343258 1000076 343398 1000156
rect 340978 997600 343178 1000076
rect 343478 997600 348258 1002770
rect 333500 997598 333579 997600
rect 333513 997595 333579 997598
rect 45921 996570 45987 996573
rect 341014 996570 341074 997600
rect 383862 997338 399714 1037600
rect 472862 997338 488714 1037600
rect 524262 997338 540114 1037600
rect 575648 1005032 590458 1036620
rect 575648 1004183 585598 1005032
rect 575699 997600 580479 1004103
rect 580559 1000165 585598 1004183
rect 580559 1000076 580699 1000165
rect 583059 1000156 585598 1000165
rect 580779 997600 582979 1000085
rect 583059 1000076 583098 1000156
rect 585458 1000076 585598 1000156
rect 583178 997600 585378 1000076
rect 585678 997600 590458 1004952
rect 580796 997598 581746 997600
rect 581686 997522 581746 997598
rect 585734 997522 585794 997600
rect 581686 997462 585794 997522
rect 585734 997114 585794 997462
rect 626062 997338 641914 1037600
rect 585734 997054 585978 997114
rect 45921 996568 341074 996570
rect 45921 996512 45926 996568
rect 45982 996512 341074 996568
rect 45921 996510 341074 996512
rect 585918 996570 585978 997054
rect 672625 996570 672691 996573
rect 585918 996568 672691 996570
rect 585918 996512 672630 996568
rect 672686 996512 672691 996568
rect 585918 996510 672691 996512
rect 45921 996507 45987 996510
rect 672625 996507 672691 996510
rect 585685 996434 585751 996437
rect 672441 996434 672507 996437
rect 585685 996432 672507 996434
rect 585685 996376 585690 996432
rect 585746 996376 672446 996432
rect 672502 996376 672507 996432
rect 585685 996374 672507 996376
rect 585685 996371 585751 996374
rect 672441 996371 672507 996374
rect 537845 995482 537911 995485
rect 538029 995482 538095 995485
rect 537845 995480 538095 995482
rect 537845 995424 537850 995480
rect 537906 995424 538034 995480
rect 538090 995424 538095 995480
rect 537845 995422 538095 995424
rect 537845 995419 537911 995422
rect 538029 995419 538095 995422
rect 193213 990586 193279 990589
rect 212441 990586 212507 990589
rect 193213 990584 212507 990586
rect 193213 990528 193218 990584
rect 193274 990528 212446 990584
rect 212502 990528 212507 990584
rect 193213 990526 212507 990528
rect 193213 990523 193279 990526
rect 212441 990523 212507 990526
rect 576853 990586 576919 990589
rect 596081 990586 596147 990589
rect 576853 990584 596147 990586
rect 576853 990528 576858 990584
rect 576914 990528 596086 990584
rect 596142 990528 596147 990584
rect 576853 990526 596147 990528
rect 576853 990523 576919 990526
rect 596081 990523 596147 990526
rect 540973 990450 541039 990453
rect 560201 990450 560267 990453
rect 540973 990448 560267 990450
rect 540973 990392 540978 990448
rect 541034 990392 560206 990448
rect 560262 990392 560267 990448
rect 540973 990390 560267 990392
rect 540973 990387 541039 990390
rect 560201 990387 560267 990390
rect 45461 990178 45527 990181
rect 676254 990178 676260 990180
rect 45461 990176 676260 990178
rect 45461 990120 45466 990176
rect 45522 990120 676260 990176
rect 45461 990118 676260 990120
rect 45461 990115 45527 990118
rect 676254 990116 676260 990118
rect 676324 990116 676330 990180
rect 0 954262 40262 970114
rect 677338 951686 717600 967538
rect 1697 922071 38140 926940
rect 38220 922314 39600 926940
rect 38220 922254 39866 922314
rect 38220 922151 39600 922254
rect 1697 921931 39593 922071
rect 1697 919596 34940 921931
rect 35020 921770 39600 921851
rect 39806 921770 39866 922254
rect 35020 921710 39866 921770
rect 35020 919730 39600 921710
rect 35020 919676 39866 919730
rect 39468 919670 39866 919676
rect 1697 919456 39593 919596
rect 1697 917120 35476 919456
rect 35556 919322 39600 919376
rect 39806 919322 39866 919670
rect 35556 919262 39866 919322
rect 35556 917282 39600 919262
rect 677542 918580 677548 918644
rect 677612 918642 677618 918644
rect 677869 918642 677935 918645
rect 677612 918640 677935 918642
rect 677612 918584 677874 918640
rect 677930 918584 677935 918640
rect 677612 918582 677935 918584
rect 677612 918580 677618 918582
rect 677869 918579 677935 918582
rect 678000 917700 679380 922500
rect 679460 917620 715903 922502
rect 678007 917480 715903 917620
rect 44357 917282 44423 917285
rect 35556 917280 44423 917282
rect 35556 917224 44362 917280
rect 44418 917224 44423 917280
rect 35556 917222 44423 917224
rect 35556 917200 39600 917222
rect 44357 917219 44423 917222
rect 1697 916980 39593 917120
rect 1697 912098 38140 916980
rect 38220 912100 39600 916900
rect 677593 915378 677659 915381
rect 678000 915378 682044 917400
rect 677593 915376 682044 915378
rect 677593 915320 677598 915376
rect 677654 915320 682044 915376
rect 677593 915318 682044 915320
rect 677593 915315 677659 915318
rect 678000 915224 682044 915318
rect 682124 915144 715903 917480
rect 678007 915004 715903 915144
rect 677593 912794 677659 912797
rect 677869 912794 677935 912797
rect 678000 912794 682580 914924
rect 677593 912792 682580 912794
rect 677593 912736 677598 912792
rect 677654 912736 677874 912792
rect 677930 912749 682580 912792
rect 677930 912736 678132 912749
rect 677593 912734 678132 912736
rect 677593 912731 677659 912734
rect 677869 912731 677935 912734
rect 682660 912669 715903 915004
rect 678007 912529 715903 912669
rect 39665 908170 39731 908173
rect 40534 908170 40540 908172
rect 39665 908168 40540 908170
rect 39665 908112 39670 908168
rect 39726 908112 40540 908168
rect 39665 908110 40540 908112
rect 39665 908107 39731 908110
rect 40534 908108 40540 908110
rect 40604 908108 40610 908172
rect 673361 908170 673427 908173
rect 677869 908170 677935 908173
rect 678000 908170 679380 912449
rect 673361 908168 679380 908170
rect 673361 908112 673366 908168
rect 673422 908112 677874 908168
rect 677930 908112 679380 908168
rect 673361 908110 679380 908112
rect 673361 908107 673427 908110
rect 677869 908107 677935 908110
rect 40401 908034 40467 908037
rect 40534 908034 40540 908036
rect 40401 908032 40540 908034
rect 40401 907976 40406 908032
rect 40462 907976 40540 908032
rect 40401 907974 40540 907976
rect 40401 907971 40467 907974
rect 40534 907972 40540 907974
rect 40604 907972 40610 908036
rect 676254 907700 676260 907764
rect 676324 907762 676330 907764
rect 677777 907762 677843 907765
rect 676324 907760 677843 907762
rect 676324 907704 677782 907760
rect 677838 907704 677843 907760
rect 676324 907702 677843 907704
rect 676324 907700 676330 907702
rect 677777 907699 677843 907702
rect 678000 907660 679380 908110
rect 679460 907660 715903 912529
rect 40401 888994 40467 888997
rect 40358 888992 40467 888994
rect 40358 888936 40406 888992
rect 40462 888936 40467 888992
rect 40358 888931 40467 888936
rect 40358 888860 40418 888931
rect 40350 888796 40356 888860
rect 40420 888796 40426 888860
rect 0 879798 35960 884658
rect 36040 880018 40000 884658
rect 40125 880018 40191 880021
rect 36040 880016 40191 880018
rect 36040 879960 40130 880016
rect 40186 879960 40191 880016
rect 36040 879958 40191 879960
rect 36040 879878 40000 879958
rect 40125 879955 40191 879958
rect 0 879658 39455 879798
rect 0 877298 37654 879658
rect 37734 877378 40000 879578
rect 0 877259 39455 877298
rect 0 874899 39375 877259
rect 39455 875122 40000 877179
rect 41413 875122 41479 875125
rect 39455 875120 41479 875122
rect 39455 875064 41418 875120
rect 41474 875064 41479 875120
rect 39455 875062 41479 875064
rect 39455 874979 40000 875062
rect 41413 875059 41479 875062
rect 0 874759 39455 874899
rect 0 869848 35960 874759
rect 36040 869899 40000 874679
rect 677338 862486 717600 878338
rect 39982 855810 39988 855812
rect 39806 855750 39988 855810
rect 39806 855540 39866 855750
rect 39982 855748 39988 855750
rect 40052 855748 40058 855812
rect 39798 855476 39804 855540
rect 39868 855476 39874 855540
rect 980 837598 32568 842458
rect 32648 837678 40000 842458
rect 980 837458 37524 837598
rect 39849 837588 39915 837589
rect 39798 837586 39804 837588
rect 39758 837526 39804 837586
rect 39868 837584 39915 837588
rect 39910 837528 39915 837584
rect 39798 837524 39804 837526
rect 39868 837524 39915 837528
rect 39849 837523 39915 837524
rect 980 835098 37444 837458
rect 37524 835274 40000 837378
rect 44449 835274 44515 835277
rect 37524 835272 44515 835274
rect 37524 835216 44454 835272
rect 44510 835216 44515 835272
rect 37524 835214 44515 835216
rect 37524 835178 40000 835214
rect 44449 835211 44515 835214
rect 980 835059 37524 835098
rect 980 832699 37435 835059
rect 37515 832779 40000 834979
rect 980 832559 37524 832699
rect 39849 832690 39915 832693
rect 39982 832690 39988 832692
rect 39849 832688 39988 832690
rect 39849 832632 39854 832688
rect 39910 832632 39988 832688
rect 39849 832630 39988 832632
rect 39849 832627 39915 832630
rect 39982 832628 39988 832630
rect 40052 832628 40058 832692
rect 980 827648 33417 832559
rect 33497 828066 40000 832479
rect 672533 828746 672599 828749
rect 676121 828746 676187 828749
rect 677600 828746 680592 833301
rect 672533 828744 680592 828746
rect 672533 828688 672538 828744
rect 672594 828688 676126 828744
rect 676182 828688 680592 828744
rect 672533 828686 680592 828688
rect 672533 828683 672599 828686
rect 676121 828683 676187 828686
rect 677600 828521 680592 828686
rect 680672 828441 717600 833352
rect 678145 828301 717600 828441
rect 44725 828066 44791 828069
rect 33497 828064 44791 828066
rect 33497 828008 44730 828064
rect 44786 828008 44791 828064
rect 33497 828006 44791 828008
rect 33497 827699 40000 828006
rect 44725 828003 44791 828006
rect 39665 827522 39731 827525
rect 39806 827522 39866 827699
rect 39665 827520 39866 827522
rect 39665 827464 39670 827520
rect 39726 827464 39866 827520
rect 39665 827462 39866 827464
rect 39665 827459 39731 827462
rect 672625 826162 672691 826165
rect 673269 826162 673335 826165
rect 677600 826162 678145 828221
rect 672625 826160 678145 826162
rect 672625 826104 672630 826160
rect 672686 826104 673274 826160
rect 673330 826104 678145 826160
rect 672625 826102 678145 826104
rect 672625 826099 672691 826102
rect 673269 826099 673335 826102
rect 677600 826021 678145 826102
rect 678225 825941 717600 828301
rect 678145 825902 717600 825941
rect 673177 823714 673243 823717
rect 676121 823714 676187 823717
rect 677600 823714 679866 825822
rect 673177 823712 679866 823714
rect 673177 823656 673182 823712
rect 673238 823656 676126 823712
rect 676182 823656 679866 823712
rect 673177 823654 679866 823656
rect 673177 823651 673243 823654
rect 676121 823651 676187 823654
rect 677600 823622 679866 823654
rect 679946 823542 717600 825902
rect 678145 823402 717600 823542
rect 677600 818542 680592 823322
rect 680672 818469 717600 823402
rect 0 784462 40262 800314
rect 40350 797676 40356 797740
rect 40420 797676 40426 797740
rect 40358 797604 40418 797676
rect 40350 797540 40356 797604
rect 40420 797540 40426 797604
rect 40350 792100 40356 792164
rect 40420 792162 40426 792164
rect 40534 792162 40540 792164
rect 40420 792102 40540 792162
rect 40420 792100 40426 792102
rect 40534 792100 40540 792102
rect 40604 792100 40610 792164
rect 672993 792162 673059 792165
rect 673177 792162 673243 792165
rect 672993 792160 673243 792162
rect 672993 792104 672998 792160
rect 673054 792104 673182 792160
rect 673238 792104 673243 792160
rect 672993 792102 673243 792104
rect 672993 792099 673059 792102
rect 673177 792099 673243 792102
rect 40534 778562 40540 778564
rect 40358 778502 40540 778562
rect 40358 778292 40418 778502
rect 40534 778500 40540 778502
rect 40604 778500 40610 778564
rect 40350 778228 40356 778292
rect 40420 778228 40426 778292
rect 677338 773286 717600 789138
rect 40350 763132 40356 763196
rect 40420 763194 40426 763196
rect 40718 763194 40724 763196
rect 40420 763134 40724 763194
rect 40420 763132 40426 763134
rect 40718 763132 40724 763134
rect 40788 763132 40794 763196
rect 0 741262 40262 757114
rect 40350 753476 40356 753540
rect 40420 753538 40426 753540
rect 40718 753538 40724 753540
rect 40420 753478 40724 753538
rect 40420 753476 40426 753478
rect 40718 753476 40724 753478
rect 40788 753476 40794 753540
rect 672809 753538 672875 753541
rect 672993 753538 673059 753541
rect 672809 753536 673059 753538
rect 672809 753480 672814 753536
rect 672870 753480 672998 753536
rect 673054 753480 673059 753536
rect 672809 753478 673059 753480
rect 672809 753475 672875 753478
rect 672993 753475 673059 753478
rect 40350 750620 40356 750684
rect 40420 750682 40426 750684
rect 40420 750622 40602 750682
rect 40420 750620 40426 750622
rect 40350 750348 40356 750412
rect 40420 750410 40426 750412
rect 40542 750410 40602 750622
rect 40420 750350 40602 750410
rect 40420 750348 40426 750350
rect 40166 731308 40172 731372
rect 40236 731308 40242 731372
rect 40174 731234 40234 731308
rect 40718 731234 40724 731236
rect 40174 731174 40724 731234
rect 40718 731172 40724 731174
rect 40788 731172 40794 731236
rect 677338 728286 717600 744138
rect 0 698062 40262 713914
rect 40350 712268 40356 712332
rect 40420 712330 40426 712332
rect 40718 712330 40724 712332
rect 40420 712270 40724 712330
rect 40420 712268 40426 712270
rect 40718 712268 40724 712270
rect 40788 712268 40794 712332
rect 40350 702068 40356 702132
rect 40420 702130 40426 702132
rect 40902 702130 40908 702132
rect 40420 702070 40908 702130
rect 40420 702068 40426 702070
rect 40902 702068 40908 702070
rect 40972 702068 40978 702132
rect 40534 695268 40540 695332
rect 40604 695330 40610 695332
rect 40902 695330 40908 695332
rect 40604 695270 40908 695330
rect 40604 695268 40610 695270
rect 40902 695268 40908 695270
rect 40972 695268 40978 695332
rect 673453 685402 673519 685405
rect 675385 685402 675451 685405
rect 673453 685400 675451 685402
rect 673453 685344 673458 685400
rect 673514 685344 675390 685400
rect 675446 685344 675451 685400
rect 673453 685342 675451 685344
rect 673453 685339 673519 685342
rect 675385 685339 675451 685342
rect 677338 683286 717600 699138
rect 40166 673372 40172 673436
rect 40236 673434 40242 673436
rect 40534 673434 40540 673436
rect 40236 673374 40540 673434
rect 40236 673372 40242 673374
rect 40534 673372 40540 673374
rect 40604 673372 40610 673436
rect 0 654862 40262 670714
rect 40534 654394 40540 654396
rect 40174 654334 40540 654394
rect 40174 654260 40234 654334
rect 40534 654332 40540 654334
rect 40604 654332 40610 654396
rect 40166 654196 40172 654260
rect 40236 654196 40242 654260
rect 677338 638086 717600 653938
rect 40350 634748 40356 634812
rect 40420 634810 40426 634812
rect 40902 634810 40908 634812
rect 40420 634750 40908 634810
rect 40420 634748 40426 634750
rect 40902 634748 40908 634750
rect 40972 634748 40978 634812
rect 0 611662 40262 627514
rect 672993 618218 673059 618221
rect 672993 618216 673194 618218
rect 672993 618160 672998 618216
rect 673054 618160 673194 618216
rect 672993 618158 673194 618160
rect 672993 618155 673059 618158
rect 672809 618082 672875 618085
rect 673134 618082 673194 618158
rect 672809 618080 673194 618082
rect 672809 618024 672814 618080
rect 672870 618024 673194 618080
rect 672809 618022 673194 618024
rect 672809 618019 672875 618022
rect 40534 598980 40540 599044
rect 40604 599042 40610 599044
rect 40902 599042 40908 599044
rect 40604 598982 40908 599042
rect 40604 598980 40610 598982
rect 40902 598980 40908 598982
rect 40972 598980 40978 599044
rect 677338 593086 717600 608938
rect 0 568462 40262 584314
rect 40166 565932 40172 565996
rect 40236 565932 40242 565996
rect 40174 565724 40234 565932
rect 40166 565660 40172 565724
rect 40236 565660 40242 565724
rect 44541 560282 44607 560285
rect 44909 560282 44975 560285
rect 44541 560280 44975 560282
rect 44541 560224 44546 560280
rect 44602 560224 44914 560280
rect 44970 560224 44975 560280
rect 44541 560222 44975 560224
rect 44541 560219 44607 560222
rect 44909 560219 44975 560222
rect 40166 550564 40172 550628
rect 40236 550626 40242 550628
rect 40534 550626 40540 550628
rect 40236 550566 40540 550626
rect 40236 550564 40242 550566
rect 40534 550564 40540 550566
rect 40604 550564 40610 550628
rect 677338 547886 717600 563738
rect 0 525262 40262 541114
rect 40534 540908 40540 540972
rect 40604 540970 40610 540972
rect 40902 540970 40908 540972
rect 40604 540910 40908 540970
rect 40604 540908 40610 540910
rect 40902 540908 40908 540910
rect 40972 540908 40978 540972
rect 40902 521930 40908 521932
rect 40174 521870 40908 521930
rect 40174 521796 40234 521870
rect 40902 521868 40908 521870
rect 40972 521868 40978 521932
rect 40166 521732 40172 521796
rect 40236 521732 40242 521796
rect 676121 514178 676187 514181
rect 677600 514178 680592 518701
rect 676121 514176 680592 514178
rect 676121 514120 676126 514176
rect 676182 514120 680592 514176
rect 676121 514118 680592 514120
rect 676121 514115 676187 514118
rect 677600 513921 680592 514118
rect 680672 513841 717600 518752
rect 678145 513701 717600 513841
rect 673085 511458 673151 511461
rect 673269 511458 673335 511461
rect 677600 511458 678145 513621
rect 673085 511456 678145 511458
rect 673085 511400 673090 511456
rect 673146 511400 673274 511456
rect 673330 511421 678145 511456
rect 673330 511400 677764 511421
rect 673085 511398 677764 511400
rect 673085 511395 673151 511398
rect 673269 511395 673335 511398
rect 678225 511341 717600 513701
rect 678145 511302 717600 511341
rect 672993 509146 673059 509149
rect 676121 509146 676187 509149
rect 677600 509146 679866 511222
rect 672993 509144 679866 509146
rect 672993 509088 672998 509144
rect 673054 509088 676126 509144
rect 676182 509088 679866 509144
rect 672993 509086 679866 509088
rect 672993 509083 673059 509086
rect 676121 509083 676187 509086
rect 677600 509022 679866 509086
rect 679946 508942 717600 511302
rect 678145 508802 717600 508942
rect 40166 508058 40172 508060
rect 39990 507998 40172 508058
rect 39990 507788 40050 507998
rect 40166 507996 40172 507998
rect 40236 507996 40242 508060
rect 39982 507724 39988 507788
rect 40052 507724 40058 507788
rect 677600 503942 680592 508722
rect 680672 503869 717600 508802
rect 673269 502346 673335 502349
rect 673637 502346 673703 502349
rect 673269 502344 673703 502346
rect 673269 502288 673274 502344
rect 673330 502288 673642 502344
rect 673698 502288 673703 502344
rect 673269 502286 673703 502288
rect 673269 502283 673335 502286
rect 673637 502283 673703 502286
rect 0 492998 36928 497931
rect 37008 493234 40000 497858
rect 44449 493234 44515 493237
rect 37008 493232 44515 493234
rect 37008 493176 44454 493232
rect 44510 493176 44515 493232
rect 37008 493174 44515 493176
rect 37008 493078 40000 493174
rect 44449 493171 44515 493174
rect 0 492858 39455 492998
rect 39806 492965 39866 493078
rect 39757 492960 39866 492965
rect 39757 492904 39762 492960
rect 39818 492904 39866 492960
rect 39757 492902 39866 492904
rect 39757 492899 39823 492902
rect 0 490498 37654 492858
rect 37734 490578 40000 492778
rect 0 490459 39455 490498
rect 0 488099 39375 490459
rect 39455 488610 40000 490379
rect 44541 488610 44607 488613
rect 39455 488608 44607 488610
rect 39455 488552 44546 488608
rect 44602 488552 44607 488608
rect 39455 488550 44607 488552
rect 39455 488179 40000 488550
rect 44541 488547 44607 488550
rect 0 487959 39455 488099
rect 0 483048 36928 487959
rect 37008 483099 40000 487879
rect 673361 483170 673427 483173
rect 673318 483168 673427 483170
rect 673318 483112 673366 483168
rect 673422 483112 673427 483168
rect 673318 483107 673427 483112
rect 673318 483037 673378 483107
rect 673318 483032 673427 483037
rect 673318 482976 673366 483032
rect 673422 482976 673427 483032
rect 673318 482974 673427 482976
rect 673361 482971 673427 482974
rect 677542 477532 677548 477596
rect 677612 477594 677618 477596
rect 678053 477594 678119 477597
rect 677612 477592 678119 477594
rect 677612 477536 678058 477592
rect 678114 477536 678119 477592
rect 677612 477534 678119 477536
rect 677612 477532 677618 477534
rect 678053 477531 678119 477534
rect 677869 469978 677935 469981
rect 678000 469978 685920 474700
rect 677869 469976 685920 469978
rect 677869 469920 677874 469976
rect 677930 469920 685920 469976
rect 677869 469918 685920 469920
rect 677869 469915 677935 469918
rect 678000 469900 685920 469918
rect 686000 469820 715903 474700
rect 681558 469680 715903 469820
rect 673361 467530 673427 467533
rect 678000 467530 682044 469600
rect 673361 467528 682044 467530
rect 673361 467472 673366 467528
rect 673422 467472 682044 467528
rect 673361 467470 682044 467472
rect 673361 467467 673427 467470
rect 678000 467424 682044 467470
rect 678102 467124 678162 467424
rect 682124 467344 715903 469680
rect 681558 467204 715903 467344
rect 678000 464949 682580 467124
rect 682660 464869 715903 467204
rect 681558 464729 715903 464869
rect 673269 463722 673335 463725
rect 673453 463722 673519 463725
rect 673269 463720 673519 463722
rect 673269 463664 673274 463720
rect 673330 463664 673458 463720
rect 673514 463664 673519 463720
rect 673269 463662 673519 463664
rect 673269 463659 673335 463662
rect 673453 463659 673519 463662
rect 673453 463586 673519 463589
rect 673729 463586 673795 463589
rect 673453 463584 673795 463586
rect 673453 463528 673458 463584
rect 673514 463528 673734 463584
rect 673790 463528 673795 463584
rect 673453 463526 673795 463528
rect 673453 463523 673519 463526
rect 673729 463523 673795 463526
rect 678000 459860 685920 464649
rect 686000 459860 715903 464729
rect 1697 450871 31600 455740
rect 31680 450951 39600 455740
rect 39941 455426 40007 455429
rect 40166 455426 40172 455428
rect 39941 455424 40172 455426
rect 39941 455368 39946 455424
rect 40002 455368 40172 455424
rect 39941 455366 40172 455368
rect 39941 455363 40007 455366
rect 40166 455364 40172 455366
rect 40236 455364 40242 455428
rect 39665 451890 39731 451893
rect 40166 451890 40172 451892
rect 39665 451888 40172 451890
rect 39665 451832 39670 451888
rect 39726 451832 40172 451888
rect 39665 451830 40172 451832
rect 39665 451827 39731 451830
rect 40166 451828 40172 451830
rect 40236 451828 40242 451892
rect 1697 450731 36042 450871
rect 1697 448396 34940 450731
rect 35020 448626 39600 450651
rect 44357 448626 44423 448629
rect 35020 448624 44423 448626
rect 35020 448568 44362 448624
rect 44418 448568 44423 448624
rect 35020 448566 44423 448568
rect 35020 448476 39600 448566
rect 44357 448563 44423 448566
rect 1697 448256 36042 448396
rect 1697 445920 35476 448256
rect 39438 448176 39498 448476
rect 35556 446000 39600 448176
rect 1697 445780 36042 445920
rect 1697 440900 31600 445780
rect 31680 441010 39600 445700
rect 673545 444410 673611 444413
rect 673729 444410 673795 444413
rect 673545 444408 673795 444410
rect 673545 444352 673550 444408
rect 673606 444352 673734 444408
rect 673790 444352 673795 444408
rect 673545 444350 673795 444352
rect 673545 444347 673611 444350
rect 673729 444347 673795 444350
rect 39665 441010 39731 441013
rect 31680 441008 39731 441010
rect 31680 440952 39670 441008
rect 39726 440952 39731 441008
rect 31680 440950 39731 440952
rect 31680 440900 39600 440950
rect 39665 440947 39731 440950
rect 673085 427954 673151 427957
rect 677409 427954 677475 427957
rect 673085 427952 677475 427954
rect 673085 427896 673090 427952
rect 673146 427896 677414 427952
rect 677470 427896 677475 427952
rect 673085 427894 677475 427896
rect 673085 427891 673151 427894
rect 677409 427891 677475 427894
rect 677600 425781 684103 430501
rect 677593 425776 684103 425781
rect 677593 425720 677598 425776
rect 677654 425721 684103 425776
rect 677654 425720 677764 425721
rect 677593 425718 677764 425720
rect 677593 425715 677659 425718
rect 684183 425641 716620 430552
rect 680076 425501 716620 425641
rect 677600 423221 680085 425421
rect 680165 423141 716620 425501
rect 680076 423102 716620 423141
rect 673361 420882 673427 420885
rect 677600 420882 680076 423022
rect 673361 420880 680076 420882
rect 673361 420824 673366 420880
rect 673422 420824 680076 420880
rect 673361 420822 680076 420824
rect 673361 420819 673427 420822
rect 680156 420742 716620 423102
rect 680076 420602 716620 420742
rect 677600 415742 684952 420522
rect 685032 415742 716620 420602
rect 0 397662 40262 413514
rect 42241 400210 42307 400213
rect 42609 400210 42675 400213
rect 42241 400208 42675 400210
rect 42241 400152 42246 400208
rect 42302 400152 42614 400208
rect 42670 400152 42675 400208
rect 42241 400150 42675 400152
rect 42241 400147 42307 400150
rect 42609 400147 42675 400150
rect 677338 370686 717600 386538
rect 0 354462 40262 370314
rect 0 311262 40262 327114
rect 677338 325486 717600 341338
rect 672533 314802 672599 314805
rect 672533 314800 672642 314802
rect 672533 314744 672538 314800
rect 672594 314744 672642 314800
rect 672533 314739 672642 314744
rect 672582 314533 672642 314739
rect 672533 314528 672642 314533
rect 672533 314472 672538 314528
rect 672594 314472 672642 314528
rect 672533 314470 672642 314472
rect 672533 314467 672599 314470
rect 675017 293042 675083 293045
rect 675201 293042 675267 293045
rect 675385 293042 675451 293045
rect 675017 293040 675451 293042
rect 675017 292984 675022 293040
rect 675078 292984 675206 293040
rect 675262 292984 675390 293040
rect 675446 292984 675451 293040
rect 675017 292982 675451 292984
rect 675017 292979 675083 292982
rect 675201 292979 675267 292982
rect 675385 292979 675451 292982
rect 0 268062 40262 283914
rect 677338 280486 717600 296338
rect 0 224862 40262 240714
rect 677338 235486 717600 251338
rect 672533 231842 672599 231845
rect 672901 231842 672967 231845
rect 672533 231840 672967 231842
rect 672533 231784 672538 231840
rect 672594 231784 672906 231840
rect 672962 231784 672967 231840
rect 672533 231782 672967 231784
rect 672533 231779 672599 231782
rect 672901 231779 672967 231782
rect 0 181662 40262 197514
rect 44449 193218 44515 193221
rect 44633 193218 44699 193221
rect 44449 193216 44699 193218
rect 44449 193160 44454 193216
rect 44510 193160 44638 193216
rect 44694 193160 44699 193216
rect 44449 193158 44699 193160
rect 44449 193155 44515 193158
rect 44633 193155 44699 193158
rect 672533 193218 672599 193221
rect 672901 193218 672967 193221
rect 672533 193216 672967 193218
rect 672533 193160 672538 193216
rect 672594 193160 672906 193216
rect 672962 193160 672967 193216
rect 672533 193158 672967 193160
rect 672533 193155 672599 193158
rect 672901 193155 672967 193158
rect 673729 192402 673795 192405
rect 675385 192402 675451 192405
rect 673729 192400 675451 192402
rect 673729 192344 673734 192400
rect 673790 192344 675390 192400
rect 675446 192344 675451 192400
rect 673729 192342 675451 192344
rect 673729 192339 673795 192342
rect 675385 192339 675451 192342
rect 677338 190286 717600 206138
rect 677338 145286 717600 161138
rect 0 120198 35960 125058
rect 36040 120278 40000 125058
rect 0 120058 39455 120198
rect 39757 120186 39823 120189
rect 44173 120186 44239 120189
rect 39757 120184 44239 120186
rect 39757 120128 39762 120184
rect 39818 120128 44178 120184
rect 44234 120128 44239 120184
rect 39757 120126 44239 120128
rect 39757 120123 39823 120126
rect 44173 120123 44239 120126
rect 0 117698 37654 120058
rect 37734 117778 40000 119978
rect 0 117659 39455 117698
rect 0 115299 39375 117659
rect 39455 115970 40000 117579
rect 41413 115970 41479 115973
rect 42333 115970 42399 115973
rect 39455 115968 42399 115970
rect 39455 115912 41418 115968
rect 41474 115912 42338 115968
rect 42394 115912 42399 115968
rect 39455 115910 42399 115912
rect 39455 115379 40000 115910
rect 41413 115907 41479 115910
rect 42333 115907 42399 115910
rect 0 115159 39455 115299
rect 0 110248 35960 115159
rect 36040 110530 40000 115079
rect 44173 110530 44239 110533
rect 45461 110530 45527 110533
rect 36040 110528 45527 110530
rect 36040 110472 44178 110528
rect 44234 110472 45466 110528
rect 45522 110472 45527 110528
rect 36040 110470 45527 110472
rect 36040 110299 40000 110470
rect 44173 110467 44239 110470
rect 45461 110467 45527 110470
rect 677338 100086 717600 115938
rect 39389 84282 39455 84285
rect 40166 84282 40172 84284
rect 39389 84280 40172 84282
rect 39389 84224 39394 84280
rect 39450 84224 40172 84280
rect 39389 84222 40172 84224
rect 39389 84219 39455 84222
rect 40166 84220 40172 84222
rect 40236 84220 40242 84284
rect 1697 78071 38140 82940
rect 38220 78151 39600 82940
rect 1697 77931 39593 78071
rect 1697 75596 34940 77931
rect 35020 75850 39600 77851
rect 44265 75850 44331 75853
rect 35020 75848 44331 75850
rect 35020 75792 44270 75848
rect 44326 75792 44331 75848
rect 35020 75790 44331 75792
rect 35020 75676 39600 75790
rect 44265 75787 44331 75790
rect 1697 75456 39593 75596
rect 1697 73120 35476 75456
rect 35556 73266 39600 75376
rect 44265 73266 44331 73269
rect 35556 73264 44331 73266
rect 35556 73208 44270 73264
rect 44326 73208 44331 73264
rect 35556 73206 44331 73208
rect 35556 73200 39600 73206
rect 44265 73203 44331 73206
rect 1697 72980 39593 73120
rect 1697 68098 38140 72980
rect 38220 68234 39600 72900
rect 44265 68234 44331 68237
rect 45553 68234 45619 68237
rect 38220 68232 45619 68234
rect 38220 68176 44270 68232
rect 44326 68176 45558 68232
rect 45614 68176 45619 68232
rect 38220 68174 45619 68176
rect 38220 68100 39600 68174
rect 44265 68171 44331 68174
rect 45553 68171 45619 68174
rect 212533 47698 212599 47701
rect 231577 47698 231643 47701
rect 212533 47696 231643 47698
rect 212533 47640 212538 47696
rect 212594 47640 231582 47696
rect 231638 47640 231643 47696
rect 212533 47638 231643 47640
rect 212533 47635 212599 47638
rect 231577 47635 231643 47638
rect 270493 47698 270559 47701
rect 289629 47698 289695 47701
rect 270493 47696 289695 47698
rect 270493 47640 270498 47696
rect 270554 47640 289634 47696
rect 289690 47640 289695 47696
rect 270493 47638 289695 47640
rect 270493 47635 270559 47638
rect 289629 47635 289695 47638
rect 154573 47154 154639 47157
rect 173801 47154 173867 47157
rect 154573 47152 173867 47154
rect 154573 47096 154578 47152
rect 154634 47096 173806 47152
rect 173862 47096 173867 47152
rect 154573 47094 173867 47096
rect 154573 47091 154639 47094
rect 173801 47091 173867 47094
rect 622945 40490 623011 40493
rect 84334 40488 623011 40490
rect 84334 40432 622950 40488
rect 623006 40432 623011 40488
rect 84334 40430 623011 40432
rect 84334 40218 84394 40430
rect 622945 40427 623011 40430
rect 149053 40354 149119 40357
rect 145838 40352 149119 40354
rect 145838 40296 149058 40352
rect 149114 40296 149119 40352
rect 145838 40294 149119 40296
rect 84150 40158 84394 40218
rect 86309 40218 86375 40221
rect 86309 40216 86602 40218
rect 86309 40160 86314 40216
rect 86370 40160 86602 40216
rect 86309 40158 86602 40160
rect 84150 40000 84210 40158
rect 86309 40155 86375 40158
rect 86542 40000 86602 40158
rect 145838 40000 145898 40294
rect 149053 40291 149119 40294
rect 47600 35977 51202 36017
rect 47600 35175 47646 35977
rect 51144 35175 51202 35977
rect 47600 33577 51202 35175
rect 47600 32987 47652 33577
rect 51182 32987 51202 33577
rect 47600 32953 51202 32987
rect 51600 35977 55202 36017
rect 51600 35175 51646 35977
rect 55144 35175 55202 35977
rect 51600 33577 55202 35175
rect 51600 32987 51652 33577
rect 55182 32987 55202 33577
rect 51600 32953 55202 32987
rect 55600 35977 59202 36017
rect 55600 35175 55646 35977
rect 59144 35175 59202 35977
rect 55600 33577 59202 35175
rect 55600 32987 55652 33577
rect 59182 32987 59202 33577
rect 55600 32953 59202 32987
rect 59600 35977 63202 36017
rect 59600 35175 59646 35977
rect 63144 35175 63202 35977
rect 59600 33577 63202 35175
rect 59600 32987 59652 33577
rect 63182 32987 63202 33577
rect 59600 32953 63202 32987
rect 63600 35977 67202 36017
rect 63600 35175 63646 35977
rect 67144 35175 67202 35977
rect 63600 33577 67202 35175
rect 63600 32987 63652 33577
rect 67182 32987 67202 33577
rect 63600 32953 67202 32987
rect 67600 35977 71202 36017
rect 67600 35175 67646 35977
rect 71144 35175 71202 35977
rect 67600 33577 71202 35175
rect 67600 32987 67652 33577
rect 71182 32987 71202 33577
rect 67600 32953 71202 32987
rect 78942 32648 83722 40000
rect 84022 37524 86222 40000
rect 86421 39810 88621 40000
rect 88921 39810 93701 40000
rect 86421 39750 93701 39810
rect 83802 37444 83942 37524
rect 86302 37444 86341 37524
rect 86421 37515 88621 39750
rect 83802 37435 86341 37444
rect 88701 37435 88841 37524
rect 83802 33417 88841 37435
rect 88921 33497 93701 39750
rect 101400 35977 105002 36017
rect 101400 35175 101446 35977
rect 104944 35175 105002 35977
rect 101400 33577 105002 35175
rect 83802 32568 93752 33417
rect 101400 32987 101452 33577
rect 104982 32987 105002 33577
rect 101400 32953 105002 32987
rect 105400 35977 109002 36017
rect 105400 35175 105446 35977
rect 108944 35175 109002 35977
rect 105400 33577 109002 35175
rect 105400 32987 105452 33577
rect 108982 32987 109002 33577
rect 105400 32953 109002 32987
rect 109400 35977 113002 36017
rect 109400 35175 109446 35977
rect 112944 35175 113002 35977
rect 109400 33577 113002 35175
rect 109400 32987 109452 33577
rect 112982 32987 113002 33577
rect 109400 32953 113002 32987
rect 113400 35977 117002 36017
rect 113400 35175 113446 35977
rect 116944 35175 117002 35977
rect 113400 33577 117002 35175
rect 113400 32987 113452 33577
rect 116982 32987 117002 33577
rect 113400 32953 117002 32987
rect 117400 35977 121002 36017
rect 117400 35175 117446 35977
rect 120944 35175 121002 35977
rect 117400 33577 121002 35175
rect 117400 32987 117452 33577
rect 120982 32987 121002 33577
rect 117400 32953 121002 32987
rect 121400 35977 125002 36017
rect 121400 35175 121446 35977
rect 124944 35175 125002 35977
rect 121400 33577 125002 35175
rect 121400 32987 121452 33577
rect 124982 32987 125002 33577
rect 121400 32953 125002 32987
rect 78942 980 93752 32568
rect 132660 30216 132868 39875
rect 132660 26680 132735 30216
rect 132948 30136 133162 40000
rect 132815 30016 133162 30136
rect 133242 37738 141587 39875
rect 141893 38746 143275 39875
rect 141893 38453 142982 38746
rect 143355 38666 143585 40000
rect 141893 38397 142926 38453
rect 143062 38420 143585 38666
rect 141893 38111 142710 38397
rect 143062 38373 143355 38420
rect 143388 38373 143585 38420
rect 143665 39293 143738 39875
rect 143818 39373 144151 40000
rect 144231 39293 145736 39875
rect 143006 38317 143062 38373
rect 143332 38317 143388 38373
rect 141953 38051 142710 38111
rect 133242 36966 141740 37738
rect 142046 37467 142710 38051
rect 142790 38300 143006 38317
rect 143019 38300 143332 38317
rect 142790 38120 143332 38300
rect 143665 38293 145736 39293
rect 143468 38237 145736 38293
rect 142790 38101 143006 38120
rect 143019 38101 143332 38120
rect 142790 38004 143332 38101
rect 142790 37547 143019 38004
rect 143412 37924 145736 38237
rect 143099 37467 145736 37924
rect 142046 36966 145736 37467
rect 133242 36603 145736 36966
rect 145816 36843 145920 40000
rect 146000 36923 147407 39875
rect 146042 36881 147407 36923
rect 145816 36801 145962 36843
rect 145816 36741 145934 36801
rect 145962 36741 146052 36801
rect 146132 36791 147407 36881
rect 145816 36711 146052 36741
rect 145816 36683 145934 36711
rect 145934 36651 146026 36683
rect 146052 36651 146142 36711
rect 146222 36701 147407 36791
rect 145934 36621 146142 36651
rect 133242 36511 145854 36603
rect 145934 36591 146245 36621
rect 146026 36531 146141 36591
rect 146142 36531 146245 36591
rect 133242 36396 145946 36511
rect 146026 36476 146245 36531
rect 133242 33821 146061 36396
rect 133242 33704 145944 33821
rect 146141 33741 146245 36476
rect 133242 33561 145801 33704
rect 146024 33669 146245 33741
rect 146024 33624 146141 33669
rect 146170 33624 146245 33669
rect 145881 33609 146024 33624
rect 146027 33609 146170 33624
rect 133242 33444 145684 33561
rect 145881 33519 146170 33609
rect 146325 33544 147407 36701
rect 145881 33481 146024 33519
rect 146027 33481 146170 33519
rect 145764 33459 145881 33481
rect 145910 33459 146027 33481
rect 133242 33401 145641 33444
rect 133242 33095 143065 33401
rect 145764 33399 146027 33459
rect 146250 33401 147407 33544
rect 145764 33364 145881 33399
rect 145910 33364 146027 33399
rect 145721 33321 145764 33364
rect 145806 33321 145910 33364
rect 143145 33291 145910 33321
rect 143145 33260 145777 33261
rect 145806 33260 145910 33291
rect 146107 33284 147407 33401
rect 143145 33231 145806 33260
rect 145721 33201 145806 33231
rect 143145 33175 145806 33201
rect 145990 33180 147407 33284
rect 145886 33095 147407 33180
rect 132815 30003 132948 30016
rect 132815 27080 133162 30003
rect 133242 27160 147407 33095
rect 155200 35977 158802 36017
rect 155200 35175 155246 35977
rect 158744 35175 158802 35977
rect 155200 33577 158802 35175
rect 155200 32987 155252 33577
rect 158782 32987 158802 33577
rect 155200 32953 158802 32987
rect 159200 35977 162802 36017
rect 159200 35175 159246 35977
rect 162744 35175 162802 35977
rect 159200 33577 162802 35175
rect 159200 32987 159252 33577
rect 162782 32987 162802 33577
rect 159200 32953 162802 32987
rect 163200 35977 166802 36017
rect 163200 35175 163246 35977
rect 166744 35175 166802 35977
rect 163200 33577 166802 35175
rect 163200 32987 163252 33577
rect 166782 32987 166802 33577
rect 163200 32953 166802 32987
rect 167200 35977 170802 36017
rect 167200 35175 167246 35977
rect 170744 35175 170802 35977
rect 167200 33577 170802 35175
rect 167200 32987 167252 33577
rect 170782 32987 170802 33577
rect 167200 32953 170802 32987
rect 171200 35977 174802 36017
rect 171200 35175 171246 35977
rect 174744 35175 174802 35977
rect 171200 33577 174802 35175
rect 171200 32987 171252 33577
rect 174782 32987 174802 33577
rect 171200 32953 174802 32987
rect 175200 35977 178802 36017
rect 175200 35175 175246 35977
rect 178744 35175 178802 35977
rect 175200 33577 178802 35175
rect 175200 32987 175252 33577
rect 178782 32987 178802 33577
rect 175200 32953 178802 32987
rect 132815 26760 133482 27080
rect 133562 26840 147407 27160
rect 132660 26360 133082 26680
rect 133162 26480 133762 26760
rect 133842 26560 147407 26840
rect 133162 26450 133949 26480
rect 133162 26440 133482 26450
rect 133482 26390 133739 26440
rect 133762 26390 133949 26450
rect 132660 26103 133402 26360
rect 133482 26293 133949 26390
rect 134029 26373 147407 26560
rect 133482 26270 133942 26293
rect 133482 26240 133739 26270
rect 133949 26240 134122 26293
rect 133482 26210 134122 26240
rect 133482 26183 133739 26210
rect 133739 26180 133929 26183
rect 133949 26180 134122 26210
rect 134202 26200 147407 26373
rect 133739 26120 134122 26180
rect 132660 25913 133659 26103
rect 133739 26090 134392 26120
rect 133739 26060 133929 26090
rect 134122 26060 134392 26090
rect 133739 26000 134392 26060
rect 133739 25993 133929 26000
rect 134122 25993 134392 26000
rect 132660 25720 133849 25913
rect 133929 25850 134392 25993
rect 134472 25930 147407 26200
rect 133929 25820 134628 25850
rect 133929 25800 134122 25820
rect 134122 25760 134364 25800
rect 134392 25760 134628 25820
rect 132660 25478 134042 25720
rect 134122 25584 134628 25760
rect 134122 25558 134364 25584
rect 134368 25558 134628 25584
rect 134364 25520 134628 25558
rect 132660 25440 134284 25478
rect 132660 20991 134322 25440
rect 134402 21071 134628 25520
rect 134708 20991 147407 25930
rect 132660 0 147407 20991
rect 186486 0 202338 40262
rect 240133 39946 240199 39949
rect 253933 39946 253999 39949
rect 240133 39944 246498 39946
rect 240133 39888 240138 39944
rect 240194 39888 246498 39944
rect 240133 39886 246498 39888
rect 240133 39883 240199 39886
rect 241237 39810 241303 39813
rect 242893 39810 242959 39813
rect 241156 39808 242959 39810
rect 241156 39752 241242 39808
rect 241298 39752 242898 39808
rect 242954 39752 242959 39808
rect 241156 39750 242959 39752
rect 241237 39747 241346 39750
rect 242893 39747 242959 39750
rect 241286 39600 241346 39747
rect 246438 39600 246498 39886
rect 248830 39944 253999 39946
rect 248830 39888 253938 39944
rect 253994 39888 253999 39944
rect 248830 39886 253999 39888
rect 248830 39600 248890 39886
rect 253933 39883 253999 39886
rect 210000 35977 213602 36017
rect 210000 35175 210046 35977
rect 213544 35175 213602 35977
rect 210000 33577 213602 35175
rect 210000 32987 210052 33577
rect 213582 32987 213602 33577
rect 210000 32953 213602 32987
rect 214000 35977 217602 36017
rect 214000 35175 214046 35977
rect 217544 35175 217602 35977
rect 214000 33577 217602 35175
rect 214000 32987 214052 33577
rect 217582 32987 217602 33577
rect 214000 32953 217602 32987
rect 218000 35977 221602 36017
rect 218000 35175 218046 35977
rect 221544 35175 221602 35977
rect 218000 33577 221602 35175
rect 218000 32987 218052 33577
rect 221582 32987 221602 33577
rect 218000 32953 221602 32987
rect 222000 35977 225602 36017
rect 222000 35175 222046 35977
rect 225544 35175 225602 35977
rect 222000 33577 225602 35175
rect 222000 32987 222052 33577
rect 225582 32987 225602 33577
rect 222000 32953 225602 32987
rect 226000 35977 229602 36017
rect 226000 35175 226046 35977
rect 229544 35175 229602 35977
rect 226000 33577 229602 35175
rect 226000 32987 226052 33577
rect 229582 32987 229602 33577
rect 226000 32953 229602 32987
rect 230000 35977 233602 36017
rect 230000 35175 230046 35977
rect 233544 35175 233602 35977
rect 230000 33577 233602 35175
rect 230000 32987 230052 33577
rect 233582 32987 233602 33577
rect 230000 32953 233602 32987
rect 241260 31680 246049 39600
rect 246349 39538 248524 39600
rect 248824 39538 251000 39600
rect 246349 39478 251000 39538
rect 246129 34940 246269 36042
rect 246349 35020 248524 39478
rect 248604 35476 248744 36042
rect 248824 35556 251000 39478
rect 251080 35476 251220 36042
rect 248604 34940 251220 35476
rect 246129 31600 251220 34940
rect 251300 31680 256100 39600
rect 263800 35977 267402 36017
rect 263800 35175 263846 35977
rect 267344 35175 267402 35977
rect 263800 33577 267402 35175
rect 263800 32987 263852 33577
rect 267382 32987 267402 33577
rect 263800 32953 267402 32987
rect 267800 35977 271402 36017
rect 267800 35175 267846 35977
rect 271344 35175 271402 35977
rect 267800 33577 271402 35175
rect 267800 32987 267852 33577
rect 271382 32987 271402 33577
rect 267800 32953 271402 32987
rect 271800 35977 275402 36017
rect 271800 35175 271846 35977
rect 275344 35175 275402 35977
rect 271800 33577 275402 35175
rect 271800 32987 271852 33577
rect 275382 32987 275402 33577
rect 271800 32953 275402 32987
rect 275800 35977 279402 36017
rect 275800 35175 275846 35977
rect 279344 35175 279402 35977
rect 275800 33577 279402 35175
rect 275800 32987 275852 33577
rect 279382 32987 279402 33577
rect 275800 32953 279402 32987
rect 279800 35977 283402 36017
rect 279800 35175 279846 35977
rect 283344 35175 283402 35977
rect 279800 33577 283402 35175
rect 279800 32987 279852 33577
rect 283382 32987 283402 33577
rect 279800 32953 283402 32987
rect 283800 35977 287402 36017
rect 283800 35175 283846 35977
rect 287344 35175 287402 35977
rect 283800 33577 287402 35175
rect 283800 32987 283852 33577
rect 287382 32987 287402 33577
rect 283800 32953 287402 32987
rect 241260 1697 256100 31600
rect 295086 0 310938 40262
rect 318600 35977 322202 36017
rect 318600 35175 318646 35977
rect 322144 35175 322202 35977
rect 318600 33577 322202 35175
rect 318600 32987 318652 33577
rect 322182 32987 322202 33577
rect 318600 32953 322202 32987
rect 322600 35977 326202 36017
rect 322600 35175 322646 35977
rect 326144 35175 326202 35977
rect 322600 33577 326202 35175
rect 322600 32987 322652 33577
rect 326182 32987 326202 33577
rect 322600 32953 326202 32987
rect 326600 35977 330202 36017
rect 326600 35175 326646 35977
rect 330144 35175 330202 35977
rect 326600 33577 330202 35175
rect 326600 32987 326652 33577
rect 330182 32987 330202 33577
rect 326600 32953 330202 32987
rect 330600 35977 334202 36017
rect 330600 35175 330646 35977
rect 334144 35175 334202 35977
rect 330600 33577 334202 35175
rect 330600 32987 330652 33577
rect 334182 32987 334202 33577
rect 330600 32953 334202 32987
rect 334600 35977 338202 36017
rect 334600 35175 334646 35977
rect 338144 35175 338202 35977
rect 334600 33577 338202 35175
rect 334600 32987 334652 33577
rect 338182 32987 338202 33577
rect 334600 32953 338202 32987
rect 338600 35977 342202 36017
rect 338600 35175 338646 35977
rect 342144 35175 342202 35977
rect 338600 33577 342202 35175
rect 338600 32987 338652 33577
rect 342182 32987 342202 33577
rect 338600 32953 342202 32987
rect 349886 0 365738 40262
rect 373400 35977 377002 36017
rect 373400 35175 373446 35977
rect 376944 35175 377002 35977
rect 373400 33577 377002 35175
rect 373400 32987 373452 33577
rect 376982 32987 377002 33577
rect 373400 32953 377002 32987
rect 377400 35977 381002 36017
rect 377400 35175 377446 35977
rect 380944 35175 381002 35977
rect 377400 33577 381002 35175
rect 377400 32987 377452 33577
rect 380982 32987 381002 33577
rect 377400 32953 381002 32987
rect 381400 35977 385002 36017
rect 381400 35175 381446 35977
rect 384944 35175 385002 35977
rect 381400 33577 385002 35175
rect 381400 32987 381452 33577
rect 384982 32987 385002 33577
rect 381400 32953 385002 32987
rect 385400 35977 389002 36017
rect 385400 35175 385446 35977
rect 388944 35175 389002 35977
rect 385400 33577 389002 35175
rect 385400 32987 385452 33577
rect 388982 32987 389002 33577
rect 385400 32953 389002 32987
rect 389400 35977 393002 36017
rect 389400 35175 389446 35977
rect 392944 35175 393002 35977
rect 389400 33577 393002 35175
rect 389400 32987 389452 33577
rect 392982 32987 393002 33577
rect 389400 32953 393002 32987
rect 393400 35977 397002 36017
rect 393400 35175 393446 35977
rect 396944 35175 397002 35977
rect 393400 33577 397002 35175
rect 393400 32987 393452 33577
rect 396982 32987 397002 33577
rect 393400 32953 397002 32987
rect 404686 0 420538 40262
rect 428200 35977 431802 36017
rect 428200 35175 428246 35977
rect 431744 35175 431802 35977
rect 428200 33577 431802 35175
rect 428200 32987 428252 33577
rect 431782 32987 431802 33577
rect 428200 32953 431802 32987
rect 432200 35977 435802 36017
rect 432200 35175 432246 35977
rect 435744 35175 435802 35977
rect 432200 33577 435802 35175
rect 432200 32987 432252 33577
rect 435782 32987 435802 33577
rect 432200 32953 435802 32987
rect 436200 35977 439802 36017
rect 436200 35175 436246 35977
rect 439744 35175 439802 35977
rect 436200 33577 439802 35175
rect 436200 32987 436252 33577
rect 439782 32987 439802 33577
rect 436200 32953 439802 32987
rect 440200 35977 443802 36017
rect 440200 35175 440246 35977
rect 443744 35175 443802 35977
rect 440200 33577 443802 35175
rect 440200 32987 440252 33577
rect 443782 32987 443802 33577
rect 440200 32953 443802 32987
rect 444200 35977 447802 36017
rect 444200 35175 444246 35977
rect 447744 35175 447802 35977
rect 444200 33577 447802 35175
rect 444200 32987 444252 33577
rect 447782 32987 447802 33577
rect 444200 32953 447802 32987
rect 448200 35977 451802 36017
rect 448200 35175 448246 35977
rect 451744 35175 451802 35977
rect 448200 33577 451802 35175
rect 448200 32987 448252 33577
rect 451782 32987 451802 33577
rect 448200 32953 451802 32987
rect 459486 0 475338 40262
rect 483000 35977 486602 36017
rect 483000 35175 483046 35977
rect 486544 35175 486602 35977
rect 483000 33577 486602 35175
rect 483000 32987 483052 33577
rect 486582 32987 486602 33577
rect 483000 32953 486602 32987
rect 487000 35977 490602 36017
rect 487000 35175 487046 35977
rect 490544 35175 490602 35977
rect 487000 33577 490602 35175
rect 487000 32987 487052 33577
rect 490582 32987 490602 33577
rect 487000 32953 490602 32987
rect 491000 35977 494602 36017
rect 491000 35175 491046 35977
rect 494544 35175 494602 35977
rect 491000 33577 494602 35175
rect 491000 32987 491052 33577
rect 494582 32987 494602 33577
rect 491000 32953 494602 32987
rect 495000 35977 498602 36017
rect 495000 35175 495046 35977
rect 498544 35175 498602 35977
rect 495000 33577 498602 35175
rect 495000 32987 495052 33577
rect 498582 32987 498602 33577
rect 495000 32953 498602 32987
rect 499000 35977 502602 36017
rect 499000 35175 499046 35977
rect 502544 35175 502602 35977
rect 499000 33577 502602 35175
rect 499000 32987 499052 33577
rect 502582 32987 502602 33577
rect 499000 32953 502602 32987
rect 503000 35977 506602 36017
rect 503000 35175 503046 35977
rect 506544 35175 506602 35977
rect 503000 33577 506602 35175
rect 503000 32987 503052 33577
rect 506582 32987 506602 33577
rect 503000 32953 506602 32987
rect 514286 0 530138 40262
rect 569217 40218 569283 40221
rect 579153 40218 579219 40221
rect 569174 40216 579219 40218
rect 569174 40160 569222 40216
rect 569278 40160 579158 40216
rect 579214 40160 579219 40216
rect 569174 40158 579219 40160
rect 569174 40155 569283 40158
rect 579153 40155 579219 40158
rect 632973 40218 633039 40221
rect 634813 40218 634879 40221
rect 632973 40216 634879 40218
rect 632973 40160 632978 40216
rect 633034 40160 634818 40216
rect 634874 40160 634879 40216
rect 632973 40158 634879 40160
rect 632973 40155 633039 40158
rect 634813 40155 634879 40158
rect 569174 40000 569234 40155
rect 537800 35977 541402 36017
rect 537800 35175 537846 35977
rect 541344 35175 541402 35977
rect 537800 33577 541402 35175
rect 537800 32987 537852 33577
rect 541382 32987 541402 33577
rect 537800 32953 541402 32987
rect 541800 35977 545402 36017
rect 541800 35175 541846 35977
rect 545344 35175 545402 35977
rect 541800 33577 545402 35175
rect 541800 32987 541852 33577
rect 545382 32987 545402 33577
rect 541800 32953 545402 32987
rect 545800 35977 549402 36017
rect 545800 35175 545846 35977
rect 549344 35175 549402 35977
rect 545800 33577 549402 35175
rect 545800 32987 545852 33577
rect 549382 32987 549402 33577
rect 545800 32953 549402 32987
rect 549800 35977 553402 36017
rect 549800 35175 549846 35977
rect 553344 35175 553402 35977
rect 549800 33577 553402 35175
rect 549800 32987 549852 33577
rect 553382 32987 553402 33577
rect 549800 32953 553402 32987
rect 553800 35977 557402 36017
rect 553800 35175 553846 35977
rect 557344 35175 557402 35977
rect 553800 33577 557402 35175
rect 553800 32987 553852 33577
rect 557382 32987 557402 33577
rect 553800 32953 557402 32987
rect 557800 35977 561402 36017
rect 557800 35175 557846 35977
rect 561344 35175 561402 35977
rect 557800 33577 561402 35175
rect 569142 34830 573922 40000
rect 574222 37524 576422 40000
rect 574002 37444 574142 37524
rect 576502 37444 576541 37524
rect 576621 37515 578821 40000
rect 574002 37435 576541 37444
rect 578901 37435 579041 37524
rect 574002 34750 579041 37435
rect 579121 34830 583901 40000
rect 622942 39672 627722 40000
rect 622942 39616 622950 39672
rect 623006 39616 627722 39672
rect 622942 37008 627722 39616
rect 627802 37654 627942 39455
rect 628022 37734 630222 40000
rect 630421 39455 632621 40000
rect 630302 39375 630341 39455
rect 632701 39375 632841 39455
rect 630302 37654 632841 39375
rect 627802 36928 632841 37654
rect 632921 37008 637701 40000
rect 591600 35977 595202 36017
rect 591600 35175 591646 35977
rect 595144 35175 595202 35977
rect 557800 32987 557852 33577
rect 561382 32987 561402 33577
rect 557800 32953 561402 32987
rect 569142 0 583952 34750
rect 591600 33577 595202 35175
rect 591600 32987 591652 33577
rect 595182 32987 595202 33577
rect 591600 32953 595202 32987
rect 595600 35977 599202 36017
rect 595600 35175 595646 35977
rect 599144 35175 599202 35977
rect 595600 33577 599202 35175
rect 595600 32987 595652 33577
rect 599182 32987 599202 33577
rect 595600 32953 599202 32987
rect 599600 35977 603202 36017
rect 599600 35175 599646 35977
rect 603144 35175 603202 35977
rect 599600 33577 603202 35175
rect 599600 32987 599652 33577
rect 603182 32987 603202 33577
rect 599600 32953 603202 32987
rect 603600 35977 607202 36017
rect 603600 35175 603646 35977
rect 607144 35175 607202 35977
rect 603600 33577 607202 35175
rect 603600 32987 603652 33577
rect 607182 32987 607202 33577
rect 603600 32953 607202 32987
rect 607600 35977 611202 36017
rect 607600 35175 607646 35977
rect 611144 35175 611202 35977
rect 607600 33577 611202 35175
rect 607600 32987 607652 33577
rect 611182 32987 611202 33577
rect 607600 32953 611202 32987
rect 611600 35977 615202 36017
rect 611600 35175 611646 35977
rect 615144 35175 615202 35977
rect 611600 33577 615202 35175
rect 611600 32987 611652 33577
rect 615182 32987 615202 33577
rect 611600 32953 615202 32987
rect 622869 0 637752 36928
rect 645400 35977 649002 36017
rect 645400 35175 645446 35977
rect 648944 35175 649002 35977
rect 645400 33577 649002 35175
rect 645400 32987 645452 33577
rect 648982 32987 649002 33577
rect 645400 32953 649002 32987
rect 649400 35977 653002 36017
rect 649400 35175 649446 35977
rect 652944 35175 653002 35977
rect 649400 33577 653002 35175
rect 649400 32987 649452 33577
rect 652982 32987 653002 33577
rect 649400 32953 653002 32987
rect 653400 35977 657002 36017
rect 653400 35175 653446 35977
rect 656944 35175 657002 35977
rect 653400 33577 657002 35175
rect 653400 32987 653452 33577
rect 656982 32987 657002 33577
rect 653400 32953 657002 32987
rect 657400 35977 661002 36017
rect 657400 35175 657446 35977
rect 660944 35175 661002 35977
rect 657400 33577 661002 35175
rect 657400 32987 657452 33577
rect 660982 32987 661002 33577
rect 657400 32953 661002 32987
rect 661400 35977 665002 36017
rect 661400 35175 661446 35977
rect 664944 35175 665002 35977
rect 661400 33577 665002 35175
rect 661400 32987 661452 33577
rect 664982 32987 665002 33577
rect 661400 32953 665002 32987
rect 665400 35977 669002 36017
rect 665400 35175 665446 35977
rect 668944 35175 669002 35977
rect 665400 33577 669002 35175
rect 665400 32987 665452 33577
rect 668982 32987 669002 33577
rect 665400 32953 669002 32987
<< via3 >>
rect 39854 837528 39868 837584
<< obsm4 >>
rect 0 1032677 40466 1037600
rect 40546 1032757 76454 1037600
rect 0 1016680 40549 1032677
rect 0 1011527 40349 1016680
rect 40800 1016600 76200 1032757
rect 76534 1032677 91866 1037600
rect 91946 1032757 127854 1037600
rect 76393 1016680 91994 1032677
rect 40429 1011607 76454 1016600
rect 0 1011387 40549 1011527
rect 40800 1011387 76200 1011607
rect 76534 1011527 91866 1016680
rect 92200 1016600 127600 1032757
rect 127934 1032677 143266 1037600
rect 143346 1032757 179254 1037600
rect 127793 1016680 143394 1032677
rect 91946 1011607 127854 1016600
rect 76393 1011387 91994 1011527
rect 92200 1011387 127600 1011607
rect 127934 1011527 143266 1016680
rect 143600 1016600 179000 1032757
rect 179334 1032677 194666 1037600
rect 194746 1032757 230654 1037600
rect 179193 1016680 194794 1032677
rect 143346 1011607 179254 1016600
rect 127793 1011387 143394 1011527
rect 143600 1011387 179000 1011607
rect 179334 1011527 194666 1016680
rect 195000 1016600 230400 1032757
rect 230734 1032677 246066 1037600
rect 246146 1032757 282254 1037600
rect 230593 1016680 246194 1032677
rect 194746 1011607 230654 1016600
rect 179193 1011387 194794 1011527
rect 195000 1011387 230400 1011607
rect 230734 1011527 246066 1016680
rect 246400 1016600 282000 1032757
rect 282334 1032677 297666 1037600
rect 297746 1032757 333654 1037600
rect 282193 1016680 297794 1032677
rect 246146 1011607 282254 1016600
rect 230593 1011387 246194 1011527
rect 246400 1011387 282000 1011607
rect 282334 1011527 297666 1016680
rect 298000 1016600 333400 1032757
rect 333734 1032677 348066 1037600
rect 348146 1032757 384054 1037600
rect 333593 1016680 348207 1032677
rect 297746 1011607 333654 1016600
rect 282193 1011387 297794 1011527
rect 298000 1011387 333400 1011607
rect 333734 1011527 348066 1016680
rect 348400 1016600 383800 1032757
rect 384134 1032677 399466 1037600
rect 399546 1032757 473054 1037600
rect 383993 1016680 399594 1032677
rect 348146 1011607 384054 1016600
rect 333593 1011387 348207 1011527
rect 348400 1011387 383800 1011607
rect 384134 1011527 399466 1016680
rect 399800 1016600 472800 1032757
rect 473134 1032677 488466 1037600
rect 488546 1032757 524454 1037600
rect 472993 1016680 488594 1032677
rect 399546 1011607 473054 1016600
rect 383993 1011387 399594 1011527
rect 399800 1011387 435200 1011607
rect 436200 1011387 472800 1011607
rect 473134 1011527 488466 1016680
rect 488800 1016600 524200 1032757
rect 524534 1032677 539866 1037600
rect 539946 1032757 575854 1037600
rect 524393 1016680 539994 1032677
rect 488546 1011607 524454 1016600
rect 472993 1011387 488594 1011527
rect 488800 1011387 524200 1011607
rect 524534 1011527 539866 1016680
rect 540200 1016600 575600 1032757
rect 575934 1032677 590266 1037600
rect 590346 1032757 626254 1037600
rect 575793 1016680 590407 1032677
rect 539946 1011607 575854 1016600
rect 524393 1011387 539994 1011527
rect 540200 1011387 575600 1011607
rect 575934 1011527 590266 1016680
rect 590600 1016600 626000 1032757
rect 626334 1032677 641666 1037600
rect 641746 1032757 677887 1037600
rect 642000 1032677 677600 1032757
rect 677967 1032677 717600 1037600
rect 626193 1016680 641794 1032677
rect 642000 1016680 717600 1032677
rect 590346 1011607 626254 1016600
rect 575793 1011387 590407 1011527
rect 590600 1011387 626000 1011607
rect 626334 1011527 641666 1016680
rect 642000 1016600 677600 1016680
rect 641746 1011607 678129 1016600
rect 642000 1011527 677600 1011607
rect 678209 1011527 717600 1016680
rect 626193 1011387 641794 1011527
rect 642000 1011387 717600 1011527
rect 0 1010337 40466 1011387
rect 40546 1010417 76454 1011307
rect 76534 1010337 91866 1011387
rect 91946 1010417 127854 1011307
rect 127934 1010337 143266 1011387
rect 143346 1010417 179254 1011307
rect 179334 1010337 194666 1011387
rect 194746 1010417 230654 1011307
rect 230734 1010337 246066 1011387
rect 246146 1010417 282254 1011307
rect 282334 1010337 297666 1011387
rect 297746 1010417 333654 1011307
rect 333734 1010337 348066 1011387
rect 348146 1010417 384054 1011307
rect 384134 1010337 399466 1011387
rect 399546 1010417 473054 1011307
rect 473134 1010337 488466 1011387
rect 488546 1010417 524454 1011307
rect 524534 1010337 539866 1011387
rect 539946 1010417 575854 1011307
rect 575934 1010337 590266 1011387
rect 590346 1010417 626254 1011307
rect 626334 1010337 641666 1011387
rect 641746 1010417 677896 1011307
rect 677976 1010337 717600 1011387
rect 0 1010217 40549 1010337
rect 40800 1010217 76200 1010337
rect 76393 1010217 91994 1010337
rect 92200 1010217 127600 1010337
rect 127793 1010217 143394 1010337
rect 143600 1010217 179000 1010337
rect 179193 1010217 194794 1010337
rect 195000 1010217 230400 1010337
rect 230593 1010217 246194 1010337
rect 246400 1010217 282000 1010337
rect 282193 1010217 297794 1010337
rect 298000 1010217 333400 1010337
rect 333593 1010217 348207 1010337
rect 348400 1010217 383800 1010337
rect 383993 1010217 399594 1010337
rect 399800 1010217 435200 1010337
rect 436200 1010217 472800 1010337
rect 472993 1010217 488594 1010337
rect 488800 1010217 524200 1010337
rect 524393 1010217 539994 1010337
rect 540200 1010217 575600 1010337
rect 575793 1010217 590407 1010337
rect 590600 1010217 626000 1010337
rect 626193 1010217 641794 1010337
rect 642000 1010217 717600 1010337
rect 0 1009167 40466 1010217
rect 40546 1009247 76454 1010137
rect 76534 1009167 91866 1010217
rect 91946 1009247 127854 1010137
rect 127934 1009167 143266 1010217
rect 143346 1009247 179254 1010137
rect 179334 1009167 194666 1010217
rect 194746 1009247 230654 1010137
rect 230734 1009167 246066 1010217
rect 246146 1009247 282254 1010137
rect 282334 1009167 297666 1010217
rect 297746 1009247 333654 1010137
rect 333734 1009167 348066 1010217
rect 348146 1009247 384054 1010137
rect 384134 1009167 399466 1010217
rect 399546 1009247 473054 1010137
rect 473134 1009167 488466 1010217
rect 488546 1009247 524454 1010137
rect 524534 1009167 539866 1010217
rect 539946 1009247 575854 1010137
rect 575934 1009167 590266 1010217
rect 590346 1009247 626254 1010137
rect 626334 1009167 641666 1010217
rect 641746 1009247 677925 1010137
rect 678005 1009167 717600 1010217
rect 0 1009027 40549 1009167
rect 40800 1009027 76200 1009167
rect 76393 1009027 91994 1009167
rect 92200 1009027 127600 1009167
rect 127793 1009027 143394 1009167
rect 143600 1009027 179000 1009167
rect 179193 1009027 194794 1009167
rect 195000 1009027 230400 1009167
rect 230593 1009027 246194 1009167
rect 246400 1009027 282000 1009167
rect 282193 1009027 297794 1009167
rect 298000 1009027 333400 1009167
rect 333593 1009027 348207 1009167
rect 348400 1009027 383800 1009167
rect 383993 1009027 399594 1009167
rect 399800 1009027 435200 1009167
rect 436200 1009027 472800 1009167
rect 472993 1009027 488594 1009167
rect 488800 1009027 524200 1009167
rect 524393 1009027 539994 1009167
rect 540200 1009027 575600 1009167
rect 575793 1009027 590407 1009167
rect 590600 1009027 626000 1009167
rect 626193 1009027 641794 1009167
rect 642000 1009027 717600 1009167
rect 0 1008801 35285 1009027
rect 35365 1008881 76722 1008947
rect 76802 1008901 85538 1009027
rect 0 1008145 35338 1008801
rect 35418 1008225 83488 1008821
rect 36489 1008145 40800 1008165
rect 76200 1008145 76454 1008165
rect 83568 1008145 83872 1008901
rect 85618 1008881 128122 1008947
rect 128202 1008901 136938 1009027
rect 83952 1008225 134888 1008821
rect 91946 1008145 92200 1008165
rect 127600 1008145 127854 1008165
rect 134968 1008145 135272 1008901
rect 137018 1008881 179522 1008947
rect 179602 1008901 188338 1009027
rect 135352 1008225 186288 1008821
rect 143346 1008145 143600 1008165
rect 179000 1008145 179254 1008165
rect 186368 1008145 186672 1008901
rect 188418 1008881 230922 1008947
rect 231002 1008901 239738 1009027
rect 186752 1008225 237688 1008821
rect 194746 1008145 195000 1008165
rect 230400 1008145 230654 1008165
rect 237768 1008145 238072 1008901
rect 239818 1008881 282522 1008947
rect 282602 1008901 291338 1009027
rect 238152 1008225 289288 1008821
rect 246146 1008145 246400 1008165
rect 282000 1008145 282254 1008165
rect 289368 1008145 289672 1008901
rect 291418 1008881 384322 1008947
rect 384402 1008901 393138 1009027
rect 289752 1008225 391088 1008821
rect 297746 1008145 298000 1008165
rect 333400 1008145 333654 1008165
rect 348146 1008145 348400 1008165
rect 383800 1008145 384054 1008165
rect 391168 1008145 391472 1008901
rect 393218 1008881 435200 1008947
rect 436200 1008881 473322 1008947
rect 473402 1008901 482138 1009027
rect 391552 1008225 480088 1008821
rect 399546 1008145 399800 1008165
rect 472800 1008145 473054 1008165
rect 480168 1008145 480472 1008901
rect 482218 1008881 524722 1008947
rect 524802 1008901 533538 1009027
rect 480552 1008225 531488 1008821
rect 488546 1008145 488800 1008165
rect 524200 1008145 524454 1008165
rect 531568 1008145 531872 1008901
rect 533618 1008881 575854 1008947
rect 575934 1008901 590266 1009027
rect 590346 1008881 626522 1008947
rect 626602 1008901 635338 1009027
rect 531952 1008225 633288 1008821
rect 539946 1008145 540200 1008165
rect 575600 1008145 575854 1008165
rect 590346 1008145 590600 1008165
rect 626000 1008145 626254 1008165
rect 633368 1008145 633672 1008901
rect 635418 1008881 682235 1008947
rect 633752 1008225 682182 1008821
rect 682315 1008801 717600 1009027
rect 641746 1008145 642000 1008165
rect 677600 1008145 681910 1008165
rect 682262 1008145 717600 1008801
rect 0 1007849 36409 1008145
rect 36489 1007949 76454 1008145
rect 76534 1007949 91866 1008145
rect 91946 1007949 127854 1008145
rect 127934 1007949 143266 1008145
rect 143346 1007949 179254 1008145
rect 179334 1007949 194666 1008145
rect 194746 1007949 230654 1008145
rect 230734 1007949 246066 1008145
rect 246146 1007949 282254 1008145
rect 282334 1007949 297666 1008145
rect 297746 1007949 333654 1008145
rect 333734 1007949 348066 1008145
rect 348146 1007949 384054 1008145
rect 384134 1007949 399466 1008145
rect 399546 1007949 435200 1008145
rect 436200 1007949 473054 1008145
rect 473134 1007949 488466 1008145
rect 488546 1007949 524454 1008145
rect 524534 1007949 539866 1008145
rect 539946 1007949 575854 1008145
rect 575934 1007949 590266 1008145
rect 590346 1007949 626254 1008145
rect 626334 1007949 641666 1008145
rect 641746 1007949 681910 1008145
rect 36489 1007929 40800 1007949
rect 76200 1007929 76454 1007949
rect 0 1007293 36545 1007849
rect 0 1007067 36005 1007293
rect 36625 1007273 86629 1007869
rect 86709 1007293 87013 1007949
rect 91946 1007929 92200 1007949
rect 127600 1007929 127854 1007949
rect 87093 1007273 138029 1007869
rect 138109 1007293 138413 1007949
rect 143346 1007929 143600 1007949
rect 179000 1007929 179254 1007949
rect 138493 1007273 189429 1007869
rect 189509 1007293 189813 1007949
rect 194746 1007929 195000 1007949
rect 230400 1007929 230654 1007949
rect 189893 1007273 240829 1007869
rect 240909 1007293 241213 1007949
rect 246146 1007929 246400 1007949
rect 282000 1007929 282254 1007949
rect 241293 1007273 292429 1007869
rect 292509 1007293 292813 1007949
rect 297746 1007929 298000 1007949
rect 333400 1007929 333654 1007949
rect 348146 1007929 348400 1007949
rect 383800 1007929 384054 1007949
rect 292893 1007273 394229 1007869
rect 394309 1007293 394613 1007949
rect 399546 1007929 399800 1007949
rect 472800 1007929 473054 1007949
rect 394693 1007273 483229 1007869
rect 483309 1007293 483613 1007949
rect 488546 1007929 488800 1007949
rect 524200 1007929 524454 1007949
rect 483693 1007273 534629 1007869
rect 534709 1007293 535013 1007949
rect 539946 1007929 540200 1007949
rect 575600 1007929 575854 1007949
rect 590346 1007929 590600 1007949
rect 626000 1007929 626254 1007949
rect 535093 1007273 636429 1007869
rect 636509 1007293 636813 1007949
rect 641746 1007929 642000 1007949
rect 677600 1007929 681910 1007949
rect 636893 1007273 681787 1007869
rect 681990 1007849 717600 1008145
rect 36085 1007147 76722 1007213
rect 76802 1007067 85538 1007193
rect 85618 1007147 128122 1007213
rect 128202 1007067 136938 1007193
rect 137018 1007147 179522 1007213
rect 179602 1007067 188338 1007193
rect 188418 1007147 230922 1007213
rect 231002 1007067 239738 1007193
rect 239818 1007147 282522 1007213
rect 282602 1007067 291338 1007193
rect 291418 1007147 384322 1007213
rect 384402 1007067 393138 1007193
rect 393218 1007147 435200 1007213
rect 436200 1007147 473322 1007213
rect 473402 1007067 482138 1007193
rect 482218 1007147 524722 1007213
rect 524802 1007067 533538 1007193
rect 533618 1007147 575854 1007213
rect 575934 1007067 590266 1007193
rect 590346 1007147 626522 1007213
rect 626602 1007067 635338 1007193
rect 635418 1007147 681515 1007213
rect 681867 1007193 717600 1007849
rect 681595 1007067 717600 1007193
rect 0 1006927 40549 1007067
rect 76393 1006927 91994 1007067
rect 127793 1006927 143394 1007067
rect 179193 1006927 194794 1007067
rect 230593 1006927 246194 1007067
rect 282193 1006927 297794 1007067
rect 333593 1006927 348207 1007067
rect 383993 1006927 399594 1007067
rect 472993 1006927 488594 1007067
rect 524393 1006927 539994 1007067
rect 575793 1006927 590407 1007067
rect 626193 1006927 641794 1007067
rect 677600 1006927 717600 1007067
rect 0 1005837 40466 1006927
rect 40546 1005917 76454 1006847
rect 76534 1005837 91866 1006927
rect 91946 1005917 127854 1006847
rect 127934 1005837 143266 1006927
rect 143346 1005917 179254 1006847
rect 179334 1005837 194666 1006927
rect 194746 1005917 230654 1006847
rect 230734 1005837 246066 1006927
rect 246146 1005917 282254 1006847
rect 282334 1005837 297666 1006927
rect 297746 1005917 333654 1006847
rect 333734 1005837 348066 1006927
rect 348146 1005917 384054 1006847
rect 384134 1005837 399466 1006927
rect 399546 1005917 436200 1006847
rect 437200 1005917 473054 1006847
rect 473134 1005837 488466 1006927
rect 488546 1005917 524454 1006847
rect 524534 1005837 539866 1006927
rect 539946 1005917 575854 1006847
rect 575934 1005837 590266 1006927
rect 590346 1005917 626254 1006847
rect 626334 1005837 641666 1006927
rect 641746 1005917 677895 1006847
rect 677975 1005837 717600 1006927
rect 0 1005717 40549 1005837
rect 76393 1005717 91994 1005837
rect 127793 1005717 143394 1005837
rect 179193 1005717 194794 1005837
rect 230593 1005717 246194 1005837
rect 282193 1005717 297794 1005837
rect 333593 1005717 348207 1005837
rect 383993 1005717 399594 1005837
rect 472993 1005717 488594 1005837
rect 524393 1005717 539994 1005837
rect 575793 1005717 590407 1005837
rect 626193 1005717 641794 1005837
rect 677600 1005717 717600 1005837
rect 0 1004867 40466 1005717
rect 40546 1004947 76454 1005637
rect 76534 1004867 91866 1005717
rect 91946 1004947 127854 1005637
rect 127934 1004867 143266 1005717
rect 143346 1004947 179254 1005637
rect 179334 1004867 194666 1005717
rect 194746 1004947 230654 1005637
rect 230734 1004867 246066 1005717
rect 246146 1004947 282254 1005637
rect 282334 1004867 297666 1005717
rect 297746 1004947 333654 1005637
rect 333734 1004867 348066 1005717
rect 348146 1004947 384054 1005637
rect 384134 1004867 399466 1005717
rect 399546 1004947 435200 1005637
rect 436200 1004947 473054 1005637
rect 473134 1004867 488466 1005717
rect 488546 1004947 524454 1005637
rect 524534 1004867 539866 1005717
rect 539946 1004947 575854 1005637
rect 575934 1004867 590266 1005717
rect 590346 1004947 626254 1005637
rect 626334 1004867 641666 1005717
rect 641746 1004947 677867 1005637
rect 677947 1004867 717600 1005717
rect 0 1004747 40549 1004867
rect 76393 1004747 91994 1004867
rect 127793 1004747 143394 1004867
rect 179193 1004747 194794 1004867
rect 230593 1004747 246194 1004867
rect 282193 1004747 297794 1004867
rect 333593 1004747 348207 1004867
rect 383993 1004747 399594 1004867
rect 472993 1004747 488594 1004867
rect 524393 1004747 539994 1004867
rect 575793 1004747 590407 1004867
rect 626193 1004747 641794 1004867
rect 677600 1004747 717600 1004867
rect 0 1003897 40466 1004747
rect 40546 1003977 76454 1004667
rect 76534 1003897 91866 1004747
rect 91946 1003977 127854 1004667
rect 127934 1003897 143266 1004747
rect 143346 1003977 179254 1004667
rect 179334 1003897 194666 1004747
rect 194746 1003977 230654 1004667
rect 230734 1003897 246066 1004747
rect 246146 1003977 282254 1004667
rect 282334 1003897 297666 1004747
rect 297746 1003977 333654 1004667
rect 333734 1003897 348066 1004747
rect 348146 1003977 384054 1004667
rect 384134 1003897 399466 1004747
rect 399546 1003977 473054 1004667
rect 473134 1003897 488466 1004747
rect 488546 1003977 524454 1004667
rect 524534 1003897 539866 1004747
rect 539946 1003977 575854 1004667
rect 575934 1003897 590266 1004747
rect 590346 1003977 626254 1004667
rect 626334 1003897 641666 1004747
rect 641746 1003977 677877 1004667
rect 677957 1003897 717600 1004747
rect 0 1003777 40549 1003897
rect 76393 1003777 91994 1003897
rect 127793 1003777 143394 1003897
rect 179193 1003777 194794 1003897
rect 230593 1003777 246194 1003897
rect 282193 1003777 297794 1003897
rect 333593 1003777 348207 1003897
rect 383993 1003777 399594 1003897
rect 472993 1003777 488594 1003897
rect 524393 1003777 539994 1003897
rect 575793 1003777 590407 1003897
rect 626193 1003777 641794 1003897
rect 677600 1003777 717600 1003897
rect 0 1002687 40466 1003777
rect 40546 1002767 76454 1003697
rect 76534 1002687 91866 1003777
rect 91946 1002767 127854 1003697
rect 127934 1002687 143266 1003777
rect 143346 1002767 179254 1003697
rect 179334 1002687 194666 1003777
rect 194746 1002767 230654 1003697
rect 230734 1002687 246066 1003777
rect 246146 1002767 282254 1003697
rect 282334 1002687 297666 1003777
rect 297746 1002767 333654 1003697
rect 333734 1002687 348066 1003777
rect 348146 1002767 384054 1003697
rect 384134 1002687 399466 1003777
rect 399546 1002767 473054 1003697
rect 473134 1002687 488466 1003777
rect 488546 1002767 524454 1003697
rect 524534 1002687 539866 1003777
rect 539946 1002767 575854 1003697
rect 575934 1002687 590266 1003777
rect 590346 1002767 626254 1003697
rect 626334 1002687 641666 1003777
rect 641746 1002767 677920 1003697
rect 678000 1002687 717600 1003777
rect 0 1002567 40549 1002687
rect 76393 1002567 91994 1002687
rect 127793 1002567 143394 1002687
rect 179193 1002567 194794 1002687
rect 230593 1002567 246194 1002687
rect 282193 1002567 297794 1002687
rect 333593 1002567 348207 1002687
rect 383993 1002567 399594 1002687
rect 472993 1002567 488594 1002687
rect 524393 1002567 539994 1002687
rect 575793 1002567 590407 1002687
rect 626193 1002567 641794 1002687
rect 677600 1002567 717600 1002687
rect 0 1002315 40466 1002567
rect 0 998209 28573 1002315
rect 28799 1002262 40466 1002315
rect 0 997967 20920 998209
rect 0 997600 4843 997887
rect 4923 997600 20920 997967
rect 21000 997600 25993 998129
rect 26073 998005 28573 998209
rect 26073 997976 27383 998005
rect 26073 997600 26213 997976
rect 0 970200 26213 997600
rect 0 969946 4843 970200
rect 4923 969866 20920 969994
rect 21000 969946 25993 970200
rect 26073 969866 26213 969994
rect 26293 969946 27183 997896
rect 27263 970200 27383 997976
rect 27263 969866 27383 969994
rect 27463 969946 28353 997925
rect 28433 970200 28573 998005
rect 28433 969866 28573 969994
rect 0 963538 28573 969866
rect 28653 963618 28719 1002235
rect 0 961872 28699 963538
rect 28779 961952 29375 1002182
rect 29455 1001990 40466 1002262
rect 29435 997600 29671 1001910
rect 29751 1001867 40466 1001990
rect 29455 970200 29651 997600
rect 29435 969946 29671 970200
rect 29455 965013 29651 969866
rect 29731 965093 30327 1001787
rect 30407 1001595 40466 1001867
rect 29455 964709 30307 965013
rect 29455 961872 29651 964709
rect 0 961568 29651 961872
rect 0 954802 28699 961568
rect 0 954534 28573 954802
rect 0 954200 4843 954454
rect 4923 954393 20920 954534
rect 21000 954200 25993 954454
rect 26073 954393 26213 954534
rect 0 927000 26213 954200
rect 0 926746 4843 927000
rect 4923 926666 20920 926807
rect 21000 926746 25993 927000
rect 26073 926666 26213 926807
rect 26293 926746 27183 954454
rect 27263 954393 27383 954534
rect 27263 927000 27383 954200
rect 27263 926666 27383 926807
rect 27463 926746 28353 954454
rect 28433 954393 28573 954534
rect 28433 927000 28573 954200
rect 28433 926666 28573 926807
rect 0 912334 28573 926666
rect 0 912000 4843 912254
rect 4923 912193 20920 912334
rect 21000 912000 25993 912254
rect 26073 912193 26213 912334
rect 0 884800 26213 912000
rect 0 884546 4843 884800
rect 4923 884466 20920 884607
rect 21000 884546 25993 884800
rect 26073 884466 26213 884607
rect 26293 884546 27183 912254
rect 27263 912193 27383 912334
rect 27263 884800 27383 912000
rect 27263 884466 27383 884607
rect 27463 884546 28353 912254
rect 28433 912193 28573 912334
rect 28433 884800 28573 912000
rect 28433 884466 28573 884607
rect 0 870134 28573 884466
rect 0 869800 4843 870054
rect 4923 869993 20920 870134
rect 21000 869800 25993 870054
rect 26073 869993 26213 870134
rect 0 842600 26213 869800
rect 0 842346 4843 842600
rect 4923 842266 20920 842407
rect 21000 842346 25993 842600
rect 26073 842266 26213 842407
rect 26293 842346 27183 870054
rect 27263 869993 27383 870134
rect 27263 842600 27383 869800
rect 27263 842266 27383 842407
rect 27463 842346 28353 870054
rect 28433 869993 28573 870134
rect 28433 842600 28573 869800
rect 28433 842266 28573 842407
rect 28653 842346 28719 954722
rect 0 827934 28699 842266
rect 0 827600 4843 827854
rect 4923 827793 20920 827934
rect 21000 827600 25993 827854
rect 26073 827793 26213 827934
rect 0 800400 26213 827600
rect 0 800146 4843 800400
rect 4923 800066 20920 800194
rect 21000 800146 25993 800400
rect 26073 800066 26213 800194
rect 26293 800146 27183 827854
rect 27263 827793 27383 827934
rect 27263 800400 27383 827600
rect 27263 800066 27383 800194
rect 27463 800146 28353 827854
rect 28433 827793 28573 827934
rect 28433 800400 28573 827600
rect 28433 800066 28573 800194
rect 0 793738 28573 800066
rect 28653 793818 28719 827854
rect 0 792072 28699 793738
rect 28779 792152 29375 961488
rect 29455 954534 29651 961568
rect 29435 954200 29671 954454
rect 29455 927000 29651 954200
rect 29435 926746 29671 927000
rect 29455 912334 29651 926666
rect 29435 912000 29671 912254
rect 29455 884800 29651 912000
rect 29435 884546 29671 884800
rect 29455 870134 29651 884466
rect 29435 869800 29671 870054
rect 29455 842600 29651 869800
rect 29435 842346 29671 842600
rect 29455 827934 29651 842266
rect 29435 827600 29671 827854
rect 29455 800400 29651 827600
rect 29435 800146 29671 800400
rect 29455 795213 29651 800066
rect 29731 795293 30327 964629
rect 30387 963618 30453 1001515
rect 30533 1001477 40466 1001595
rect 40546 1001557 76454 1002487
rect 76534 1001477 91866 1002567
rect 91946 1001557 127854 1002487
rect 127934 1001477 143266 1002567
rect 143346 1001557 179254 1002487
rect 179334 1001477 194666 1002567
rect 194746 1001557 230654 1002487
rect 230734 1001477 246066 1002567
rect 246146 1001557 282254 1002487
rect 282334 1001477 297666 1002567
rect 297746 1001557 333654 1002487
rect 333734 1001477 348066 1002567
rect 348146 1001557 384054 1002487
rect 384134 1001477 399466 1002567
rect 399546 1001557 473054 1002487
rect 473134 1001477 488466 1002567
rect 488546 1001557 524454 1002487
rect 524534 1001477 539866 1002567
rect 539946 1001557 575854 1002487
rect 575934 1001477 590266 1002567
rect 590346 1001557 626254 1002487
rect 626334 1001477 641666 1002567
rect 641746 1001557 677905 1002487
rect 677985 1002315 717600 1002567
rect 677985 1002262 688801 1002315
rect 677985 1001595 688145 1002262
rect 677985 1001477 687067 1001595
rect 30533 1001357 40549 1001477
rect 76393 1001357 91994 1001477
rect 127793 1001357 143394 1001477
rect 179193 1001357 194794 1001477
rect 230593 1001357 246194 1001477
rect 282193 1001357 297794 1001477
rect 333593 1001357 348207 1001477
rect 383993 1001357 399594 1001477
rect 472993 1001357 488594 1001477
rect 524393 1001357 539994 1001477
rect 575793 1001357 590407 1001477
rect 626193 1001357 641794 1001477
rect 677600 1001357 687067 1001477
rect 30533 1000507 40469 1001357
rect 40549 1000587 76393 1001277
rect 76473 1000507 91914 1001357
rect 91994 1000587 127793 1001277
rect 127873 1000507 143314 1001357
rect 143394 1000587 179193 1001277
rect 179273 1000507 194714 1001357
rect 194794 1000587 230593 1001277
rect 230673 1000507 246114 1001357
rect 246194 1000587 282193 1001277
rect 282273 1000507 297714 1001357
rect 297794 1000587 333593 1001277
rect 333673 1000507 348127 1001357
rect 348207 1000587 383993 1001277
rect 384073 1000507 399514 1001357
rect 399594 1000587 435200 1001277
rect 436200 1000587 472993 1001277
rect 473073 1000507 488514 1001357
rect 488594 1000587 524393 1001277
rect 524473 1000507 539914 1001357
rect 539994 1000587 575793 1001277
rect 575873 1000507 590327 1001357
rect 590407 1000587 626193 1001277
rect 626273 1000507 641714 1001357
rect 641794 1000587 677894 1001277
rect 677974 1000507 687067 1001357
rect 30533 1000387 40549 1000507
rect 76393 1000387 91994 1000507
rect 127793 1000387 143394 1000507
rect 179193 1000387 194794 1000507
rect 230593 1000387 246194 1000507
rect 282193 1000387 297794 1000507
rect 333593 1000387 348207 1000507
rect 383993 1000387 399594 1000507
rect 472993 1000387 488594 1000507
rect 524393 1000387 539994 1000507
rect 575793 1000387 590407 1000507
rect 626193 1000387 641794 1000507
rect 677600 1000387 687067 1000507
rect 30533 999297 40466 1000387
rect 40546 999377 76454 1000307
rect 76534 999297 91866 1000387
rect 91946 999377 127854 1000307
rect 127934 999297 143266 1000387
rect 143346 999377 179254 1000307
rect 179334 999297 194666 1000387
rect 194746 999377 230654 1000307
rect 230734 999297 246066 1000387
rect 246146 999377 282254 1000307
rect 282334 999297 297666 1000387
rect 297746 999377 333654 1000307
rect 333734 999297 348066 1000387
rect 348146 999377 384054 1000307
rect 384134 999297 399466 1000387
rect 399546 999377 436200 1000307
rect 437200 999377 473054 1000307
rect 473134 999297 488466 1000387
rect 488546 999377 524454 1000307
rect 524534 999297 539866 1000387
rect 539946 999377 575854 1000307
rect 575934 999297 590266 1000387
rect 590346 999377 626254 1000307
rect 626334 999297 641666 1000387
rect 641746 999377 678357 1000307
rect 678437 999297 687067 1000387
rect 30533 999177 40549 999297
rect 76393 999177 91994 999297
rect 127793 999177 143394 999297
rect 179193 999177 194794 999297
rect 230593 999177 246194 999297
rect 282193 999177 297794 999297
rect 333593 999177 348207 999297
rect 383993 999177 399594 999297
rect 472993 999177 488594 999297
rect 524393 999177 539994 999297
rect 575793 999177 590407 999297
rect 626193 999177 641794 999297
rect 677600 999177 687067 999297
rect 30533 998437 40466 999177
rect 30533 998000 37213 998437
rect 30533 997975 33823 998000
rect 30533 997600 30673 997975
rect 31763 997957 33823 997975
rect 31763 997947 32853 997957
rect 30533 969866 30673 969994
rect 30753 969946 31683 997895
rect 31763 997600 31883 997947
rect 31763 969866 31883 969994
rect 31963 969946 32653 997867
rect 32733 997600 32853 997947
rect 32733 969866 32853 969994
rect 32933 969946 33623 997877
rect 33703 997600 33823 997957
rect 34913 997985 37213 998000
rect 33703 969866 33823 969994
rect 33903 969946 34833 997920
rect 34913 997600 35033 997985
rect 36123 997974 37213 997985
rect 34913 969866 35033 969994
rect 35113 969946 36043 997905
rect 36123 997600 36243 997974
rect 36323 969994 37013 997894
rect 37093 997600 37213 997974
rect 36123 969914 36243 969994
rect 37093 969914 37213 969994
rect 37293 969946 38223 998357
rect 38303 998150 40466 998437
rect 38303 997600 38423 998150
rect 36123 969866 37213 969914
rect 38303 969866 38423 969994
rect 38503 969946 39593 998070
rect 39673 997927 40466 998150
rect 40546 998007 76454 999097
rect 76534 997927 91866 999177
rect 91946 998007 127854 999097
rect 127934 997927 143266 999177
rect 143346 998007 179254 999097
rect 179334 997927 194666 999177
rect 194746 998007 230654 999097
rect 230734 997927 246066 999177
rect 246146 998007 282254 999097
rect 282334 997927 297666 999177
rect 297746 998007 333654 999097
rect 333734 998007 348066 999177
rect 348146 998007 384054 999097
rect 384134 997927 399466 999177
rect 399546 998007 473054 999097
rect 473134 997927 488466 999177
rect 488546 998007 524454 999097
rect 524534 997927 539866 999177
rect 539946 998007 575854 999097
rect 575934 998007 590266 999177
rect 590346 998007 626254 999097
rect 626334 997927 641666 999177
rect 641746 998007 678070 999097
rect 678150 997927 687067 999177
rect 39673 997600 40549 997927
rect 76393 997707 91994 997927
rect 127793 997707 143394 997927
rect 179193 997707 194794 997927
rect 230593 997707 246194 997927
rect 282193 997707 297794 997927
rect 383993 997707 399594 997927
rect 472993 997707 488594 997927
rect 524393 997707 539994 997927
rect 626193 997707 641794 997927
rect 677600 997134 687067 997927
rect 677600 997051 677927 997134
rect 676259 990180 676325 990181
rect 676259 990116 676260 990180
rect 676324 990116 676325 990180
rect 676259 990115 676325 990116
rect 39673 969866 39893 969994
rect 30533 963538 39893 969866
rect 30407 954802 39893 963538
rect 30387 842346 30453 954722
rect 30533 954534 39893 954802
rect 30533 954393 30673 954534
rect 30533 926666 30673 926807
rect 30753 926746 31683 954454
rect 31763 954393 31883 954534
rect 31763 926666 31883 926807
rect 31963 926746 32653 954454
rect 32733 954393 32853 954534
rect 32733 926666 32853 926807
rect 32933 926746 33623 954454
rect 33703 954393 33823 954534
rect 33703 926666 33823 926807
rect 33903 926746 34833 954454
rect 34913 954393 35033 954534
rect 36123 954473 37213 954534
rect 34913 926666 35033 926807
rect 35113 926746 36043 954454
rect 36123 954393 36243 954473
rect 37093 954393 37213 954473
rect 36323 926807 37013 954393
rect 36123 926727 36243 926807
rect 37093 926727 37213 926807
rect 37293 926746 38223 954454
rect 38303 954393 38423 954534
rect 36123 926666 37213 926727
rect 38303 926666 38423 926807
rect 38503 926746 39593 954454
rect 39673 954393 39893 954534
rect 30533 912334 39593 926666
rect 30533 912193 30673 912334
rect 30533 884466 30673 884607
rect 30753 884546 31683 912254
rect 31763 912193 31883 912334
rect 31763 884466 31883 884607
rect 31963 884546 32653 912254
rect 32733 912193 32853 912334
rect 32733 884466 32853 884607
rect 32933 884546 33623 912254
rect 33703 912193 33823 912334
rect 33703 884466 33823 884607
rect 33903 884546 34833 912254
rect 34913 912193 35033 912334
rect 36123 912273 37213 912334
rect 34913 884466 35033 884607
rect 35113 884546 36043 912254
rect 36123 912193 36243 912273
rect 37093 912193 37213 912273
rect 36323 884607 37013 912193
rect 36123 884527 36243 884607
rect 37093 884527 37213 884607
rect 37293 884546 38223 912254
rect 38303 912193 38423 912334
rect 36123 884466 37213 884527
rect 38303 884466 38423 884607
rect 38503 884546 39593 912254
rect 40539 908172 40605 908173
rect 40539 908108 40540 908172
rect 40604 908108 40605 908172
rect 40539 908107 40605 908108
rect 40542 908037 40602 908107
rect 40539 908036 40605 908037
rect 40539 907972 40540 908036
rect 40604 907972 40605 908036
rect 40539 907971 40605 907972
rect 676262 907765 676322 990115
rect 677707 967266 677927 967407
rect 678007 967346 679097 997054
rect 679177 997051 679297 997134
rect 680387 997131 681477 997134
rect 679177 967266 679297 967407
rect 679377 967346 680307 997054
rect 680387 997051 680507 997131
rect 681357 997051 681477 997131
rect 680587 967407 681277 997051
rect 680387 967327 680507 967407
rect 681357 967327 681477 967407
rect 681557 967346 682487 997054
rect 682567 997051 682687 997134
rect 680387 967266 681477 967327
rect 682567 967266 682687 967407
rect 682767 967346 683697 997054
rect 683777 997051 683897 997134
rect 683777 967266 683897 967407
rect 683977 967346 684667 997054
rect 684747 997051 684867 997134
rect 684747 967266 684867 967407
rect 684947 967346 685637 997054
rect 685717 997051 685837 997134
rect 685717 967266 685837 967407
rect 685917 967346 686847 997054
rect 686927 997051 687067 997134
rect 686927 967266 687067 967407
rect 677707 966998 687067 967266
rect 687147 967078 687213 1001515
rect 687293 1001191 688145 1001595
rect 687293 1001055 687849 1001191
rect 677707 958262 687193 966998
rect 677707 951934 687067 958262
rect 677707 951806 677927 951934
rect 678007 922346 679097 951854
rect 679177 951806 679297 951934
rect 680387 951886 681477 951934
rect 679177 922266 679297 922407
rect 679377 922346 680307 951854
rect 680387 951806 680507 951886
rect 681357 951806 681477 951886
rect 680587 922407 681277 951806
rect 680387 922327 680507 922407
rect 681357 922327 681477 922407
rect 681557 922346 682487 951854
rect 682567 951806 682687 951934
rect 680387 922266 681477 922327
rect 682567 922266 682687 922407
rect 682767 922346 683697 951854
rect 683777 951806 683897 951934
rect 683777 922266 683897 922407
rect 683977 922346 684667 951854
rect 684747 951806 684867 951934
rect 684747 922266 684867 922407
rect 684947 922346 685637 951854
rect 685717 951806 685837 951934
rect 685717 922266 685837 922407
rect 685917 922346 686847 951854
rect 686927 951806 687067 951934
rect 686927 922266 687067 922407
rect 677547 918644 677613 918645
rect 677547 918580 677548 918644
rect 677612 918580 677613 918644
rect 677547 918579 677613 918580
rect 676259 907764 676325 907765
rect 676259 907700 676260 907764
rect 676324 907700 676325 907764
rect 676259 907699 676325 907700
rect 40355 888860 40421 888861
rect 40355 888796 40356 888860
rect 40420 888796 40421 888860
rect 40355 888795 40421 888796
rect 30533 870134 39593 884466
rect 40358 874850 40418 888795
rect 39990 874790 40418 874850
rect 30533 869993 30673 870134
rect 30533 842266 30673 842407
rect 30753 842346 31683 870054
rect 31763 869993 31883 870134
rect 31763 842266 31883 842407
rect 31963 842346 32653 870054
rect 32733 869993 32853 870134
rect 32733 842266 32853 842407
rect 32933 842346 33623 870054
rect 33703 869993 33823 870134
rect 33703 842266 33823 842407
rect 33903 842346 34833 870054
rect 34913 869993 35033 870134
rect 36123 870073 37213 870134
rect 34913 842266 35033 842407
rect 35113 842346 36043 870054
rect 36123 869993 36243 870073
rect 37093 869993 37213 870073
rect 36323 842407 37013 869993
rect 36123 842327 36243 842407
rect 37093 842327 37213 842407
rect 37293 842346 38223 870054
rect 38303 869993 38423 870134
rect 36123 842266 37213 842327
rect 38303 842266 38423 842407
rect 38503 842346 39593 870054
rect 39990 855813 40050 874790
rect 39987 855812 40053 855813
rect 39987 855748 39988 855812
rect 40052 855748 40053 855812
rect 39987 855747 40053 855748
rect 39803 855540 39869 855541
rect 39803 855476 39804 855540
rect 39868 855476 39869 855540
rect 39803 855475 39869 855476
rect 30407 827934 39593 842266
rect 39806 837589 39866 855475
rect 39803 837588 39869 837589
rect 39803 837524 39804 837588
rect 39868 837524 39869 837588
rect 39803 837523 39869 837524
rect 39987 832692 40053 832693
rect 39987 832628 39988 832692
rect 40052 832628 40053 832692
rect 39987 832627 40053 832628
rect 29455 794909 30307 795213
rect 29455 792072 29651 794909
rect 0 791768 29651 792072
rect 0 785002 28699 791768
rect 0 784734 28573 785002
rect 0 784400 4843 784654
rect 4923 784593 20920 784734
rect 21000 784400 25993 784654
rect 26073 784593 26213 784734
rect 0 757200 26213 784400
rect 0 756946 4843 757200
rect 4923 756866 20920 756994
rect 21000 756946 25993 757200
rect 26073 756866 26213 756994
rect 26293 756946 27183 784654
rect 27263 784593 27383 784734
rect 27263 757200 27383 784400
rect 27263 756866 27383 756994
rect 27463 756946 28353 784654
rect 28433 784593 28573 784734
rect 28433 757200 28573 784400
rect 28433 756866 28573 756994
rect 0 750538 28573 756866
rect 28653 750618 28719 784922
rect 0 748872 28699 750538
rect 28779 748952 29375 791688
rect 29455 784734 29651 791768
rect 29435 784400 29671 784654
rect 29455 757200 29651 784400
rect 29435 756946 29671 757200
rect 29455 752013 29651 756866
rect 29731 752093 30327 794829
rect 30387 793818 30453 827854
rect 30533 827793 30673 827934
rect 30533 800066 30673 800194
rect 30753 800146 31683 827854
rect 31763 827793 31883 827934
rect 31763 800066 31883 800194
rect 31963 800146 32653 827854
rect 32733 827793 32853 827934
rect 32733 800066 32853 800194
rect 32933 800146 33623 827854
rect 33703 827793 33823 827934
rect 33703 800066 33823 800194
rect 33903 800146 34833 827854
rect 34913 827793 35033 827934
rect 36123 827873 37213 827934
rect 34913 800066 35033 800194
rect 35113 800146 36043 827854
rect 36123 827793 36243 827873
rect 37093 827793 37213 827873
rect 36323 800194 37013 827793
rect 36123 800114 36243 800194
rect 37093 800114 37213 800194
rect 37293 800146 38223 827854
rect 38303 827793 38423 827934
rect 36123 800066 37213 800114
rect 38303 800066 38423 800194
rect 38503 800146 39593 827854
rect 39990 817050 40050 832627
rect 39990 816990 40418 817050
rect 39673 800066 39893 800194
rect 30533 793738 39893 800066
rect 40358 797741 40418 816990
rect 40355 797740 40421 797741
rect 40355 797676 40356 797740
rect 40420 797676 40421 797740
rect 40355 797675 40421 797676
rect 40355 797604 40421 797605
rect 40355 797540 40356 797604
rect 40420 797540 40421 797604
rect 40355 797539 40421 797540
rect 30407 785002 39893 793738
rect 40358 792165 40418 797539
rect 40355 792164 40421 792165
rect 40355 792100 40356 792164
rect 40420 792100 40421 792164
rect 40355 792099 40421 792100
rect 40539 792164 40605 792165
rect 40539 792100 40540 792164
rect 40604 792100 40605 792164
rect 40539 792099 40605 792100
rect 29455 751709 30307 752013
rect 29455 748872 29651 751709
rect 0 748568 29651 748872
rect 0 741802 28699 748568
rect 0 741534 28573 741802
rect 0 741200 4843 741454
rect 4923 741393 20920 741534
rect 21000 741200 25993 741454
rect 26073 741393 26213 741534
rect 0 714000 26213 741200
rect 0 713746 4843 714000
rect 4923 713666 20920 713794
rect 21000 713746 25993 714000
rect 26073 713666 26213 713794
rect 26293 713746 27183 741454
rect 27263 741393 27383 741534
rect 27263 714000 27383 741200
rect 27263 713666 27383 713794
rect 27463 713746 28353 741454
rect 28433 741393 28573 741534
rect 28433 714000 28573 741200
rect 28433 713666 28573 713794
rect 0 707338 28573 713666
rect 28653 707418 28719 741722
rect 0 705672 28699 707338
rect 28779 705752 29375 748488
rect 29455 741534 29651 748568
rect 29435 741200 29671 741454
rect 29455 714000 29651 741200
rect 29435 713746 29671 714000
rect 29455 708813 29651 713666
rect 29731 708893 30327 751629
rect 30387 750618 30453 784922
rect 30533 784734 39893 785002
rect 30533 784593 30673 784734
rect 30533 756866 30673 756994
rect 30753 756946 31683 784654
rect 31763 784593 31883 784734
rect 31763 756866 31883 756994
rect 31963 756946 32653 784654
rect 32733 784593 32853 784734
rect 32733 756866 32853 756994
rect 32933 756946 33623 784654
rect 33703 784593 33823 784734
rect 33703 756866 33823 756994
rect 33903 756946 34833 784654
rect 34913 784593 35033 784734
rect 36123 784673 37213 784734
rect 34913 756866 35033 756994
rect 35113 756946 36043 784654
rect 36123 784593 36243 784673
rect 37093 784593 37213 784673
rect 36323 756994 37013 784593
rect 36123 756914 36243 756994
rect 37093 756914 37213 756994
rect 37293 756946 38223 784654
rect 38303 784593 38423 784734
rect 36123 756866 37213 756914
rect 38303 756866 38423 756994
rect 38503 756946 39593 784654
rect 39673 784593 39893 784734
rect 40542 778565 40602 792099
rect 40539 778564 40605 778565
rect 40539 778500 40540 778564
rect 40604 778500 40605 778564
rect 40539 778499 40605 778500
rect 40355 778292 40421 778293
rect 40355 778228 40356 778292
rect 40420 778228 40421 778292
rect 40355 778227 40421 778228
rect 40358 763197 40418 778227
rect 40355 763196 40421 763197
rect 40355 763132 40356 763196
rect 40420 763132 40421 763196
rect 40355 763131 40421 763132
rect 40723 763196 40789 763197
rect 40723 763132 40724 763196
rect 40788 763132 40789 763196
rect 40723 763131 40789 763132
rect 39673 756866 39893 756994
rect 30533 750538 39893 756866
rect 40726 753541 40786 763131
rect 40355 753540 40421 753541
rect 40355 753476 40356 753540
rect 40420 753476 40421 753540
rect 40355 753475 40421 753476
rect 40723 753540 40789 753541
rect 40723 753476 40724 753540
rect 40788 753476 40789 753540
rect 40723 753475 40789 753476
rect 40358 750685 40418 753475
rect 40355 750684 40421 750685
rect 40355 750620 40356 750684
rect 40420 750620 40421 750684
rect 40355 750619 40421 750620
rect 30407 741802 39893 750538
rect 40355 750412 40421 750413
rect 40355 750410 40356 750412
rect 29455 708509 30307 708813
rect 29455 705672 29651 708509
rect 0 705368 29651 705672
rect 0 698602 28699 705368
rect 0 698334 28573 698602
rect 0 698000 4843 698254
rect 4923 698193 20920 698334
rect 21000 698000 25993 698254
rect 26073 698193 26213 698334
rect 0 670800 26213 698000
rect 0 670546 4843 670800
rect 4923 670466 20920 670594
rect 21000 670546 25993 670800
rect 26073 670466 26213 670594
rect 26293 670546 27183 698254
rect 27263 698193 27383 698334
rect 27263 670800 27383 698000
rect 27263 670466 27383 670594
rect 27463 670546 28353 698254
rect 28433 698193 28573 698334
rect 28433 670800 28573 698000
rect 28433 670466 28573 670594
rect 0 664138 28573 670466
rect 28653 664218 28719 698522
rect 0 662472 28699 664138
rect 28779 662552 29375 705288
rect 29455 698334 29651 705368
rect 29435 698000 29671 698254
rect 29455 670800 29651 698000
rect 29435 670546 29671 670800
rect 29455 665613 29651 670466
rect 29731 665693 30327 708429
rect 30387 707418 30453 741722
rect 30533 741534 39893 741802
rect 30533 741393 30673 741534
rect 30533 713666 30673 713794
rect 30753 713746 31683 741454
rect 31763 741393 31883 741534
rect 31763 713666 31883 713794
rect 31963 713746 32653 741454
rect 32733 741393 32853 741534
rect 32733 713666 32853 713794
rect 32933 713746 33623 741454
rect 33703 741393 33823 741534
rect 33703 713666 33823 713794
rect 33903 713746 34833 741454
rect 34913 741393 35033 741534
rect 36123 741473 37213 741534
rect 34913 713666 35033 713794
rect 35113 713746 36043 741454
rect 36123 741393 36243 741473
rect 37093 741393 37213 741473
rect 36323 713794 37013 741393
rect 36123 713714 36243 713794
rect 37093 713714 37213 713794
rect 37293 713746 38223 741454
rect 38303 741393 38423 741534
rect 36123 713666 37213 713714
rect 38303 713666 38423 713794
rect 38503 713746 39593 741454
rect 39673 741393 39893 741534
rect 40174 750350 40356 750410
rect 40174 731373 40234 750350
rect 40355 750348 40356 750350
rect 40420 750348 40421 750412
rect 40355 750347 40421 750348
rect 40171 731372 40237 731373
rect 40171 731308 40172 731372
rect 40236 731308 40237 731372
rect 40171 731307 40237 731308
rect 40723 731236 40789 731237
rect 40723 731172 40724 731236
rect 40788 731172 40789 731236
rect 40723 731171 40789 731172
rect 39673 713666 39893 713794
rect 30533 707338 39893 713666
rect 40726 712333 40786 731171
rect 40355 712332 40421 712333
rect 40355 712330 40356 712332
rect 30407 698602 39893 707338
rect 40174 712270 40356 712330
rect 40174 702130 40234 712270
rect 40355 712268 40356 712270
rect 40420 712268 40421 712332
rect 40355 712267 40421 712268
rect 40723 712332 40789 712333
rect 40723 712268 40724 712332
rect 40788 712268 40789 712332
rect 40723 712267 40789 712268
rect 40355 702132 40421 702133
rect 40355 702130 40356 702132
rect 40174 702070 40356 702130
rect 40355 702068 40356 702070
rect 40420 702068 40421 702132
rect 40355 702067 40421 702068
rect 40907 702132 40973 702133
rect 40907 702068 40908 702132
rect 40972 702068 40973 702132
rect 40907 702067 40973 702068
rect 29455 665309 30307 665613
rect 29455 662472 29651 665309
rect 0 662168 29651 662472
rect 0 655402 28699 662168
rect 0 655134 28573 655402
rect 0 654800 4843 655054
rect 4923 654993 20920 655134
rect 21000 654800 25993 655054
rect 26073 654993 26213 655134
rect 0 627600 26213 654800
rect 0 627346 4843 627600
rect 4923 627266 20920 627394
rect 21000 627346 25993 627600
rect 26073 627266 26213 627394
rect 26293 627346 27183 655054
rect 27263 654993 27383 655134
rect 27263 627600 27383 654800
rect 27263 627266 27383 627394
rect 27463 627346 28353 655054
rect 28433 654993 28573 655134
rect 28433 627600 28573 654800
rect 28433 627266 28573 627394
rect 0 620938 28573 627266
rect 28653 621018 28719 655322
rect 0 619272 28699 620938
rect 28779 619352 29375 662088
rect 29455 655134 29651 662168
rect 29435 654800 29671 655054
rect 29455 627600 29651 654800
rect 29435 627346 29671 627600
rect 29455 622413 29651 627266
rect 29731 622493 30327 665229
rect 30387 664218 30453 698522
rect 30533 698334 39893 698602
rect 30533 698193 30673 698334
rect 30533 670466 30673 670594
rect 30753 670546 31683 698254
rect 31763 698193 31883 698334
rect 31763 670466 31883 670594
rect 31963 670546 32653 698254
rect 32733 698193 32853 698334
rect 32733 670466 32853 670594
rect 32933 670546 33623 698254
rect 33703 698193 33823 698334
rect 33703 670466 33823 670594
rect 33903 670546 34833 698254
rect 34913 698193 35033 698334
rect 36123 698273 37213 698334
rect 34913 670466 35033 670594
rect 35113 670546 36043 698254
rect 36123 698193 36243 698273
rect 37093 698193 37213 698273
rect 36323 670594 37013 698193
rect 36123 670514 36243 670594
rect 37093 670514 37213 670594
rect 37293 670546 38223 698254
rect 38303 698193 38423 698334
rect 36123 670466 37213 670514
rect 38303 670466 38423 670594
rect 38503 670546 39593 698254
rect 39673 698193 39893 698334
rect 40910 695333 40970 702067
rect 40539 695332 40605 695333
rect 40539 695268 40540 695332
rect 40604 695268 40605 695332
rect 40539 695267 40605 695268
rect 40907 695332 40973 695333
rect 40907 695268 40908 695332
rect 40972 695268 40973 695332
rect 40907 695267 40973 695268
rect 40542 676290 40602 695267
rect 40174 676230 40602 676290
rect 40174 673437 40234 676230
rect 40171 673436 40237 673437
rect 40171 673372 40172 673436
rect 40236 673372 40237 673436
rect 40171 673371 40237 673372
rect 40539 673436 40605 673437
rect 40539 673372 40540 673436
rect 40604 673372 40605 673436
rect 40539 673371 40605 673372
rect 39673 670466 39893 670594
rect 30533 664138 39893 670466
rect 30407 655402 39893 664138
rect 29455 622109 30307 622413
rect 29455 619272 29651 622109
rect 0 618968 29651 619272
rect 0 612202 28699 618968
rect 0 611934 28573 612202
rect 0 611600 4843 611854
rect 4923 611793 20920 611934
rect 21000 611600 25993 611854
rect 26073 611793 26213 611934
rect 0 584400 26213 611600
rect 0 584146 4843 584400
rect 4923 584066 20920 584194
rect 21000 584146 25993 584400
rect 26073 584066 26213 584194
rect 26293 584146 27183 611854
rect 27263 611793 27383 611934
rect 27263 584400 27383 611600
rect 27263 584066 27383 584194
rect 27463 584146 28353 611854
rect 28433 611793 28573 611934
rect 28433 584400 28573 611600
rect 28433 584066 28573 584194
rect 0 577738 28573 584066
rect 28653 577818 28719 612122
rect 0 576072 28699 577738
rect 28779 576152 29375 618888
rect 29455 611934 29651 618968
rect 29435 611600 29671 611854
rect 29455 584400 29651 611600
rect 29435 584146 29671 584400
rect 29455 579213 29651 584066
rect 29731 579293 30327 622029
rect 30387 621018 30453 655322
rect 30533 655134 39893 655402
rect 30533 654993 30673 655134
rect 30533 627266 30673 627394
rect 30753 627346 31683 655054
rect 31763 654993 31883 655134
rect 31763 627266 31883 627394
rect 31963 627346 32653 655054
rect 32733 654993 32853 655134
rect 32733 627266 32853 627394
rect 32933 627346 33623 655054
rect 33703 654993 33823 655134
rect 33703 627266 33823 627394
rect 33903 627346 34833 655054
rect 34913 654993 35033 655134
rect 36123 655073 37213 655134
rect 34913 627266 35033 627394
rect 35113 627346 36043 655054
rect 36123 654993 36243 655073
rect 37093 654993 37213 655073
rect 36323 627394 37013 654993
rect 36123 627314 36243 627394
rect 37093 627314 37213 627394
rect 37293 627346 38223 655054
rect 38303 654993 38423 655134
rect 36123 627266 37213 627314
rect 38303 627266 38423 627394
rect 38503 627346 39593 655054
rect 39673 654993 39893 655134
rect 40542 654397 40602 673371
rect 40539 654396 40605 654397
rect 40539 654332 40540 654396
rect 40604 654332 40605 654396
rect 40539 654331 40605 654332
rect 40171 654260 40237 654261
rect 40171 654196 40172 654260
rect 40236 654196 40237 654260
rect 40171 654195 40237 654196
rect 40174 642970 40234 654195
rect 39990 642910 40234 642970
rect 39990 637530 40050 642910
rect 39990 637470 40418 637530
rect 40358 634813 40418 637470
rect 40355 634812 40421 634813
rect 40355 634748 40356 634812
rect 40420 634748 40421 634812
rect 40355 634747 40421 634748
rect 40907 634812 40973 634813
rect 40907 634748 40908 634812
rect 40972 634748 40973 634812
rect 40907 634747 40973 634748
rect 39673 627266 39893 627394
rect 30533 620938 39893 627266
rect 30407 612202 39893 620938
rect 29455 578909 30307 579213
rect 29455 576072 29651 578909
rect 0 575768 29651 576072
rect 0 569002 28699 575768
rect 0 568734 28573 569002
rect 0 568400 4843 568654
rect 4923 568593 20920 568734
rect 21000 568400 25993 568654
rect 26073 568593 26213 568734
rect 0 541200 26213 568400
rect 0 540946 4843 541200
rect 4923 540866 20920 540994
rect 21000 540946 25993 541200
rect 26073 540866 26213 540994
rect 26293 540946 27183 568654
rect 27263 568593 27383 568734
rect 27263 541200 27383 568400
rect 27263 540866 27383 540994
rect 27463 540946 28353 568654
rect 28433 568593 28573 568734
rect 28433 541200 28573 568400
rect 28433 540866 28573 540994
rect 0 534538 28573 540866
rect 28653 534618 28719 568922
rect 0 532872 28699 534538
rect 28779 532952 29375 575688
rect 29455 568734 29651 575768
rect 29435 568400 29671 568654
rect 29455 541200 29651 568400
rect 29435 540946 29671 541200
rect 29455 536013 29651 540866
rect 29731 536093 30327 578829
rect 30387 577818 30453 612122
rect 30533 611934 39893 612202
rect 30533 611793 30673 611934
rect 30533 584066 30673 584194
rect 30753 584146 31683 611854
rect 31763 611793 31883 611934
rect 31763 584066 31883 584194
rect 31963 584146 32653 611854
rect 32733 611793 32853 611934
rect 32733 584066 32853 584194
rect 32933 584146 33623 611854
rect 33703 611793 33823 611934
rect 33703 584066 33823 584194
rect 33903 584146 34833 611854
rect 34913 611793 35033 611934
rect 36123 611873 37213 611934
rect 34913 584066 35033 584194
rect 35113 584146 36043 611854
rect 36123 611793 36243 611873
rect 37093 611793 37213 611873
rect 36323 584194 37013 611793
rect 36123 584114 36243 584194
rect 37093 584114 37213 584194
rect 37293 584146 38223 611854
rect 38303 611793 38423 611934
rect 36123 584066 37213 584114
rect 38303 584066 38423 584194
rect 38503 584146 39593 611854
rect 39673 611793 39893 611934
rect 40910 599045 40970 634747
rect 40539 599044 40605 599045
rect 40539 598980 40540 599044
rect 40604 598980 40605 599044
rect 40539 598979 40605 598980
rect 40907 599044 40973 599045
rect 40907 598980 40908 599044
rect 40972 598980 40973 599044
rect 40907 598979 40973 598980
rect 40542 585170 40602 598979
rect 40174 585110 40602 585170
rect 39673 584066 39893 584194
rect 30533 577738 39893 584066
rect 30407 569002 39893 577738
rect 29455 535709 30307 536013
rect 29455 532872 29651 535709
rect 0 532568 29651 532872
rect 0 525802 28699 532568
rect 0 525534 28573 525802
rect 0 525200 4843 525454
rect 4923 525393 20920 525534
rect 21000 525200 25993 525454
rect 26073 525393 26213 525534
rect 0 498000 26213 525200
rect 0 497746 4843 498000
rect 4923 497666 20920 497807
rect 21000 497746 25993 498000
rect 26073 497666 26213 497807
rect 26293 497746 27183 525454
rect 27263 525393 27383 525534
rect 27263 498000 27383 525200
rect 27263 497666 27383 497807
rect 27463 497746 28353 525454
rect 28433 525393 28573 525534
rect 28433 498000 28573 525200
rect 28433 497666 28573 497807
rect 0 483334 28573 497666
rect 0 483000 4843 483254
rect 4923 483193 20920 483334
rect 21000 483000 25993 483254
rect 26073 483193 26213 483334
rect 0 455800 26213 483000
rect 0 455546 4843 455800
rect 4923 455466 20920 455607
rect 21000 455546 25993 455800
rect 26073 455466 26213 455607
rect 26293 455546 27183 483254
rect 27263 483193 27383 483334
rect 27263 455800 27383 483000
rect 27263 455466 27383 455607
rect 27463 455546 28353 483254
rect 28433 483193 28573 483334
rect 28433 455800 28573 483000
rect 28433 455466 28573 455607
rect 0 441134 28573 455466
rect 0 440800 4843 441054
rect 4923 440993 20920 441134
rect 21000 440800 25993 441054
rect 26073 440993 26213 441134
rect 0 413600 26213 440800
rect 0 413346 4843 413600
rect 4923 413266 20920 413394
rect 21000 413346 25993 413600
rect 26073 413266 26213 413394
rect 26293 413346 27183 441054
rect 27263 440993 27383 441134
rect 27263 413600 27383 440800
rect 27263 413266 27383 413394
rect 27463 413346 28353 441054
rect 28433 440993 28573 441134
rect 28433 413600 28573 440800
rect 28433 413266 28573 413394
rect 0 406938 28573 413266
rect 28653 407018 28719 525722
rect 0 405272 28699 406938
rect 28779 405352 29375 532488
rect 29455 525534 29651 532568
rect 29435 525200 29671 525454
rect 29455 498000 29651 525200
rect 29435 497746 29671 498000
rect 29455 483334 29651 497666
rect 29435 483000 29671 483254
rect 29455 455800 29651 483000
rect 29435 455546 29671 455800
rect 29455 441134 29651 455466
rect 29435 440800 29671 441054
rect 29455 413600 29651 440800
rect 29435 413346 29671 413600
rect 29455 408413 29651 413266
rect 29731 408493 30327 535629
rect 30387 534618 30453 568922
rect 30533 568734 39893 569002
rect 30533 568593 30673 568734
rect 30533 540866 30673 540994
rect 30753 540946 31683 568654
rect 31763 568593 31883 568734
rect 31763 540866 31883 540994
rect 31963 540946 32653 568654
rect 32733 568593 32853 568734
rect 32733 540866 32853 540994
rect 32933 540946 33623 568654
rect 33703 568593 33823 568734
rect 33703 540866 33823 540994
rect 33903 540946 34833 568654
rect 34913 568593 35033 568734
rect 36123 568673 37213 568734
rect 34913 540866 35033 540994
rect 35113 540946 36043 568654
rect 36123 568593 36243 568673
rect 37093 568593 37213 568673
rect 36323 540994 37013 568593
rect 36123 540914 36243 540994
rect 37093 540914 37213 540994
rect 37293 540946 38223 568654
rect 38303 568593 38423 568734
rect 36123 540866 37213 540914
rect 38303 540866 38423 540994
rect 38503 540946 39593 568654
rect 39673 568593 39893 568734
rect 40174 565997 40234 585110
rect 40171 565996 40237 565997
rect 40171 565932 40172 565996
rect 40236 565932 40237 565996
rect 40171 565931 40237 565932
rect 40171 565724 40237 565725
rect 40171 565660 40172 565724
rect 40236 565660 40237 565724
rect 40171 565659 40237 565660
rect 40174 550629 40234 565659
rect 40171 550628 40237 550629
rect 40171 550564 40172 550628
rect 40236 550564 40237 550628
rect 40171 550563 40237 550564
rect 40539 550628 40605 550629
rect 40539 550564 40540 550628
rect 40604 550564 40605 550628
rect 40539 550563 40605 550564
rect 39673 540866 39893 540994
rect 40542 540973 40602 550563
rect 40539 540972 40605 540973
rect 40539 540908 40540 540972
rect 40604 540908 40605 540972
rect 40539 540907 40605 540908
rect 40907 540972 40973 540973
rect 40907 540908 40908 540972
rect 40972 540908 40973 540972
rect 40907 540907 40973 540908
rect 30533 534538 39893 540866
rect 30407 525802 39893 534538
rect 29455 408109 30307 408413
rect 29455 405272 29651 408109
rect 0 404968 29651 405272
rect 0 398202 28699 404968
rect 0 397934 28573 398202
rect 0 397600 4843 397854
rect 4923 397793 20920 397934
rect 21000 397600 25993 397854
rect 26073 397793 26213 397934
rect 0 370400 26213 397600
rect 0 370146 4843 370400
rect 4923 370066 20920 370194
rect 21000 370146 25993 370400
rect 26073 370066 26213 370194
rect 26293 370146 27183 397854
rect 27263 397793 27383 397934
rect 27263 370400 27383 397600
rect 27263 370066 27383 370194
rect 27463 370146 28353 397854
rect 28433 397793 28573 397934
rect 28433 370400 28573 397600
rect 28433 370066 28573 370194
rect 0 363738 28573 370066
rect 28653 363818 28719 398122
rect 0 362072 28699 363738
rect 28779 362152 29375 404888
rect 29455 397934 29651 404968
rect 29435 397600 29671 397854
rect 29455 370400 29651 397600
rect 29435 370146 29671 370400
rect 29455 365213 29651 370066
rect 29731 365293 30327 408029
rect 30387 407018 30453 525722
rect 30533 525534 39893 525802
rect 30533 525393 30673 525534
rect 30533 497666 30673 497807
rect 30753 497746 31683 525454
rect 31763 525393 31883 525534
rect 31763 497666 31883 497807
rect 31963 497746 32653 525454
rect 32733 525393 32853 525534
rect 32733 497666 32853 497807
rect 32933 497746 33623 525454
rect 33703 525393 33823 525534
rect 33703 497666 33823 497807
rect 33903 497746 34833 525454
rect 34913 525393 35033 525534
rect 36123 525473 37213 525534
rect 34913 497666 35033 497807
rect 35113 497746 36043 525454
rect 36123 525393 36243 525473
rect 37093 525393 37213 525473
rect 36323 497807 37013 525393
rect 36123 497727 36243 497807
rect 37093 497727 37213 497807
rect 37293 497746 38223 525454
rect 38303 525393 38423 525534
rect 36123 497666 37213 497727
rect 38303 497666 38423 497807
rect 38503 497746 39593 525454
rect 39673 525393 39893 525534
rect 40910 521933 40970 540907
rect 40907 521932 40973 521933
rect 40907 521868 40908 521932
rect 40972 521868 40973 521932
rect 40907 521867 40973 521868
rect 40171 521796 40237 521797
rect 40171 521732 40172 521796
rect 40236 521732 40237 521796
rect 40171 521731 40237 521732
rect 40174 508061 40234 521731
rect 40171 508060 40237 508061
rect 40171 507996 40172 508060
rect 40236 507996 40237 508060
rect 40171 507995 40237 507996
rect 39987 507788 40053 507789
rect 39987 507724 39988 507788
rect 40052 507724 40053 507788
rect 39987 507723 40053 507724
rect 30533 483334 39593 497666
rect 39990 488610 40050 507723
rect 39990 488550 40234 488610
rect 30533 483193 30673 483334
rect 30533 455466 30673 455607
rect 30753 455546 31683 483254
rect 31763 483193 31883 483334
rect 31763 455466 31883 455607
rect 31963 455546 32653 483254
rect 32733 483193 32853 483334
rect 32733 455466 32853 455607
rect 32933 455546 33623 483254
rect 33703 483193 33823 483334
rect 33703 455466 33823 455607
rect 33903 455546 34833 483254
rect 34913 483193 35033 483334
rect 36123 483273 37213 483334
rect 34913 455466 35033 455607
rect 35113 455546 36043 483254
rect 36123 483193 36243 483273
rect 37093 483193 37213 483273
rect 36323 455607 37013 483193
rect 36123 455527 36243 455607
rect 37093 455527 37213 455607
rect 37293 455546 38223 483254
rect 38303 483193 38423 483334
rect 36123 455466 37213 455527
rect 38303 455466 38423 455607
rect 38503 455546 39593 483254
rect 30533 441134 39593 455466
rect 40174 455429 40234 488550
rect 677550 477597 677610 918579
rect 678007 907934 687067 922266
rect 677707 878066 677927 878207
rect 678007 878146 679097 907854
rect 679177 907793 679297 907934
rect 680387 907873 681477 907934
rect 679177 878066 679297 878207
rect 679377 878146 680307 907854
rect 680387 907793 680507 907873
rect 681357 907793 681477 907873
rect 680587 878207 681277 907793
rect 680387 878127 680507 878207
rect 681357 878127 681477 878207
rect 681557 878146 682487 907854
rect 682567 907793 682687 907934
rect 680387 878066 681477 878127
rect 682567 878066 682687 878207
rect 682767 878146 683697 907854
rect 683777 907793 683897 907934
rect 683777 878066 683897 878207
rect 683977 878146 684667 907854
rect 684747 907793 684867 907934
rect 684747 878066 684867 878207
rect 684947 878146 685637 907854
rect 685717 907793 685837 907934
rect 685717 878066 685837 878207
rect 685917 878146 686847 907854
rect 686927 907793 687067 907934
rect 686927 878066 687067 878207
rect 677707 877798 687067 878066
rect 687147 877878 687213 958182
rect 687273 957171 687869 1000975
rect 687929 996800 688165 1001111
rect 687949 967600 688145 996800
rect 687929 967346 688165 967600
rect 687949 960232 688145 967266
rect 688225 960312 688821 1002182
rect 688881 967078 688947 1002235
rect 689027 997251 717600 1002315
rect 689027 997134 691527 997251
rect 689027 997051 689167 997134
rect 689027 967600 689167 996800
rect 689027 967266 689167 967407
rect 689247 967346 690137 997054
rect 690217 997051 690337 997134
rect 690217 967600 690337 996800
rect 690217 967266 690337 967407
rect 690417 967346 691307 997054
rect 691387 997051 691527 997134
rect 691607 996800 696600 997171
rect 696680 997134 717600 997251
rect 696680 997051 712677 997134
rect 712757 996800 717600 997054
rect 691387 967600 717600 996800
rect 691387 967266 691527 967407
rect 691607 967346 696600 967600
rect 696680 967266 712677 967407
rect 712757 967346 717600 967600
rect 689027 966998 717600 967266
rect 688901 960232 717600 966998
rect 687949 959928 717600 960232
rect 687949 957091 688145 959928
rect 687293 956787 688145 957091
rect 677707 869062 687193 877798
rect 677707 862734 687067 869062
rect 677707 862606 677927 862734
rect 678007 833146 679097 862654
rect 679177 862606 679297 862734
rect 680387 862686 681477 862734
rect 679177 833066 679297 833207
rect 679377 833146 680307 862654
rect 680387 862606 680507 862686
rect 681357 862606 681477 862686
rect 680587 833207 681277 862606
rect 680387 833127 680507 833207
rect 681357 833127 681477 833207
rect 681557 833146 682487 862654
rect 682567 862606 682687 862734
rect 680387 833066 681477 833127
rect 682567 833066 682687 833207
rect 682767 833146 683697 862654
rect 683777 862606 683897 862734
rect 683777 833066 683897 833207
rect 683977 833146 684667 862654
rect 684747 862606 684867 862734
rect 684747 833066 684867 833207
rect 684947 833146 685637 862654
rect 685717 862606 685837 862734
rect 685717 833066 685837 833207
rect 685917 833146 686847 862654
rect 686927 862606 687067 862734
rect 686927 833066 687067 833207
rect 678007 818734 687067 833066
rect 677707 788866 677927 789007
rect 678007 788946 679097 818654
rect 679177 818593 679297 818734
rect 680387 818673 681477 818734
rect 679177 788866 679297 789007
rect 679377 788946 680307 818654
rect 680387 818593 680507 818673
rect 681357 818593 681477 818673
rect 680587 789007 681277 818593
rect 680387 788927 680507 789007
rect 681357 788927 681477 789007
rect 681557 788946 682487 818654
rect 682567 818593 682687 818734
rect 680387 788866 681477 788927
rect 682567 788866 682687 789007
rect 682767 788946 683697 818654
rect 683777 818593 683897 818734
rect 683777 788866 683897 789007
rect 683977 788946 684667 818654
rect 684747 818593 684867 818734
rect 684747 788866 684867 789007
rect 684947 788946 685637 818654
rect 685717 818593 685837 818734
rect 685717 788866 685837 789007
rect 685917 788946 686847 818654
rect 686927 818593 687067 818734
rect 686927 788866 687067 789007
rect 677707 788598 687067 788866
rect 687147 788678 687213 868982
rect 687273 867971 687869 956707
rect 687949 951934 688145 956787
rect 687929 951600 688165 951854
rect 687949 922600 688145 951600
rect 687929 922346 688165 922600
rect 687949 907934 688145 922266
rect 687929 907600 688165 907854
rect 687949 878400 688145 907600
rect 687929 878146 688165 878400
rect 687949 871032 688145 878066
rect 688225 871112 688821 959848
rect 688901 958262 717600 959928
rect 688881 877878 688947 958182
rect 689027 951934 717600 958262
rect 689027 951806 689167 951934
rect 689027 922600 689167 951600
rect 689027 922266 689167 922407
rect 689247 922346 690137 951854
rect 690217 951806 690337 951934
rect 690217 922600 690337 951600
rect 690217 922266 690337 922407
rect 690417 922346 691307 951854
rect 691387 951806 691527 951934
rect 691607 951600 696600 951854
rect 696680 951806 712677 951934
rect 712757 951600 717600 951854
rect 691387 922600 717600 951600
rect 691387 922266 691527 922407
rect 691607 922346 696600 922600
rect 696680 922266 712677 922407
rect 712757 922346 717600 922600
rect 689027 907934 717600 922266
rect 689027 907793 689167 907934
rect 689027 878400 689167 907600
rect 689027 878066 689167 878207
rect 689247 878146 690137 907854
rect 690217 907793 690337 907934
rect 690217 878400 690337 907600
rect 690217 878066 690337 878207
rect 690417 878146 691307 907854
rect 691387 907793 691527 907934
rect 691607 907600 696600 907854
rect 696680 907793 712677 907934
rect 712757 907600 717600 907854
rect 691387 878400 717600 907600
rect 691387 878066 691527 878207
rect 691607 878146 696600 878400
rect 696680 878066 712677 878207
rect 712757 878146 717600 878400
rect 689027 877798 717600 878066
rect 688901 871032 717600 877798
rect 687949 870728 717600 871032
rect 687949 867891 688145 870728
rect 687293 867587 688145 867891
rect 677707 779862 687193 788598
rect 677707 773534 687067 779862
rect 677707 773406 677927 773534
rect 677707 743866 677927 744007
rect 678007 743946 679097 773454
rect 679177 773406 679297 773534
rect 680387 773486 681477 773534
rect 679177 743866 679297 744007
rect 679377 743946 680307 773454
rect 680387 773406 680507 773486
rect 681357 773406 681477 773486
rect 680587 744007 681277 773406
rect 680387 743927 680507 744007
rect 681357 743927 681477 744007
rect 681557 743946 682487 773454
rect 682567 773406 682687 773534
rect 680387 743866 681477 743927
rect 682567 743866 682687 744007
rect 682767 743946 683697 773454
rect 683777 773406 683897 773534
rect 683777 743866 683897 744007
rect 683977 743946 684667 773454
rect 684747 773406 684867 773534
rect 684747 743866 684867 744007
rect 684947 743946 685637 773454
rect 685717 773406 685837 773534
rect 685717 743866 685837 744007
rect 685917 743946 686847 773454
rect 686927 773406 687067 773534
rect 686927 743866 687067 744007
rect 677707 743598 687067 743866
rect 687147 743678 687213 779782
rect 687273 778771 687869 867507
rect 687949 862734 688145 867587
rect 687929 862400 688165 862654
rect 687949 833400 688145 862400
rect 687929 833146 688165 833400
rect 687949 818734 688145 833066
rect 687929 818400 688165 818654
rect 687949 789200 688145 818400
rect 687929 788946 688165 789200
rect 687949 781832 688145 788866
rect 688225 781912 688821 870648
rect 688901 869062 717600 870728
rect 688881 788678 688947 868982
rect 689027 862734 717600 869062
rect 689027 862606 689167 862734
rect 689027 833400 689167 862400
rect 689027 833066 689167 833207
rect 689247 833146 690137 862654
rect 690217 862606 690337 862734
rect 690217 833400 690337 862400
rect 690217 833066 690337 833207
rect 690417 833146 691307 862654
rect 691387 862606 691527 862734
rect 691607 862400 696600 862654
rect 696680 862606 712677 862734
rect 712757 862400 717600 862654
rect 691387 833400 717600 862400
rect 691387 833066 691527 833207
rect 691607 833146 696600 833400
rect 696680 833066 712677 833207
rect 712757 833146 717600 833400
rect 689027 818734 717600 833066
rect 689027 818593 689167 818734
rect 689027 789200 689167 818400
rect 689027 788866 689167 789007
rect 689247 788946 690137 818654
rect 690217 818593 690337 818734
rect 690217 789200 690337 818400
rect 690217 788866 690337 789007
rect 690417 788946 691307 818654
rect 691387 818593 691527 818734
rect 691607 818400 696600 818654
rect 696680 818593 712677 818734
rect 712757 818400 717600 818654
rect 691387 789200 717600 818400
rect 691387 788866 691527 789007
rect 691607 788946 696600 789200
rect 696680 788866 712677 789007
rect 712757 788946 717600 789200
rect 689027 788598 717600 788866
rect 688901 781832 717600 788598
rect 687949 781528 717600 781832
rect 687949 778691 688145 781528
rect 687293 778387 688145 778691
rect 677707 734862 687193 743598
rect 677707 728534 687067 734862
rect 677707 728406 677927 728534
rect 677707 698866 677927 699007
rect 678007 698946 679097 728454
rect 679177 728406 679297 728534
rect 680387 728486 681477 728534
rect 679177 698866 679297 699007
rect 679377 698946 680307 728454
rect 680387 728406 680507 728486
rect 681357 728406 681477 728486
rect 680587 699007 681277 728406
rect 680387 698927 680507 699007
rect 681357 698927 681477 699007
rect 681557 698946 682487 728454
rect 682567 728406 682687 728534
rect 680387 698866 681477 698927
rect 682567 698866 682687 699007
rect 682767 698946 683697 728454
rect 683777 728406 683897 728534
rect 683777 698866 683897 699007
rect 683977 698946 684667 728454
rect 684747 728406 684867 728534
rect 684747 698866 684867 699007
rect 684947 698946 685637 728454
rect 685717 728406 685837 728534
rect 685717 698866 685837 699007
rect 685917 698946 686847 728454
rect 686927 728406 687067 728534
rect 686927 698866 687067 699007
rect 677707 698598 687067 698866
rect 687147 698678 687213 734782
rect 687273 733771 687869 778307
rect 687949 773534 688145 778387
rect 687929 773200 688165 773454
rect 687949 744200 688145 773200
rect 687929 743946 688165 744200
rect 687949 736832 688145 743866
rect 688225 736912 688821 781448
rect 688901 779862 717600 781528
rect 688881 743678 688947 779782
rect 689027 773534 717600 779862
rect 689027 773406 689167 773534
rect 689027 744200 689167 773200
rect 689027 743866 689167 744007
rect 689247 743946 690137 773454
rect 690217 773406 690337 773534
rect 690217 744200 690337 773200
rect 690217 743866 690337 744007
rect 690417 743946 691307 773454
rect 691387 773406 691527 773534
rect 691607 773200 696600 773454
rect 696680 773406 712677 773534
rect 712757 773200 717600 773454
rect 691387 744200 717600 773200
rect 691387 743866 691527 744007
rect 691607 743946 696600 744200
rect 696680 743866 712677 744007
rect 712757 743946 717600 744200
rect 689027 743598 717600 743866
rect 688901 736832 717600 743598
rect 687949 736528 717600 736832
rect 687949 733691 688145 736528
rect 687293 733387 688145 733691
rect 677707 689862 687193 698598
rect 677707 683534 687067 689862
rect 677707 683406 677927 683534
rect 677707 653666 677927 653807
rect 678007 653746 679097 683454
rect 679177 683406 679297 683534
rect 680387 683486 681477 683534
rect 679177 653666 679297 653807
rect 679377 653746 680307 683454
rect 680387 683406 680507 683486
rect 681357 683406 681477 683486
rect 680587 653807 681277 683406
rect 680387 653727 680507 653807
rect 681357 653727 681477 653807
rect 681557 653746 682487 683454
rect 682567 683406 682687 683534
rect 680387 653666 681477 653727
rect 682567 653666 682687 653807
rect 682767 653746 683697 683454
rect 683777 683406 683897 683534
rect 683777 653666 683897 653807
rect 683977 653746 684667 683454
rect 684747 683406 684867 683534
rect 684747 653666 684867 653807
rect 684947 653746 685637 683454
rect 685717 683406 685837 683534
rect 685717 653666 685837 653807
rect 685917 653746 686847 683454
rect 686927 683406 687067 683534
rect 686927 653666 687067 653807
rect 677707 653398 687067 653666
rect 687147 653478 687213 689782
rect 687273 688771 687869 733307
rect 687949 728534 688145 733387
rect 687929 728200 688165 728454
rect 687949 699200 688145 728200
rect 687929 698946 688165 699200
rect 687949 691832 688145 698866
rect 688225 691912 688821 736448
rect 688901 734862 717600 736528
rect 688881 698678 688947 734782
rect 689027 728534 717600 734862
rect 689027 728406 689167 728534
rect 689027 699200 689167 728200
rect 689027 698866 689167 699007
rect 689247 698946 690137 728454
rect 690217 728406 690337 728534
rect 690217 699200 690337 728200
rect 690217 698866 690337 699007
rect 690417 698946 691307 728454
rect 691387 728406 691527 728534
rect 691607 728200 696600 728454
rect 696680 728406 712677 728534
rect 712757 728200 717600 728454
rect 691387 699200 717600 728200
rect 691387 698866 691527 699007
rect 691607 698946 696600 699200
rect 696680 698866 712677 699007
rect 712757 698946 717600 699200
rect 689027 698598 717600 698866
rect 688901 691832 717600 698598
rect 687949 691528 717600 691832
rect 687949 688691 688145 691528
rect 687293 688387 688145 688691
rect 677707 644662 687193 653398
rect 677707 638334 687067 644662
rect 677707 638206 677927 638334
rect 677707 608666 677927 608807
rect 678007 608746 679097 638254
rect 679177 638206 679297 638334
rect 680387 638286 681477 638334
rect 679177 608666 679297 608807
rect 679377 608746 680307 638254
rect 680387 638206 680507 638286
rect 681357 638206 681477 638286
rect 680587 608807 681277 638206
rect 680387 608727 680507 608807
rect 681357 608727 681477 608807
rect 681557 608746 682487 638254
rect 682567 638206 682687 638334
rect 680387 608666 681477 608727
rect 682567 608666 682687 608807
rect 682767 608746 683697 638254
rect 683777 638206 683897 638334
rect 683777 608666 683897 608807
rect 683977 608746 684667 638254
rect 684747 638206 684867 638334
rect 684747 608666 684867 608807
rect 684947 608746 685637 638254
rect 685717 638206 685837 638334
rect 685717 608666 685837 608807
rect 685917 608746 686847 638254
rect 686927 638206 687067 638334
rect 686927 608666 687067 608807
rect 677707 608398 687067 608666
rect 687147 608478 687213 644582
rect 687273 643571 687869 688307
rect 687949 683534 688145 688387
rect 687929 683200 688165 683454
rect 687949 654000 688145 683200
rect 687929 653746 688165 654000
rect 687949 646632 688145 653666
rect 688225 646712 688821 691448
rect 688901 689862 717600 691528
rect 688881 653478 688947 689782
rect 689027 683534 717600 689862
rect 689027 683406 689167 683534
rect 689027 654000 689167 683200
rect 689027 653666 689167 653807
rect 689247 653746 690137 683454
rect 690217 683406 690337 683534
rect 690217 654000 690337 683200
rect 690217 653666 690337 653807
rect 690417 653746 691307 683454
rect 691387 683406 691527 683534
rect 691607 683200 696600 683454
rect 696680 683406 712677 683534
rect 712757 683200 717600 683454
rect 691387 654000 717600 683200
rect 691387 653666 691527 653807
rect 691607 653746 696600 654000
rect 696680 653666 712677 653807
rect 712757 653746 717600 654000
rect 689027 653398 717600 653666
rect 688901 646632 717600 653398
rect 687949 646328 717600 646632
rect 687949 643491 688145 646328
rect 687293 643187 688145 643491
rect 677707 599662 687193 608398
rect 677707 593334 687067 599662
rect 677707 593206 677927 593334
rect 677707 563466 677927 563607
rect 678007 563546 679097 593254
rect 679177 593206 679297 593334
rect 680387 593286 681477 593334
rect 679177 563466 679297 563607
rect 679377 563546 680307 593254
rect 680387 593206 680507 593286
rect 681357 593206 681477 593286
rect 680587 563607 681277 593206
rect 680387 563527 680507 563607
rect 681357 563527 681477 563607
rect 681557 563546 682487 593254
rect 682567 593206 682687 593334
rect 680387 563466 681477 563527
rect 682567 563466 682687 563607
rect 682767 563546 683697 593254
rect 683777 593206 683897 593334
rect 683777 563466 683897 563607
rect 683977 563546 684667 593254
rect 684747 593206 684867 593334
rect 684747 563466 684867 563607
rect 684947 563546 685637 593254
rect 685717 593206 685837 593334
rect 685717 563466 685837 563607
rect 685917 563546 686847 593254
rect 686927 593206 687067 593334
rect 686927 563466 687067 563607
rect 677707 563198 687067 563466
rect 687147 563278 687213 599582
rect 687273 598571 687869 643107
rect 687949 638334 688145 643187
rect 687929 638000 688165 638254
rect 687949 609000 688145 638000
rect 687929 608746 688165 609000
rect 687949 601632 688145 608666
rect 688225 601712 688821 646248
rect 688901 644662 717600 646328
rect 688881 608478 688947 644582
rect 689027 638334 717600 644662
rect 689027 638206 689167 638334
rect 689027 609000 689167 638000
rect 689027 608666 689167 608807
rect 689247 608746 690137 638254
rect 690217 638206 690337 638334
rect 690217 609000 690337 638000
rect 690217 608666 690337 608807
rect 690417 608746 691307 638254
rect 691387 638206 691527 638334
rect 691607 638000 696600 638254
rect 696680 638206 712677 638334
rect 712757 638000 717600 638254
rect 691387 609000 717600 638000
rect 691387 608666 691527 608807
rect 691607 608746 696600 609000
rect 696680 608666 712677 608807
rect 712757 608746 717600 609000
rect 689027 608398 717600 608666
rect 688901 601632 717600 608398
rect 687949 601328 717600 601632
rect 687949 598491 688145 601328
rect 687293 598187 688145 598491
rect 677707 554462 687193 563198
rect 677707 548134 687067 554462
rect 677707 548006 677927 548134
rect 678007 518546 679097 548054
rect 679177 548006 679297 548134
rect 680387 548086 681477 548134
rect 679177 518466 679297 518607
rect 679377 518546 680307 548054
rect 680387 548006 680507 548086
rect 681357 548006 681477 548086
rect 680587 518607 681277 548006
rect 680387 518527 680507 518607
rect 681357 518527 681477 518607
rect 681557 518546 682487 548054
rect 682567 548006 682687 548134
rect 680387 518466 681477 518527
rect 682567 518466 682687 518607
rect 682767 518546 683697 548054
rect 683777 548006 683897 548134
rect 683777 518466 683897 518607
rect 683977 518546 684667 548054
rect 684747 548006 684867 548134
rect 684747 518466 684867 518607
rect 684947 518546 685637 548054
rect 685717 548006 685837 548134
rect 685717 518466 685837 518607
rect 685917 518546 686847 548054
rect 686927 548006 687067 548134
rect 686927 518466 687067 518607
rect 678007 504134 687067 518466
rect 677547 477596 677613 477597
rect 677547 477532 677548 477596
rect 677612 477532 677613 477596
rect 677547 477531 677613 477532
rect 678007 474546 679097 504054
rect 679177 503993 679297 504134
rect 680387 504073 681477 504134
rect 679177 474466 679297 474607
rect 679377 474546 680307 504054
rect 680387 503993 680507 504073
rect 681357 503993 681477 504073
rect 680587 474607 681277 503993
rect 680387 474527 680507 474607
rect 681357 474527 681477 474607
rect 681557 474546 682487 504054
rect 682567 503993 682687 504134
rect 680387 474466 681477 474527
rect 682567 474466 682687 474607
rect 682767 474546 683697 504054
rect 683777 503993 683897 504134
rect 683777 474466 683897 474607
rect 683977 474546 684667 504054
rect 684747 503993 684867 504134
rect 684747 474466 684867 474607
rect 684947 474546 685637 504054
rect 685717 503993 685837 504134
rect 685717 474466 685837 474607
rect 685917 474546 686847 504054
rect 686927 503993 687067 504134
rect 686927 474466 687067 474607
rect 678007 460134 687067 474466
rect 40171 455428 40237 455429
rect 40171 455364 40172 455428
rect 40236 455364 40237 455428
rect 40171 455363 40237 455364
rect 40171 451892 40237 451893
rect 40171 451828 40172 451892
rect 40236 451828 40237 451892
rect 40171 451827 40237 451828
rect 30533 440993 30673 441134
rect 30533 413266 30673 413394
rect 30753 413346 31683 441054
rect 31763 440993 31883 441134
rect 31763 413266 31883 413394
rect 31963 413346 32653 441054
rect 32733 440993 32853 441134
rect 32733 413266 32853 413394
rect 32933 413346 33623 441054
rect 33703 440993 33823 441134
rect 33703 413266 33823 413394
rect 33903 413346 34833 441054
rect 34913 440993 35033 441134
rect 36123 441073 37213 441134
rect 34913 413266 35033 413394
rect 35113 413346 36043 441054
rect 36123 440993 36243 441073
rect 37093 440993 37213 441073
rect 36323 413394 37013 440993
rect 36123 413314 36243 413394
rect 37093 413314 37213 413394
rect 37293 413346 38223 441054
rect 38303 440993 38423 441134
rect 36123 413266 37213 413314
rect 38303 413266 38423 413394
rect 38503 413346 39593 441054
rect 39673 413266 39893 413394
rect 30533 406938 39893 413266
rect 30407 398202 39893 406938
rect 29455 364909 30307 365213
rect 29455 362072 29651 364909
rect 0 361768 29651 362072
rect 0 355002 28699 361768
rect 0 354734 28573 355002
rect 0 354400 4843 354654
rect 4923 354593 20920 354734
rect 21000 354400 25993 354654
rect 26073 354593 26213 354734
rect 0 327200 26213 354400
rect 0 326946 4843 327200
rect 4923 326866 20920 326994
rect 21000 326946 25993 327200
rect 26073 326866 26213 326994
rect 26293 326946 27183 354654
rect 27263 354593 27383 354734
rect 27263 327200 27383 354400
rect 27263 326866 27383 326994
rect 27463 326946 28353 354654
rect 28433 354593 28573 354734
rect 28433 327200 28573 354400
rect 28433 326866 28573 326994
rect 0 320538 28573 326866
rect 28653 320618 28719 354922
rect 0 318872 28699 320538
rect 28779 318952 29375 361688
rect 29455 354734 29651 361768
rect 29435 354400 29671 354654
rect 29455 327200 29651 354400
rect 29435 326946 29671 327200
rect 29455 322013 29651 326866
rect 29731 322093 30327 364829
rect 30387 363818 30453 398122
rect 30533 397934 39893 398202
rect 30533 397793 30673 397934
rect 30533 370066 30673 370194
rect 30753 370146 31683 397854
rect 31763 397793 31883 397934
rect 31763 370066 31883 370194
rect 31963 370146 32653 397854
rect 32733 397793 32853 397934
rect 32733 370066 32853 370194
rect 32933 370146 33623 397854
rect 33703 397793 33823 397934
rect 33703 370066 33823 370194
rect 33903 370146 34833 397854
rect 34913 397793 35033 397934
rect 36123 397873 37213 397934
rect 34913 370066 35033 370194
rect 35113 370146 36043 397854
rect 36123 397793 36243 397873
rect 37093 397793 37213 397873
rect 36323 370194 37013 397793
rect 36123 370114 36243 370194
rect 37093 370114 37213 370194
rect 37293 370146 38223 397854
rect 38303 397793 38423 397934
rect 36123 370066 37213 370114
rect 38303 370066 38423 370194
rect 38503 370146 39593 397854
rect 39673 397793 39893 397934
rect 39673 370066 39893 370194
rect 30533 363738 39893 370066
rect 30407 355002 39893 363738
rect 29455 321709 30307 322013
rect 29455 318872 29651 321709
rect 0 318568 29651 318872
rect 0 311802 28699 318568
rect 0 311534 28573 311802
rect 0 311200 4843 311454
rect 4923 311393 20920 311534
rect 21000 311200 25993 311454
rect 26073 311393 26213 311534
rect 0 284000 26213 311200
rect 0 283746 4843 284000
rect 4923 283666 20920 283794
rect 21000 283746 25993 284000
rect 26073 283666 26213 283794
rect 26293 283746 27183 311454
rect 27263 311393 27383 311534
rect 27263 284000 27383 311200
rect 27263 283666 27383 283794
rect 27463 283746 28353 311454
rect 28433 311393 28573 311534
rect 28433 284000 28573 311200
rect 28433 283666 28573 283794
rect 0 277338 28573 283666
rect 28653 277418 28719 311722
rect 0 275672 28699 277338
rect 28779 275752 29375 318488
rect 29455 311534 29651 318568
rect 29435 311200 29671 311454
rect 29455 284000 29651 311200
rect 29435 283746 29671 284000
rect 29455 278813 29651 283666
rect 29731 278893 30327 321629
rect 30387 320618 30453 354922
rect 30533 354734 39893 355002
rect 30533 354593 30673 354734
rect 30533 326866 30673 326994
rect 30753 326946 31683 354654
rect 31763 354593 31883 354734
rect 31763 326866 31883 326994
rect 31963 326946 32653 354654
rect 32733 354593 32853 354734
rect 32733 326866 32853 326994
rect 32933 326946 33623 354654
rect 33703 354593 33823 354734
rect 33703 326866 33823 326994
rect 33903 326946 34833 354654
rect 34913 354593 35033 354734
rect 36123 354673 37213 354734
rect 34913 326866 35033 326994
rect 35113 326946 36043 354654
rect 36123 354593 36243 354673
rect 37093 354593 37213 354673
rect 36323 326994 37013 354593
rect 36123 326914 36243 326994
rect 37093 326914 37213 326994
rect 37293 326946 38223 354654
rect 38303 354593 38423 354734
rect 36123 326866 37213 326914
rect 38303 326866 38423 326994
rect 38503 326946 39593 354654
rect 39673 354593 39893 354734
rect 39673 326866 39893 326994
rect 30533 320538 39893 326866
rect 30407 311802 39893 320538
rect 29455 278509 30307 278813
rect 29455 275672 29651 278509
rect 0 275368 29651 275672
rect 0 268602 28699 275368
rect 0 268334 28573 268602
rect 0 268000 4843 268254
rect 4923 268193 20920 268334
rect 21000 268000 25993 268254
rect 26073 268193 26213 268334
rect 0 240800 26213 268000
rect 0 240546 4843 240800
rect 4923 240466 20920 240594
rect 21000 240546 25993 240800
rect 26073 240466 26213 240594
rect 26293 240546 27183 268254
rect 27263 268193 27383 268334
rect 27263 240800 27383 268000
rect 27263 240466 27383 240594
rect 27463 240546 28353 268254
rect 28433 268193 28573 268334
rect 28433 240800 28573 268000
rect 28433 240466 28573 240594
rect 0 234138 28573 240466
rect 28653 234218 28719 268522
rect 0 232472 28699 234138
rect 28779 232552 29375 275288
rect 29455 268334 29651 275368
rect 29435 268000 29671 268254
rect 29455 240800 29651 268000
rect 29435 240546 29671 240800
rect 29455 235613 29651 240466
rect 29731 235693 30327 278429
rect 30387 277418 30453 311722
rect 30533 311534 39893 311802
rect 30533 311393 30673 311534
rect 30533 283666 30673 283794
rect 30753 283746 31683 311454
rect 31763 311393 31883 311534
rect 31763 283666 31883 283794
rect 31963 283746 32653 311454
rect 32733 311393 32853 311534
rect 32733 283666 32853 283794
rect 32933 283746 33623 311454
rect 33703 311393 33823 311534
rect 33703 283666 33823 283794
rect 33903 283746 34833 311454
rect 34913 311393 35033 311534
rect 36123 311473 37213 311534
rect 34913 283666 35033 283794
rect 35113 283746 36043 311454
rect 36123 311393 36243 311473
rect 37093 311393 37213 311473
rect 36323 283794 37013 311393
rect 36123 283714 36243 283794
rect 37093 283714 37213 283794
rect 37293 283746 38223 311454
rect 38303 311393 38423 311534
rect 36123 283666 37213 283714
rect 38303 283666 38423 283794
rect 38503 283746 39593 311454
rect 39673 311393 39893 311534
rect 39673 283666 39893 283794
rect 30533 277338 39893 283666
rect 30407 268602 39893 277338
rect 29455 235309 30307 235613
rect 29455 232472 29651 235309
rect 0 232168 29651 232472
rect 0 225402 28699 232168
rect 0 225134 28573 225402
rect 0 224800 4843 225054
rect 4923 224993 20920 225134
rect 21000 224800 25993 225054
rect 26073 224993 26213 225134
rect 0 197600 26213 224800
rect 0 197346 4843 197600
rect 4923 197266 20920 197394
rect 21000 197346 25993 197600
rect 26073 197266 26213 197394
rect 26293 197346 27183 225054
rect 27263 224993 27383 225134
rect 27263 197600 27383 224800
rect 27263 197266 27383 197394
rect 27463 197346 28353 225054
rect 28433 224993 28573 225134
rect 28433 197600 28573 224800
rect 28433 197266 28573 197394
rect 0 190938 28573 197266
rect 28653 191018 28719 225322
rect 0 189272 28699 190938
rect 28779 189352 29375 232088
rect 29455 225134 29651 232168
rect 29435 224800 29671 225054
rect 29455 197600 29651 224800
rect 29435 197346 29671 197600
rect 29455 192413 29651 197266
rect 29731 192493 30327 235229
rect 30387 234218 30453 268522
rect 30533 268334 39893 268602
rect 30533 268193 30673 268334
rect 30533 240466 30673 240594
rect 30753 240546 31683 268254
rect 31763 268193 31883 268334
rect 31763 240466 31883 240594
rect 31963 240546 32653 268254
rect 32733 268193 32853 268334
rect 32733 240466 32853 240594
rect 32933 240546 33623 268254
rect 33703 268193 33823 268334
rect 33703 240466 33823 240594
rect 33903 240546 34833 268254
rect 34913 268193 35033 268334
rect 36123 268273 37213 268334
rect 34913 240466 35033 240594
rect 35113 240546 36043 268254
rect 36123 268193 36243 268273
rect 37093 268193 37213 268273
rect 36323 240594 37013 268193
rect 36123 240514 36243 240594
rect 37093 240514 37213 240594
rect 37293 240546 38223 268254
rect 38303 268193 38423 268334
rect 36123 240466 37213 240514
rect 38303 240466 38423 240594
rect 38503 240546 39593 268254
rect 39673 268193 39893 268334
rect 39673 240466 39893 240594
rect 30533 234138 39893 240466
rect 30407 225402 39893 234138
rect 29455 192109 30307 192413
rect 29455 189272 29651 192109
rect 0 188968 29651 189272
rect 0 182202 28699 188968
rect 0 181934 28573 182202
rect 0 181600 4843 181854
rect 4923 181793 20920 181934
rect 21000 181600 25993 181854
rect 26073 181793 26213 181934
rect 0 153400 26213 181600
rect 0 152400 25993 153400
rect 0 125200 26213 152400
rect 0 124946 4843 125200
rect 4923 124866 20920 125007
rect 21000 124946 25993 125200
rect 26073 124866 26213 125007
rect 26293 124946 27183 181854
rect 27263 181793 27383 181934
rect 27263 153400 27383 181600
rect 27263 125200 27383 152400
rect 27263 124866 27383 125007
rect 27463 124946 28353 181854
rect 28433 181793 28573 181934
rect 28433 153400 28573 181600
rect 28653 153400 28719 182122
rect 28433 125200 28573 152400
rect 28433 124866 28573 125007
rect 0 110534 28573 124866
rect 0 110200 4843 110454
rect 4923 110393 20920 110534
rect 21000 110200 25993 110454
rect 26073 110393 26213 110534
rect 0 83000 26213 110200
rect 0 82746 4843 83000
rect 4923 82666 20920 82807
rect 21000 82746 25993 83000
rect 26073 82666 26213 82807
rect 26293 82746 27183 110454
rect 27263 110393 27383 110534
rect 27263 83000 27383 110200
rect 27263 82666 27383 82807
rect 27463 82746 28353 110454
rect 28433 110393 28573 110534
rect 28433 83000 28573 110200
rect 28433 82666 28573 82807
rect 0 68334 28573 82666
rect 0 68000 4843 68254
rect 4923 68193 20920 68334
rect 21000 68000 25993 68254
rect 26073 68193 26213 68334
rect 0 40800 26213 68000
rect 0 40546 4843 40800
rect 4923 40466 20920 40549
rect 0 40349 20920 40466
rect 21000 40429 25993 40800
rect 26073 40466 26213 40549
rect 26293 40546 27183 68254
rect 27263 68193 27383 68334
rect 27263 40800 27383 68000
rect 27263 40466 27383 40549
rect 27463 40546 28353 68254
rect 28433 68193 28573 68334
rect 28433 40800 28573 68000
rect 28433 40466 28573 40549
rect 26073 40349 28573 40466
rect 0 35285 28573 40349
rect 28653 35365 28719 152400
rect 28779 35418 29375 188888
rect 29455 181934 29651 188968
rect 29435 181600 29671 181854
rect 29455 153400 29651 181600
rect 29455 125200 29651 152400
rect 29435 124946 29671 125200
rect 29455 110534 29651 124866
rect 29435 110200 29671 110454
rect 29455 83000 29651 110200
rect 29435 82746 29671 83000
rect 29455 68334 29651 82666
rect 29435 68000 29671 68254
rect 29455 40800 29651 68000
rect 29435 36489 29671 40800
rect 29731 36625 30327 192029
rect 30387 191018 30453 225322
rect 30533 225134 39893 225402
rect 30533 224993 30673 225134
rect 30533 197266 30673 197394
rect 30753 197346 31683 225054
rect 31763 224993 31883 225134
rect 31763 197266 31883 197394
rect 31963 197346 32653 225054
rect 32733 224993 32853 225134
rect 32733 197266 32853 197394
rect 32933 197346 33623 225054
rect 33703 224993 33823 225134
rect 33703 197266 33823 197394
rect 33903 197346 34833 225054
rect 34913 224993 35033 225134
rect 36123 225073 37213 225134
rect 34913 197266 35033 197394
rect 35113 197346 36043 225054
rect 36123 224993 36243 225073
rect 37093 224993 37213 225073
rect 36323 197394 37013 224993
rect 36123 197314 36243 197394
rect 37093 197314 37213 197394
rect 37293 197346 38223 225054
rect 38303 224993 38423 225134
rect 36123 197266 37213 197314
rect 38303 197266 38423 197394
rect 38503 197346 39593 225054
rect 39673 224993 39893 225134
rect 39673 197266 39893 197394
rect 30533 190938 39893 197266
rect 30407 182202 39893 190938
rect 30387 153400 30453 182122
rect 30533 181934 39893 182202
rect 30533 181793 30673 181934
rect 30753 154400 31683 181854
rect 31763 181793 31883 181934
rect 31963 153400 32653 181854
rect 32733 181793 32853 181934
rect 29751 36409 30307 36545
rect 29455 36005 30307 36409
rect 30387 36085 30453 152400
rect 30533 124866 30673 125007
rect 30753 124946 31683 153400
rect 31763 124866 31883 125007
rect 31963 124946 32653 152400
rect 32733 124866 32853 125007
rect 32933 124946 33623 181854
rect 33703 181793 33823 181934
rect 33703 124866 33823 125007
rect 33903 124946 34833 181854
rect 34913 181793 35033 181934
rect 36123 181873 37213 181934
rect 34913 124866 35033 125007
rect 35113 124946 36043 181854
rect 36123 181793 36243 181873
rect 37093 181793 37213 181873
rect 36323 153400 37013 181793
rect 37293 154400 38223 181854
rect 38303 181793 38423 181934
rect 36323 125007 37013 152400
rect 36123 124927 36243 125007
rect 37093 124927 37213 125007
rect 37293 124946 38223 153400
rect 36123 124866 37213 124927
rect 38303 124866 38423 125007
rect 38503 124946 39593 181854
rect 39673 181793 39893 181934
rect 30533 110534 39593 124866
rect 30533 110393 30673 110534
rect 30533 82666 30673 82807
rect 30753 82746 31683 110454
rect 31763 110393 31883 110534
rect 31763 82666 31883 82807
rect 31963 82746 32653 110454
rect 32733 110393 32853 110534
rect 32733 82666 32853 82807
rect 32933 82746 33623 110454
rect 33703 110393 33823 110534
rect 33703 82666 33823 82807
rect 33903 82746 34833 110454
rect 34913 110393 35033 110534
rect 36123 110473 37213 110534
rect 34913 82666 35033 82807
rect 35113 82746 36043 110454
rect 36123 110393 36243 110473
rect 37093 110393 37213 110473
rect 36323 82807 37013 110393
rect 36123 82727 36243 82807
rect 37093 82727 37213 82807
rect 37293 82746 38223 110454
rect 38303 110393 38423 110534
rect 36123 82666 37213 82727
rect 38303 82666 38423 82807
rect 38503 82746 39593 110454
rect 40174 84285 40234 451827
rect 678007 430346 679097 460054
rect 679177 459993 679297 460134
rect 680387 460073 681477 460134
rect 679177 430266 679297 430407
rect 679377 430346 680307 460054
rect 680387 459993 680507 460073
rect 681357 459993 681477 460073
rect 680587 430407 681277 459993
rect 680387 430327 680507 430407
rect 681357 430327 681477 430407
rect 681557 430346 682487 460054
rect 682567 459993 682687 460134
rect 680387 430266 681477 430327
rect 682567 430266 682687 430407
rect 682767 430346 683697 460054
rect 683777 459993 683897 460134
rect 683777 430266 683897 430407
rect 683977 430346 684667 460054
rect 684747 459993 684867 460134
rect 684747 430266 684867 430407
rect 684947 430346 685637 460054
rect 685717 459993 685837 460134
rect 685717 430266 685837 430407
rect 685917 430346 686847 460054
rect 686927 459993 687067 460134
rect 686927 430266 687067 430407
rect 687147 430346 687213 554382
rect 687273 553371 687869 598107
rect 687949 593334 688145 598187
rect 687929 593000 688165 593254
rect 687949 563800 688145 593000
rect 687929 563546 688165 563800
rect 687949 556432 688145 563466
rect 688225 556512 688821 601248
rect 688901 599662 717600 601328
rect 688881 563278 688947 599582
rect 689027 593334 717600 599662
rect 689027 593206 689167 593334
rect 689027 563800 689167 593000
rect 689027 563466 689167 563607
rect 689247 563546 690137 593254
rect 690217 593206 690337 593334
rect 690217 563800 690337 593000
rect 690217 563466 690337 563607
rect 690417 563546 691307 593254
rect 691387 593206 691527 593334
rect 691607 593000 696600 593254
rect 696680 593206 712677 593334
rect 712757 593000 717600 593254
rect 691387 563800 717600 593000
rect 691387 563466 691527 563607
rect 691607 563546 696600 563800
rect 696680 563466 712677 563607
rect 712757 563546 717600 563800
rect 689027 563198 717600 563466
rect 688901 556432 717600 563198
rect 687949 556128 717600 556432
rect 687949 553291 688145 556128
rect 687293 552987 688145 553291
rect 678007 415934 687193 430266
rect 677707 386266 677927 386407
rect 678007 386346 679097 415854
rect 679177 415793 679297 415934
rect 680387 415873 681477 415934
rect 679177 386266 679297 386407
rect 679377 386346 680307 415854
rect 680387 415793 680507 415873
rect 681357 415793 681477 415873
rect 680587 386407 681277 415793
rect 680387 386327 680507 386407
rect 681357 386327 681477 386407
rect 681557 386346 682487 415854
rect 682567 415793 682687 415934
rect 680387 386266 681477 386327
rect 682567 386266 682687 386407
rect 682767 386346 683697 415854
rect 683777 415793 683897 415934
rect 683777 386266 683897 386407
rect 683977 386346 684667 415854
rect 684747 415793 684867 415934
rect 684747 386266 684867 386407
rect 684947 386346 685637 415854
rect 685717 415793 685837 415934
rect 685717 386266 685837 386407
rect 685917 386346 686847 415854
rect 686927 415793 687067 415934
rect 686927 386266 687067 386407
rect 677707 385998 687067 386266
rect 687147 386078 687213 415854
rect 677707 377262 687193 385998
rect 677707 370934 687067 377262
rect 677707 370806 677927 370934
rect 677707 341066 677927 341207
rect 678007 341146 679097 370854
rect 679177 370806 679297 370934
rect 680387 370886 681477 370934
rect 679177 341066 679297 341207
rect 679377 341146 680307 370854
rect 680387 370806 680507 370886
rect 681357 370806 681477 370886
rect 680587 341207 681277 370806
rect 680387 341127 680507 341207
rect 681357 341127 681477 341207
rect 681557 341146 682487 370854
rect 682567 370806 682687 370934
rect 680387 341066 681477 341127
rect 682567 341066 682687 341207
rect 682767 341146 683697 370854
rect 683777 370806 683897 370934
rect 683777 341066 683897 341207
rect 683977 341146 684667 370854
rect 684747 370806 684867 370934
rect 684747 341066 684867 341207
rect 684947 341146 685637 370854
rect 685717 370806 685837 370934
rect 685717 341066 685837 341207
rect 685917 341146 686847 370854
rect 686927 370806 687067 370934
rect 686927 341066 687067 341207
rect 677707 340798 687067 341066
rect 687147 340878 687213 377182
rect 687273 376171 687869 552907
rect 687949 548134 688145 552987
rect 687929 547800 688165 548054
rect 687949 518800 688145 547800
rect 687929 518546 688165 518800
rect 687949 504134 688145 518466
rect 687929 503800 688165 504054
rect 687949 474800 688145 503800
rect 687929 474546 688165 474800
rect 687949 460134 688145 474466
rect 687929 459800 688165 460054
rect 687949 430600 688145 459800
rect 687929 430346 688165 430600
rect 687949 415934 688145 430266
rect 687929 415600 688165 415854
rect 687949 386600 688145 415600
rect 687929 386346 688165 386600
rect 687949 379232 688145 386266
rect 688225 379312 688821 556048
rect 688901 554462 717600 556128
rect 688881 430346 688947 554382
rect 689027 548134 717600 554462
rect 689027 548006 689167 548134
rect 689027 518800 689167 547800
rect 689027 518466 689167 518607
rect 689247 518546 690137 548054
rect 690217 548006 690337 548134
rect 690217 518800 690337 547800
rect 690217 518466 690337 518607
rect 690417 518546 691307 548054
rect 691387 548006 691527 548134
rect 691607 547800 696600 548054
rect 696680 548006 712677 548134
rect 712757 547800 717600 548054
rect 691387 518800 717600 547800
rect 691387 518466 691527 518607
rect 691607 518546 696600 518800
rect 696680 518466 712677 518607
rect 712757 518546 717600 518800
rect 689027 504134 717600 518466
rect 689027 503993 689167 504134
rect 689027 474800 689167 503800
rect 689027 474466 689167 474607
rect 689247 474546 690137 504054
rect 690217 503993 690337 504134
rect 690217 474800 690337 503800
rect 690217 474466 690337 474607
rect 690417 474546 691307 504054
rect 691387 503993 691527 504134
rect 691607 503800 696600 504054
rect 696680 503993 712677 504134
rect 712757 503800 717600 504054
rect 691387 474800 717600 503800
rect 691387 474466 691527 474607
rect 691607 474546 696600 474800
rect 696680 474466 712677 474607
rect 712757 474546 717600 474800
rect 689027 460134 717600 474466
rect 689027 459993 689167 460134
rect 689027 430600 689167 459800
rect 689027 430266 689167 430407
rect 689247 430346 690137 460054
rect 690217 459993 690337 460134
rect 690217 430600 690337 459800
rect 690217 430266 690337 430407
rect 690417 430346 691307 460054
rect 691387 459993 691527 460134
rect 691607 459800 696600 460054
rect 696680 459993 712677 460134
rect 712757 459800 717600 460054
rect 691387 430600 717600 459800
rect 691387 430266 691527 430407
rect 691607 430346 696600 430600
rect 696680 430266 712677 430407
rect 712757 430346 717600 430600
rect 688901 415934 717600 430266
rect 688881 386078 688947 415854
rect 689027 415793 689167 415934
rect 689027 386600 689167 415600
rect 689027 386266 689167 386407
rect 689247 386346 690137 415854
rect 690217 415793 690337 415934
rect 690217 386600 690337 415600
rect 690217 386266 690337 386407
rect 690417 386346 691307 415854
rect 691387 415793 691527 415934
rect 691607 415600 696600 415854
rect 696680 415793 712677 415934
rect 712757 415600 717600 415854
rect 691387 386600 717600 415600
rect 691387 386266 691527 386407
rect 691607 386346 696600 386600
rect 696680 386266 712677 386407
rect 712757 386346 717600 386600
rect 689027 385998 717600 386266
rect 688901 379232 717600 385998
rect 687949 378928 717600 379232
rect 687949 376091 688145 378928
rect 687293 375787 688145 376091
rect 677707 332062 687193 340798
rect 677707 325734 687067 332062
rect 677707 325606 677927 325734
rect 677707 296066 677927 296207
rect 678007 296146 679097 325654
rect 679177 325606 679297 325734
rect 680387 325686 681477 325734
rect 679177 296066 679297 296207
rect 679377 296146 680307 325654
rect 680387 325606 680507 325686
rect 681357 325606 681477 325686
rect 680587 296207 681277 325606
rect 680387 296127 680507 296207
rect 681357 296127 681477 296207
rect 681557 296146 682487 325654
rect 682567 325606 682687 325734
rect 680387 296066 681477 296127
rect 682567 296066 682687 296207
rect 682767 296146 683697 325654
rect 683777 325606 683897 325734
rect 683777 296066 683897 296207
rect 683977 296146 684667 325654
rect 684747 325606 684867 325734
rect 684747 296066 684867 296207
rect 684947 296146 685637 325654
rect 685717 325606 685837 325734
rect 685717 296066 685837 296207
rect 685917 296146 686847 325654
rect 686927 325606 687067 325734
rect 686927 296066 687067 296207
rect 677707 295798 687067 296066
rect 687147 295878 687213 331982
rect 687273 330971 687869 375707
rect 687949 370934 688145 375787
rect 687929 370600 688165 370854
rect 687949 341400 688145 370600
rect 687929 341146 688165 341400
rect 687949 334032 688145 341066
rect 688225 334112 688821 378848
rect 688901 377262 717600 378928
rect 688881 340878 688947 377182
rect 689027 370934 717600 377262
rect 689027 370806 689167 370934
rect 689027 341400 689167 370600
rect 689027 341066 689167 341207
rect 689247 341146 690137 370854
rect 690217 370806 690337 370934
rect 690217 341400 690337 370600
rect 690217 341066 690337 341207
rect 690417 341146 691307 370854
rect 691387 370806 691527 370934
rect 691607 370600 696600 370854
rect 696680 370806 712677 370934
rect 712757 370600 717600 370854
rect 691387 341400 717600 370600
rect 691387 341066 691527 341207
rect 691607 341146 696600 341400
rect 696680 341066 712677 341207
rect 712757 341146 717600 341400
rect 689027 340798 717600 341066
rect 688901 334032 717600 340798
rect 687949 333728 717600 334032
rect 687949 330891 688145 333728
rect 687293 330587 688145 330891
rect 677707 287062 687193 295798
rect 677707 280734 687067 287062
rect 677707 280606 677927 280734
rect 677707 251066 677927 251207
rect 678007 251146 679097 280654
rect 679177 280606 679297 280734
rect 680387 280686 681477 280734
rect 679177 251066 679297 251207
rect 679377 251146 680307 280654
rect 680387 280606 680507 280686
rect 681357 280606 681477 280686
rect 680587 251207 681277 280606
rect 680387 251127 680507 251207
rect 681357 251127 681477 251207
rect 681557 251146 682487 280654
rect 682567 280606 682687 280734
rect 680387 251066 681477 251127
rect 682567 251066 682687 251207
rect 682767 251146 683697 280654
rect 683777 280606 683897 280734
rect 683777 251066 683897 251207
rect 683977 251146 684667 280654
rect 684747 280606 684867 280734
rect 684747 251066 684867 251207
rect 684947 251146 685637 280654
rect 685717 280606 685837 280734
rect 685717 251066 685837 251207
rect 685917 251146 686847 280654
rect 686927 280606 687067 280734
rect 686927 251066 687067 251207
rect 677707 250798 687067 251066
rect 687147 250878 687213 286982
rect 687273 285971 687869 330507
rect 687949 325734 688145 330587
rect 687929 325400 688165 325654
rect 687949 296400 688145 325400
rect 687929 296146 688165 296400
rect 687949 289032 688145 296066
rect 688225 289112 688821 333648
rect 688901 332062 717600 333728
rect 688881 295878 688947 331982
rect 689027 325734 717600 332062
rect 689027 325606 689167 325734
rect 689027 296400 689167 325400
rect 689027 296066 689167 296207
rect 689247 296146 690137 325654
rect 690217 325606 690337 325734
rect 690217 296400 690337 325400
rect 690217 296066 690337 296207
rect 690417 296146 691307 325654
rect 691387 325606 691527 325734
rect 691607 325400 696600 325654
rect 696680 325606 712677 325734
rect 712757 325400 717600 325654
rect 691387 296400 717600 325400
rect 691387 296066 691527 296207
rect 691607 296146 696600 296400
rect 696680 296066 712677 296207
rect 712757 296146 717600 296400
rect 689027 295798 717600 296066
rect 688901 289032 717600 295798
rect 687949 288728 717600 289032
rect 687949 285891 688145 288728
rect 687293 285587 688145 285891
rect 677707 242062 687193 250798
rect 677707 235734 687067 242062
rect 677707 235606 677927 235734
rect 677707 205866 677927 206007
rect 678007 205946 679097 235654
rect 679177 235606 679297 235734
rect 680387 235686 681477 235734
rect 679177 205866 679297 206007
rect 679377 205946 680307 235654
rect 680387 235606 680507 235686
rect 681357 235606 681477 235686
rect 680587 206007 681277 235606
rect 680387 205927 680507 206007
rect 681357 205927 681477 206007
rect 681557 205946 682487 235654
rect 682567 235606 682687 235734
rect 680387 205866 681477 205927
rect 682567 205866 682687 206007
rect 682767 205946 683697 235654
rect 683777 235606 683897 235734
rect 683777 205866 683897 206007
rect 683977 205946 684667 235654
rect 684747 235606 684867 235734
rect 684747 205866 684867 206007
rect 684947 205946 685637 235654
rect 685717 235606 685837 235734
rect 685717 205866 685837 206007
rect 685917 205946 686847 235654
rect 686927 235606 687067 235734
rect 686927 205866 687067 206007
rect 677707 205598 687067 205866
rect 687147 205678 687213 241982
rect 687273 240971 687869 285507
rect 687949 280734 688145 285587
rect 687929 280400 688165 280654
rect 687949 251400 688145 280400
rect 687929 251146 688165 251400
rect 687949 244032 688145 251066
rect 688225 244112 688821 288648
rect 688901 287062 717600 288728
rect 688881 250878 688947 286982
rect 689027 280734 717600 287062
rect 689027 280606 689167 280734
rect 689027 251400 689167 280400
rect 689027 251066 689167 251207
rect 689247 251146 690137 280654
rect 690217 280606 690337 280734
rect 690217 251400 690337 280400
rect 690217 251066 690337 251207
rect 690417 251146 691307 280654
rect 691387 280606 691527 280734
rect 691607 280400 696600 280654
rect 696680 280606 712677 280734
rect 712757 280400 717600 280654
rect 691387 251400 717600 280400
rect 691387 251066 691527 251207
rect 691607 251146 696600 251400
rect 696680 251066 712677 251207
rect 712757 251146 717600 251400
rect 689027 250798 717600 251066
rect 688901 244032 717600 250798
rect 687949 243728 717600 244032
rect 687949 240891 688145 243728
rect 687293 240587 688145 240891
rect 677707 196862 687193 205598
rect 677707 190534 687067 196862
rect 677707 190406 677927 190534
rect 677707 160866 677927 161007
rect 678007 160946 679097 190454
rect 679177 190406 679297 190534
rect 680387 190486 681477 190534
rect 679177 160866 679297 161007
rect 679377 160946 680307 190454
rect 680387 190406 680507 190486
rect 681357 190406 681477 190486
rect 680587 161007 681277 190406
rect 680387 160927 680507 161007
rect 681357 160927 681477 161007
rect 681557 160946 682487 190454
rect 682567 190406 682687 190534
rect 680387 160866 681477 160927
rect 682567 160866 682687 161007
rect 682767 160946 683697 190454
rect 683777 190406 683897 190534
rect 683777 160866 683897 161007
rect 683977 160946 684667 190454
rect 684747 190406 684867 190534
rect 684747 160866 684867 161007
rect 684947 160946 685637 190454
rect 685717 190406 685837 190534
rect 685717 160866 685837 161007
rect 685917 160946 686847 190454
rect 686927 190406 687067 190534
rect 686927 160866 687067 161007
rect 677707 160598 687067 160866
rect 687147 160678 687213 196782
rect 687273 195771 687869 240507
rect 687949 235734 688145 240587
rect 687929 235400 688165 235654
rect 687949 206200 688145 235400
rect 687929 205946 688165 206200
rect 687949 198832 688145 205866
rect 688225 198912 688821 243648
rect 688901 242062 717600 243728
rect 688881 205678 688947 241982
rect 689027 235734 717600 242062
rect 689027 235606 689167 235734
rect 689027 206200 689167 235400
rect 689027 205866 689167 206007
rect 689247 205946 690137 235654
rect 690217 235606 690337 235734
rect 690217 206200 690337 235400
rect 690217 205866 690337 206007
rect 690417 205946 691307 235654
rect 691387 235606 691527 235734
rect 691607 235400 696600 235654
rect 696680 235606 712677 235734
rect 712757 235400 717600 235654
rect 691387 206200 717600 235400
rect 691387 205866 691527 206007
rect 691607 205946 696600 206200
rect 696680 205866 712677 206007
rect 712757 205946 717600 206200
rect 689027 205598 717600 205866
rect 688901 198832 717600 205598
rect 687949 198528 717600 198832
rect 687949 195691 688145 198528
rect 687293 195387 688145 195691
rect 677707 151862 687193 160598
rect 677707 145534 687067 151862
rect 677707 145406 677927 145534
rect 677707 115666 677927 115807
rect 678007 115746 679097 145454
rect 679177 145406 679297 145534
rect 680387 145486 681477 145534
rect 679177 115666 679297 115807
rect 679377 115746 680307 145454
rect 680387 145406 680507 145486
rect 681357 145406 681477 145486
rect 680587 115807 681277 145406
rect 680387 115727 680507 115807
rect 681357 115727 681477 115807
rect 681557 115746 682487 145454
rect 682567 145406 682687 145534
rect 680387 115666 681477 115727
rect 682567 115666 682687 115807
rect 682767 115746 683697 145454
rect 683777 145406 683897 145534
rect 683777 115666 683897 115807
rect 683977 115746 684667 145454
rect 684747 145406 684867 145534
rect 684747 115666 684867 115807
rect 684947 115746 685637 145454
rect 685717 145406 685837 145534
rect 685717 115666 685837 115807
rect 685917 115746 686847 145454
rect 686927 145406 687067 145534
rect 686927 115666 687067 115807
rect 677707 115398 687067 115666
rect 687147 115478 687213 151782
rect 687273 150771 687869 195307
rect 687949 190534 688145 195387
rect 687929 190200 688165 190454
rect 687949 161200 688145 190200
rect 687929 160946 688165 161200
rect 687949 153832 688145 160866
rect 688225 153912 688821 198448
rect 688901 196862 717600 198528
rect 688881 160678 688947 196782
rect 689027 190534 717600 196862
rect 689027 190406 689167 190534
rect 689027 161200 689167 190200
rect 689027 160866 689167 161007
rect 689247 160946 690137 190454
rect 690217 190406 690337 190534
rect 690217 161200 690337 190200
rect 690217 160866 690337 161007
rect 690417 160946 691307 190454
rect 691387 190406 691527 190534
rect 691607 190200 696600 190454
rect 696680 190406 712677 190534
rect 712757 190200 717600 190454
rect 691387 161200 717600 190200
rect 691387 160866 691527 161007
rect 691607 160946 696600 161200
rect 696680 160866 712677 161007
rect 712757 160946 717600 161200
rect 689027 160598 717600 160866
rect 688901 153832 717600 160598
rect 687949 153528 717600 153832
rect 687949 150691 688145 153528
rect 687293 150387 688145 150691
rect 677707 106662 687193 115398
rect 677707 100334 687067 106662
rect 677707 100206 677927 100334
rect 40171 84284 40237 84285
rect 40171 84220 40172 84284
rect 40236 84220 40237 84284
rect 40171 84219 40237 84220
rect 30533 68334 39593 82666
rect 30533 68193 30673 68334
rect 30533 40466 30673 40549
rect 30753 40546 31683 68254
rect 31763 68193 31883 68334
rect 31763 40466 31883 40549
rect 31963 40546 32653 68254
rect 32733 68193 32853 68334
rect 32733 40466 32853 40549
rect 32933 40546 33623 68254
rect 33703 68193 33823 68334
rect 33703 40466 33823 40549
rect 33903 40546 34833 68254
rect 34913 68193 35033 68334
rect 36123 68273 37213 68334
rect 34913 40466 35033 40549
rect 35113 40546 36043 68254
rect 36123 68193 36243 68273
rect 37093 68193 37213 68273
rect 36323 40549 37013 68193
rect 36123 40469 36243 40549
rect 37093 40469 37213 40549
rect 37293 40546 38223 68254
rect 38303 68193 38423 68334
rect 36123 40466 37213 40469
rect 38303 40466 38423 40549
rect 38503 40546 39593 68254
rect 39673 40466 40000 40549
rect 30533 39673 40000 40466
rect 186606 39673 202207 39893
rect 295206 39673 310807 39893
rect 350006 39673 365607 39893
rect 404806 39673 420407 39893
rect 459606 39673 475207 39893
rect 514406 39673 530007 39893
rect 677051 39673 677927 40000
rect 30533 38423 39450 39673
rect 39530 38503 79054 39593
rect 79134 38423 93466 39593
rect 93546 38503 186654 39593
rect 30533 38303 40000 38423
rect 78993 38303 93607 38423
rect 30533 37213 39163 38303
rect 39243 37293 79054 38223
rect 79134 37213 93466 38303
rect 132600 38223 147600 38503
rect 186734 38423 202066 39673
rect 202146 38503 241454 39593
rect 241534 38423 255866 39593
rect 255946 38503 295254 39593
rect 295334 38423 310666 39673
rect 310746 38503 350054 39593
rect 350134 38423 365466 39673
rect 365546 38503 404854 39593
rect 404934 38423 420266 39673
rect 420346 38503 459654 39593
rect 459734 38423 475066 39673
rect 475146 38503 514454 39593
rect 514534 38423 529866 39673
rect 529946 38503 569254 39593
rect 569334 38423 583666 39593
rect 583746 38503 623054 39593
rect 623134 38423 637466 39593
rect 637546 38503 677054 39593
rect 677134 39450 677927 39673
rect 678007 39530 679097 100254
rect 679177 100206 679297 100334
rect 680387 100286 681477 100334
rect 679377 71000 680307 100254
rect 680387 100206 680507 100286
rect 681357 100206 681477 100286
rect 680587 70000 681277 100206
rect 679177 39450 679297 40000
rect 677134 39163 679297 39450
rect 679377 39243 680307 70000
rect 680387 39626 680507 40000
rect 680587 39706 681277 69000
rect 681357 39626 681477 40000
rect 681557 39695 682487 100254
rect 682567 100206 682687 100334
rect 680387 39615 681477 39626
rect 682567 39615 682687 40000
rect 682767 39680 683697 100254
rect 683777 100206 683897 100334
rect 680387 39600 682687 39615
rect 683777 39643 683897 40000
rect 683977 39723 684667 100254
rect 684747 100206 684867 100334
rect 684947 70000 685637 100254
rect 685717 100206 685837 100334
rect 685917 71000 686847 100254
rect 686927 100206 687067 100334
rect 687147 70000 687213 106582
rect 687273 105571 687869 150307
rect 687949 145534 688145 150387
rect 687929 145200 688165 145454
rect 687949 116000 688145 145200
rect 687929 115746 688165 116000
rect 687949 108632 688145 115666
rect 688225 108712 688821 153448
rect 688901 151862 717600 153528
rect 688881 115478 688947 151782
rect 689027 145534 717600 151862
rect 689027 145406 689167 145534
rect 689027 116000 689167 145200
rect 689027 115666 689167 115807
rect 689247 115746 690137 145454
rect 690217 145406 690337 145534
rect 690217 116000 690337 145200
rect 690217 115666 690337 115807
rect 690417 115746 691307 145454
rect 691387 145406 691527 145534
rect 691607 145200 696600 145454
rect 696680 145406 712677 145534
rect 712757 145200 717600 145454
rect 691387 116000 717600 145200
rect 691387 115666 691527 115807
rect 691607 115746 696600 116000
rect 696680 115666 712677 115807
rect 712757 115746 717600 116000
rect 689027 115398 717600 115666
rect 688901 108632 717600 115398
rect 687949 108328 717600 108632
rect 687949 105491 688145 108328
rect 687293 105187 688145 105491
rect 684747 39653 684867 40000
rect 684947 39733 685637 69000
rect 685717 39653 685837 40000
rect 685917 39705 686847 70000
rect 684747 39643 685837 39653
rect 683777 39625 685837 39643
rect 686927 39625 687067 40000
rect 683777 39600 687067 39625
rect 680387 39163 687067 39600
rect 677134 38423 687067 39163
rect 186606 38303 202207 38423
rect 241393 38303 256007 38423
rect 295206 38303 310807 38423
rect 350006 38303 365607 38423
rect 404806 38303 420407 38423
rect 459606 38303 475207 38423
rect 514406 38303 530007 38423
rect 569193 38303 583807 38423
rect 622993 38303 637607 38423
rect 677051 38303 687067 38423
rect 93546 37293 186654 38223
rect 30533 37093 40000 37213
rect 78993 37093 93607 37213
rect 30533 36243 39626 37093
rect 39706 36323 78993 37013
rect 79073 36243 93527 37093
rect 132600 37013 147600 37293
rect 186734 37213 202066 38303
rect 202146 37293 241454 38223
rect 241534 37213 255866 38303
rect 255946 37293 295254 38223
rect 295334 37213 310666 38303
rect 310746 37293 350054 38223
rect 350134 37213 365466 38303
rect 365546 37293 404854 38223
rect 404934 37213 420266 38303
rect 420346 37293 459654 38223
rect 459734 37213 475066 38303
rect 475146 37293 514454 38223
rect 514534 37213 529866 38303
rect 529946 37293 569254 38223
rect 569334 37213 583666 38303
rect 583746 37293 623054 38223
rect 623134 37213 637466 38303
rect 637546 37293 677054 38223
rect 677134 37213 687067 38303
rect 186606 37093 202207 37213
rect 241393 37093 256007 37213
rect 295206 37093 310807 37213
rect 350006 37093 365607 37213
rect 404806 37093 420407 37213
rect 459606 37093 475207 37213
rect 514406 37093 530007 37213
rect 569193 37093 583807 37213
rect 622993 37093 637607 37213
rect 677051 37093 687067 37213
rect 93607 36323 186606 37013
rect 30533 36123 40000 36243
rect 78993 36123 93607 36243
rect 30533 36005 39615 36123
rect 29455 35338 39615 36005
rect 28799 35285 39615 35338
rect 0 35033 39615 35285
rect 39695 35977 79054 36043
rect 39695 35175 47646 35977
rect 51144 35175 51646 35977
rect 55144 35175 55646 35977
rect 59144 35175 59646 35977
rect 63144 35175 63646 35977
rect 67144 35175 67646 35977
rect 71144 35175 79054 35977
rect 39695 35113 79054 35175
rect 79134 35033 93466 36123
rect 132600 36043 147600 36323
rect 186686 36243 202127 37093
rect 202207 36323 241393 37013
rect 241473 36243 255927 37093
rect 256007 36323 295206 37013
rect 295286 36243 310727 37093
rect 310807 36323 350006 37013
rect 350086 36243 365527 37093
rect 365607 36323 404806 37013
rect 404886 36243 420327 37093
rect 420407 36323 459606 37013
rect 459686 36243 475127 37093
rect 475207 36323 514406 37013
rect 514486 36243 529927 37093
rect 530007 36323 569193 37013
rect 569273 36243 583727 37093
rect 583807 36323 622993 37013
rect 623073 36243 637527 37093
rect 637607 36323 677051 37013
rect 677131 36243 687067 37093
rect 186606 36123 202207 36243
rect 241393 36123 256007 36243
rect 295206 36123 310807 36243
rect 350006 36123 365607 36243
rect 404806 36123 420407 36243
rect 459606 36123 475207 36243
rect 514406 36123 530007 36243
rect 569193 36123 583807 36243
rect 622993 36123 637607 36243
rect 677051 36123 687067 36243
rect 93546 35977 186654 36043
rect 93546 35175 101446 35977
rect 104944 35175 105446 35977
rect 108944 35175 109446 35977
rect 112944 35175 113446 35977
rect 116944 35175 117446 35977
rect 120944 35175 121446 35977
rect 124944 35175 155246 35977
rect 158744 35175 159246 35977
rect 162744 35175 163246 35977
rect 166744 35175 167246 35977
rect 170744 35175 171246 35977
rect 174744 35175 175246 35977
rect 178744 35175 186654 35977
rect 93546 35113 186654 35175
rect 0 34913 40000 35033
rect 78993 34913 93607 35033
rect 0 33823 39600 34913
rect 39680 33903 79054 34833
rect 79134 33823 93466 34913
rect 132600 34833 147600 35113
rect 186734 35033 202066 36123
rect 202146 35977 241454 36043
rect 202146 35175 210046 35977
rect 213544 35175 214046 35977
rect 217544 35175 218046 35977
rect 221544 35175 222046 35977
rect 225544 35175 226046 35977
rect 229544 35175 230046 35977
rect 233544 35175 241454 35977
rect 202146 35113 241454 35175
rect 241534 35033 255866 36123
rect 255946 35977 295254 36043
rect 255946 35175 263846 35977
rect 267344 35175 267846 35977
rect 271344 35175 271846 35977
rect 275344 35175 275846 35977
rect 279344 35175 279846 35977
rect 283344 35175 283846 35977
rect 287344 35175 295254 35977
rect 255946 35113 295254 35175
rect 295334 35033 310666 36123
rect 310746 35977 350054 36043
rect 310746 35175 318646 35977
rect 322144 35175 322646 35977
rect 326144 35175 326646 35977
rect 330144 35175 330646 35977
rect 334144 35175 334646 35977
rect 338144 35175 338646 35977
rect 342144 35175 350054 35977
rect 310746 35113 350054 35175
rect 350134 35033 365466 36123
rect 365546 35977 404854 36043
rect 365546 35175 373446 35977
rect 376944 35175 377446 35977
rect 380944 35175 381446 35977
rect 384944 35175 385446 35977
rect 388944 35175 389446 35977
rect 392944 35175 393446 35977
rect 396944 35175 404854 35977
rect 365546 35113 404854 35175
rect 404934 35033 420266 36123
rect 420346 35977 459654 36043
rect 420346 35175 428246 35977
rect 431744 35175 432246 35977
rect 435744 35175 436246 35977
rect 439744 35175 440246 35977
rect 443744 35175 444246 35977
rect 447744 35175 448246 35977
rect 451744 35175 459654 35977
rect 420346 35113 459654 35175
rect 459734 35033 475066 36123
rect 475146 35977 514454 36043
rect 475146 35175 483046 35977
rect 486544 35175 487046 35977
rect 490544 35175 491046 35977
rect 494544 35175 495046 35977
rect 498544 35175 499046 35977
rect 502544 35175 503046 35977
rect 506544 35175 514454 35977
rect 475146 35113 514454 35175
rect 514534 35033 529866 36123
rect 529946 35977 569254 36043
rect 529946 35175 537846 35977
rect 541344 35175 541846 35977
rect 545344 35175 545846 35977
rect 549344 35175 549846 35977
rect 553344 35175 553846 35977
rect 557344 35175 557846 35977
rect 561344 35175 569254 35977
rect 529946 35113 569254 35175
rect 569334 35033 583666 36123
rect 583746 35977 623054 36043
rect 583746 35175 591646 35977
rect 595144 35175 595646 35977
rect 599144 35175 599646 35977
rect 603144 35175 603646 35977
rect 607144 35175 607646 35977
rect 611144 35175 611646 35977
rect 615144 35175 623054 35977
rect 583746 35113 623054 35175
rect 623134 35033 637466 36123
rect 637546 35977 677054 36043
rect 637546 35175 645446 35977
rect 648944 35175 649446 35977
rect 652944 35175 653446 35977
rect 656944 35175 657446 35977
rect 660944 35175 661446 35977
rect 664944 35175 665446 35977
rect 668944 35175 677054 35977
rect 637546 35113 677054 35175
rect 677134 36005 687067 36123
rect 687147 36085 687213 69000
rect 677134 35733 687193 36005
rect 687273 35813 687869 105107
rect 687949 100334 688145 105187
rect 687929 100000 688165 100254
rect 687949 70000 688145 100000
rect 687949 40000 688145 69000
rect 677134 35610 687849 35733
rect 687929 35690 688165 40000
rect 677134 35338 688145 35610
rect 688225 35418 688821 108248
rect 688901 106662 717600 108328
rect 688881 70000 688947 106582
rect 689027 100334 717600 106662
rect 689027 100206 689167 100334
rect 689027 70000 689167 100000
rect 688881 35365 688947 69000
rect 689027 39595 689167 69000
rect 689247 39675 690137 100254
rect 690217 100206 690337 100334
rect 690217 70000 690337 100000
rect 690217 39624 690337 69000
rect 690417 39704 691307 100254
rect 691387 100206 691527 100334
rect 691607 100000 696600 100254
rect 696680 100206 712677 100334
rect 712757 100000 717600 100254
rect 691387 70000 717600 100000
rect 691607 69000 717600 70000
rect 691387 40000 717600 69000
rect 691387 39624 691527 40000
rect 690217 39595 691527 39624
rect 689027 39391 691527 39595
rect 691607 39471 696600 40000
rect 696680 39633 712677 40000
rect 712757 39713 717600 40000
rect 696680 39391 717600 39633
rect 677134 35285 688801 35338
rect 689027 35285 717600 39391
rect 677134 35033 717600 35285
rect 186606 34913 202207 35033
rect 241393 34913 256007 35033
rect 295206 34913 310807 35033
rect 350006 34913 365607 35033
rect 404806 34913 420407 35033
rect 459606 34913 475207 35033
rect 514406 34913 530007 35033
rect 569193 34913 583807 35033
rect 622993 34913 637607 35033
rect 677051 34913 717600 35033
rect 93546 33903 186654 34833
rect 0 33703 40000 33823
rect 78993 33703 93607 33823
rect 0 32853 39643 33703
rect 39723 33577 79054 33623
rect 39723 32987 47652 33577
rect 51182 32987 51652 33577
rect 55182 32987 55652 33577
rect 59182 32987 59652 33577
rect 63182 32987 63652 33577
rect 67182 32987 67652 33577
rect 71182 32987 79054 33577
rect 39723 32933 79054 32987
rect 79134 32853 93466 33703
rect 132600 33623 147600 33903
rect 186734 33823 202066 34913
rect 202146 33903 241454 34833
rect 241534 33823 255866 34913
rect 255946 33903 295254 34833
rect 295334 33823 310666 34913
rect 310746 33903 350054 34833
rect 350134 33823 365466 34913
rect 365546 33903 404854 34833
rect 404934 33823 420266 34913
rect 420346 33903 459654 34833
rect 459734 33823 475066 34913
rect 475146 33903 514454 34833
rect 514534 33823 529866 34913
rect 529946 33903 569254 34833
rect 569334 33823 583666 34913
rect 583746 33903 623054 34833
rect 623134 33823 637466 34913
rect 637546 33903 677054 34833
rect 677134 33823 717600 34913
rect 186606 33703 202207 33823
rect 241393 33703 256007 33823
rect 295206 33703 310807 33823
rect 350006 33703 365607 33823
rect 404806 33703 420407 33823
rect 459606 33703 475207 33823
rect 514406 33703 530007 33823
rect 569193 33703 583807 33823
rect 622993 33703 637607 33823
rect 677051 33703 717600 33823
rect 93546 33577 186654 33623
rect 93546 32987 101452 33577
rect 104982 32987 105452 33577
rect 108982 32987 109452 33577
rect 112982 32987 113452 33577
rect 116982 32987 117452 33577
rect 120982 32987 121452 33577
rect 124982 32987 155252 33577
rect 158782 32987 159252 33577
rect 162782 32987 163252 33577
rect 166782 32987 167252 33577
rect 170782 32987 171252 33577
rect 174782 32987 175252 33577
rect 178782 32987 186654 33577
rect 93546 32933 186654 32987
rect 0 32733 40000 32853
rect 78993 32733 93607 32853
rect 0 31883 39653 32733
rect 39733 31963 79054 32653
rect 79134 31883 93466 32733
rect 132600 32653 147600 32933
rect 186734 32853 202066 33703
rect 202146 33577 241454 33623
rect 202146 32987 210052 33577
rect 213582 32987 214052 33577
rect 217582 32987 218052 33577
rect 221582 32987 222052 33577
rect 225582 32987 226052 33577
rect 229582 32987 230052 33577
rect 233582 32987 241454 33577
rect 202146 32933 241454 32987
rect 241534 32853 255866 33703
rect 255946 33577 295254 33623
rect 255946 32987 263852 33577
rect 267382 32987 267852 33577
rect 271382 32987 271852 33577
rect 275382 32987 275852 33577
rect 279382 32987 279852 33577
rect 283382 32987 283852 33577
rect 287382 32987 295254 33577
rect 255946 32933 295254 32987
rect 295334 32853 310666 33703
rect 310746 33577 350054 33623
rect 310746 32987 318652 33577
rect 322182 32987 322652 33577
rect 326182 32987 326652 33577
rect 330182 32987 330652 33577
rect 334182 32987 334652 33577
rect 338182 32987 338652 33577
rect 342182 32987 350054 33577
rect 310746 32933 350054 32987
rect 350134 32853 365466 33703
rect 365546 33577 404854 33623
rect 365546 32987 373452 33577
rect 376982 32987 377452 33577
rect 380982 32987 381452 33577
rect 384982 32987 385452 33577
rect 388982 32987 389452 33577
rect 392982 32987 393452 33577
rect 396982 32987 404854 33577
rect 365546 32933 404854 32987
rect 404934 32853 420266 33703
rect 420346 33577 459654 33623
rect 420346 32987 428252 33577
rect 431782 32987 432252 33577
rect 435782 32987 436252 33577
rect 439782 32987 440252 33577
rect 443782 32987 444252 33577
rect 447782 32987 448252 33577
rect 451782 32987 459654 33577
rect 420346 32933 459654 32987
rect 459734 32853 475066 33703
rect 475146 33577 514454 33623
rect 475146 32987 483052 33577
rect 486582 32987 487052 33577
rect 490582 32987 491052 33577
rect 494582 32987 495052 33577
rect 498582 32987 499052 33577
rect 502582 32987 503052 33577
rect 506582 32987 514454 33577
rect 475146 32933 514454 32987
rect 514534 32853 529866 33703
rect 529946 33577 569254 33623
rect 529946 32987 537852 33577
rect 541382 32987 541852 33577
rect 545382 32987 545852 33577
rect 549382 32987 549852 33577
rect 553382 32987 553852 33577
rect 557382 32987 557852 33577
rect 561382 32987 569254 33577
rect 529946 32933 569254 32987
rect 569334 32853 583666 33703
rect 583746 33577 623054 33623
rect 583746 32987 591652 33577
rect 595182 32987 595652 33577
rect 599182 32987 599652 33577
rect 603182 32987 603652 33577
rect 607182 32987 607652 33577
rect 611182 32987 611652 33577
rect 615182 32987 623054 33577
rect 583746 32933 623054 32987
rect 623134 32853 637466 33703
rect 637546 33577 677054 33623
rect 637546 32987 645452 33577
rect 648982 32987 649452 33577
rect 652982 32987 653452 33577
rect 656982 32987 657452 33577
rect 660982 32987 661452 33577
rect 664982 32987 665452 33577
rect 668982 32987 677054 33577
rect 637546 32933 677054 32987
rect 677134 32853 717600 33703
rect 186606 32733 202207 32853
rect 241393 32733 256007 32853
rect 295206 32733 310807 32853
rect 350006 32733 365607 32853
rect 404806 32733 420407 32853
rect 459606 32733 475207 32853
rect 514406 32733 530007 32853
rect 569193 32733 583807 32853
rect 622993 32733 637607 32853
rect 677051 32733 717600 32853
rect 93546 31963 186654 32653
rect 0 31763 40000 31883
rect 78993 31763 93607 31883
rect 0 30673 39625 31763
rect 39705 30753 79054 31683
rect 79134 30673 93466 31763
rect 132600 31683 147600 31963
rect 186734 31883 202066 32733
rect 202146 31963 241454 32653
rect 241534 31883 255866 32733
rect 255946 31963 295254 32653
rect 295334 31883 310666 32733
rect 310746 31963 350054 32653
rect 350134 31883 365466 32733
rect 365546 31963 404854 32653
rect 404934 31883 420266 32733
rect 420346 31963 459654 32653
rect 459734 31883 475066 32733
rect 475146 31963 514454 32653
rect 514534 31883 529866 32733
rect 529946 31963 569254 32653
rect 569334 31883 583666 32733
rect 583746 31963 623054 32653
rect 623134 31883 637466 32733
rect 637546 31963 677054 32653
rect 677134 31883 717600 32733
rect 186606 31763 202207 31883
rect 241393 31763 256007 31883
rect 295206 31763 310807 31883
rect 350006 31763 365607 31883
rect 404806 31763 420407 31883
rect 459606 31763 475207 31883
rect 514406 31763 530007 31883
rect 569193 31763 583807 31883
rect 622993 31763 637607 31883
rect 677051 31763 717600 31883
rect 93546 30753 186654 31683
rect 0 30533 40000 30673
rect 78993 30533 93607 30673
rect 0 30407 36005 30533
rect 0 29751 35733 30407
rect 36085 30387 79054 30453
rect 79134 30407 93466 30533
rect 132600 30453 147600 30753
rect 186734 30673 202066 31763
rect 202146 30753 241454 31683
rect 241534 30673 255866 31763
rect 255946 30753 295254 31683
rect 295334 30673 310666 31763
rect 310746 30753 350054 31683
rect 350134 30673 365466 31763
rect 365546 30753 404854 31683
rect 404934 30673 420266 31763
rect 420346 30753 459654 31683
rect 459734 30673 475066 31763
rect 475146 30753 514454 31683
rect 514534 30673 529866 31763
rect 529946 30753 569254 31683
rect 569334 30673 583666 31763
rect 583746 30753 623054 31683
rect 623134 30673 637466 31763
rect 637546 30753 677054 31683
rect 677134 30673 717600 31763
rect 186606 30533 202207 30673
rect 241393 30533 256007 30673
rect 295206 30533 310807 30673
rect 350006 30533 365607 30673
rect 404806 30533 420407 30673
rect 459606 30533 475207 30673
rect 514406 30533 530007 30673
rect 569193 30533 583807 30673
rect 622993 30533 637607 30673
rect 677051 30533 717600 30673
rect 93546 30407 192982 30453
rect 193062 30407 201798 30533
rect 93546 30387 132600 30407
rect 147600 30387 192982 30407
rect 201878 30387 301582 30453
rect 301662 30407 310398 30533
rect 310478 30387 356382 30453
rect 356462 30407 365198 30533
rect 365278 30387 411182 30453
rect 411262 30407 419998 30533
rect 420078 30387 465982 30453
rect 466062 30407 474798 30533
rect 474878 30387 520782 30453
rect 520862 30407 529598 30533
rect 529678 30387 681515 30453
rect 0 29455 35610 29751
rect 35813 29731 191507 30327
rect 35690 29651 40000 29671
rect 47400 29651 71400 29671
rect 78800 29651 79054 29671
rect 93546 29651 93800 29671
rect 101200 29651 125200 29671
rect 155000 29651 179000 29671
rect 186400 29651 186654 29671
rect 191587 29651 191891 30307
rect 191971 29731 300107 30327
rect 202146 29651 202400 29671
rect 209800 29651 233800 29671
rect 241200 29651 241454 29671
rect 255946 29651 256200 29671
rect 263600 29651 287600 29671
rect 295000 29651 295254 29671
rect 300187 29651 300491 30307
rect 300571 29731 354907 30327
rect 310746 29651 311000 29671
rect 318400 29651 342400 29671
rect 349800 29651 350054 29671
rect 354987 29651 355291 30307
rect 355371 29731 409707 30327
rect 365546 29651 365800 29671
rect 373200 29651 397200 29671
rect 404600 29651 404854 29671
rect 409787 29651 410091 30307
rect 410171 29731 464507 30327
rect 420346 29651 420600 29671
rect 428000 29651 452000 29671
rect 459400 29651 459654 29671
rect 464587 29651 464891 30307
rect 464971 29731 519307 30327
rect 475146 29651 475400 29671
rect 482800 29651 506800 29671
rect 514200 29651 514454 29671
rect 519387 29651 519691 30307
rect 519771 29731 680975 30327
rect 681595 30307 717600 30533
rect 681055 29751 717600 30307
rect 529946 29651 530200 29671
rect 537600 29651 561600 29671
rect 569000 29651 569254 29671
rect 583746 29651 584000 29671
rect 591400 29651 615400 29671
rect 622800 29651 623054 29671
rect 637546 29651 637800 29671
rect 645200 29651 669200 29671
rect 676800 29651 681111 29671
rect 35690 29455 79054 29651
rect 79134 29455 93466 29651
rect 93546 29455 186654 29651
rect 186734 29455 202066 29651
rect 202146 29455 241454 29651
rect 241534 29455 255866 29651
rect 255946 29455 295254 29651
rect 295334 29455 310666 29651
rect 310746 29455 350054 29651
rect 350134 29455 365466 29651
rect 365546 29455 404854 29651
rect 404934 29455 420266 29651
rect 420346 29455 459654 29651
rect 459734 29455 475066 29651
rect 475146 29455 514454 29651
rect 514534 29455 529866 29651
rect 529946 29455 569254 29651
rect 569334 29455 583666 29651
rect 583746 29455 623054 29651
rect 623134 29455 637466 29651
rect 637546 29455 681111 29651
rect 681191 29455 717600 29751
rect 0 28799 35338 29455
rect 35690 29435 40000 29455
rect 47400 29435 71400 29455
rect 78800 29435 79054 29455
rect 93546 29435 93800 29455
rect 101200 29435 125200 29455
rect 155000 29435 179000 29455
rect 186400 29435 186654 29455
rect 0 28573 35285 28799
rect 35418 28779 194648 29375
rect 35365 28653 79054 28719
rect 93546 28699 132600 28719
rect 147600 28699 192982 28719
rect 194728 28699 195032 29455
rect 202146 29435 202400 29455
rect 209800 29435 233800 29455
rect 241200 29435 241454 29455
rect 255946 29435 256200 29455
rect 263600 29435 287600 29455
rect 295000 29435 295254 29455
rect 195112 28779 303248 29375
rect 79134 28573 93466 28699
rect 93546 28653 192982 28699
rect 132600 28573 147600 28653
rect 193062 28573 201798 28699
rect 201878 28653 301582 28719
rect 303328 28699 303632 29455
rect 310746 29435 311000 29455
rect 318400 29435 342400 29455
rect 349800 29435 350054 29455
rect 303712 28779 358048 29375
rect 301662 28573 310398 28699
rect 310478 28653 356382 28719
rect 358128 28699 358432 29455
rect 365546 29435 365800 29455
rect 373200 29435 397200 29455
rect 404600 29435 404854 29455
rect 358512 28779 412848 29375
rect 356462 28573 365198 28699
rect 365278 28653 411182 28719
rect 412928 28699 413232 29455
rect 420346 29435 420600 29455
rect 428000 29435 452000 29455
rect 459400 29435 459654 29455
rect 413312 28779 467648 29375
rect 411262 28573 419998 28699
rect 420078 28653 465982 28719
rect 467728 28699 468032 29455
rect 475146 29435 475400 29455
rect 482800 29435 506800 29455
rect 514200 29435 514454 29455
rect 468112 28779 522448 29375
rect 466062 28573 474798 28699
rect 474878 28653 520782 28719
rect 522528 28699 522832 29455
rect 529946 29435 530200 29455
rect 537600 29435 561600 29455
rect 569000 29435 569254 29455
rect 583746 29435 584000 29455
rect 591400 29435 615400 29455
rect 622800 29435 623054 29455
rect 637546 29435 637800 29455
rect 645200 29435 669200 29455
rect 676800 29435 681111 29455
rect 522912 28779 682182 29375
rect 682262 28799 717600 29455
rect 520862 28573 529598 28699
rect 529678 28653 682235 28719
rect 682315 28573 717600 28799
rect 0 28433 47400 28573
rect 71400 28433 78800 28573
rect 78993 28433 93607 28573
rect 93800 28433 101200 28573
rect 125200 28433 155000 28573
rect 179000 28433 186400 28573
rect 186606 28433 202207 28573
rect 202400 28433 209800 28573
rect 233800 28433 241200 28573
rect 241393 28433 256007 28573
rect 256200 28433 263600 28573
rect 287600 28433 295000 28573
rect 295206 28433 310807 28573
rect 311000 28433 318400 28573
rect 342400 28433 349800 28573
rect 350006 28433 365607 28573
rect 365800 28433 373200 28573
rect 397200 28433 404600 28573
rect 404806 28433 420407 28573
rect 420600 28433 428000 28573
rect 452000 28433 459400 28573
rect 459606 28433 475207 28573
rect 475400 28433 482800 28573
rect 506800 28433 514200 28573
rect 514406 28433 530007 28573
rect 530200 28433 537600 28573
rect 561600 28433 569000 28573
rect 569193 28433 583807 28573
rect 584000 28433 591400 28573
rect 615400 28433 622800 28573
rect 622993 28433 637607 28573
rect 637800 28433 645200 28573
rect 669200 28433 676800 28573
rect 677051 28433 717600 28573
rect 0 27383 39595 28433
rect 39675 27463 79054 28353
rect 79134 27383 93466 28433
rect 132600 28353 147600 28433
rect 93546 27463 186654 28353
rect 132600 27383 147600 27463
rect 186734 27383 202066 28433
rect 202146 27463 241454 28353
rect 241534 27383 255866 28433
rect 255946 27463 295254 28353
rect 295334 27383 310666 28433
rect 310746 27463 350054 28353
rect 350134 27383 365466 28433
rect 365546 27463 404854 28353
rect 404934 27383 420266 28433
rect 420346 27463 459654 28353
rect 459734 27383 475066 28433
rect 475146 27463 514454 28353
rect 514534 27383 529866 28433
rect 529946 27463 569254 28353
rect 569334 27383 583666 28433
rect 583746 27463 623054 28353
rect 623134 27383 637466 28433
rect 637546 27463 677054 28353
rect 677134 27383 717600 28433
rect 0 27263 47400 27383
rect 71400 27263 78800 27383
rect 78993 27263 93607 27383
rect 93800 27263 101200 27383
rect 125200 27263 155000 27383
rect 179000 27263 186400 27383
rect 186606 27263 202207 27383
rect 202400 27263 209800 27383
rect 233800 27263 241200 27383
rect 241393 27263 256007 27383
rect 256200 27263 263600 27383
rect 287600 27263 295000 27383
rect 295206 27263 310807 27383
rect 311000 27263 318400 27383
rect 342400 27263 349800 27383
rect 350006 27263 365607 27383
rect 365800 27263 373200 27383
rect 397200 27263 404600 27383
rect 404806 27263 420407 27383
rect 420600 27263 428000 27383
rect 452000 27263 459400 27383
rect 459606 27263 475207 27383
rect 475400 27263 482800 27383
rect 506800 27263 514200 27383
rect 514406 27263 530007 27383
rect 530200 27263 537600 27383
rect 561600 27263 569000 27383
rect 569193 27263 583807 27383
rect 584000 27263 591400 27383
rect 615400 27263 622800 27383
rect 622993 27263 637607 27383
rect 637800 27263 645200 27383
rect 669200 27263 676800 27383
rect 677051 27263 717600 27383
rect 0 26213 39624 27263
rect 39704 26293 79054 27183
rect 79134 26213 93466 27263
rect 132600 27183 147600 27263
rect 93546 26293 186654 27183
rect 132600 26213 147600 26293
rect 186734 26213 202066 27263
rect 202146 26293 241454 27183
rect 241534 26213 255866 27263
rect 255946 26293 295254 27183
rect 295334 26213 310666 27263
rect 310746 26293 350054 27183
rect 350134 26213 365466 27263
rect 365546 26293 404854 27183
rect 404934 26213 420266 27263
rect 420346 26293 459654 27183
rect 459734 26213 475066 27263
rect 475146 26293 514454 27183
rect 514534 26213 529866 27263
rect 529946 26293 569254 27183
rect 569334 26213 583666 27263
rect 583746 26293 623054 27183
rect 623134 26213 637466 27263
rect 637546 26293 677054 27183
rect 677134 26213 717600 27263
rect 0 26073 47400 26213
rect 0 20920 39391 26073
rect 40000 25993 47400 26073
rect 71400 25993 78800 26213
rect 78993 26073 93607 26213
rect 39471 21000 79054 25993
rect 40000 20920 47400 21000
rect 0 4923 47400 20920
rect 0 0 39633 4923
rect 40000 4843 47400 4923
rect 71400 4843 78800 21000
rect 79134 20920 93466 26073
rect 93800 25993 101200 26213
rect 125200 25993 155000 26213
rect 179000 25993 186400 26213
rect 186606 26073 202207 26213
rect 93546 21000 186654 25993
rect 78993 4923 93607 20920
rect 39713 0 79054 4843
rect 79134 0 93466 4923
rect 93800 4843 101200 21000
rect 125200 4843 155000 21000
rect 179000 4843 186400 21000
rect 186734 20920 202066 26073
rect 202400 25993 209800 26213
rect 233800 25993 241200 26213
rect 241393 26073 256007 26213
rect 202146 21000 241454 25993
rect 186606 4923 202207 20920
rect 93546 0 186654 4843
rect 186734 0 202066 4923
rect 202400 4843 209800 21000
rect 233800 4843 241200 21000
rect 241534 20920 255866 26073
rect 256200 25993 263600 26213
rect 287600 25993 295000 26213
rect 295206 26073 310807 26213
rect 255946 21000 295254 25993
rect 241393 4923 256007 20920
rect 202146 0 241454 4843
rect 241534 0 255866 4923
rect 256200 4843 263600 21000
rect 287600 4843 295000 21000
rect 295334 20920 310666 26073
rect 311000 25993 318400 26213
rect 342400 25993 349800 26213
rect 350006 26073 365607 26213
rect 310746 21000 350054 25993
rect 295206 4923 310807 20920
rect 255946 0 295254 4843
rect 295334 0 310666 4923
rect 311000 4843 318400 21000
rect 342400 4843 349800 21000
rect 350134 20920 365466 26073
rect 365800 25993 373200 26213
rect 397200 25993 404600 26213
rect 404806 26073 420407 26213
rect 365546 21000 404854 25993
rect 350006 4923 365607 20920
rect 310746 0 350054 4843
rect 350134 0 365466 4923
rect 365800 4843 373200 21000
rect 397200 4843 404600 21000
rect 404934 20920 420266 26073
rect 420600 25993 428000 26213
rect 452000 25993 459400 26213
rect 459606 26073 475207 26213
rect 420346 21000 459654 25993
rect 404806 4923 420407 20920
rect 365546 0 404854 4843
rect 404934 0 420266 4923
rect 420600 4843 428000 21000
rect 452000 4843 459400 21000
rect 459734 20920 475066 26073
rect 475400 25993 482800 26213
rect 506800 25993 514200 26213
rect 514406 26073 530007 26213
rect 475146 21000 514454 25993
rect 459606 4923 475207 20920
rect 420346 0 459654 4843
rect 459734 0 475066 4923
rect 475400 4843 482800 21000
rect 506800 4843 514200 21000
rect 514534 20920 529866 26073
rect 530200 25993 537600 26213
rect 561600 25993 569000 26213
rect 569193 26073 583807 26213
rect 529946 21000 569254 25993
rect 514406 4923 530007 20920
rect 475146 0 514454 4843
rect 514534 0 529866 4923
rect 530200 4843 537600 21000
rect 561600 4843 569000 21000
rect 569334 20920 583666 26073
rect 584000 25993 591400 26213
rect 615400 25993 622800 26213
rect 622993 26073 637607 26213
rect 583746 21000 623054 25993
rect 569193 4923 583807 20920
rect 529946 0 569254 4843
rect 569334 0 583666 4923
rect 584000 4843 591400 21000
rect 615400 4843 622800 21000
rect 623134 20920 637466 26073
rect 637800 25993 645200 26213
rect 669200 25993 676800 26213
rect 677051 26073 717600 26213
rect 637546 21000 677171 25993
rect 622993 4923 637607 20920
rect 583746 0 623054 4843
rect 623134 0 637466 4923
rect 637800 4843 645200 21000
rect 669200 4843 676800 21000
rect 677251 20920 717600 26073
rect 677051 4923 717600 20920
rect 637546 0 677054 4843
rect 677134 0 717600 4923
<< metal5 >>
rect 78440 1018512 90960 1031002
rect 129840 1018512 142360 1031002
rect 181240 1018512 193760 1031002
rect 232640 1018512 245160 1031002
rect 284240 1018512 296760 1031002
rect 334620 1018402 347160 1030925
rect 386040 1018512 398560 1031002
rect 475040 1018512 487560 1031002
rect 526440 1018512 538960 1031002
rect 576820 1018402 589360 1030925
rect 628240 1018512 640760 1031002
rect 6598 956440 19088 968960
rect 698512 952840 711002 965360
rect 6086 913863 19572 925191
rect 698028 909409 711514 920737
rect 698512 863640 711002 876160
rect 6675 828820 19198 841360
rect 698402 819640 710925 832180
rect 6598 786640 19088 799160
rect 698512 774440 711002 786960
rect 6598 743440 19088 755960
rect 698512 729440 711002 741960
rect 6598 700240 19088 712760
rect 698512 684440 711002 696960
rect 6598 657040 19088 669560
rect 698512 639240 711002 651760
rect 6598 613840 19088 626360
rect 698512 594240 711002 606760
rect 6598 570640 19088 583160
rect 698512 549040 711002 561560
rect 6598 527440 19088 539960
rect 6675 484220 19198 496760
rect 698028 461609 711514 472937
rect 6086 442663 19572 453991
rect 6598 399840 19088 412360
rect 698512 371840 711002 384360
rect 6598 356640 19088 369160
rect 6598 313440 19088 325960
rect 698512 326640 711002 339160
rect 6598 270240 19088 282760
rect 698512 281640 711002 294160
rect 6598 227040 19088 239560
rect 698512 236640 711002 249160
rect 6598 183840 19088 196360
rect 698512 191440 711002 203960
rect 698512 146440 711002 158960
rect 6675 111420 19198 123960
rect 698512 101240 711002 113760
rect 6086 69863 19572 81191
rect 80040 6675 92580 19198
rect 133840 6675 146380 19198
rect 187640 6598 200160 19088
rect 243009 6086 254337 19572
rect 296240 6598 308760 19088
rect 351040 6598 363560 19088
rect 405840 6598 418360 19088
rect 460640 6598 473160 19088
rect 515440 6598 527960 19088
rect 624040 6675 636580 19198
<< obsm5 >>
rect 0 1032757 717600 1037600
rect 0 1016917 40800 1032757
rect 76200 1031322 92200 1032757
rect 76200 1018192 78120 1031322
rect 91280 1018192 92200 1031322
rect 76200 1016917 92200 1018192
rect 127600 1031322 143600 1032757
rect 127600 1018192 129520 1031322
rect 142680 1018192 143600 1031322
rect 127600 1016917 143600 1018192
rect 179000 1031322 195000 1032757
rect 179000 1018192 180920 1031322
rect 194080 1018192 195000 1031322
rect 179000 1016917 195000 1018192
rect 230400 1031322 246400 1032757
rect 230400 1018192 232320 1031322
rect 245480 1018192 246400 1031322
rect 230400 1016917 246400 1018192
rect 282000 1031322 298000 1032757
rect 282000 1018192 283920 1031322
rect 297080 1018192 298000 1031322
rect 282000 1016917 298000 1018192
rect 333400 1031245 348400 1032757
rect 333400 1018082 334300 1031245
rect 347480 1018082 348400 1031245
rect 333400 1016917 348400 1018082
rect 383800 1031322 399800 1032757
rect 383800 1018192 385720 1031322
rect 398880 1018192 399800 1031322
rect 383800 1016917 399800 1018192
rect 472800 1031322 488800 1032757
rect 472800 1018192 474720 1031322
rect 487880 1018192 488800 1031322
rect 472800 1016917 488800 1018192
rect 524200 1031322 540200 1032757
rect 524200 1018192 526120 1031322
rect 539280 1018192 540200 1031322
rect 524200 1016917 540200 1018192
rect 575600 1031245 590600 1032757
rect 575600 1018082 576500 1031245
rect 589680 1018082 590600 1031245
rect 575600 1016917 590600 1018082
rect 626000 1031322 642000 1032757
rect 626000 1018192 627920 1031322
rect 641080 1018192 642000 1031322
rect 626000 1016917 642000 1018192
rect 677600 1016917 717600 1032757
rect 0 1011287 40109 1016917
rect 40800 1016597 41000 1016600
rect 40429 1011607 41000 1016597
rect 41320 1011607 44280 1016597
rect 44600 1011607 45000 1016600
rect 45320 1011607 48280 1016597
rect 48600 1011607 49000 1016600
rect 49320 1011607 52280 1016597
rect 52600 1011607 53000 1016600
rect 53320 1011607 56280 1016597
rect 56600 1011607 57000 1016600
rect 57320 1011607 60280 1016597
rect 60600 1011607 61000 1016600
rect 61320 1011607 64280 1016597
rect 64600 1011607 65000 1016600
rect 65320 1011607 68280 1016597
rect 68600 1011607 69000 1016600
rect 69320 1011607 72280 1016597
rect 72600 1011607 73000 1016600
rect 73320 1011607 74280 1016597
rect 74600 1011607 75000 1016600
rect 75600 1016597 76200 1016600
rect 75600 1011607 76454 1016597
rect 0 1009267 40226 1011287
rect 40546 1010437 76454 1011287
rect 40546 1009267 76454 1010117
rect 0 1006827 35049 1009267
rect 35369 1007147 76454 1008947
rect 0 1002551 40226 1006827
rect 40546 1005937 76454 1006827
rect 40546 1004968 76454 1005617
rect 40800 1004967 76200 1004968
rect 40546 1003997 76454 1004647
rect 40546 1002787 76454 1003677
rect 0 998449 28333 1002551
rect 0 997600 20683 998449
rect 26313 998245 28333 998449
rect 26313 998216 27163 998245
rect 21003 997600 25993 998129
rect 0 970200 4843 997600
rect 21000 997000 25993 997600
rect 21000 996000 25993 996400
rect 21003 994720 25993 995680
rect 21000 994000 25993 994400
rect 21003 990720 25993 993680
rect 21000 990000 25993 990400
rect 21003 986720 25993 989680
rect 21000 986000 25993 986400
rect 21003 982720 25993 985680
rect 21000 982000 25993 982400
rect 21003 978720 25993 981680
rect 21000 978000 25993 978400
rect 21003 974720 25993 977680
rect 21000 974000 25993 974400
rect 21003 970720 25993 973680
rect 21000 970200 25993 970400
rect 0 969626 20683 970200
rect 21003 969946 25993 970200
rect 26313 969946 27163 997896
rect 27483 969946 28333 997925
rect 28653 969946 30453 1002231
rect 30773 1001257 40226 1002551
rect 40546 1001577 76454 1002467
rect 76774 1001257 91626 1016917
rect 92200 1016597 92400 1016600
rect 91946 1011607 92400 1016597
rect 92720 1011607 95680 1016597
rect 96000 1011607 96400 1016600
rect 96720 1011607 99680 1016597
rect 100000 1011607 100400 1016600
rect 100720 1011607 103680 1016597
rect 104000 1011607 104400 1016600
rect 104720 1011607 107680 1016597
rect 108000 1011607 108400 1016600
rect 108720 1011607 111680 1016597
rect 112000 1011607 112400 1016600
rect 112720 1011607 115680 1016597
rect 116000 1011607 116400 1016600
rect 116720 1011607 119680 1016597
rect 120000 1011607 120400 1016600
rect 120720 1011607 123680 1016597
rect 124000 1011607 124400 1016600
rect 124720 1011607 125680 1016597
rect 126000 1011607 126400 1016600
rect 127000 1016597 127600 1016600
rect 127000 1011607 127854 1016597
rect 91946 1010437 127854 1011287
rect 91946 1009267 127854 1010117
rect 91946 1007147 127854 1008947
rect 91946 1005937 127854 1006827
rect 91946 1004968 127854 1005617
rect 92200 1004967 127600 1004968
rect 91946 1003997 127854 1004647
rect 91946 1002787 127854 1003677
rect 91946 1001577 127854 1002467
rect 128174 1001257 143026 1016917
rect 143600 1016597 143800 1016600
rect 143346 1011607 143800 1016597
rect 144120 1011607 147080 1016597
rect 147400 1011607 147800 1016600
rect 148120 1011607 151080 1016597
rect 151400 1011607 151800 1016600
rect 152120 1011607 155080 1016597
rect 155400 1011607 155800 1016600
rect 156120 1011607 159080 1016597
rect 159400 1011607 159800 1016600
rect 160120 1011607 163080 1016597
rect 163400 1011607 163800 1016600
rect 164120 1011607 167080 1016597
rect 167400 1011607 167800 1016600
rect 168120 1011607 171080 1016597
rect 171400 1011607 171800 1016600
rect 172120 1011607 175080 1016597
rect 175400 1011607 175800 1016600
rect 176120 1011607 177080 1016597
rect 177400 1011607 177800 1016600
rect 178400 1016597 179000 1016600
rect 178400 1011607 179254 1016597
rect 143346 1010437 179254 1011287
rect 143346 1009267 179254 1010117
rect 143346 1007147 179254 1008947
rect 143346 1005937 179254 1006827
rect 143346 1004968 179254 1005617
rect 143600 1004967 179000 1004968
rect 143346 1003997 179254 1004647
rect 143346 1002787 179254 1003677
rect 143346 1001577 179254 1002467
rect 179574 1001257 194426 1016917
rect 195000 1016597 195200 1016600
rect 194746 1011607 195200 1016597
rect 195520 1011607 198480 1016597
rect 198800 1011607 199200 1016600
rect 199520 1011607 202480 1016597
rect 202800 1011607 203200 1016600
rect 203520 1011607 206480 1016597
rect 206800 1011607 207200 1016600
rect 207520 1011607 210480 1016597
rect 210800 1011607 211200 1016600
rect 211520 1011607 214480 1016597
rect 214800 1011607 215200 1016600
rect 215520 1011607 218480 1016597
rect 218800 1011607 219200 1016600
rect 219520 1011607 222480 1016597
rect 222800 1011607 223200 1016600
rect 223520 1011607 226480 1016597
rect 226800 1011607 227200 1016600
rect 227520 1011607 228480 1016597
rect 228800 1011607 229200 1016600
rect 229800 1016597 230400 1016600
rect 229800 1011607 230654 1016597
rect 194746 1010437 230654 1011287
rect 194746 1009267 230654 1010117
rect 194746 1007147 230654 1008947
rect 194746 1005937 230654 1006827
rect 194746 1004968 230654 1005617
rect 195000 1004967 230400 1004968
rect 194746 1003997 230654 1004647
rect 194746 1002787 230654 1003677
rect 194746 1001577 230654 1002467
rect 230974 1001257 245826 1016917
rect 246400 1016597 246600 1016600
rect 246146 1011607 246600 1016597
rect 246920 1011607 249880 1016597
rect 250200 1011607 250600 1016600
rect 250920 1011607 253880 1016597
rect 254200 1011607 254600 1016600
rect 254920 1011607 257880 1016597
rect 258200 1011607 258600 1016600
rect 258920 1011607 261880 1016597
rect 262200 1011607 262600 1016600
rect 262920 1011607 265880 1016597
rect 266200 1011607 266600 1016600
rect 266920 1011607 269880 1016597
rect 270200 1011607 270600 1016600
rect 270920 1011607 273880 1016597
rect 274200 1011607 274600 1016600
rect 274920 1011607 277880 1016597
rect 278200 1011607 278600 1016600
rect 278920 1011607 279880 1016597
rect 280200 1011607 280600 1016600
rect 281200 1016597 282000 1016600
rect 281200 1011607 282254 1016597
rect 246146 1010437 282254 1011287
rect 246146 1009267 282254 1010117
rect 246146 1007147 282254 1008947
rect 246146 1005937 282254 1006827
rect 246146 1004968 282254 1005617
rect 246400 1004967 282000 1004968
rect 246146 1003997 282254 1004647
rect 246146 1002787 282254 1003677
rect 246146 1001577 282254 1002467
rect 282574 1001257 297426 1016917
rect 298000 1016597 298200 1016600
rect 297746 1011607 298200 1016597
rect 298520 1011607 301480 1016597
rect 301800 1011607 302200 1016600
rect 302520 1011607 305480 1016597
rect 305800 1011607 306200 1016600
rect 306520 1011607 309480 1016597
rect 309800 1011607 310200 1016600
rect 310520 1011607 313480 1016597
rect 313800 1011607 314200 1016600
rect 314520 1011607 317480 1016597
rect 317800 1011607 318200 1016600
rect 318520 1011607 321480 1016597
rect 321800 1011607 322200 1016600
rect 322520 1011607 325480 1016597
rect 325800 1011607 326200 1016600
rect 326520 1011607 329480 1016597
rect 329800 1011607 330200 1016600
rect 330520 1011607 331480 1016597
rect 331800 1011607 332200 1016600
rect 332800 1016597 333400 1016600
rect 332800 1011607 333654 1016597
rect 297746 1010437 333654 1011287
rect 297746 1009267 333654 1010117
rect 297746 1007147 333654 1008947
rect 297746 1005937 333654 1006827
rect 297746 1004968 333654 1005617
rect 298000 1004967 333400 1004968
rect 297746 1003997 333654 1004647
rect 297746 1002787 333654 1003677
rect 297746 1001577 333654 1002467
rect 333974 1001257 347826 1016917
rect 348400 1016597 348600 1016600
rect 348146 1011607 348600 1016597
rect 348920 1011607 351880 1016597
rect 352200 1011607 352600 1016600
rect 352920 1011607 355880 1016597
rect 356200 1011607 356600 1016600
rect 356920 1011607 359880 1016597
rect 360200 1011607 360600 1016600
rect 360920 1011607 363880 1016597
rect 364200 1011607 364600 1016600
rect 364920 1011607 367880 1016597
rect 368200 1011607 368600 1016600
rect 368920 1011607 371880 1016597
rect 372200 1011607 372600 1016600
rect 372920 1011607 375880 1016597
rect 376200 1011607 376600 1016600
rect 376920 1011607 379880 1016597
rect 380200 1011607 380600 1016600
rect 380920 1011607 381880 1016597
rect 382200 1011607 382600 1016600
rect 383200 1016597 383800 1016600
rect 383200 1011607 384054 1016597
rect 348146 1010437 384054 1011287
rect 348146 1009267 384054 1010117
rect 348146 1007147 384054 1008947
rect 348146 1005937 384054 1006827
rect 348146 1004968 384054 1005617
rect 348400 1004967 383800 1004968
rect 348146 1003997 384054 1004647
rect 348146 1002787 384054 1003677
rect 348146 1001577 384054 1002467
rect 384374 1001257 399226 1016917
rect 399800 1016597 400000 1016600
rect 399546 1011607 400000 1016597
rect 400320 1011607 403280 1016597
rect 403600 1011607 404000 1016600
rect 404320 1011607 407280 1016597
rect 407600 1011607 408000 1016600
rect 408320 1011607 411280 1016597
rect 411600 1011607 412000 1016600
rect 412320 1011607 415280 1016597
rect 415600 1011607 416000 1016600
rect 416320 1011607 419280 1016597
rect 419600 1011607 420000 1016600
rect 420320 1011607 423280 1016597
rect 423600 1011607 424000 1016600
rect 424320 1011607 427280 1016597
rect 427600 1011607 428000 1016600
rect 428320 1011607 431280 1016597
rect 431600 1011607 432000 1016600
rect 432320 1011607 433280 1016597
rect 433600 1011607 434000 1016600
rect 434600 1011607 435400 1016600
rect 436000 1011607 436400 1016600
rect 437000 1011607 437400 1016600
rect 437720 1011607 440680 1016597
rect 441000 1011607 441400 1016600
rect 441720 1011607 444680 1016597
rect 445000 1011607 445400 1016600
rect 445720 1011607 448680 1016597
rect 449000 1011607 449400 1016600
rect 449720 1011607 452680 1016597
rect 453000 1011607 453400 1016600
rect 453720 1011607 456680 1016597
rect 457000 1011607 457400 1016600
rect 457720 1011607 460680 1016597
rect 461000 1011607 461400 1016600
rect 461720 1011607 464680 1016597
rect 465000 1011607 465400 1016600
rect 465720 1011607 468680 1016597
rect 469000 1011607 469400 1016600
rect 469720 1011607 470680 1016597
rect 471000 1011607 471400 1016600
rect 472000 1016597 472800 1016600
rect 472000 1011607 473054 1016597
rect 399546 1010437 473054 1011287
rect 399546 1009267 473054 1010117
rect 399546 1007147 435200 1008947
rect 436200 1007147 473054 1008947
rect 399546 1005937 436200 1006827
rect 437200 1005937 473054 1006827
rect 399546 1004968 435200 1005617
rect 399800 1004967 435200 1004968
rect 436200 1004968 473054 1005617
rect 436200 1004967 472800 1004968
rect 399546 1003997 473054 1004647
rect 399546 1002787 473054 1003677
rect 399546 1001577 473054 1002467
rect 473374 1001257 488226 1016917
rect 488800 1016597 489000 1016600
rect 488546 1011607 489000 1016597
rect 489320 1011607 492280 1016597
rect 492600 1011607 493000 1016600
rect 493320 1011607 496280 1016597
rect 496600 1011607 497000 1016600
rect 497320 1011607 500280 1016597
rect 500600 1011607 501000 1016600
rect 501320 1011607 504280 1016597
rect 504600 1011607 505000 1016600
rect 505320 1011607 508280 1016597
rect 508600 1011607 509000 1016600
rect 509320 1011607 512280 1016597
rect 512600 1011607 513000 1016600
rect 513320 1011607 516280 1016597
rect 516600 1011607 517000 1016600
rect 517320 1011607 520280 1016597
rect 520600 1011607 521000 1016600
rect 521320 1011607 522280 1016597
rect 522600 1011607 523000 1016600
rect 523600 1016597 524200 1016600
rect 523600 1011607 524454 1016597
rect 488546 1010437 524454 1011287
rect 488546 1009267 524454 1010117
rect 488546 1007147 524454 1008947
rect 488546 1005937 524454 1006827
rect 488546 1004968 524454 1005617
rect 488800 1004967 524200 1004968
rect 488546 1003997 524454 1004647
rect 488546 1002787 524454 1003677
rect 488546 1001577 524454 1002467
rect 524774 1001257 539626 1016917
rect 540200 1016597 540400 1016600
rect 539946 1011607 540400 1016597
rect 540720 1011607 543680 1016597
rect 544000 1011607 544400 1016600
rect 544720 1011607 547680 1016597
rect 548000 1011607 548400 1016600
rect 548720 1011607 551680 1016597
rect 552000 1011607 552400 1016600
rect 552720 1011607 555680 1016597
rect 556000 1011607 556400 1016600
rect 556720 1011607 559680 1016597
rect 560000 1011607 560400 1016600
rect 560720 1011607 563680 1016597
rect 564000 1011607 564400 1016600
rect 564720 1011607 567680 1016597
rect 568000 1011607 568400 1016600
rect 568720 1011607 571680 1016597
rect 572000 1011607 572400 1016600
rect 572720 1011607 573680 1016597
rect 574000 1011607 574400 1016600
rect 575000 1016597 575600 1016600
rect 575000 1011607 575854 1016597
rect 539946 1010437 575854 1011287
rect 539946 1009267 575854 1010117
rect 539946 1007147 575854 1008947
rect 539946 1005937 575854 1006827
rect 539946 1004968 575854 1005617
rect 540200 1004967 575600 1004968
rect 539946 1003997 575854 1004647
rect 539946 1002787 575854 1003677
rect 539946 1001577 575854 1002467
rect 576174 1001257 590026 1016917
rect 590600 1016597 590800 1016600
rect 590346 1011607 590800 1016597
rect 591120 1011607 594080 1016597
rect 594400 1011607 594800 1016600
rect 595120 1011607 598080 1016597
rect 598400 1011607 598800 1016600
rect 599120 1011607 602080 1016597
rect 602400 1011607 602800 1016600
rect 603120 1011607 606080 1016597
rect 606400 1011607 606800 1016600
rect 607120 1011607 610080 1016597
rect 610400 1011607 610800 1016600
rect 611120 1011607 614080 1016597
rect 614400 1011607 614800 1016600
rect 615120 1011607 618080 1016597
rect 618400 1011607 618800 1016600
rect 619120 1011607 622080 1016597
rect 622400 1011607 622800 1016600
rect 623120 1011607 624080 1016597
rect 624400 1011607 624800 1016600
rect 625400 1016597 626000 1016600
rect 625400 1011607 626254 1016597
rect 590346 1010437 626254 1011287
rect 590346 1009267 626254 1010117
rect 590346 1007147 626254 1008947
rect 590346 1005937 626254 1006827
rect 590346 1004968 626254 1005617
rect 590600 1004967 626000 1004968
rect 590346 1003997 626254 1004647
rect 590346 1002787 626254 1003677
rect 590346 1001577 626254 1002467
rect 626574 1001257 641426 1016917
rect 642000 1016597 642200 1016600
rect 641746 1011607 642200 1016597
rect 642520 1011607 645480 1016597
rect 645800 1011607 646200 1016600
rect 646520 1011607 649480 1016597
rect 649800 1011607 650200 1016600
rect 650520 1011607 653480 1016597
rect 653800 1011607 654200 1016600
rect 654520 1011607 657480 1016597
rect 657800 1011607 658200 1016600
rect 658520 1011607 661480 1016597
rect 661800 1011607 662200 1016600
rect 662520 1011607 665480 1016597
rect 665800 1011607 666200 1016600
rect 666520 1011607 669480 1016597
rect 669800 1011607 670200 1016600
rect 670520 1011607 673480 1016597
rect 673800 1011607 674200 1016600
rect 674520 1011607 675480 1016597
rect 675800 1011607 676200 1016600
rect 676800 1016597 677600 1016600
rect 676800 1011607 678129 1016597
rect 678449 1011287 717600 1016917
rect 641746 1010437 677896 1011287
rect 678216 1010437 717600 1011287
rect 641746 1009267 677925 1010117
rect 678245 1009267 717600 1010437
rect 641746 1007147 682231 1008947
rect 682551 1006827 717600 1009267
rect 641746 1005937 677895 1006827
rect 678215 1005617 717600 1006827
rect 641746 1004968 677867 1005617
rect 642000 1004967 677867 1004968
rect 678187 1004967 717600 1005617
rect 641746 1003997 677877 1004647
rect 678197 1003997 717600 1004967
rect 641746 1002787 677920 1003677
rect 678240 1002551 717600 1003997
rect 678240 1002467 686827 1002551
rect 641746 1001577 677905 1002467
rect 678225 1001257 686827 1002467
rect 30773 1000607 40229 1001257
rect 40549 1000607 76393 1001257
rect 76713 1000607 91674 1001257
rect 91994 1000607 127793 1001257
rect 128113 1000607 143074 1001257
rect 143394 1000607 179193 1001257
rect 179513 1000607 194474 1001257
rect 194794 1000607 230593 1001257
rect 230913 1000607 245874 1001257
rect 246194 1000607 282193 1001257
rect 282513 1000607 297474 1001257
rect 297794 1000607 333593 1001257
rect 333913 1000607 347887 1001257
rect 348207 1000607 383993 1001257
rect 384313 1000607 399274 1001257
rect 399594 1000607 435200 1001257
rect 436200 1000607 472993 1001257
rect 473313 1000607 488274 1001257
rect 488594 1000607 524393 1001257
rect 524713 1000607 539674 1001257
rect 539994 1000607 575793 1001257
rect 576113 1000607 590087 1001257
rect 590407 1000607 626193 1001257
rect 626513 1000607 641474 1001257
rect 641794 1000607 677894 1001257
rect 678214 1000607 686827 1001257
rect 30773 998677 40226 1000607
rect 40546 999397 76454 1000287
rect 30773 998240 36993 998677
rect 38523 998390 40226 998677
rect 30773 998215 33603 998240
rect 35133 998225 36993 998240
rect 31983 998197 33603 998215
rect 36343 998214 36993 998225
rect 31983 998187 32633 998197
rect 30773 969946 31663 997895
rect 31983 970200 32633 997867
rect 31983 969946 32632 970200
rect 32953 969946 33603 997877
rect 33923 969946 34813 997920
rect 35133 969946 36023 997905
rect 36343 969994 36993 997894
rect 37313 969946 38203 998357
rect 38523 969946 39573 998070
rect 39893 997707 40226 998390
rect 40546 998027 76454 999077
rect 76774 998027 91626 1000607
rect 91946 999397 127854 1000287
rect 91946 998027 127854 999077
rect 128174 998027 143026 1000607
rect 143346 999397 179254 1000287
rect 143346 998027 179254 999077
rect 179574 998027 194426 1000607
rect 194746 999397 230654 1000287
rect 194746 998027 230654 999077
rect 230974 998027 245826 1000607
rect 246146 999397 282254 1000287
rect 246146 998027 282254 999077
rect 282574 998027 297426 1000607
rect 297746 999397 333654 1000287
rect 297746 998027 333654 999077
rect 333974 998027 347826 1000607
rect 348146 999397 384054 1000287
rect 348146 998027 384054 999077
rect 384374 998027 399226 1000607
rect 399546 999397 436200 1000287
rect 437200 999397 473054 1000287
rect 399546 998027 473054 999077
rect 473374 998027 488226 1000607
rect 488546 999397 524454 1000287
rect 488546 998027 524454 999077
rect 524774 998027 539626 1000607
rect 539946 999397 575854 1000287
rect 539946 998027 575854 999077
rect 576174 998027 590026 1000607
rect 590346 999397 626254 1000287
rect 590346 998027 626254 999077
rect 626574 998027 641426 1000607
rect 641746 999397 678357 1000287
rect 678677 999077 686827 1000607
rect 641746 998027 678070 999077
rect 678390 997707 686827 999077
rect 39893 997600 40800 997707
rect 677600 997374 686827 997707
rect 677600 996800 677707 997374
rect 680607 997371 681257 997374
rect 36343 969626 36993 969674
rect 0 969280 39573 969626
rect 0 956120 6278 969280
rect 19408 956120 39573 969280
rect 678027 967346 679077 997054
rect 679397 967346 680287 997054
rect 680607 967407 681257 997051
rect 681577 967346 682467 997054
rect 682787 967346 683677 997054
rect 683997 967346 684647 997054
rect 684968 996800 685617 997054
rect 684967 967600 685617 996800
rect 684968 967346 685617 967600
rect 685937 967346 686827 997054
rect 687147 967346 688947 1002231
rect 689267 997491 717600 1002551
rect 689267 997374 691287 997491
rect 689267 967346 690117 997054
rect 690437 967346 691287 997054
rect 691607 996800 696597 997171
rect 696917 996800 717600 997491
rect 691607 996400 696600 996800
rect 691607 995400 696600 995800
rect 691607 992120 696597 995080
rect 691607 991400 696600 991800
rect 691607 988120 696597 991080
rect 691607 987400 696600 987800
rect 691607 984120 696597 987080
rect 691607 983400 696600 983800
rect 691607 980120 696597 983080
rect 691607 979400 696600 979800
rect 691607 976120 696597 979080
rect 691607 975400 696600 975800
rect 691607 972120 696597 975080
rect 691607 971400 696600 971800
rect 691607 968120 696597 971080
rect 691607 967600 696600 967800
rect 712757 967600 717600 996800
rect 691607 967346 696597 967600
rect 680607 967026 681257 967087
rect 696917 967026 717600 967600
rect 0 954774 39573 956120
rect 678027 965680 717600 967026
rect 0 954200 20683 954774
rect 36343 954713 36993 954774
rect 21003 954200 25993 954454
rect 0 927000 4843 954200
rect 21000 953800 25993 954200
rect 21000 952800 25993 953200
rect 21003 951520 25993 952480
rect 21000 950800 25993 951200
rect 21003 947520 25993 950480
rect 21000 946800 25993 947200
rect 21003 943520 25993 946480
rect 21000 942800 25993 943200
rect 21003 939520 25993 942480
rect 21000 938800 25993 939200
rect 21003 935520 25993 938480
rect 21000 934800 25993 935200
rect 21003 931520 25993 934480
rect 21000 930800 25993 931200
rect 21003 927520 25993 930480
rect 21000 927000 25993 927200
rect 0 926426 20683 927000
rect 21003 926746 25993 927000
rect 26313 926746 27163 954454
rect 27483 926746 28333 954454
rect 28653 926746 30453 954454
rect 30773 926746 31663 954454
rect 31983 954200 32632 954454
rect 31983 927000 32633 954200
rect 31983 926746 32632 927000
rect 32953 926746 33603 954454
rect 33923 926746 34813 954454
rect 35133 926746 36023 954454
rect 36343 926807 36993 954393
rect 37313 926746 38203 954454
rect 38523 926746 39573 954454
rect 678027 952520 698192 965680
rect 711322 952520 717600 965680
rect 678027 952174 717600 952520
rect 680607 952126 681257 952174
rect 36343 926426 36993 926487
rect 0 925511 39573 926426
rect 0 913543 5766 925511
rect 19892 913543 39573 925511
rect 678027 922346 679077 951854
rect 679397 922346 680287 951854
rect 680607 922407 681257 951806
rect 681577 922346 682467 951854
rect 682787 922346 683677 951854
rect 683997 922346 684647 951854
rect 684968 951600 685617 951854
rect 684967 922600 685617 951600
rect 684968 922346 685617 922600
rect 685937 922346 686827 951854
rect 687147 922346 688947 951854
rect 689267 922346 690117 951854
rect 690437 922346 691287 951854
rect 691607 951600 696597 951854
rect 696917 951600 717600 952174
rect 691607 951400 696600 951600
rect 691607 950400 696600 950800
rect 691607 947120 696597 950080
rect 691607 946400 696600 946800
rect 691607 943120 696597 946080
rect 691607 942400 696600 942800
rect 691607 939120 696597 942080
rect 691607 938400 696600 938800
rect 691607 935120 696597 938080
rect 691607 934400 696600 934800
rect 691607 931120 696597 934080
rect 691607 930400 696600 930800
rect 691607 927120 696597 930080
rect 691607 926400 696600 926800
rect 691607 923120 696597 926080
rect 691607 922600 696600 922800
rect 712757 922600 717600 951600
rect 691607 922346 696597 922600
rect 680607 922026 681257 922087
rect 696917 922026 717600 922600
rect 0 912574 39573 913543
rect 678027 921057 717600 922026
rect 0 912000 20683 912574
rect 36343 912513 36993 912574
rect 21003 912000 25993 912254
rect 0 884800 4843 912000
rect 21000 911600 25993 912000
rect 21000 910600 25993 911000
rect 21003 909320 25993 910280
rect 21000 908600 25993 909000
rect 21003 905320 25993 908280
rect 21000 904600 25993 905000
rect 21003 901320 25993 904280
rect 21000 900600 25993 901000
rect 21003 897320 25993 900280
rect 21000 896600 25993 897000
rect 21003 893320 25993 896280
rect 21000 892600 25993 893000
rect 21003 889320 25993 892280
rect 21000 888600 25993 889000
rect 21003 885320 25993 888280
rect 21000 884800 25993 885000
rect 0 884226 20683 884800
rect 21003 884546 25993 884800
rect 26313 884546 27163 912254
rect 27483 884546 28333 912254
rect 28653 884546 30453 912254
rect 30773 884546 31663 912254
rect 31983 912000 32632 912254
rect 31983 884800 32633 912000
rect 31983 884546 32632 884800
rect 32953 884546 33603 912254
rect 33923 884546 34813 912254
rect 35133 884546 36023 912254
rect 36343 884607 36993 912193
rect 37313 884546 38203 912254
rect 38523 884546 39573 912254
rect 678027 909089 697708 921057
rect 711834 909089 717600 921057
rect 678027 908174 717600 909089
rect 680607 908113 681257 908174
rect 36343 884226 36993 884287
rect 0 883880 39573 884226
rect 0 870700 6355 883880
rect 6675 871020 19198 883560
rect 19518 870700 39573 883880
rect 678027 878146 679077 907854
rect 679397 878146 680287 907854
rect 680607 878207 681257 907793
rect 681577 878146 682467 907854
rect 682787 878146 683677 907854
rect 683997 878146 684647 907854
rect 684968 907600 685617 907854
rect 684967 878400 685617 907600
rect 684968 878146 685617 878400
rect 685937 878146 686827 907854
rect 687147 878146 688947 907854
rect 689267 878146 690117 907854
rect 690437 878146 691287 907854
rect 691607 907600 696597 907854
rect 696917 907600 717600 908174
rect 691607 907200 696600 907600
rect 691607 906200 696600 906600
rect 691607 902920 696597 905880
rect 691607 902200 696600 902600
rect 691607 898920 696597 901880
rect 691607 898200 696600 898600
rect 691607 894920 696597 897880
rect 691607 894200 696600 894600
rect 691607 890920 696597 893880
rect 691607 890200 696600 890600
rect 691607 886920 696597 889880
rect 691607 886200 696600 886600
rect 691607 882920 696597 885880
rect 691607 882200 696600 882600
rect 691607 878920 696597 881880
rect 691607 878400 696600 878600
rect 712757 878400 717600 907600
rect 691607 878146 696597 878400
rect 680607 877826 681257 877887
rect 696917 877826 717600 878400
rect 0 870374 39573 870700
rect 678027 876480 717600 877826
rect 0 869800 20683 870374
rect 36343 870313 36993 870374
rect 21003 869800 25993 870054
rect 0 842600 4843 869800
rect 21000 869400 25993 869800
rect 21000 868400 25993 868800
rect 21003 867120 25993 868080
rect 21000 866400 25993 866800
rect 21003 863120 25993 866080
rect 21000 862400 25993 862800
rect 21003 859120 25993 862080
rect 21000 858400 25993 858800
rect 21003 855120 25993 858080
rect 21000 854400 25993 854800
rect 21003 851120 25993 854080
rect 21000 850400 25993 850800
rect 21003 847120 25993 850080
rect 21000 846400 25993 846800
rect 21003 843120 25993 846080
rect 21000 842600 25993 842800
rect 0 842026 20683 842600
rect 21003 842346 25993 842600
rect 26313 842346 27163 870054
rect 27483 842346 28333 870054
rect 28653 842346 30453 870054
rect 30773 842346 31663 870054
rect 31983 869800 32632 870054
rect 31983 842600 32633 869800
rect 31983 842346 32632 842600
rect 32953 842346 33603 870054
rect 33923 842346 34813 870054
rect 35133 842346 36023 870054
rect 36343 842407 36993 869993
rect 37313 842346 38203 870054
rect 38523 842346 39573 870054
rect 678027 863320 698192 876480
rect 711322 863320 717600 876480
rect 678027 862974 717600 863320
rect 680607 862926 681257 862974
rect 36343 842026 36993 842087
rect 0 841680 39573 842026
rect 0 828500 6355 841680
rect 19518 828500 39573 841680
rect 678027 833146 679077 862654
rect 679397 833146 680287 862654
rect 680607 833207 681257 862606
rect 681577 833146 682467 862654
rect 682787 833146 683677 862654
rect 683997 833146 684647 862654
rect 684968 862400 685617 862654
rect 684967 833400 685617 862400
rect 684968 833146 685617 833400
rect 685937 833146 686827 862654
rect 687147 833146 688947 862654
rect 689267 833146 690117 862654
rect 690437 833146 691287 862654
rect 691607 862400 696597 862654
rect 696917 862400 717600 862974
rect 691607 862200 696600 862400
rect 691607 861200 696600 861600
rect 691607 857920 696597 860880
rect 691607 857200 696600 857600
rect 691607 853920 696597 856880
rect 691607 853200 696600 853600
rect 691607 849920 696597 852880
rect 691607 849200 696600 849600
rect 691607 845920 696597 848880
rect 691607 845200 696600 845600
rect 691607 841920 696597 844880
rect 691607 841200 696600 841600
rect 691607 837920 696597 840880
rect 691607 837200 696600 837600
rect 691607 833920 696597 836880
rect 691607 833400 696600 833600
rect 712757 833400 717600 862400
rect 691607 833146 696597 833400
rect 680607 832826 681257 832887
rect 696917 832826 717600 833400
rect 0 828174 39573 828500
rect 678027 832500 717600 832826
rect 0 827600 20683 828174
rect 36343 828113 36993 828174
rect 21003 827600 25993 827854
rect 0 800400 4843 827600
rect 21000 827200 25993 827600
rect 21000 826200 25993 826600
rect 21003 824920 25993 825880
rect 21000 824200 25993 824600
rect 21003 820920 25993 823880
rect 21000 820200 25993 820600
rect 21003 816920 25993 819880
rect 21000 816200 25993 816600
rect 21003 812920 25993 815880
rect 21000 812200 25993 812600
rect 21003 808920 25993 811880
rect 21000 808200 25993 808600
rect 21003 804920 25993 807880
rect 21000 804200 25993 804600
rect 21003 800920 25993 803880
rect 21000 800400 25993 800600
rect 0 799826 20683 800400
rect 21003 800146 25993 800400
rect 26313 800146 27163 827854
rect 27483 800146 28333 827854
rect 28653 800146 30453 827854
rect 30773 800146 31663 827854
rect 31983 827600 32632 827854
rect 31983 800400 32633 827600
rect 31983 800146 32632 800400
rect 32953 800146 33603 827854
rect 33923 800146 34813 827854
rect 35133 800146 36023 827854
rect 36343 800194 36993 827793
rect 37313 800146 38203 827854
rect 38523 800146 39573 827854
rect 678027 819320 698082 832500
rect 711245 819320 717600 832500
rect 678027 818974 717600 819320
rect 680607 818913 681257 818974
rect 36343 799826 36993 799874
rect 0 799480 39573 799826
rect 0 786320 6278 799480
rect 19408 786320 39573 799480
rect 678027 788946 679077 818654
rect 679397 788946 680287 818654
rect 680607 789007 681257 818593
rect 681577 788946 682467 818654
rect 682787 788946 683677 818654
rect 683997 788946 684647 818654
rect 684968 818400 685617 818654
rect 684967 789200 685617 818400
rect 684968 788946 685617 789200
rect 685937 788946 686827 818654
rect 687147 788946 688947 818654
rect 689267 788946 690117 818654
rect 690437 788946 691287 818654
rect 691607 818400 696597 818654
rect 696917 818400 717600 818974
rect 691607 818000 696600 818400
rect 691607 817000 696600 817400
rect 691607 813720 696597 816680
rect 691607 813000 696600 813400
rect 691607 809720 696597 812680
rect 691607 809000 696600 809400
rect 691607 805720 696597 808680
rect 691607 805000 696600 805400
rect 691607 801720 696597 804680
rect 691607 801000 696600 801400
rect 691607 797720 696597 800680
rect 691607 797000 696600 797400
rect 691607 793720 696597 796680
rect 691607 793000 696600 793400
rect 691607 789720 696597 792680
rect 691607 789200 696600 789400
rect 712757 789200 717600 818400
rect 691607 788946 696597 789200
rect 680607 788626 681257 788687
rect 696917 788626 717600 789200
rect 0 784974 39573 786320
rect 678027 787280 717600 788626
rect 0 784400 20683 784974
rect 36343 784913 36993 784974
rect 21003 784400 25993 784654
rect 0 757200 4843 784400
rect 21000 784000 25993 784400
rect 21000 783000 25993 783400
rect 21003 781720 25993 782680
rect 21000 781000 25993 781400
rect 21003 777720 25993 780680
rect 21000 777000 25993 777400
rect 21003 773720 25993 776680
rect 21000 773000 25993 773400
rect 21003 769720 25993 772680
rect 21000 769000 25993 769400
rect 21003 765720 25993 768680
rect 21000 765000 25993 765400
rect 21003 761720 25993 764680
rect 21000 761000 25993 761400
rect 21003 757720 25993 760680
rect 21000 757200 25993 757400
rect 0 756626 20683 757200
rect 21003 756946 25993 757200
rect 26313 756946 27163 784654
rect 27483 756946 28333 784654
rect 28653 756946 30453 784654
rect 30773 756946 31663 784654
rect 31983 784400 32632 784654
rect 31983 757200 32633 784400
rect 31983 756946 32632 757200
rect 32953 756946 33603 784654
rect 33923 756946 34813 784654
rect 35133 756946 36023 784654
rect 36343 756994 36993 784593
rect 37313 756946 38203 784654
rect 38523 756946 39573 784654
rect 678027 774120 698192 787280
rect 711322 774120 717600 787280
rect 678027 773774 717600 774120
rect 680607 773726 681257 773774
rect 36343 756626 36993 756674
rect 0 756280 39573 756626
rect 0 743120 6278 756280
rect 19408 743120 39573 756280
rect 678027 743946 679077 773454
rect 679397 743946 680287 773454
rect 680607 744007 681257 773406
rect 681577 743946 682467 773454
rect 682787 743946 683677 773454
rect 683997 743946 684647 773454
rect 684968 773200 685617 773454
rect 684967 744200 685617 773200
rect 684968 743946 685617 744200
rect 685937 743946 686827 773454
rect 687147 743946 688947 773454
rect 689267 743946 690117 773454
rect 690437 743946 691287 773454
rect 691607 773200 696597 773454
rect 696917 773200 717600 773774
rect 691607 773000 696600 773200
rect 691607 772000 696600 772400
rect 691607 768720 696597 771680
rect 691607 768000 696600 768400
rect 691607 764720 696597 767680
rect 691607 764000 696600 764400
rect 691607 760720 696597 763680
rect 691607 760000 696600 760400
rect 691607 756720 696597 759680
rect 691607 756000 696600 756400
rect 691607 752720 696597 755680
rect 691607 752000 696600 752400
rect 691607 748720 696597 751680
rect 691607 748000 696600 748400
rect 691607 744720 696597 747680
rect 691607 744200 696600 744400
rect 712757 744200 717600 773200
rect 691607 743946 696597 744200
rect 680607 743626 681257 743687
rect 696917 743626 717600 744200
rect 0 741774 39573 743120
rect 678027 742280 717600 743626
rect 0 741200 20683 741774
rect 36343 741713 36993 741774
rect 21003 741200 25993 741454
rect 0 714000 4843 741200
rect 21000 740800 25993 741200
rect 21000 739800 25993 740200
rect 21003 738520 25993 739480
rect 21000 737800 25993 738200
rect 21003 734520 25993 737480
rect 21000 733800 25993 734200
rect 21003 730520 25993 733480
rect 21000 729800 25993 730200
rect 21003 726520 25993 729480
rect 21000 725800 25993 726200
rect 21003 722520 25993 725480
rect 21000 721800 25993 722200
rect 21003 718520 25993 721480
rect 21000 717800 25993 718200
rect 21003 714520 25993 717480
rect 21000 714000 25993 714200
rect 0 713426 20683 714000
rect 21003 713746 25993 714000
rect 26313 713746 27163 741454
rect 27483 713746 28333 741454
rect 28653 713746 30453 741454
rect 30773 713746 31663 741454
rect 31983 741200 32632 741454
rect 31983 714000 32633 741200
rect 31983 713746 32632 714000
rect 32953 713746 33603 741454
rect 33923 713746 34813 741454
rect 35133 713746 36023 741454
rect 36343 713794 36993 741393
rect 37313 713746 38203 741454
rect 38523 713746 39573 741454
rect 678027 729120 698192 742280
rect 711322 729120 717600 742280
rect 678027 728774 717600 729120
rect 680607 728726 681257 728774
rect 36343 713426 36993 713474
rect 0 713080 39573 713426
rect 0 699920 6278 713080
rect 19408 699920 39573 713080
rect 0 698574 39573 699920
rect 678027 698946 679077 728454
rect 679397 698946 680287 728454
rect 680607 699007 681257 728406
rect 681577 698946 682467 728454
rect 682787 698946 683677 728454
rect 683997 698946 684647 728454
rect 684968 728200 685617 728454
rect 684967 699200 685617 728200
rect 684968 698946 685617 699200
rect 685937 698946 686827 728454
rect 687147 698946 688947 728454
rect 689267 698946 690117 728454
rect 690437 698946 691287 728454
rect 691607 728200 696597 728454
rect 696917 728200 717600 728774
rect 691607 728000 696600 728200
rect 691607 727000 696600 727400
rect 691607 723720 696597 726680
rect 691607 723000 696600 723400
rect 691607 719720 696597 722680
rect 691607 719000 696600 719400
rect 691607 715720 696597 718680
rect 691607 715000 696600 715400
rect 691607 711720 696597 714680
rect 691607 711000 696600 711400
rect 691607 707720 696597 710680
rect 691607 707000 696600 707400
rect 691607 703720 696597 706680
rect 691607 703000 696600 703400
rect 691607 699720 696597 702680
rect 691607 699200 696600 699400
rect 712757 699200 717600 728200
rect 691607 698946 696597 699200
rect 680607 698626 681257 698687
rect 696917 698626 717600 699200
rect 0 698000 20683 698574
rect 36343 698513 36993 698574
rect 21003 698000 25993 698254
rect 0 670800 4843 698000
rect 21000 697600 25993 698000
rect 21000 696600 25993 697000
rect 21003 695320 25993 696280
rect 21000 694600 25993 695000
rect 21003 691320 25993 694280
rect 21000 690600 25993 691000
rect 21003 687320 25993 690280
rect 21000 686600 25993 687000
rect 21003 683320 25993 686280
rect 21000 682600 25993 683000
rect 21003 679320 25993 682280
rect 21000 678600 25993 679000
rect 21003 675320 25993 678280
rect 21000 674600 25993 675000
rect 21003 671320 25993 674280
rect 21000 670800 25993 671000
rect 0 670226 20683 670800
rect 21003 670546 25993 670800
rect 26313 670546 27163 698254
rect 27483 670546 28333 698254
rect 28653 670546 30453 698254
rect 30773 670546 31663 698254
rect 31983 698000 32632 698254
rect 31983 670800 32633 698000
rect 31983 670546 32632 670800
rect 32953 670546 33603 698254
rect 33923 670546 34813 698254
rect 35133 670546 36023 698254
rect 36343 670594 36993 698193
rect 37313 670546 38203 698254
rect 38523 670546 39573 698254
rect 678027 697280 717600 698626
rect 678027 684120 698192 697280
rect 711322 684120 717600 697280
rect 678027 683774 717600 684120
rect 680607 683726 681257 683774
rect 36343 670226 36993 670274
rect 0 669880 39573 670226
rect 0 656720 6278 669880
rect 19408 656720 39573 669880
rect 0 655374 39573 656720
rect 0 654800 20683 655374
rect 36343 655313 36993 655374
rect 21003 654800 25993 655054
rect 0 627600 4843 654800
rect 21000 654400 25993 654800
rect 21000 653400 25993 653800
rect 21003 652120 25993 653080
rect 21000 651400 25993 651800
rect 21003 648120 25993 651080
rect 21000 647400 25993 647800
rect 21003 644120 25993 647080
rect 21000 643400 25993 643800
rect 21003 640120 25993 643080
rect 21000 639400 25993 639800
rect 21003 636120 25993 639080
rect 21000 635400 25993 635800
rect 21003 632120 25993 635080
rect 21000 631400 25993 631800
rect 21003 628120 25993 631080
rect 21000 627600 25993 627800
rect 0 627026 20683 627600
rect 21003 627346 25993 627600
rect 26313 627346 27163 655054
rect 27483 627346 28333 655054
rect 28653 627346 30453 655054
rect 30773 627346 31663 655054
rect 31983 654800 32632 655054
rect 31983 627600 32633 654800
rect 31983 627346 32632 627600
rect 32953 627346 33603 655054
rect 33923 627346 34813 655054
rect 35133 627346 36023 655054
rect 36343 627394 36993 654993
rect 37313 627346 38203 655054
rect 38523 627346 39573 655054
rect 678027 653746 679077 683454
rect 679397 653746 680287 683454
rect 680607 653807 681257 683406
rect 681577 653746 682467 683454
rect 682787 653746 683677 683454
rect 683997 653746 684647 683454
rect 684968 683200 685617 683454
rect 684967 654000 685617 683200
rect 684968 653746 685617 654000
rect 685937 653746 686827 683454
rect 687147 653746 688947 683454
rect 689267 653746 690117 683454
rect 690437 653746 691287 683454
rect 691607 683200 696597 683454
rect 696917 683200 717600 683774
rect 691607 682800 696600 683200
rect 691607 681800 696600 682200
rect 691607 678520 696597 681480
rect 691607 677800 696600 678200
rect 691607 674520 696597 677480
rect 691607 673800 696600 674200
rect 691607 670520 696597 673480
rect 691607 669800 696600 670200
rect 691607 666520 696597 669480
rect 691607 665800 696600 666200
rect 691607 662520 696597 665480
rect 691607 661800 696600 662200
rect 691607 658520 696597 661480
rect 691607 657800 696600 658200
rect 691607 654520 696597 657480
rect 691607 654000 696600 654200
rect 712757 654000 717600 683200
rect 691607 653746 696597 654000
rect 680607 653426 681257 653487
rect 696917 653426 717600 654000
rect 678027 652080 717600 653426
rect 678027 638920 698192 652080
rect 711322 638920 717600 652080
rect 678027 638574 717600 638920
rect 680607 638526 681257 638574
rect 36343 627026 36993 627074
rect 0 626680 39573 627026
rect 0 613520 6278 626680
rect 19408 613520 39573 626680
rect 0 612174 39573 613520
rect 0 611600 20683 612174
rect 36343 612113 36993 612174
rect 21003 611600 25993 611854
rect 0 584400 4843 611600
rect 21000 611200 25993 611600
rect 21000 610200 25993 610600
rect 21003 608920 25993 609880
rect 21000 608200 25993 608600
rect 21003 604920 25993 607880
rect 21000 604200 25993 604600
rect 21003 600920 25993 603880
rect 21000 600200 25993 600600
rect 21003 596920 25993 599880
rect 21000 596200 25993 596600
rect 21003 592920 25993 595880
rect 21000 592200 25993 592600
rect 21003 588920 25993 591880
rect 21000 588200 25993 588600
rect 21003 584920 25993 587880
rect 21000 584400 25993 584600
rect 0 583826 20683 584400
rect 21003 584146 25993 584400
rect 26313 584146 27163 611854
rect 27483 584146 28333 611854
rect 28653 584146 30453 611854
rect 30773 584146 31663 611854
rect 31983 611600 32632 611854
rect 31983 584400 32633 611600
rect 31983 584146 32632 584400
rect 32953 584146 33603 611854
rect 33923 584146 34813 611854
rect 35133 584146 36023 611854
rect 36343 584194 36993 611793
rect 37313 584146 38203 611854
rect 38523 584146 39573 611854
rect 678027 608746 679077 638254
rect 679397 608746 680287 638254
rect 680607 608807 681257 638206
rect 681577 608746 682467 638254
rect 682787 608746 683677 638254
rect 683997 608746 684647 638254
rect 684968 638000 685617 638254
rect 684967 609000 685617 638000
rect 684968 608746 685617 609000
rect 685937 608746 686827 638254
rect 687147 608746 688947 638254
rect 689267 608746 690117 638254
rect 690437 608746 691287 638254
rect 691607 638000 696597 638254
rect 696917 638000 717600 638574
rect 691607 637800 696600 638000
rect 691607 636800 696600 637200
rect 691607 633520 696597 636480
rect 691607 632800 696600 633200
rect 691607 629520 696597 632480
rect 691607 628800 696600 629200
rect 691607 625520 696597 628480
rect 691607 624800 696600 625200
rect 691607 621520 696597 624480
rect 691607 620800 696600 621200
rect 691607 617520 696597 620480
rect 691607 616800 696600 617200
rect 691607 613520 696597 616480
rect 691607 612800 696600 613200
rect 691607 609520 696597 612480
rect 691607 609000 696600 609200
rect 712757 609000 717600 638000
rect 691607 608746 696597 609000
rect 680607 608426 681257 608487
rect 696917 608426 717600 609000
rect 678027 607080 717600 608426
rect 678027 593920 698192 607080
rect 711322 593920 717600 607080
rect 678027 593574 717600 593920
rect 680607 593526 681257 593574
rect 36343 583826 36993 583874
rect 0 583480 39573 583826
rect 0 570320 6278 583480
rect 19408 570320 39573 583480
rect 0 568974 39573 570320
rect 0 568400 20683 568974
rect 36343 568913 36993 568974
rect 21003 568400 25993 568654
rect 0 541200 4843 568400
rect 21000 568000 25993 568400
rect 21000 567000 25993 567400
rect 21003 565720 25993 566680
rect 21000 565000 25993 565400
rect 21003 561720 25993 564680
rect 21000 561000 25993 561400
rect 21003 557720 25993 560680
rect 21000 557000 25993 557400
rect 21003 553720 25993 556680
rect 21000 553000 25993 553400
rect 21003 549720 25993 552680
rect 21000 549000 25993 549400
rect 21003 545720 25993 548680
rect 21000 545000 25993 545400
rect 21003 541720 25993 544680
rect 21000 541200 25993 541400
rect 0 540626 20683 541200
rect 21003 540946 25993 541200
rect 26313 540946 27163 568654
rect 27483 540946 28333 568654
rect 28653 540946 30453 568654
rect 30773 540946 31663 568654
rect 31983 568400 32632 568654
rect 31983 541200 32633 568400
rect 31983 540946 32632 541200
rect 32953 540946 33603 568654
rect 33923 540946 34813 568654
rect 35133 540946 36023 568654
rect 36343 540994 36993 568593
rect 37313 540946 38203 568654
rect 38523 540946 39573 568654
rect 678027 563546 679077 593254
rect 679397 563546 680287 593254
rect 680607 563607 681257 593206
rect 681577 563546 682467 593254
rect 682787 563546 683677 593254
rect 683997 563546 684647 593254
rect 684968 593000 685617 593254
rect 684967 563800 685617 593000
rect 684968 563546 685617 563800
rect 685937 563546 686827 593254
rect 687147 563546 688947 593254
rect 689267 563546 690117 593254
rect 690437 563546 691287 593254
rect 691607 593000 696597 593254
rect 696917 593000 717600 593574
rect 691607 592600 696600 593000
rect 691607 591600 696600 592000
rect 691607 588320 696597 591280
rect 691607 587600 696600 588000
rect 691607 584320 696597 587280
rect 691607 583600 696600 584000
rect 691607 580320 696597 583280
rect 691607 579600 696600 580000
rect 691607 576320 696597 579280
rect 691607 575600 696600 576000
rect 691607 572320 696597 575280
rect 691607 571600 696600 572000
rect 691607 568320 696597 571280
rect 691607 567600 696600 568000
rect 691607 564320 696597 567280
rect 691607 563800 696600 564000
rect 712757 563800 717600 593000
rect 691607 563546 696597 563800
rect 680607 563226 681257 563287
rect 696917 563226 717600 563800
rect 678027 561880 717600 563226
rect 678027 548720 698192 561880
rect 711322 548720 717600 561880
rect 678027 548374 717600 548720
rect 680607 548326 681257 548374
rect 36343 540626 36993 540674
rect 0 540280 39573 540626
rect 0 527120 6278 540280
rect 19408 527120 39573 540280
rect 0 525774 39573 527120
rect 0 525200 20683 525774
rect 36343 525713 36993 525774
rect 21003 525200 25993 525454
rect 0 498000 4843 525200
rect 21000 524800 25993 525200
rect 21000 523800 25993 524200
rect 21003 522520 25993 523480
rect 21000 521800 25993 522200
rect 21003 518520 25993 521480
rect 21000 517800 25993 518200
rect 21003 514520 25993 517480
rect 21000 513800 25993 514200
rect 21003 510520 25993 513480
rect 21000 509800 25993 510200
rect 21003 506520 25993 509480
rect 21000 505800 25993 506200
rect 21003 502520 25993 505480
rect 21000 501800 25993 502200
rect 21003 498520 25993 501480
rect 21000 498000 25993 498200
rect 0 497426 20683 498000
rect 21003 497746 25993 498000
rect 26313 497746 27163 525454
rect 27483 497746 28333 525454
rect 28653 497746 30453 525454
rect 30773 497746 31663 525454
rect 31983 525200 32632 525454
rect 31983 498000 32633 525200
rect 31983 497746 32632 498000
rect 32953 497746 33603 525454
rect 33923 497746 34813 525454
rect 35133 497746 36023 525454
rect 36343 497807 36993 525393
rect 37313 497746 38203 525454
rect 38523 497746 39573 525454
rect 678027 518546 679077 548054
rect 679397 518546 680287 548054
rect 680607 518607 681257 548006
rect 681577 518546 682467 548054
rect 682787 518546 683677 548054
rect 683997 518546 684647 548054
rect 684968 547800 685617 548054
rect 684967 518800 685617 547800
rect 684968 518546 685617 518800
rect 685937 518546 686827 548054
rect 687147 518546 688947 548054
rect 689267 518546 690117 548054
rect 690437 518546 691287 548054
rect 691607 547800 696597 548054
rect 696917 547800 717600 548374
rect 691607 547600 696600 547800
rect 691607 546600 696600 547000
rect 691607 543320 696597 546280
rect 691607 542600 696600 543000
rect 691607 539320 696597 542280
rect 691607 538600 696600 539000
rect 691607 535320 696597 538280
rect 691607 534600 696600 535000
rect 691607 531320 696597 534280
rect 691607 530600 696600 531000
rect 691607 527320 696597 530280
rect 691607 526600 696600 527000
rect 691607 523320 696597 526280
rect 691607 522600 696600 523000
rect 691607 519320 696597 522280
rect 691607 518800 696600 519000
rect 712757 518800 717600 547800
rect 691607 518546 696597 518800
rect 680607 518226 681257 518287
rect 696917 518226 717600 518800
rect 678027 517900 717600 518226
rect 678027 504720 698082 517900
rect 698402 505040 710925 517580
rect 711245 504720 717600 517900
rect 678027 504374 717600 504720
rect 680607 504313 681257 504374
rect 36343 497426 36993 497487
rect 0 497080 39573 497426
rect 0 483900 6355 497080
rect 19518 483900 39573 497080
rect 0 483574 39573 483900
rect 0 483000 20683 483574
rect 36343 483513 36993 483574
rect 21003 483000 25993 483254
rect 0 455800 4843 483000
rect 21000 482600 25993 483000
rect 21000 481600 25993 482000
rect 21003 480320 25993 481280
rect 21000 479600 25993 480000
rect 21003 476320 25993 479280
rect 21000 475600 25993 476000
rect 21003 472320 25993 475280
rect 21000 471600 25993 472000
rect 21003 468320 25993 471280
rect 21000 467600 25993 468000
rect 21003 464320 25993 467280
rect 21000 463600 25993 464000
rect 21003 460320 25993 463280
rect 21000 459600 25993 460000
rect 21003 456320 25993 459280
rect 21000 455800 25993 456000
rect 0 455226 20683 455800
rect 21003 455546 25993 455800
rect 26313 455546 27163 483254
rect 27483 455546 28333 483254
rect 28653 455546 30453 483254
rect 30773 455546 31663 483254
rect 31983 483000 32632 483254
rect 31983 455800 32633 483000
rect 31983 455546 32632 455800
rect 32953 455546 33603 483254
rect 33923 455546 34813 483254
rect 35133 455546 36023 483254
rect 36343 455607 36993 483193
rect 37313 455546 38203 483254
rect 38523 455546 39573 483254
rect 678027 474546 679077 504054
rect 679397 474546 680287 504054
rect 680607 474607 681257 503993
rect 681577 474546 682467 504054
rect 682787 474546 683677 504054
rect 683997 474546 684647 504054
rect 684968 503800 685617 504054
rect 684967 474800 685617 503800
rect 684968 474546 685617 474800
rect 685937 474546 686827 504054
rect 687147 474546 688947 504054
rect 689267 474546 690117 504054
rect 690437 474546 691287 504054
rect 691607 503800 696597 504054
rect 696917 503800 717600 504374
rect 691607 503600 696600 503800
rect 691607 502600 696600 503000
rect 691607 499320 696597 502280
rect 691607 498600 696600 499000
rect 691607 495320 696597 498280
rect 691607 494600 696600 495000
rect 691607 491320 696597 494280
rect 691607 490600 696600 491000
rect 691607 487320 696597 490280
rect 691607 486600 696600 487000
rect 691607 483320 696597 486280
rect 691607 482600 696600 483000
rect 691607 479320 696597 482280
rect 691607 478600 696600 479000
rect 691607 475320 696597 478280
rect 691607 474800 696600 475000
rect 712757 474800 717600 503800
rect 691607 474546 696597 474800
rect 680607 474226 681257 474287
rect 696917 474226 717600 474800
rect 678027 473257 717600 474226
rect 678027 461289 697708 473257
rect 711834 461289 717600 473257
rect 678027 460374 717600 461289
rect 680607 460313 681257 460374
rect 36343 455226 36993 455287
rect 0 454311 39573 455226
rect 0 442343 5766 454311
rect 19892 442343 39573 454311
rect 0 441374 39573 442343
rect 0 440800 20683 441374
rect 36343 441313 36993 441374
rect 21003 440800 25993 441054
rect 0 413600 4843 440800
rect 21000 440400 25993 440800
rect 21000 439400 25993 439800
rect 21003 438120 25993 439080
rect 21000 437400 25993 437800
rect 21003 434120 25993 437080
rect 21000 433400 25993 433800
rect 21003 430120 25993 433080
rect 21000 429400 25993 429800
rect 21003 426120 25993 429080
rect 21000 425400 25993 425800
rect 21003 422120 25993 425080
rect 21000 421400 25993 421800
rect 21003 418120 25993 421080
rect 21000 417400 25993 417800
rect 21003 414120 25993 417080
rect 21000 413600 25993 413800
rect 0 413026 20683 413600
rect 21003 413346 25993 413600
rect 26313 413346 27163 441054
rect 27483 413346 28333 441054
rect 28653 413346 30453 441054
rect 30773 413346 31663 441054
rect 31983 440800 32632 441054
rect 31983 413600 32633 440800
rect 31983 413346 32632 413600
rect 32953 413346 33603 441054
rect 33923 413346 34813 441054
rect 35133 413346 36023 441054
rect 36343 413394 36993 440993
rect 37313 413346 38203 441054
rect 38523 413346 39573 441054
rect 678027 430346 679077 460054
rect 679397 430346 680287 460054
rect 680607 430407 681257 459993
rect 681577 430346 682467 460054
rect 682787 430346 683677 460054
rect 683997 430346 684647 460054
rect 684968 459800 685617 460054
rect 684967 430600 685617 459800
rect 684968 430346 685617 430600
rect 685937 430346 686827 460054
rect 687147 430346 688947 460054
rect 689267 430346 690117 460054
rect 690437 430346 691287 460054
rect 691607 459800 696597 460054
rect 696917 459800 717600 460374
rect 691607 459400 696600 459800
rect 691607 458400 696600 458800
rect 691607 455120 696597 458080
rect 691607 454400 696600 454800
rect 691607 451120 696597 454080
rect 691607 450400 696600 450800
rect 691607 447120 696597 450080
rect 691607 446400 696600 446800
rect 691607 443120 696597 446080
rect 691607 442400 696600 442800
rect 691607 439120 696597 442080
rect 691607 438400 696600 438800
rect 691607 435120 696597 438080
rect 691607 434400 696600 434800
rect 691607 431120 696597 434080
rect 691607 430600 696600 430800
rect 712757 430600 717600 459800
rect 691607 430346 696597 430600
rect 680607 430026 681257 430087
rect 696917 430026 717600 430600
rect 678027 429700 717600 430026
rect 678027 416520 698082 429700
rect 698402 416840 710925 429380
rect 711245 416520 717600 429700
rect 678027 416174 717600 416520
rect 680607 416113 681257 416174
rect 36343 413026 36993 413074
rect 0 412680 39573 413026
rect 0 399520 6278 412680
rect 19408 399520 39573 412680
rect 0 398174 39573 399520
rect 0 397600 20683 398174
rect 36343 398113 36993 398174
rect 21003 397600 25993 397854
rect 0 370400 4843 397600
rect 21000 397200 25993 397600
rect 21000 396200 25993 396600
rect 21003 394920 25993 395880
rect 21000 394200 25993 394600
rect 21003 390920 25993 393880
rect 21000 390200 25993 390600
rect 21003 386920 25993 389880
rect 21000 386200 25993 386600
rect 21003 382920 25993 385880
rect 21000 382200 25993 382600
rect 21003 378920 25993 381880
rect 21000 378200 25993 378600
rect 21003 374920 25993 377880
rect 21000 374200 25993 374600
rect 21003 370920 25993 373880
rect 21000 370400 25993 370600
rect 0 369826 20683 370400
rect 21003 370146 25993 370400
rect 26313 370146 27163 397854
rect 27483 370146 28333 397854
rect 28653 370146 30453 397854
rect 30773 370146 31663 397854
rect 31983 397600 32632 397854
rect 31983 370400 32633 397600
rect 31983 370146 32632 370400
rect 32953 370146 33603 397854
rect 33923 370146 34813 397854
rect 35133 370146 36023 397854
rect 36343 370194 36993 397793
rect 37313 370146 38203 397854
rect 38523 370146 39573 397854
rect 678027 386346 679077 415854
rect 679397 386346 680287 415854
rect 680607 386407 681257 415793
rect 681577 386346 682467 415854
rect 682787 386346 683677 415854
rect 683997 386346 684647 415854
rect 684968 415600 685617 415854
rect 684967 386600 685617 415600
rect 684968 386346 685617 386600
rect 685937 386346 686827 415854
rect 687147 386346 688947 415854
rect 689267 386346 690117 415854
rect 690437 386346 691287 415854
rect 691607 415600 696597 415854
rect 696917 415600 717600 416174
rect 691607 415400 696600 415600
rect 691607 414400 696600 414800
rect 691607 411120 696597 414080
rect 691607 410400 696600 410800
rect 691607 407120 696597 410080
rect 691607 406400 696600 406800
rect 691607 403120 696597 406080
rect 691607 402400 696600 402800
rect 691607 399120 696597 402080
rect 691607 398400 696600 398800
rect 691607 395120 696597 398080
rect 691607 394400 696600 394800
rect 691607 391120 696597 394080
rect 691607 390400 696600 390800
rect 691607 387120 696597 390080
rect 691607 386600 696600 386800
rect 712757 386600 717600 415600
rect 691607 386346 696597 386600
rect 680607 386026 681257 386087
rect 696917 386026 717600 386600
rect 678027 384680 717600 386026
rect 678027 371520 698192 384680
rect 711322 371520 717600 384680
rect 678027 371174 717600 371520
rect 680607 371126 681257 371174
rect 36343 369826 36993 369874
rect 0 369480 39573 369826
rect 0 356320 6278 369480
rect 19408 356320 39573 369480
rect 0 354974 39573 356320
rect 0 354400 20683 354974
rect 36343 354913 36993 354974
rect 21003 354400 25993 354654
rect 0 327200 4843 354400
rect 21000 354000 25993 354400
rect 21000 353000 25993 353400
rect 21003 351720 25993 352680
rect 21000 351000 25993 351400
rect 21003 347720 25993 350680
rect 21000 347000 25993 347400
rect 21003 343720 25993 346680
rect 21000 343000 25993 343400
rect 21003 339720 25993 342680
rect 21000 339000 25993 339400
rect 21003 335720 25993 338680
rect 21000 335000 25993 335400
rect 21003 331720 25993 334680
rect 21000 331000 25993 331400
rect 21003 327720 25993 330680
rect 21000 327200 25993 327400
rect 0 326626 20683 327200
rect 21003 326946 25993 327200
rect 26313 326946 27163 354654
rect 27483 326946 28333 354654
rect 28653 326946 30453 354654
rect 30773 326946 31663 354654
rect 31983 354400 32632 354654
rect 31983 327200 32633 354400
rect 31983 326946 32632 327200
rect 32953 326946 33603 354654
rect 33923 326946 34813 354654
rect 35133 326946 36023 354654
rect 36343 326994 36993 354593
rect 37313 326946 38203 354654
rect 38523 326946 39573 354654
rect 678027 341146 679077 370854
rect 679397 341146 680287 370854
rect 680607 341207 681257 370806
rect 681577 341146 682467 370854
rect 682787 341146 683677 370854
rect 683997 341146 684647 370854
rect 684968 370600 685617 370854
rect 684967 341400 685617 370600
rect 684968 341146 685617 341400
rect 685937 341146 686827 370854
rect 687147 341146 688947 370854
rect 689267 341146 690117 370854
rect 690437 341146 691287 370854
rect 691607 370600 696597 370854
rect 696917 370600 717600 371174
rect 691607 370200 696600 370600
rect 691607 369200 696600 369600
rect 691607 365920 696597 368880
rect 691607 365200 696600 365600
rect 691607 361920 696597 364880
rect 691607 361200 696600 361600
rect 691607 357920 696597 360880
rect 691607 357200 696600 357600
rect 691607 353920 696597 356880
rect 691607 353200 696600 353600
rect 691607 349920 696597 352880
rect 691607 349200 696600 349600
rect 691607 345920 696597 348880
rect 691607 345200 696600 345600
rect 691607 341920 696597 344880
rect 691607 341400 696600 341600
rect 712757 341400 717600 370600
rect 691607 341146 696597 341400
rect 680607 340826 681257 340887
rect 696917 340826 717600 341400
rect 678027 339480 717600 340826
rect 36343 326626 36993 326674
rect 0 326280 39573 326626
rect 0 313120 6278 326280
rect 19408 313120 39573 326280
rect 678027 326320 698192 339480
rect 711322 326320 717600 339480
rect 678027 325974 717600 326320
rect 680607 325926 681257 325974
rect 0 311774 39573 313120
rect 0 311200 20683 311774
rect 36343 311713 36993 311774
rect 21003 311200 25993 311454
rect 0 284000 4843 311200
rect 21000 310800 25993 311200
rect 21000 309800 25993 310200
rect 21003 308520 25993 309480
rect 21000 307800 25993 308200
rect 21003 304520 25993 307480
rect 21000 303800 25993 304200
rect 21003 300520 25993 303480
rect 21000 299800 25993 300200
rect 21003 296520 25993 299480
rect 21000 295800 25993 296200
rect 21003 292520 25993 295480
rect 21000 291800 25993 292200
rect 21003 288520 25993 291480
rect 21000 287800 25993 288200
rect 21003 284520 25993 287480
rect 21000 284000 25993 284200
rect 0 283426 20683 284000
rect 21003 283746 25993 284000
rect 26313 283746 27163 311454
rect 27483 283746 28333 311454
rect 28653 283746 30453 311454
rect 30773 283746 31663 311454
rect 31983 311200 32632 311454
rect 31983 284000 32633 311200
rect 31983 283746 32632 284000
rect 32953 283746 33603 311454
rect 33923 283746 34813 311454
rect 35133 283746 36023 311454
rect 36343 283794 36993 311393
rect 37313 283746 38203 311454
rect 38523 283746 39573 311454
rect 678027 296146 679077 325654
rect 679397 296146 680287 325654
rect 680607 296207 681257 325606
rect 681577 296146 682467 325654
rect 682787 296146 683677 325654
rect 683997 296146 684647 325654
rect 684968 325400 685617 325654
rect 684967 296400 685617 325400
rect 684968 296146 685617 296400
rect 685937 296146 686827 325654
rect 687147 296146 688947 325654
rect 689267 296146 690117 325654
rect 690437 296146 691287 325654
rect 691607 325400 696597 325654
rect 696917 325400 717600 325974
rect 691607 325200 696600 325400
rect 691607 324200 696600 324600
rect 691607 320920 696597 323880
rect 691607 320200 696600 320600
rect 691607 316920 696597 319880
rect 691607 316200 696600 316600
rect 691607 312920 696597 315880
rect 691607 312200 696600 312600
rect 691607 308920 696597 311880
rect 691607 308200 696600 308600
rect 691607 304920 696597 307880
rect 691607 304200 696600 304600
rect 691607 300920 696597 303880
rect 691607 300200 696600 300600
rect 691607 296920 696597 299880
rect 691607 296400 696600 296600
rect 712757 296400 717600 325400
rect 691607 296146 696597 296400
rect 680607 295826 681257 295887
rect 696917 295826 717600 296400
rect 678027 294480 717600 295826
rect 36343 283426 36993 283474
rect 0 283080 39573 283426
rect 0 269920 6278 283080
rect 19408 269920 39573 283080
rect 678027 281320 698192 294480
rect 711322 281320 717600 294480
rect 678027 280974 717600 281320
rect 680607 280926 681257 280974
rect 0 268574 39573 269920
rect 0 268000 20683 268574
rect 36343 268513 36993 268574
rect 21003 268000 25993 268254
rect 0 240800 4843 268000
rect 21000 267600 25993 268000
rect 21000 266600 25993 267000
rect 21003 265320 25993 266280
rect 21000 264600 25993 265000
rect 21003 261320 25993 264280
rect 21000 260600 25993 261000
rect 21003 257320 25993 260280
rect 21000 256600 25993 257000
rect 21003 253320 25993 256280
rect 21000 252600 25993 253000
rect 21003 249320 25993 252280
rect 21000 248600 25993 249000
rect 21003 245320 25993 248280
rect 21000 244600 25993 245000
rect 21003 241320 25993 244280
rect 21000 240800 25993 241000
rect 0 240226 20683 240800
rect 21003 240546 25993 240800
rect 26313 240546 27163 268254
rect 27483 240546 28333 268254
rect 28653 240546 30453 268254
rect 30773 240546 31663 268254
rect 31983 268000 32632 268254
rect 31983 240800 32633 268000
rect 31983 240546 32632 240800
rect 32953 240546 33603 268254
rect 33923 240546 34813 268254
rect 35133 240546 36023 268254
rect 36343 240594 36993 268193
rect 37313 240546 38203 268254
rect 38523 240546 39573 268254
rect 678027 251146 679077 280654
rect 679397 251146 680287 280654
rect 680607 251207 681257 280606
rect 681577 251146 682467 280654
rect 682787 251146 683677 280654
rect 683997 251146 684647 280654
rect 684968 280400 685617 280654
rect 684967 251400 685617 280400
rect 684968 251146 685617 251400
rect 685937 251146 686827 280654
rect 687147 251146 688947 280654
rect 689267 251146 690117 280654
rect 690437 251146 691287 280654
rect 691607 280400 696597 280654
rect 696917 280400 717600 280974
rect 691607 280200 696600 280400
rect 691607 279200 696600 279600
rect 691607 275920 696597 278880
rect 691607 275200 696600 275600
rect 691607 271920 696597 274880
rect 691607 271200 696600 271600
rect 691607 267920 696597 270880
rect 691607 267200 696600 267600
rect 691607 263920 696597 266880
rect 691607 263200 696600 263600
rect 691607 259920 696597 262880
rect 691607 259200 696600 259600
rect 691607 255920 696597 258880
rect 691607 255200 696600 255600
rect 691607 251920 696597 254880
rect 691607 251400 696600 251600
rect 712757 251400 717600 280400
rect 691607 251146 696597 251400
rect 680607 250826 681257 250887
rect 696917 250826 717600 251400
rect 678027 249480 717600 250826
rect 36343 240226 36993 240274
rect 0 239880 39573 240226
rect 0 226720 6278 239880
rect 19408 226720 39573 239880
rect 678027 236320 698192 249480
rect 711322 236320 717600 249480
rect 678027 235974 717600 236320
rect 680607 235926 681257 235974
rect 0 225374 39573 226720
rect 0 224800 20683 225374
rect 36343 225313 36993 225374
rect 21003 224800 25993 225054
rect 0 197600 4843 224800
rect 21000 224400 25993 224800
rect 21000 223400 25993 223800
rect 21003 222120 25993 223080
rect 21000 221400 25993 221800
rect 21003 218120 25993 221080
rect 21000 217400 25993 217800
rect 21003 214120 25993 217080
rect 21000 213400 25993 213800
rect 21003 210120 25993 213080
rect 21000 209400 25993 209800
rect 21003 206120 25993 209080
rect 21000 205400 25993 205800
rect 21003 202120 25993 205080
rect 21000 201400 25993 201800
rect 21003 198120 25993 201080
rect 21000 197600 25993 197800
rect 0 197026 20683 197600
rect 21003 197346 25993 197600
rect 26313 197346 27163 225054
rect 27483 197346 28333 225054
rect 28653 197346 30453 225054
rect 30773 197346 31663 225054
rect 31983 224800 32632 225054
rect 31983 197600 32633 224800
rect 31983 197346 32632 197600
rect 32953 197346 33603 225054
rect 33923 197346 34813 225054
rect 35133 197346 36023 225054
rect 36343 197394 36993 224993
rect 37313 197346 38203 225054
rect 38523 197346 39573 225054
rect 678027 205946 679077 235654
rect 679397 205946 680287 235654
rect 680607 206007 681257 235606
rect 681577 205946 682467 235654
rect 682787 205946 683677 235654
rect 683997 205946 684647 235654
rect 684968 235400 685617 235654
rect 684967 206200 685617 235400
rect 684968 205946 685617 206200
rect 685937 205946 686827 235654
rect 687147 205946 688947 235654
rect 689267 205946 690117 235654
rect 690437 205946 691287 235654
rect 691607 235400 696597 235654
rect 696917 235400 717600 235974
rect 691607 235000 696600 235400
rect 691607 234000 696600 234400
rect 691607 230720 696597 233680
rect 691607 230000 696600 230400
rect 691607 226720 696597 229680
rect 691607 226000 696600 226400
rect 691607 222720 696597 225680
rect 691607 222000 696600 222400
rect 691607 218720 696597 221680
rect 691607 218000 696600 218400
rect 691607 214720 696597 217680
rect 691607 214000 696600 214400
rect 691607 210720 696597 213680
rect 691607 210000 696600 210400
rect 691607 206720 696597 209680
rect 691607 206200 696600 206400
rect 712757 206200 717600 235400
rect 691607 205946 696597 206200
rect 680607 205626 681257 205687
rect 696917 205626 717600 206200
rect 678027 204280 717600 205626
rect 36343 197026 36993 197074
rect 0 196680 39573 197026
rect 0 183520 6278 196680
rect 19408 183520 39573 196680
rect 678027 191120 698192 204280
rect 711322 191120 717600 204280
rect 678027 190774 717600 191120
rect 680607 190726 681257 190774
rect 0 182174 39573 183520
rect 0 181600 20683 182174
rect 36343 182113 36993 182174
rect 21003 181600 25993 181854
rect 0 125200 4843 181600
rect 21000 181200 25993 181600
rect 21000 180200 25993 180600
rect 21003 178920 25993 179880
rect 21000 178200 25993 178600
rect 21003 174920 25993 177880
rect 21000 174200 25993 174600
rect 21003 170920 25993 173880
rect 21000 170200 25993 170600
rect 21003 166920 25993 169880
rect 21000 166200 25993 166600
rect 21003 162920 25993 165880
rect 21000 162200 25993 162600
rect 21003 158920 25993 161880
rect 21000 158200 25993 158600
rect 21003 154920 25993 157880
rect 21000 154200 25993 154600
rect 21000 153200 25993 153600
rect 21000 152000 25993 152600
rect 21000 151000 25993 151400
rect 21003 149720 25993 150680
rect 21000 149000 25993 149400
rect 21003 145720 25993 148680
rect 21000 145000 25993 145400
rect 21003 141720 25993 144680
rect 21000 141000 25993 141400
rect 21003 137720 25993 140680
rect 21000 137000 25993 137400
rect 21003 133720 25993 136680
rect 21000 133000 25993 133400
rect 21003 129720 25993 132680
rect 21000 129000 25993 129400
rect 21003 125720 25993 128680
rect 21000 125200 25993 125400
rect 0 124626 20683 125200
rect 21003 124946 25993 125200
rect 26313 124946 27163 181854
rect 27483 124946 28333 181854
rect 28653 153400 30453 181854
rect 30773 154400 31663 181854
rect 31983 181600 32632 181854
rect 31983 153400 32633 181600
rect 28653 124946 30453 152400
rect 30773 124946 31663 153400
rect 31983 125200 32633 152400
rect 31983 124946 32632 125200
rect 32953 124946 33603 181854
rect 33923 124946 34813 181854
rect 35133 124946 36023 181854
rect 36343 153400 36993 181793
rect 37313 154400 38203 181854
rect 36343 125007 36993 152400
rect 37313 124946 38203 153400
rect 38523 124946 39573 181854
rect 678027 160946 679077 190454
rect 679397 160946 680287 190454
rect 680607 161007 681257 190406
rect 681577 160946 682467 190454
rect 682787 160946 683677 190454
rect 683997 160946 684647 190454
rect 684968 190200 685617 190454
rect 684967 161200 685617 190200
rect 684968 160946 685617 161200
rect 685937 160946 686827 190454
rect 687147 160946 688947 190454
rect 689267 160946 690117 190454
rect 690437 160946 691287 190454
rect 691607 190200 696597 190454
rect 696917 190200 717600 190774
rect 691607 190000 696600 190200
rect 691607 189000 696600 189400
rect 691607 185720 696597 188680
rect 691607 185000 696600 185400
rect 691607 181720 696597 184680
rect 691607 181000 696600 181400
rect 691607 177720 696597 180680
rect 691607 177000 696600 177400
rect 691607 173720 696597 176680
rect 691607 173000 696600 173400
rect 691607 169720 696597 172680
rect 691607 169000 696600 169400
rect 691607 165720 696597 168680
rect 691607 165000 696600 165400
rect 691607 161720 696597 164680
rect 691607 161200 696600 161400
rect 712757 161200 717600 190200
rect 691607 160946 696597 161200
rect 680607 160626 681257 160687
rect 696917 160626 717600 161200
rect 678027 159280 717600 160626
rect 678027 146120 698192 159280
rect 711322 146120 717600 159280
rect 678027 145774 717600 146120
rect 680607 145726 681257 145774
rect 36343 124626 36993 124687
rect 0 124280 39573 124626
rect 0 111100 6355 124280
rect 19518 111100 39573 124280
rect 678027 115746 679077 145454
rect 679397 115746 680287 145454
rect 680607 115807 681257 145406
rect 681577 115746 682467 145454
rect 682787 115746 683677 145454
rect 683997 115746 684647 145454
rect 684968 145200 685617 145454
rect 684967 116000 685617 145200
rect 684968 115746 685617 116000
rect 685937 115746 686827 145454
rect 687147 115746 688947 145454
rect 689267 115746 690117 145454
rect 690437 115746 691287 145454
rect 691607 145200 696597 145454
rect 696917 145200 717600 145774
rect 691607 144800 696600 145200
rect 691607 143800 696600 144200
rect 691607 140520 696597 143480
rect 691607 139800 696600 140200
rect 691607 136520 696597 139480
rect 691607 135800 696600 136200
rect 691607 132520 696597 135480
rect 691607 131800 696600 132200
rect 691607 128520 696597 131480
rect 691607 127800 696600 128200
rect 691607 124520 696597 127480
rect 691607 123800 696600 124200
rect 691607 120520 696597 123480
rect 691607 119800 696600 120200
rect 691607 116520 696597 119480
rect 691607 116000 696600 116200
rect 712757 116000 717600 145200
rect 691607 115746 696597 116000
rect 680607 115426 681257 115487
rect 696917 115426 717600 116000
rect 0 110774 39573 111100
rect 678027 114080 717600 115426
rect 0 110200 20683 110774
rect 36343 110713 36993 110774
rect 21003 110200 25993 110454
rect 0 83000 4843 110200
rect 21000 109800 25993 110200
rect 21000 108800 25993 109200
rect 21003 107520 25993 108480
rect 21000 106800 25993 107200
rect 21003 103520 25993 106480
rect 21000 102800 25993 103200
rect 21003 99520 25993 102480
rect 21000 98800 25993 99200
rect 21003 95520 25993 98480
rect 21000 94800 25993 95200
rect 21003 91520 25993 94480
rect 21000 90800 25993 91200
rect 21003 87520 25993 90480
rect 21000 86800 25993 87200
rect 21003 83520 25993 86480
rect 21000 83000 25993 83200
rect 0 82426 20683 83000
rect 21003 82746 25993 83000
rect 26313 82746 27163 110454
rect 27483 82746 28333 110454
rect 28653 82746 30453 110454
rect 30773 82746 31663 110454
rect 31983 110200 32632 110454
rect 31983 83000 32633 110200
rect 31983 82746 32632 83000
rect 32953 82746 33603 110454
rect 33923 82746 34813 110454
rect 35133 82746 36023 110454
rect 36343 82807 36993 110393
rect 37313 82746 38203 110454
rect 38523 82746 39573 110454
rect 678027 100920 698192 114080
rect 711322 100920 717600 114080
rect 678027 100574 717600 100920
rect 680607 100526 681257 100574
rect 36343 82426 36993 82487
rect 0 81511 39573 82426
rect 0 69543 5766 81511
rect 19892 69543 39573 81511
rect 0 68574 39573 69543
rect 0 68000 20683 68574
rect 36343 68513 36993 68574
rect 21003 68000 25993 68254
rect 0 40800 4843 68000
rect 21000 67600 25993 68000
rect 21000 66600 25993 67000
rect 21003 65320 25993 66280
rect 21000 64600 25993 65000
rect 21003 61320 25993 64280
rect 21000 60600 25993 61000
rect 21003 57320 25993 60280
rect 21000 56600 25993 57000
rect 21003 53320 25993 56280
rect 21000 52600 25993 53000
rect 21003 49320 25993 52280
rect 21000 48600 25993 49000
rect 21003 45320 25993 48280
rect 21000 44600 25993 45000
rect 21003 41320 25993 44280
rect 21000 40800 25993 41000
rect 0 40109 20683 40800
rect 21003 40429 25993 40800
rect 26313 40546 27163 68254
rect 27483 40546 28333 68254
rect 26313 40109 28333 40226
rect 0 35049 28333 40109
rect 28653 35369 30453 68254
rect 30773 40546 31663 68254
rect 31983 68000 32632 68254
rect 31983 40800 32633 68000
rect 31983 40546 32632 40800
rect 32953 40546 33603 68254
rect 33923 40546 34813 68254
rect 35133 40546 36023 68254
rect 36343 40549 36993 68193
rect 37313 40546 38203 68254
rect 38523 40546 39573 68254
rect 36343 40226 36993 40229
rect 39893 40226 40000 40800
rect 30773 39893 40000 40226
rect 676800 39893 677707 40000
rect 30773 38523 39210 39893
rect 39530 38523 79054 39573
rect 30773 36993 38923 38523
rect 47400 38203 71400 38523
rect 39243 37313 79054 38203
rect 79374 36993 93226 39573
rect 93546 38523 132854 39573
rect 133174 38523 186654 39573
rect 101200 38203 125200 38523
rect 133174 38203 147600 38523
rect 155000 38203 179000 38523
rect 93546 37313 132854 38203
rect 133174 37313 186654 38203
rect 133174 36993 147600 37313
rect 186974 36993 201826 39573
rect 202146 38523 241454 39573
rect 209800 38203 233800 38523
rect 202146 37313 241454 38203
rect 241774 36993 255626 39573
rect 255946 38523 295254 39573
rect 263600 38203 287600 38523
rect 255946 37313 295254 38203
rect 295574 36993 310426 39573
rect 310746 38523 350054 39573
rect 318400 38203 342400 38523
rect 310746 37313 350054 38203
rect 350374 36993 365226 39573
rect 365546 38523 404854 39573
rect 373200 38203 397200 38523
rect 365546 37313 404854 38203
rect 405174 36993 420026 39573
rect 420346 38523 459654 39573
rect 428000 38203 452000 38523
rect 420346 37313 459654 38203
rect 459974 36993 474826 39573
rect 475146 38523 514454 39573
rect 482800 38203 506800 38523
rect 475146 37313 514454 38203
rect 514774 36993 529626 39573
rect 529946 38523 569254 39573
rect 537600 38203 561600 38523
rect 529946 37313 569254 38203
rect 569574 36993 583426 39573
rect 583746 38523 623054 39573
rect 591400 38203 615400 38523
rect 583746 37313 623054 38203
rect 623374 36993 637226 39573
rect 637546 38523 677054 39573
rect 677374 39210 677707 39893
rect 678027 39530 679077 100254
rect 679397 71000 680287 100254
rect 680607 70000 681257 100206
rect 679397 39243 680287 70000
rect 680607 39706 681257 69000
rect 681577 39695 682467 100254
rect 682787 39680 683677 100254
rect 683997 39723 684647 100254
rect 684968 100000 685617 100254
rect 684967 70000 685617 100000
rect 685937 71000 686827 100254
rect 687147 70000 688947 100254
rect 684967 39733 685617 69000
rect 685937 39705 686827 70000
rect 684967 39403 685617 39413
rect 680607 39375 681257 39386
rect 683997 39385 685617 39403
rect 680607 39360 682467 39375
rect 683997 39360 686827 39385
rect 677374 38923 679077 39210
rect 680607 38923 686827 39360
rect 645200 38203 669200 38523
rect 637546 37313 677054 38203
rect 677374 36993 686827 38923
rect 30773 36343 39386 36993
rect 39706 36343 78993 36993
rect 79313 36343 93287 36993
rect 93607 36343 132793 36993
rect 133113 36343 186606 36993
rect 186926 36343 201887 36993
rect 202207 36343 241393 36993
rect 241713 36343 255687 36993
rect 256007 36343 295206 36993
rect 295526 36343 310487 36993
rect 310807 36343 350006 36993
rect 350326 36343 365287 36993
rect 365607 36343 404806 36993
rect 405126 36343 420087 36993
rect 420407 36343 459606 36993
rect 459926 36343 474887 36993
rect 475207 36343 514406 36993
rect 514726 36343 529687 36993
rect 530007 36343 569193 36993
rect 569513 36343 583487 36993
rect 583807 36343 622993 36993
rect 623313 36343 637287 36993
rect 637607 36343 677051 36993
rect 677371 36343 686827 36993
rect 30773 35133 39375 36343
rect 39695 35133 79054 36023
rect 30773 35049 39360 35133
rect 0 33603 39360 35049
rect 39680 33923 79054 34813
rect 0 32633 39403 33603
rect 39723 32953 79054 33603
rect 0 31983 39413 32633
rect 39733 32632 78800 32633
rect 39733 31983 79054 32632
rect 0 30773 39385 31983
rect 39705 30773 79054 31663
rect 0 28333 35049 30773
rect 35369 28653 79054 30453
rect 0 27163 39355 28333
rect 39675 27483 79054 28333
rect 0 26313 39384 27163
rect 39704 26313 79054 27163
rect 0 20683 39151 26313
rect 39471 21003 40200 25993
rect 40520 21003 43480 25993
rect 40000 21000 40200 21003
rect 43800 21000 44200 25993
rect 44520 21003 45480 25993
rect 45800 21000 46200 25993
rect 46800 21003 71600 25993
rect 71920 21003 74880 25993
rect 46800 21000 47600 21003
rect 51200 21000 51600 21003
rect 55200 21000 55600 21003
rect 59200 21000 59600 21003
rect 63200 21000 63600 21003
rect 67200 21000 67600 21003
rect 71200 21000 71600 21003
rect 75200 21000 75600 25993
rect 75920 21003 76880 25993
rect 77200 21000 77600 25993
rect 78200 21003 79054 25993
rect 78200 21000 78800 21003
rect 79374 20683 93226 36343
rect 133113 36023 147600 36343
rect 93546 35133 186654 36023
rect 133174 34813 147600 35133
rect 93546 33923 132854 34813
rect 133174 33923 186654 34813
rect 133174 33603 147600 33923
rect 93546 32953 132854 33603
rect 133174 32953 186654 33603
rect 133174 32633 147600 32953
rect 93800 32632 186400 32633
rect 93546 31983 186654 32632
rect 133174 31663 147600 31983
rect 93546 30773 132854 31663
rect 133174 30773 186654 31663
rect 133174 30453 147600 30773
rect 93546 28653 132854 30453
rect 133174 28653 186654 30453
rect 133174 28333 147600 28653
rect 93546 27483 132854 28333
rect 133174 27483 186654 28333
rect 133174 27163 147600 27483
rect 93546 26313 132854 27163
rect 133174 26313 186654 27163
rect 133174 25993 147600 26313
rect 93546 21003 94000 25993
rect 94320 21003 97280 25993
rect 93800 21000 94000 21003
rect 97600 21000 98000 25993
rect 98320 21003 99280 25993
rect 99600 21000 100000 25993
rect 100600 21003 125400 25993
rect 125720 21003 128680 25993
rect 100600 21000 101400 21003
rect 105000 21000 105400 21003
rect 109000 21000 109400 21003
rect 113000 21000 113400 21003
rect 117000 21000 117400 21003
rect 121000 21000 121400 21003
rect 125000 21000 125400 21003
rect 129000 21000 129400 25993
rect 129720 21003 130680 25993
rect 131000 21000 131400 25993
rect 132000 21003 132854 25993
rect 132000 21000 132600 21003
rect 133174 21000 147800 25993
rect 148120 21003 151080 25993
rect 151400 21000 151800 25993
rect 152120 21003 153080 25993
rect 153400 21000 153800 25993
rect 154400 21003 179200 25993
rect 179520 21003 182480 25993
rect 154400 21000 155200 21003
rect 158800 21000 159200 21003
rect 162800 21000 163200 21003
rect 166800 21000 167200 21003
rect 170800 21000 171200 21003
rect 174800 21000 175200 21003
rect 178800 21000 179200 21003
rect 182800 21000 183200 25993
rect 183520 21003 184480 25993
rect 184800 21000 185200 25993
rect 185800 21003 186654 25993
rect 185800 21000 186400 21003
rect 133174 20683 147600 21000
rect 186974 20683 201826 36343
rect 202146 35133 241454 36023
rect 202146 33923 241454 34813
rect 202146 32953 241454 33603
rect 202400 32632 241200 32633
rect 202146 31983 241454 32632
rect 202146 30773 241454 31663
rect 202146 28653 241454 30453
rect 202146 27483 241454 28333
rect 202146 26313 241454 27163
rect 202146 21003 202600 25993
rect 202920 21003 205880 25993
rect 202400 21000 202600 21003
rect 206200 21000 206600 25993
rect 206920 21003 207880 25993
rect 208200 21000 208600 25993
rect 209200 21003 234000 25993
rect 234320 21003 237280 25993
rect 209200 21000 210000 21003
rect 213600 21000 214000 21003
rect 217600 21000 218000 21003
rect 221600 21000 222000 21003
rect 225600 21000 226000 21003
rect 229600 21000 230000 21003
rect 233600 21000 234000 21003
rect 237600 21000 238000 25993
rect 238320 21003 239280 25993
rect 239600 21000 240000 25993
rect 240600 21003 241454 25993
rect 240600 21000 241200 21003
rect 241774 20683 255626 36343
rect 255946 35133 295254 36023
rect 255946 33923 295254 34813
rect 255946 32953 295254 33603
rect 256200 32632 295000 32633
rect 255946 31983 295254 32632
rect 255946 30773 295254 31663
rect 255946 28653 295254 30453
rect 255946 27483 295254 28333
rect 255946 26313 295254 27163
rect 255946 21003 256400 25993
rect 256720 21003 259680 25993
rect 256200 21000 256400 21003
rect 260000 21000 260400 25993
rect 260720 21003 261680 25993
rect 262000 21000 262400 25993
rect 263000 21003 287800 25993
rect 288120 21003 291080 25993
rect 263000 21000 263800 21003
rect 267400 21000 267800 21003
rect 271400 21000 271800 21003
rect 275400 21000 275800 21003
rect 279400 21000 279800 21003
rect 283400 21000 283800 21003
rect 287400 21000 287800 21003
rect 291400 21000 291800 25993
rect 292120 21003 293080 25993
rect 293400 21000 293800 25993
rect 294400 21003 295254 25993
rect 294400 21000 295000 21003
rect 295574 20683 310426 36343
rect 310746 35133 350054 36023
rect 310746 33923 350054 34813
rect 310746 32953 350054 33603
rect 311000 32632 349800 32633
rect 310746 31983 350054 32632
rect 310746 30773 350054 31663
rect 310746 28653 350054 30453
rect 310746 27483 350054 28333
rect 310746 26313 350054 27163
rect 310746 21003 311200 25993
rect 311520 21003 314480 25993
rect 311000 21000 311200 21003
rect 314800 21000 315200 25993
rect 315520 21003 316480 25993
rect 316800 21000 317200 25993
rect 317800 21003 342600 25993
rect 342920 21003 345880 25993
rect 317800 21000 318600 21003
rect 322200 21000 322600 21003
rect 326200 21000 326600 21003
rect 330200 21000 330600 21003
rect 334200 21000 334600 21003
rect 338200 21000 338600 21003
rect 342200 21000 342600 21003
rect 346200 21000 346600 25993
rect 346920 21003 347880 25993
rect 348200 21000 348600 25993
rect 349200 21003 350054 25993
rect 349200 21000 349800 21003
rect 350374 20683 365226 36343
rect 365546 35133 404854 36023
rect 365546 33923 404854 34813
rect 365546 32953 404854 33603
rect 365800 32632 404600 32633
rect 365546 31983 404854 32632
rect 365546 30773 404854 31663
rect 365546 28653 404854 30453
rect 365546 27483 404854 28333
rect 365546 26313 404854 27163
rect 365546 21003 366000 25993
rect 366320 21003 369280 25993
rect 365800 21000 366000 21003
rect 369600 21000 370000 25993
rect 370320 21003 371280 25993
rect 371600 21000 372000 25993
rect 372600 21003 397400 25993
rect 397720 21003 400680 25993
rect 372600 21000 373400 21003
rect 377000 21000 377400 21003
rect 381000 21000 381400 21003
rect 385000 21000 385400 21003
rect 389000 21000 389400 21003
rect 393000 21000 393400 21003
rect 397000 21000 397400 21003
rect 401000 21000 401400 25993
rect 401720 21003 402680 25993
rect 403000 21000 403400 25993
rect 404000 21003 404854 25993
rect 404000 21000 404600 21003
rect 405174 20683 420026 36343
rect 420346 35133 459654 36023
rect 420346 33923 459654 34813
rect 420346 32953 459654 33603
rect 420600 32632 459400 32633
rect 420346 31983 459654 32632
rect 420346 30773 459654 31663
rect 420346 28653 459654 30453
rect 420346 27483 459654 28333
rect 420346 26313 459654 27163
rect 420346 21003 420800 25993
rect 421120 21003 424080 25993
rect 420600 21000 420800 21003
rect 424400 21000 424800 25993
rect 425120 21003 426080 25993
rect 426400 21000 426800 25993
rect 427400 21003 452200 25993
rect 452520 21003 455480 25993
rect 427400 21000 428200 21003
rect 431800 21000 432200 21003
rect 435800 21000 436200 21003
rect 439800 21000 440200 21003
rect 443800 21000 444200 21003
rect 447800 21000 448200 21003
rect 451800 21000 452200 21003
rect 455800 21000 456200 25993
rect 456520 21003 457480 25993
rect 457800 21000 458200 25993
rect 458800 21003 459654 25993
rect 458800 21000 459400 21003
rect 459974 20683 474826 36343
rect 475146 35133 514454 36023
rect 475146 33923 514454 34813
rect 475146 32953 514454 33603
rect 475400 32632 514200 32633
rect 475146 31983 514454 32632
rect 475146 30773 514454 31663
rect 475146 28653 514454 30453
rect 475146 27483 514454 28333
rect 475146 26313 514454 27163
rect 475146 21003 475600 25993
rect 475920 21003 478880 25993
rect 475400 21000 475600 21003
rect 479200 21000 479600 25993
rect 479920 21003 480880 25993
rect 481200 21000 481600 25993
rect 482200 21003 507000 25993
rect 507320 21003 510280 25993
rect 482200 21000 483000 21003
rect 486600 21000 487000 21003
rect 490600 21000 491000 21003
rect 494600 21000 495000 21003
rect 498600 21000 499000 21003
rect 502600 21000 503000 21003
rect 506600 21000 507000 21003
rect 510600 21000 511000 25993
rect 511320 21003 512280 25993
rect 512600 21000 513000 25993
rect 513600 21003 514454 25993
rect 513600 21000 514200 21003
rect 514774 20683 529626 36343
rect 529946 35133 569254 36023
rect 529946 33923 569254 34813
rect 529946 32953 569254 33603
rect 530200 32632 569000 32633
rect 529946 31983 569254 32632
rect 529946 30773 569254 31663
rect 529946 28653 569254 30453
rect 529946 27483 569254 28333
rect 529946 26313 569254 27163
rect 529946 21003 530400 25993
rect 530720 21003 533680 25993
rect 530200 21000 530400 21003
rect 534000 21000 534400 25993
rect 534720 21003 535680 25993
rect 536000 21000 536400 25993
rect 537000 21003 561800 25993
rect 562120 21003 565080 25993
rect 537000 21000 537800 21003
rect 541400 21000 541800 21003
rect 545400 21000 545800 21003
rect 549400 21000 549800 21003
rect 553400 21000 553800 21003
rect 557400 21000 557800 21003
rect 561400 21000 561800 21003
rect 565400 21000 565800 25993
rect 566120 21003 567080 25993
rect 567400 21000 567800 25993
rect 568400 21003 569254 25993
rect 568400 21000 569000 21003
rect 569574 20683 583426 36343
rect 583746 35133 623054 36023
rect 583746 33923 623054 34813
rect 583746 32953 623054 33603
rect 584000 32632 622800 32633
rect 583746 31983 623054 32632
rect 583746 30773 623054 31663
rect 583746 28653 623054 30453
rect 583746 27483 623054 28333
rect 583746 26313 623054 27163
rect 583746 21003 584200 25993
rect 584520 21003 587480 25993
rect 584000 21000 584200 21003
rect 587800 21000 588200 25993
rect 588520 21003 589480 25993
rect 589800 21000 590200 25993
rect 590800 21003 615600 25993
rect 615920 21003 618880 25993
rect 590800 21000 591600 21003
rect 595200 21000 595600 21003
rect 599200 21000 599600 21003
rect 603200 21000 603600 21003
rect 607200 21000 607600 21003
rect 611200 21000 611600 21003
rect 615200 21000 615600 21003
rect 619200 21000 619600 25993
rect 619920 21003 620880 25993
rect 621200 21000 621600 25993
rect 622200 21003 623054 25993
rect 622200 21000 622800 21003
rect 623374 20683 637226 36343
rect 637546 35133 677054 36023
rect 677374 35049 686827 36343
rect 687147 35369 688947 69000
rect 689267 39675 690117 100254
rect 690437 39704 691287 100254
rect 691607 100000 696597 100254
rect 696917 100000 717600 100574
rect 691607 99800 696600 100000
rect 691607 98800 696600 99200
rect 691607 95520 696597 98480
rect 691607 94800 696600 95200
rect 691607 91520 696597 94480
rect 691607 90800 696600 91200
rect 691607 87520 696597 90480
rect 691607 86800 696600 87200
rect 691607 83520 696597 86480
rect 691607 82800 696600 83200
rect 691607 79520 696597 82480
rect 691607 78800 696600 79200
rect 691607 75520 696597 78480
rect 691607 74800 696600 75200
rect 691607 71520 696597 74480
rect 691607 70800 696600 71200
rect 691607 69800 696600 70200
rect 691607 68800 696600 69200
rect 691607 67800 696600 68200
rect 691607 64520 696597 67480
rect 691607 63800 696600 64200
rect 691607 60520 696597 63480
rect 691607 59800 696600 60200
rect 691607 56520 696597 59480
rect 691607 55800 696600 56200
rect 691607 52520 696597 55480
rect 691607 51800 696600 52200
rect 691607 48520 696597 51480
rect 691607 47800 696600 48200
rect 691607 44520 696597 47480
rect 691607 43800 696600 44200
rect 691607 40520 696597 43480
rect 691607 40000 696600 40200
rect 712757 40000 717600 100000
rect 691607 39471 696597 40000
rect 690437 39355 691287 39384
rect 689267 39151 691287 39355
rect 696917 39151 717600 40000
rect 689267 35049 717600 39151
rect 637546 33923 677054 34813
rect 637546 32953 677054 33603
rect 637800 32632 676800 32633
rect 637546 31983 677054 32632
rect 637546 30773 677054 31663
rect 677374 30773 717600 35049
rect 637546 28653 682231 30453
rect 682551 28333 717600 30773
rect 637546 27483 677054 28333
rect 637546 26313 677054 27163
rect 677374 26313 717600 28333
rect 637546 21003 638000 25993
rect 638320 21003 641280 25993
rect 637800 21000 638000 21003
rect 641600 21000 642000 25993
rect 642320 21003 643280 25993
rect 643600 21000 644000 25993
rect 644600 21003 669400 25993
rect 669720 21003 672680 25993
rect 644600 21000 645400 21003
rect 649000 21000 649400 21003
rect 653000 21000 653400 21003
rect 657000 21000 657400 21003
rect 661000 21000 661400 21003
rect 665000 21000 665400 21003
rect 669000 21000 669400 21003
rect 673000 21000 673400 25993
rect 673720 21003 674680 25993
rect 675000 21000 675400 25993
rect 676000 21003 677171 25993
rect 676000 21000 676800 21003
rect 677491 20683 717600 26313
rect 0 4843 40000 20683
rect 78800 19518 93800 20683
rect 78800 6355 79720 19518
rect 92900 6355 93800 19518
rect 78800 4843 93800 6355
rect 132600 19518 147600 20683
rect 132600 6355 133520 19518
rect 146700 6355 147600 19518
rect 132600 4843 147600 6355
rect 186400 19408 202400 20683
rect 186400 6278 187320 19408
rect 200480 6278 202400 19408
rect 186400 4843 202400 6278
rect 241200 19892 256200 20683
rect 241200 5766 242689 19892
rect 254657 5766 256200 19892
rect 241200 4843 256200 5766
rect 295000 19408 311000 20683
rect 295000 6278 295920 19408
rect 309080 6278 311000 19408
rect 295000 4843 311000 6278
rect 349800 19408 365800 20683
rect 349800 6278 350720 19408
rect 363880 6278 365800 19408
rect 349800 4843 365800 6278
rect 404600 19408 420600 20683
rect 404600 6278 405520 19408
rect 418680 6278 420600 19408
rect 404600 4843 420600 6278
rect 459400 19408 475400 20683
rect 459400 6278 460320 19408
rect 473480 6278 475400 19408
rect 459400 4843 475400 6278
rect 514200 19408 530200 20683
rect 514200 6278 515120 19408
rect 528280 6278 530200 19408
rect 514200 4843 530200 6278
rect 569000 19518 584000 20683
rect 569000 6355 569920 19518
rect 570240 6675 582780 19198
rect 583100 6355 584000 19518
rect 569000 4843 584000 6355
rect 622800 19518 637800 20683
rect 622800 6355 623720 19518
rect 636900 6355 637800 19518
rect 622800 4843 637800 6355
rect 676800 4843 717600 20683
rect 0 0 717600 4843
<< labels >>
rlabel metal5 s 187640 6598 200160 19088 6 clock
port 1 nsew
rlabel metal2 s 187327 41713 187383 42193 6 clock_core
port 2 nsew
rlabel metal2 s 194043 41713 194099 42193 6 por
port 3 nsew
rlabel metal5 s 351040 6598 363560 19088 6 flash_clk
port 4 nsew
rlabel metal2 s 361767 41713 361823 42193 6 flash_clk_core
port 5 nsew
rlabel metal2 s 357443 41713 357499 42193 6 flash_clk_ieb_core
port 6 nsew
rlabel metal2 s 364895 41713 364951 42193 6 flash_clk_oeb_core
port 7 nsew
rlabel metal5 s 296240 6598 308760 19088 6 flash_csb
port 8 nsew
rlabel metal2 s 306967 41713 307023 42193 6 flash_csb_core
port 9 nsew
rlabel metal2 s 302643 41713 302699 42193 6 flash_csb_ieb_core
port 10 nsew
rlabel metal2 s 310095 41713 310151 42193 6 flash_csb_oeb_core
port 11 nsew
rlabel metal5 s 405840 6598 418360 19088 6 flash_io0
port 12 nsew
rlabel metal2 s 405527 41713 405583 42193 6 flash_io0_di_core
port 13 nsew
rlabel metal2 s 416567 41713 416623 42193 6 flash_io0_do_core
port 14 nsew
rlabel metal2 s 415371 41713 415427 41806 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 412243 41713 412299 41806 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 409207 41713 409263 41806 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 415371 41806 415532 41822 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 412243 41806 412404 41822 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 409207 41806 409368 41822 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 415371 41822 415544 41834 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 415492 41834 415544 41886 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 415371 41834 415427 42193 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 412243 41822 412416 41834 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 412364 41834 412416 41886 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 412243 41834 412299 42193 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 409207 41822 409380 41834 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 409328 41834 409380 41886 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 409207 41834 409263 42193 6 flash_io0_ieb_core
port 15 nsew
rlabel via1 s 415492 41828 415544 41880 6 flash_io0_ieb_core
port 15 nsew
rlabel via1 s 412364 41828 412416 41880 6 flash_io0_ieb_core
port 15 nsew
rlabel via1 s 409328 41828 409380 41880 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 415486 41828 415550 41840 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 412358 41828 412422 41840 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 409322 41828 409386 41840 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 409322 41840 415550 41868 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 415486 41868 415550 41880 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 412358 41868 412422 41880 6 flash_io0_ieb_core
port 15 nsew
rlabel metal1 s 409322 41868 409386 41880 6 flash_io0_ieb_core
port 15 nsew
rlabel metal2 s 419695 41713 419751 41806 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 411047 41713 411103 41806 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 419552 41806 419751 41822 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 419540 41822 419751 41834 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 419695 41834 419751 42193 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 419540 41834 419592 41886 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 411047 41806 411208 41834 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 411180 41834 411208 41890 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 411168 41890 411220 41954 6 flash_io0_oeb_core
port 16 nsew
rlabel metal2 s 411047 41834 411103 42193 6 flash_io0_oeb_core
port 16 nsew
rlabel via1 s 419540 41828 419592 41880 6 flash_io0_oeb_core
port 16 nsew
rlabel via1 s 411168 41896 411220 41948 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 419534 41828 419598 41840 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 415596 41840 419598 41868 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 419534 41868 419598 41880 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 415596 41868 415624 41908 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 411162 41896 411226 41908 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 411162 41908 415624 41936 6 flash_io0_oeb_core
port 16 nsew
rlabel metal1 s 411162 41936 411226 41948 6 flash_io0_oeb_core
port 16 nsew
rlabel metal5 s 460640 6598 473160 19088 6 flash_io1
port 17 nsew
rlabel metal2 s 460327 41713 460383 42193 6 flash_io1_di_core
port 18 nsew
rlabel metal2 s 471367 41713 471423 42193 6 flash_io1_do_core
port 19 nsew
rlabel metal2 s 470171 41713 470227 41806 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 470048 41754 470100 41806 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 470048 41806 470227 41818 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 467196 41754 467248 41806 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 467043 41713 467099 41806 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 467043 41806 467248 41818 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 464160 41754 464212 41806 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 464007 41713 464063 41806 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 464007 41806 464212 41818 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 470060 41818 470227 41834 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 467043 41818 467236 41834 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 464007 41818 464200 41834 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 470171 41834 470227 42193 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 467043 41834 467099 42193 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 464007 41834 464063 42193 6 flash_io1_ieb_core
port 20 nsew
rlabel via1 s 470048 41760 470100 41812 6 flash_io1_ieb_core
port 20 nsew
rlabel via1 s 467196 41760 467248 41812 6 flash_io1_ieb_core
port 20 nsew
rlabel via1 s 464160 41760 464212 41812 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 470042 41760 470106 41772 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 467190 41760 467254 41772 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 464154 41760 464218 41772 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 464154 41772 470106 41800 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 470042 41800 470106 41812 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 467190 41800 467254 41812 6 flash_io1_ieb_core
port 20 nsew
rlabel metal1 s 464154 41800 464218 41812 6 flash_io1_ieb_core
port 20 nsew
rlabel metal2 s 474495 41713 474551 41806 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 465847 41713 465903 41806 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 474384 41806 474551 41834 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 474495 41834 474551 42193 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 474384 41834 474412 41890 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 465847 41806 466040 41834 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 466012 41834 466040 41890 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 474372 41890 474424 41954 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 466000 41890 466052 41954 6 flash_io1_oeb_core
port 21 nsew
rlabel metal2 s 465847 41834 465903 42193 6 flash_io1_oeb_core
port 21 nsew
rlabel via1 s 474372 41896 474424 41948 6 flash_io1_oeb_core
port 21 nsew
rlabel via1 s 466000 41896 466052 41948 6 flash_io1_oeb_core
port 21 nsew
rlabel metal1 s 474366 41896 474430 41908 6 flash_io1_oeb_core
port 21 nsew
rlabel metal1 s 465994 41896 466058 41908 6 flash_io1_oeb_core
port 21 nsew
rlabel metal1 s 465994 41908 474430 41936 6 flash_io1_oeb_core
port 21 nsew
rlabel metal1 s 474366 41936 474430 41948 6 flash_io1_oeb_core
port 21 nsew
rlabel metal1 s 465994 41936 466058 41948 6 flash_io1_oeb_core
port 21 nsew
rlabel metal5 s 515440 6598 527960 19088 6 gpio
port 22 nsew
rlabel metal2 s 515127 41713 515183 42193 6 gpio_in_core
port 23 nsew
rlabel metal2 s 521843 41713 521899 42193 6 gpio_inenb_core
port 24 nsew
rlabel metal2 s 520647 41713 520703 42193 6 gpio_mode0_core
port 25 nsew
rlabel metal2 s 524971 41713 525027 41806 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 518807 41713 518863 41806 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 524892 41806 525027 41822 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 518807 41806 518940 41822 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 524880 41822 525027 41834 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 524971 41834 525027 42193 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 524880 41834 524932 41886 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 518807 41822 518952 41834 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 518900 41834 518952 41886 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 518807 41834 518863 42193 6 gpio_mode1_core
port 26 nsew
rlabel via1 s 524880 41828 524932 41880 6 gpio_mode1_core
port 26 nsew
rlabel via1 s 518900 41828 518952 41880 6 gpio_mode1_core
port 26 nsew
rlabel metal1 s 524874 41828 524938 41840 6 gpio_mode1_core
port 26 nsew
rlabel metal1 s 518894 41828 518958 41840 6 gpio_mode1_core
port 26 nsew
rlabel metal1 s 518894 41840 524938 41868 6 gpio_mode1_core
port 26 nsew
rlabel metal1 s 524874 41868 524938 41880 6 gpio_mode1_core
port 26 nsew
rlabel metal1 s 518894 41868 518958 41880 6 gpio_mode1_core
port 26 nsew
rlabel metal2 s 526167 41713 526223 42193 6 gpio_out_core
port 27 nsew
rlabel metal2 s 529295 41713 529351 42193 6 gpio_outenb_core
port 28 nsew
rlabel metal5 s 6086 69863 19572 81191 6 vccd
port 29 nsew
rlabel metal5 s 624040 6675 636580 19198 6 vdda
port 30 nsew
rlabel metal5 s 6675 111420 19198 123960 6 vddio
port 31 nsew
rlabel metal5 s 80040 6675 92580 19198 6 vssa
port 32 nsew
rlabel metal5 s 243009 6086 254337 19572 6 vssd
port 33 nsew
rlabel metal5 s 334620 1018402 347160 1030925 6 vssio
port 34 nsew
rlabel metal5 s 698512 101240 711002 113760 6 mprj_io[0]
port 35 nsew
rlabel metal2 s 675407 105803 675887 105859 6 mprj_io_analog_en[0]
port 36 nsew
rlabel metal2 s 675407 107091 675887 107147 6 mprj_io_analog_pol[0]
port 37 nsew
rlabel metal2 s 675407 110127 675887 110183 6 mprj_io_analog_sel[0]
port 38 nsew
rlabel metal2 s 675407 106447 675887 106503 6 mprj_io_dm[0]
port 39 nsew
rlabel metal2 s 675407 104607 675887 104663 6 mprj_io_dm[1]
port 40 nsew
rlabel metal2 s 675407 110771 675887 110827 6 mprj_io_dm[2]
port 41 nsew
rlabel metal2 s 675407 108931 675887 108987 6 mprj_io_enh[0]
port 42 nsew
rlabel metal2 s 675407 109575 675887 109631 6 mprj_io_hldh_n[0]
port 43 nsew
rlabel metal2 s 675407 111415 675887 111471 6 mprj_io_holdover[0]
port 44 nsew
rlabel metal2 s 675407 114451 675887 114507 6 mprj_io_ib_mode_sel[0]
port 45 nsew
rlabel metal2 s 675407 107643 675887 107699 6 mprj_io_inp_dis[0]
port 46 nsew
rlabel metal2 s 675407 115095 675887 115151 6 mprj_io_oeb[0]
port 47 nsew
rlabel metal2 s 675407 111967 675887 112023 6 mprj_io_out[0]
port 48 nsew
rlabel metal2 s 675407 102767 675887 102823 6 mprj_io_slow_sel[0]
port 49 nsew
rlabel metal2 s 675407 113807 675887 113863 6 mprj_io_vtrip_sel[0]
port 50 nsew
rlabel metal2 s 675407 100927 675887 100983 6 mprj_io_in[0]
port 51 nsew
rlabel metal5 s 698512 684440 711002 696960 6 mprj_io[10]
port 52 nsew
rlabel metal2 s 675407 689003 675887 689059 6 mprj_io_analog_en[10]
port 53 nsew
rlabel metal2 s 675407 690291 675887 690347 6 mprj_io_analog_pol[10]
port 54 nsew
rlabel metal2 s 675407 693327 675887 693383 6 mprj_io_analog_sel[10]
port 55 nsew
rlabel metal2 s 675407 689647 675887 689703 6 mprj_io_dm[30]
port 56 nsew
rlabel metal2 s 675407 687807 675887 687863 6 mprj_io_dm[31]
port 57 nsew
rlabel metal2 s 675407 693971 675887 694027 6 mprj_io_dm[32]
port 58 nsew
rlabel metal2 s 675407 692131 675887 692187 6 mprj_io_enh[10]
port 59 nsew
rlabel metal2 s 675407 692775 675887 692831 6 mprj_io_hldh_n[10]
port 60 nsew
rlabel metal2 s 675407 694615 675887 694671 6 mprj_io_holdover[10]
port 61 nsew
rlabel metal2 s 675407 697651 675887 697707 6 mprj_io_ib_mode_sel[10]
port 62 nsew
rlabel metal2 s 675407 690843 675887 690899 6 mprj_io_inp_dis[10]
port 63 nsew
rlabel metal2 s 675407 698295 675887 698351 6 mprj_io_oeb[10]
port 64 nsew
rlabel metal2 s 675407 695167 675887 695223 6 mprj_io_out[10]
port 65 nsew
rlabel metal2 s 675407 685967 675887 686023 6 mprj_io_slow_sel[10]
port 66 nsew
rlabel metal2 s 675407 697007 675887 697063 6 mprj_io_vtrip_sel[10]
port 67 nsew
rlabel metal2 s 675407 684127 675887 684183 6 mprj_io_in[10]
port 68 nsew
rlabel metal5 s 698512 729440 711002 741960 6 mprj_io[11]
port 69 nsew
rlabel metal2 s 675407 734003 675887 734059 6 mprj_io_analog_en[11]
port 70 nsew
rlabel metal2 s 675407 735291 675887 735347 6 mprj_io_analog_pol[11]
port 71 nsew
rlabel metal2 s 675407 738327 675887 738383 6 mprj_io_analog_sel[11]
port 72 nsew
rlabel metal2 s 675407 734647 675887 734703 6 mprj_io_dm[33]
port 73 nsew
rlabel metal2 s 675407 732807 675887 732863 6 mprj_io_dm[34]
port 74 nsew
rlabel metal2 s 675407 738971 675887 739027 6 mprj_io_dm[35]
port 75 nsew
rlabel metal2 s 675407 737131 675887 737187 6 mprj_io_enh[11]
port 76 nsew
rlabel metal2 s 675407 737775 675887 737831 6 mprj_io_hldh_n[11]
port 77 nsew
rlabel metal2 s 675407 739615 675887 739671 6 mprj_io_holdover[11]
port 78 nsew
rlabel metal2 s 675407 742651 675887 742707 6 mprj_io_ib_mode_sel[11]
port 79 nsew
rlabel metal2 s 675407 735843 675887 735899 6 mprj_io_inp_dis[11]
port 80 nsew
rlabel metal2 s 675407 743295 675887 743351 6 mprj_io_oeb[11]
port 81 nsew
rlabel metal2 s 675407 740167 675887 740223 6 mprj_io_out[11]
port 82 nsew
rlabel metal2 s 675407 730967 675887 731023 6 mprj_io_slow_sel[11]
port 83 nsew
rlabel metal2 s 675407 742007 675887 742063 6 mprj_io_vtrip_sel[11]
port 84 nsew
rlabel metal2 s 675407 729127 675887 729183 6 mprj_io_in[11]
port 85 nsew
rlabel metal5 s 698512 774440 711002 786960 6 mprj_io[12]
port 86 nsew
rlabel metal2 s 675407 779003 675887 779059 6 mprj_io_analog_en[12]
port 87 nsew
rlabel metal2 s 675407 780291 675887 780347 6 mprj_io_analog_pol[12]
port 88 nsew
rlabel metal2 s 675407 783327 675887 783383 6 mprj_io_analog_sel[12]
port 89 nsew
rlabel metal2 s 675407 779647 675887 779703 6 mprj_io_dm[36]
port 90 nsew
rlabel metal2 s 675407 777807 675887 777863 6 mprj_io_dm[37]
port 91 nsew
rlabel metal2 s 675407 783971 675887 784027 6 mprj_io_dm[38]
port 92 nsew
rlabel metal2 s 675407 782131 675887 782187 6 mprj_io_enh[12]
port 93 nsew
rlabel metal2 s 675407 782775 675887 782831 6 mprj_io_hldh_n[12]
port 94 nsew
rlabel metal2 s 675407 784615 675887 784671 6 mprj_io_holdover[12]
port 95 nsew
rlabel metal2 s 675407 787651 675887 787707 6 mprj_io_ib_mode_sel[12]
port 96 nsew
rlabel metal2 s 675407 780843 675887 780899 6 mprj_io_inp_dis[12]
port 97 nsew
rlabel metal2 s 675407 788295 675887 788351 6 mprj_io_oeb[12]
port 98 nsew
rlabel metal2 s 675407 785167 675887 785223 6 mprj_io_out[12]
port 99 nsew
rlabel metal2 s 675407 775967 675887 776023 6 mprj_io_slow_sel[12]
port 100 nsew
rlabel metal2 s 675407 787007 675887 787063 6 mprj_io_vtrip_sel[12]
port 101 nsew
rlabel metal2 s 675407 774127 675887 774183 6 mprj_io_in[12]
port 102 nsew
rlabel metal5 s 698512 863640 711002 876160 6 mprj_io[13]
port 103 nsew
rlabel metal2 s 675407 868203 675887 868259 6 mprj_io_analog_en[13]
port 104 nsew
rlabel metal2 s 675407 869491 675887 869547 6 mprj_io_analog_pol[13]
port 105 nsew
rlabel metal2 s 675407 872527 675887 872583 6 mprj_io_analog_sel[13]
port 106 nsew
rlabel metal2 s 675407 868847 675887 868903 6 mprj_io_dm[39]
port 107 nsew
rlabel metal2 s 675407 867007 675887 867063 6 mprj_io_dm[40]
port 108 nsew
rlabel metal2 s 675407 873171 675887 873227 6 mprj_io_dm[41]
port 109 nsew
rlabel metal2 s 675407 871331 675887 871387 6 mprj_io_enh[13]
port 110 nsew
rlabel metal2 s 675407 871975 675887 872031 6 mprj_io_hldh_n[13]
port 111 nsew
rlabel metal2 s 675407 873815 675887 873871 6 mprj_io_holdover[13]
port 112 nsew
rlabel metal2 s 675407 876851 675887 876907 6 mprj_io_ib_mode_sel[13]
port 113 nsew
rlabel metal2 s 675407 870043 675887 870099 6 mprj_io_inp_dis[13]
port 114 nsew
rlabel metal2 s 675407 877495 675887 877551 6 mprj_io_oeb[13]
port 115 nsew
rlabel metal2 s 675407 874367 675887 874423 6 mprj_io_out[13]
port 116 nsew
rlabel metal2 s 675407 865167 675887 865223 6 mprj_io_slow_sel[13]
port 117 nsew
rlabel metal2 s 675407 876207 675887 876263 6 mprj_io_vtrip_sel[13]
port 118 nsew
rlabel metal2 s 675407 863327 675887 863383 6 mprj_io_in[13]
port 119 nsew
rlabel metal5 s 698512 952840 711002 965360 6 mprj_io[14]
port 120 nsew
rlabel metal2 s 675407 957403 675887 957459 6 mprj_io_analog_en[14]
port 121 nsew
rlabel metal2 s 675407 958691 675887 958747 6 mprj_io_analog_pol[14]
port 122 nsew
rlabel metal2 s 675407 961727 675887 961783 6 mprj_io_analog_sel[14]
port 123 nsew
rlabel metal2 s 675407 958047 675887 958103 6 mprj_io_dm[42]
port 124 nsew
rlabel metal2 s 675407 956207 675887 956263 6 mprj_io_dm[43]
port 125 nsew
rlabel metal2 s 675407 962371 675887 962427 6 mprj_io_dm[44]
port 126 nsew
rlabel metal2 s 675407 960531 675887 960587 6 mprj_io_enh[14]
port 127 nsew
rlabel metal2 s 675407 961175 675887 961231 6 mprj_io_hldh_n[14]
port 128 nsew
rlabel metal2 s 675407 963015 675887 963071 6 mprj_io_holdover[14]
port 129 nsew
rlabel metal2 s 675407 966051 675887 966107 6 mprj_io_ib_mode_sel[14]
port 130 nsew
rlabel metal2 s 675407 959243 675887 959299 6 mprj_io_inp_dis[14]
port 131 nsew
rlabel metal2 s 675407 966695 675887 966751 6 mprj_io_oeb[14]
port 132 nsew
rlabel metal2 s 675407 963567 675887 963623 6 mprj_io_out[14]
port 133 nsew
rlabel metal2 s 675407 954367 675887 954423 6 mprj_io_slow_sel[14]
port 134 nsew
rlabel metal2 s 675407 965407 675887 965463 6 mprj_io_vtrip_sel[14]
port 135 nsew
rlabel metal2 s 675407 952527 675887 952583 6 mprj_io_in[14]
port 136 nsew
rlabel metal5 s 628240 1018512 640760 1031002 6 mprj_io[15]
port 137 nsew
rlabel metal2 s 636141 995407 636197 995887 6 mprj_io_analog_en[15]
port 138 nsew
rlabel metal2 s 634853 995407 634909 995887 6 mprj_io_analog_pol[15]
port 139 nsew
rlabel metal2 s 631817 995407 631873 995887 6 mprj_io_analog_sel[15]
port 140 nsew
rlabel metal2 s 635497 995407 635553 995887 6 mprj_io_dm[45]
port 141 nsew
rlabel metal2 s 637337 995407 637393 995887 6 mprj_io_dm[46]
port 142 nsew
rlabel metal2 s 631173 995407 631229 995887 6 mprj_io_dm[47]
port 143 nsew
rlabel metal2 s 633013 995407 633069 995887 6 mprj_io_enh[15]
port 144 nsew
rlabel metal2 s 632369 995407 632425 995887 6 mprj_io_hldh_n[15]
port 145 nsew
rlabel metal2 s 630529 995407 630585 995887 6 mprj_io_holdover[15]
port 146 nsew
rlabel metal2 s 627493 995407 627549 995887 6 mprj_io_ib_mode_sel[15]
port 147 nsew
rlabel metal2 s 634301 995407 634357 995887 6 mprj_io_inp_dis[15]
port 148 nsew
rlabel metal2 s 626849 995407 626905 995887 6 mprj_io_oeb[15]
port 149 nsew
rlabel metal2 s 629977 995407 630033 995887 6 mprj_io_out[15]
port 150 nsew
rlabel metal2 s 639177 995407 639233 995887 6 mprj_io_slow_sel[15]
port 151 nsew
rlabel metal2 s 628137 995407 628193 995887 6 mprj_io_vtrip_sel[15]
port 152 nsew
rlabel metal2 s 641017 995407 641073 995887 6 mprj_io_in[15]
port 153 nsew
rlabel metal5 s 526440 1018512 538960 1031002 6 mprj_io[16]
port 154 nsew
rlabel metal2 s 534341 995407 534397 995887 6 mprj_io_analog_en[16]
port 155 nsew
rlabel metal2 s 533053 995407 533109 995887 6 mprj_io_analog_pol[16]
port 156 nsew
rlabel metal2 s 530017 995407 530073 995887 6 mprj_io_analog_sel[16]
port 157 nsew
rlabel metal2 s 533697 995407 533753 995887 6 mprj_io_dm[48]
port 158 nsew
rlabel metal2 s 535537 995407 535593 995887 6 mprj_io_dm[49]
port 159 nsew
rlabel metal2 s 529373 995407 529429 995887 6 mprj_io_dm[50]
port 160 nsew
rlabel metal2 s 531213 995407 531269 995887 6 mprj_io_enh[16]
port 161 nsew
rlabel metal2 s 530569 995407 530625 995887 6 mprj_io_hldh_n[16]
port 162 nsew
rlabel metal2 s 528729 995407 528785 995887 6 mprj_io_holdover[16]
port 163 nsew
rlabel metal2 s 525693 995407 525749 995887 6 mprj_io_ib_mode_sel[16]
port 164 nsew
rlabel metal2 s 532501 995407 532557 995887 6 mprj_io_inp_dis[16]
port 165 nsew
rlabel metal2 s 525049 995407 525105 995887 6 mprj_io_oeb[16]
port 166 nsew
rlabel metal2 s 528177 995407 528233 995887 6 mprj_io_out[16]
port 167 nsew
rlabel metal2 s 537377 995407 537433 995887 6 mprj_io_slow_sel[16]
port 168 nsew
rlabel metal2 s 526337 995407 526393 995887 6 mprj_io_vtrip_sel[16]
port 169 nsew
rlabel metal2 s 539217 995407 539273 995887 6 mprj_io_in[16]
port 170 nsew
rlabel metal5 s 475040 1018512 487560 1031002 6 mprj_io[17]
port 171 nsew
rlabel metal2 s 482941 995407 482997 995887 6 mprj_io_analog_en[17]
port 172 nsew
rlabel metal2 s 481653 995407 481709 995887 6 mprj_io_analog_pol[17]
port 173 nsew
rlabel metal2 s 478617 995407 478673 995887 6 mprj_io_analog_sel[17]
port 174 nsew
rlabel metal2 s 482297 995407 482353 995887 6 mprj_io_dm[51]
port 175 nsew
rlabel metal2 s 484137 995407 484193 995887 6 mprj_io_dm[52]
port 176 nsew
rlabel metal2 s 477973 995407 478029 995887 6 mprj_io_dm[53]
port 177 nsew
rlabel metal2 s 479813 995407 479869 995887 6 mprj_io_enh[17]
port 178 nsew
rlabel metal2 s 479169 995407 479225 995887 6 mprj_io_hldh_n[17]
port 179 nsew
rlabel metal2 s 477329 995407 477385 995887 6 mprj_io_holdover[17]
port 180 nsew
rlabel metal2 s 474293 995407 474349 995887 6 mprj_io_ib_mode_sel[17]
port 181 nsew
rlabel metal2 s 481101 995407 481157 995887 6 mprj_io_inp_dis[17]
port 182 nsew
rlabel metal2 s 473649 995407 473705 995887 6 mprj_io_oeb[17]
port 183 nsew
rlabel metal2 s 476777 995407 476833 995887 6 mprj_io_out[17]
port 184 nsew
rlabel metal2 s 485977 995407 486033 995887 6 mprj_io_slow_sel[17]
port 185 nsew
rlabel metal2 s 474937 995407 474993 995887 6 mprj_io_vtrip_sel[17]
port 186 nsew
rlabel metal2 s 487817 995407 487873 995887 6 mprj_io_in[17]
port 187 nsew
rlabel metal5 s 698512 146440 711002 158960 6 mprj_io[1]
port 188 nsew
rlabel metal2 s 675407 151003 675887 151059 6 mprj_io_analog_en[1]
port 189 nsew
rlabel metal2 s 675407 152291 675887 152347 6 mprj_io_analog_pol[1]
port 190 nsew
rlabel metal2 s 675407 155327 675887 155383 6 mprj_io_analog_sel[1]
port 191 nsew
rlabel metal2 s 675407 151647 675887 151703 6 mprj_io_dm[3]
port 192 nsew
rlabel metal2 s 675407 149807 675887 149863 6 mprj_io_dm[4]
port 193 nsew
rlabel metal2 s 675407 155971 675887 156027 6 mprj_io_dm[5]
port 194 nsew
rlabel metal2 s 675407 154131 675887 154187 6 mprj_io_enh[1]
port 195 nsew
rlabel metal2 s 675407 154775 675887 154831 6 mprj_io_hldh_n[1]
port 196 nsew
rlabel metal2 s 675407 156615 675887 156671 6 mprj_io_holdover[1]
port 197 nsew
rlabel metal2 s 675407 159651 675887 159707 6 mprj_io_ib_mode_sel[1]
port 198 nsew
rlabel metal2 s 675407 152843 675887 152899 6 mprj_io_inp_dis[1]
port 199 nsew
rlabel metal2 s 675407 160295 675887 160351 6 mprj_io_oeb[1]
port 200 nsew
rlabel metal2 s 675407 157167 675887 157223 6 mprj_io_out[1]
port 201 nsew
rlabel metal2 s 675407 147967 675887 148023 6 mprj_io_slow_sel[1]
port 202 nsew
rlabel metal2 s 675407 159007 675887 159063 6 mprj_io_vtrip_sel[1]
port 203 nsew
rlabel metal2 s 675407 146127 675887 146183 6 mprj_io_in[1]
port 204 nsew
rlabel metal5 s 698512 191440 711002 203960 6 mprj_io[2]
port 205 nsew
rlabel metal2 s 675407 196003 675887 196059 6 mprj_io_analog_en[2]
port 206 nsew
rlabel metal2 s 675407 197291 675887 197347 6 mprj_io_analog_pol[2]
port 207 nsew
rlabel metal2 s 675407 200327 675887 200383 6 mprj_io_analog_sel[2]
port 208 nsew
rlabel metal2 s 675407 196647 675887 196703 6 mprj_io_dm[6]
port 209 nsew
rlabel metal2 s 675407 194807 675887 194863 6 mprj_io_dm[7]
port 210 nsew
rlabel metal2 s 675407 200971 675887 201027 6 mprj_io_dm[8]
port 211 nsew
rlabel metal2 s 675407 199131 675887 199187 6 mprj_io_enh[2]
port 212 nsew
rlabel metal2 s 675407 199775 675887 199831 6 mprj_io_hldh_n[2]
port 213 nsew
rlabel metal2 s 675407 201615 675887 201671 6 mprj_io_holdover[2]
port 214 nsew
rlabel metal2 s 675407 204651 675887 204707 6 mprj_io_ib_mode_sel[2]
port 215 nsew
rlabel metal2 s 675407 197843 675887 197899 6 mprj_io_inp_dis[2]
port 216 nsew
rlabel metal2 s 675407 205295 675887 205351 6 mprj_io_oeb[2]
port 217 nsew
rlabel metal2 s 675407 202167 675887 202223 6 mprj_io_out[2]
port 218 nsew
rlabel metal2 s 675407 192967 675887 193023 6 mprj_io_slow_sel[2]
port 219 nsew
rlabel metal2 s 675407 204007 675887 204063 6 mprj_io_vtrip_sel[2]
port 220 nsew
rlabel metal2 s 675407 191127 675887 191183 6 mprj_io_in[2]
port 221 nsew
rlabel metal5 s 698512 236640 711002 249160 6 mprj_io[3]
port 222 nsew
rlabel metal2 s 675407 241203 675887 241259 6 mprj_io_analog_en[3]
port 223 nsew
rlabel metal2 s 675407 242491 675887 242547 6 mprj_io_analog_pol[3]
port 224 nsew
rlabel metal2 s 675407 245527 675887 245583 6 mprj_io_analog_sel[3]
port 225 nsew
rlabel metal2 s 675407 240007 675887 240063 6 mprj_io_dm[10]
port 226 nsew
rlabel metal2 s 675407 246171 675887 246227 6 mprj_io_dm[11]
port 227 nsew
rlabel metal2 s 675407 241847 675887 241903 6 mprj_io_dm[9]
port 228 nsew
rlabel metal2 s 675407 244331 675887 244387 6 mprj_io_enh[3]
port 229 nsew
rlabel metal2 s 675407 244975 675887 245031 6 mprj_io_hldh_n[3]
port 230 nsew
rlabel metal2 s 675407 246815 675887 246871 6 mprj_io_holdover[3]
port 231 nsew
rlabel metal2 s 675407 249851 675887 249907 6 mprj_io_ib_mode_sel[3]
port 232 nsew
rlabel metal2 s 675407 243043 675887 243099 6 mprj_io_inp_dis[3]
port 233 nsew
rlabel metal2 s 675407 250495 675887 250551 6 mprj_io_oeb[3]
port 234 nsew
rlabel metal2 s 675407 247367 675887 247423 6 mprj_io_out[3]
port 235 nsew
rlabel metal2 s 675407 238167 675887 238223 6 mprj_io_slow_sel[3]
port 236 nsew
rlabel metal2 s 675407 249207 675887 249263 6 mprj_io_vtrip_sel[3]
port 237 nsew
rlabel metal2 s 675407 236327 675887 236383 6 mprj_io_in[3]
port 238 nsew
rlabel metal5 s 698512 281640 711002 294160 6 mprj_io[4]
port 239 nsew
rlabel metal2 s 675407 286203 675887 286259 6 mprj_io_analog_en[4]
port 240 nsew
rlabel metal2 s 675407 287491 675887 287547 6 mprj_io_analog_pol[4]
port 241 nsew
rlabel metal2 s 675407 290527 675887 290583 6 mprj_io_analog_sel[4]
port 242 nsew
rlabel metal2 s 675407 286847 675887 286903 6 mprj_io_dm[12]
port 243 nsew
rlabel metal2 s 675407 285007 675887 285063 6 mprj_io_dm[13]
port 244 nsew
rlabel metal2 s 675407 291171 675887 291227 6 mprj_io_dm[14]
port 245 nsew
rlabel metal2 s 675407 289331 675887 289387 6 mprj_io_enh[4]
port 246 nsew
rlabel metal2 s 675407 289975 675887 290031 6 mprj_io_hldh_n[4]
port 247 nsew
rlabel metal2 s 675407 291815 675887 291871 6 mprj_io_holdover[4]
port 248 nsew
rlabel metal2 s 675407 294851 675887 294907 6 mprj_io_ib_mode_sel[4]
port 249 nsew
rlabel metal2 s 675407 288043 675887 288099 6 mprj_io_inp_dis[4]
port 250 nsew
rlabel metal2 s 675407 295495 675887 295551 6 mprj_io_oeb[4]
port 251 nsew
rlabel metal2 s 675407 292367 675887 292423 6 mprj_io_out[4]
port 252 nsew
rlabel metal2 s 675407 283167 675887 283223 6 mprj_io_slow_sel[4]
port 253 nsew
rlabel metal2 s 675407 294207 675887 294263 6 mprj_io_vtrip_sel[4]
port 254 nsew
rlabel metal2 s 675407 281327 675887 281383 6 mprj_io_in[4]
port 255 nsew
rlabel metal5 s 698512 326640 711002 339160 6 mprj_io[5]
port 256 nsew
rlabel metal2 s 675407 331203 675887 331259 6 mprj_io_analog_en[5]
port 257 nsew
rlabel metal2 s 675407 332491 675887 332547 6 mprj_io_analog_pol[5]
port 258 nsew
rlabel metal2 s 675407 335527 675887 335583 6 mprj_io_analog_sel[5]
port 259 nsew
rlabel metal2 s 675407 331847 675887 331903 6 mprj_io_dm[15]
port 260 nsew
rlabel metal2 s 675407 330007 675887 330063 6 mprj_io_dm[16]
port 261 nsew
rlabel metal2 s 675407 336171 675887 336227 6 mprj_io_dm[17]
port 262 nsew
rlabel metal2 s 675407 334331 675887 334387 6 mprj_io_enh[5]
port 263 nsew
rlabel metal2 s 675407 334975 675887 335031 6 mprj_io_hldh_n[5]
port 264 nsew
rlabel metal2 s 675407 336815 675887 336871 6 mprj_io_holdover[5]
port 265 nsew
rlabel metal2 s 675407 339851 675887 339907 6 mprj_io_ib_mode_sel[5]
port 266 nsew
rlabel metal2 s 675407 333043 675887 333099 6 mprj_io_inp_dis[5]
port 267 nsew
rlabel metal2 s 675407 340495 675887 340551 6 mprj_io_oeb[5]
port 268 nsew
rlabel metal2 s 675407 337367 675887 337423 6 mprj_io_out[5]
port 269 nsew
rlabel metal2 s 675407 328167 675887 328223 6 mprj_io_slow_sel[5]
port 270 nsew
rlabel metal2 s 675407 339207 675887 339263 6 mprj_io_vtrip_sel[5]
port 271 nsew
rlabel metal2 s 675407 326327 675887 326383 6 mprj_io_in[5]
port 272 nsew
rlabel metal5 s 698512 371840 711002 384360 6 mprj_io[6]
port 273 nsew
rlabel metal2 s 675407 376403 675887 376459 6 mprj_io_analog_en[6]
port 274 nsew
rlabel metal2 s 675407 377691 675887 377747 6 mprj_io_analog_pol[6]
port 275 nsew
rlabel metal2 s 675407 380727 675887 380783 6 mprj_io_analog_sel[6]
port 276 nsew
rlabel metal2 s 675407 377047 675887 377103 6 mprj_io_dm[18]
port 277 nsew
rlabel metal2 s 675407 375207 675887 375263 6 mprj_io_dm[19]
port 278 nsew
rlabel metal2 s 675407 381371 675887 381427 6 mprj_io_dm[20]
port 279 nsew
rlabel metal2 s 675407 379531 675887 379587 6 mprj_io_enh[6]
port 280 nsew
rlabel metal2 s 675407 380175 675887 380231 6 mprj_io_hldh_n[6]
port 281 nsew
rlabel metal2 s 675407 382015 675887 382071 6 mprj_io_holdover[6]
port 282 nsew
rlabel metal2 s 675407 385051 675887 385107 6 mprj_io_ib_mode_sel[6]
port 283 nsew
rlabel metal2 s 675407 378243 675887 378299 6 mprj_io_inp_dis[6]
port 284 nsew
rlabel metal2 s 675407 385695 675887 385751 6 mprj_io_oeb[6]
port 285 nsew
rlabel metal2 s 675407 382567 675887 382623 6 mprj_io_out[6]
port 286 nsew
rlabel metal2 s 675407 373367 675887 373423 6 mprj_io_slow_sel[6]
port 287 nsew
rlabel metal2 s 675407 384407 675887 384463 6 mprj_io_vtrip_sel[6]
port 288 nsew
rlabel metal2 s 675407 371527 675887 371583 6 mprj_io_in[6]
port 289 nsew
rlabel metal5 s 698512 549040 711002 561560 6 mprj_io[7]
port 290 nsew
rlabel metal2 s 675407 553603 675887 553659 6 mprj_io_analog_en[7]
port 291 nsew
rlabel metal2 s 675407 554891 675887 554947 6 mprj_io_analog_pol[7]
port 292 nsew
rlabel metal2 s 675407 557927 675887 557983 6 mprj_io_analog_sel[7]
port 293 nsew
rlabel metal2 s 675407 554247 675887 554303 6 mprj_io_dm[21]
port 294 nsew
rlabel metal2 s 675407 552407 675887 552463 6 mprj_io_dm[22]
port 295 nsew
rlabel metal2 s 675407 558571 675887 558627 6 mprj_io_dm[23]
port 296 nsew
rlabel metal2 s 675407 556731 675887 556787 6 mprj_io_enh[7]
port 297 nsew
rlabel metal2 s 675407 557375 675887 557431 6 mprj_io_hldh_n[7]
port 298 nsew
rlabel metal2 s 675407 559215 675887 559271 6 mprj_io_holdover[7]
port 299 nsew
rlabel metal2 s 675407 562251 675887 562307 6 mprj_io_ib_mode_sel[7]
port 300 nsew
rlabel metal2 s 675407 555443 675887 555499 6 mprj_io_inp_dis[7]
port 301 nsew
rlabel metal2 s 675407 562895 675887 562951 6 mprj_io_oeb[7]
port 302 nsew
rlabel metal2 s 675407 559767 675887 559823 6 mprj_io_out[7]
port 303 nsew
rlabel metal2 s 675407 550567 675887 550623 6 mprj_io_slow_sel[7]
port 304 nsew
rlabel metal2 s 675407 561607 675887 561663 6 mprj_io_vtrip_sel[7]
port 305 nsew
rlabel metal2 s 675407 548727 675887 548783 6 mprj_io_in[7]
port 306 nsew
rlabel metal5 s 698512 594240 711002 606760 6 mprj_io[8]
port 307 nsew
rlabel metal2 s 675407 598803 675887 598859 6 mprj_io_analog_en[8]
port 308 nsew
rlabel metal2 s 675407 600091 675887 600147 6 mprj_io_analog_pol[8]
port 309 nsew
rlabel metal2 s 675407 603127 675887 603183 6 mprj_io_analog_sel[8]
port 310 nsew
rlabel metal2 s 675407 599447 675887 599503 6 mprj_io_dm[24]
port 311 nsew
rlabel metal2 s 675407 597607 675887 597663 6 mprj_io_dm[25]
port 312 nsew
rlabel metal2 s 675407 603771 675887 603827 6 mprj_io_dm[26]
port 313 nsew
rlabel metal2 s 675407 601931 675887 601987 6 mprj_io_enh[8]
port 314 nsew
rlabel metal2 s 675407 602575 675887 602631 6 mprj_io_hldh_n[8]
port 315 nsew
rlabel metal2 s 675407 604415 675887 604471 6 mprj_io_holdover[8]
port 316 nsew
rlabel metal2 s 675407 607451 675887 607507 6 mprj_io_ib_mode_sel[8]
port 317 nsew
rlabel metal2 s 675407 600643 675887 600699 6 mprj_io_inp_dis[8]
port 318 nsew
rlabel metal2 s 675407 608095 675887 608151 6 mprj_io_oeb[8]
port 319 nsew
rlabel metal2 s 675407 604967 675887 605023 6 mprj_io_out[8]
port 320 nsew
rlabel metal2 s 675407 595767 675887 595823 6 mprj_io_slow_sel[8]
port 321 nsew
rlabel metal2 s 675407 606807 675887 606863 6 mprj_io_vtrip_sel[8]
port 322 nsew
rlabel metal2 s 675407 593927 675887 593983 6 mprj_io_in[8]
port 323 nsew
rlabel metal5 s 698512 639240 711002 651760 6 mprj_io[9]
port 324 nsew
rlabel metal2 s 675407 643803 675887 643859 6 mprj_io_analog_en[9]
port 325 nsew
rlabel metal2 s 675407 645091 675887 645147 6 mprj_io_analog_pol[9]
port 326 nsew
rlabel metal2 s 675407 648127 675887 648183 6 mprj_io_analog_sel[9]
port 327 nsew
rlabel metal2 s 675407 644447 675887 644503 6 mprj_io_dm[27]
port 328 nsew
rlabel metal2 s 675407 642607 675887 642663 6 mprj_io_dm[28]
port 329 nsew
rlabel metal2 s 675407 648771 675887 648827 6 mprj_io_dm[29]
port 330 nsew
rlabel metal2 s 675407 646931 675887 646987 6 mprj_io_enh[9]
port 331 nsew
rlabel metal2 s 675407 647575 675887 647631 6 mprj_io_hldh_n[9]
port 332 nsew
rlabel metal2 s 675407 649415 675887 649471 6 mprj_io_holdover[9]
port 333 nsew
rlabel metal2 s 675407 652451 675887 652507 6 mprj_io_ib_mode_sel[9]
port 334 nsew
rlabel metal2 s 675407 645643 675887 645699 6 mprj_io_inp_dis[9]
port 335 nsew
rlabel metal2 s 675407 653095 675887 653151 6 mprj_io_oeb[9]
port 336 nsew
rlabel metal2 s 675407 649967 675887 650023 6 mprj_io_out[9]
port 337 nsew
rlabel metal2 s 675407 640767 675887 640823 6 mprj_io_slow_sel[9]
port 338 nsew
rlabel metal2 s 675407 651807 675887 651863 6 mprj_io_vtrip_sel[9]
port 339 nsew
rlabel metal2 s 675407 638927 675887 638983 6 mprj_io_in[9]
port 340 nsew
rlabel metal5 s 386040 1018512 398560 1031002 6 mprj_io[18]
port 341 nsew
rlabel metal2 s 393941 995407 393997 995887 6 mprj_io_analog_en[18]
port 342 nsew
rlabel metal2 s 392653 995407 392709 995887 6 mprj_io_analog_pol[18]
port 343 nsew
rlabel metal2 s 389617 995407 389673 995887 6 mprj_io_analog_sel[18]
port 344 nsew
rlabel metal2 s 393297 995407 393353 995887 6 mprj_io_dm[54]
port 345 nsew
rlabel metal2 s 395137 995407 395193 995887 6 mprj_io_dm[55]
port 346 nsew
rlabel metal2 s 388973 995407 389029 995887 6 mprj_io_dm[56]
port 347 nsew
rlabel metal2 s 390813 995407 390869 995887 6 mprj_io_enh[18]
port 348 nsew
rlabel metal2 s 390169 995407 390225 995887 6 mprj_io_hldh_n[18]
port 349 nsew
rlabel metal2 s 388329 995407 388385 995887 6 mprj_io_holdover[18]
port 350 nsew
rlabel metal2 s 385293 995407 385349 995887 6 mprj_io_ib_mode_sel[18]
port 351 nsew
rlabel metal2 s 392101 995407 392157 995887 6 mprj_io_inp_dis[18]
port 352 nsew
rlabel metal2 s 384649 995407 384705 995887 6 mprj_io_oeb[18]
port 353 nsew
rlabel metal2 s 387777 995407 387833 995887 6 mprj_io_out[18]
port 354 nsew
rlabel metal2 s 396977 995407 397033 995887 6 mprj_io_slow_sel[18]
port 355 nsew
rlabel metal2 s 385937 995407 385993 995887 6 mprj_io_vtrip_sel[18]
port 356 nsew
rlabel metal2 s 398817 995407 398873 995887 6 mprj_io_in[18]
port 357 nsew
rlabel metal5 s 6598 657040 19088 669560 6 mprj_io[28]
port 358 nsew
rlabel metal2 s 41713 664941 42193 664997 6 mprj_io_analog_en[28]
port 359 nsew
rlabel metal2 s 41713 663653 42193 663709 6 mprj_io_analog_pol[28]
port 360 nsew
rlabel metal2 s 41713 660617 42193 660673 6 mprj_io_analog_sel[28]
port 361 nsew
rlabel metal2 s 41713 664297 42193 664353 6 mprj_io_dm[84]
port 362 nsew
rlabel metal2 s 41713 666137 42193 666193 6 mprj_io_dm[85]
port 363 nsew
rlabel metal2 s 41713 659973 42193 660029 6 mprj_io_dm[86]
port 364 nsew
rlabel metal2 s 41713 661813 42193 661869 6 mprj_io_enh[28]
port 365 nsew
rlabel metal2 s 41713 661169 42193 661225 6 mprj_io_hldh_n[28]
port 366 nsew
rlabel metal2 s 41713 659329 42193 659385 6 mprj_io_holdover[28]
port 367 nsew
rlabel metal2 s 41713 656293 42193 656349 6 mprj_io_ib_mode_sel[28]
port 368 nsew
rlabel metal2 s 41713 663101 42193 663157 6 mprj_io_inp_dis[28]
port 369 nsew
rlabel metal2 s 41713 655649 42193 655705 6 mprj_io_oeb[28]
port 370 nsew
rlabel metal2 s 41713 658777 42193 658833 6 mprj_io_out[28]
port 371 nsew
rlabel metal2 s 41713 667977 42193 668033 6 mprj_io_slow_sel[28]
port 372 nsew
rlabel metal2 s 41713 656937 42193 656993 6 mprj_io_vtrip_sel[28]
port 373 nsew
rlabel metal2 s 41713 669817 42193 669873 6 mprj_io_in[28]
port 374 nsew
rlabel metal5 s 6598 613840 19088 626360 6 mprj_io[29]
port 375 nsew
rlabel metal2 s 41713 621741 42193 621797 6 mprj_io_analog_en[29]
port 376 nsew
rlabel metal2 s 41713 620453 42193 620509 6 mprj_io_analog_pol[29]
port 377 nsew
rlabel metal2 s 41713 617417 42193 617473 6 mprj_io_analog_sel[29]
port 378 nsew
rlabel metal2 s 41713 621097 42193 621153 6 mprj_io_dm[87]
port 379 nsew
rlabel metal2 s 41713 622937 42193 622993 6 mprj_io_dm[88]
port 380 nsew
rlabel metal2 s 41713 616773 42193 616829 6 mprj_io_dm[89]
port 381 nsew
rlabel metal2 s 41713 618613 42193 618669 6 mprj_io_enh[29]
port 382 nsew
rlabel metal2 s 41713 617969 42193 618025 6 mprj_io_hldh_n[29]
port 383 nsew
rlabel metal2 s 41713 616129 42193 616185 6 mprj_io_holdover[29]
port 384 nsew
rlabel metal2 s 41713 613093 42193 613149 6 mprj_io_ib_mode_sel[29]
port 385 nsew
rlabel metal2 s 41713 619901 42193 619957 6 mprj_io_inp_dis[29]
port 386 nsew
rlabel metal2 s 41713 612449 42193 612505 6 mprj_io_oeb[29]
port 387 nsew
rlabel metal2 s 41713 615577 42193 615633 6 mprj_io_out[29]
port 388 nsew
rlabel metal2 s 41713 624777 42193 624833 6 mprj_io_slow_sel[29]
port 389 nsew
rlabel metal2 s 41713 613737 42193 613793 6 mprj_io_vtrip_sel[29]
port 390 nsew
rlabel metal2 s 41713 626617 42193 626673 6 mprj_io_in[29]
port 391 nsew
rlabel metal5 s 6598 570640 19088 583160 6 mprj_io[30]
port 392 nsew
rlabel metal2 s 41713 578541 42193 578597 6 mprj_io_analog_en[30]
port 393 nsew
rlabel metal2 s 41713 577253 42193 577309 6 mprj_io_analog_pol[30]
port 394 nsew
rlabel metal2 s 41713 574217 42193 574273 6 mprj_io_analog_sel[30]
port 395 nsew
rlabel metal2 s 41713 577897 42193 577953 6 mprj_io_dm[90]
port 396 nsew
rlabel metal2 s 41713 579737 42193 579793 6 mprj_io_dm[91]
port 397 nsew
rlabel metal2 s 41713 573573 42193 573629 6 mprj_io_dm[92]
port 398 nsew
rlabel metal2 s 41713 575413 42193 575469 6 mprj_io_enh[30]
port 399 nsew
rlabel metal2 s 41713 574769 42193 574825 6 mprj_io_hldh_n[30]
port 400 nsew
rlabel metal2 s 41713 572929 42193 572985 6 mprj_io_holdover[30]
port 401 nsew
rlabel metal2 s 41713 569893 42193 569949 6 mprj_io_ib_mode_sel[30]
port 402 nsew
rlabel metal2 s 41713 576701 42193 576757 6 mprj_io_inp_dis[30]
port 403 nsew
rlabel metal2 s 41713 569249 42193 569305 6 mprj_io_oeb[30]
port 404 nsew
rlabel metal2 s 41713 572377 42193 572433 6 mprj_io_out[30]
port 405 nsew
rlabel metal2 s 41713 581577 42193 581633 6 mprj_io_slow_sel[30]
port 406 nsew
rlabel metal2 s 41713 570537 42193 570593 6 mprj_io_vtrip_sel[30]
port 407 nsew
rlabel metal2 s 41713 583417 42193 583473 6 mprj_io_in[30]
port 408 nsew
rlabel metal5 s 6598 527440 19088 539960 6 mprj_io[31]
port 409 nsew
rlabel metal2 s 41713 535341 42193 535397 6 mprj_io_analog_en[31]
port 410 nsew
rlabel metal2 s 41713 534053 42193 534109 6 mprj_io_analog_pol[31]
port 411 nsew
rlabel metal2 s 41713 531017 42193 531073 6 mprj_io_analog_sel[31]
port 412 nsew
rlabel metal2 s 41713 534697 42193 534753 6 mprj_io_dm[93]
port 413 nsew
rlabel metal2 s 41713 536537 42193 536593 6 mprj_io_dm[94]
port 414 nsew
rlabel metal2 s 41713 530373 42193 530429 6 mprj_io_dm[95]
port 415 nsew
rlabel metal2 s 41713 532213 42193 532269 6 mprj_io_enh[31]
port 416 nsew
rlabel metal2 s 41713 531569 42193 531625 6 mprj_io_hldh_n[31]
port 417 nsew
rlabel metal2 s 41713 529729 42193 529785 6 mprj_io_holdover[31]
port 418 nsew
rlabel metal2 s 41713 526693 42193 526749 6 mprj_io_ib_mode_sel[31]
port 419 nsew
rlabel metal2 s 41713 533501 42193 533557 6 mprj_io_inp_dis[31]
port 420 nsew
rlabel metal2 s 41713 526049 42193 526105 6 mprj_io_oeb[31]
port 421 nsew
rlabel metal2 s 41713 529177 42193 529233 6 mprj_io_out[31]
port 422 nsew
rlabel metal2 s 41713 538377 42193 538433 6 mprj_io_slow_sel[31]
port 423 nsew
rlabel metal2 s 41713 527337 42193 527393 6 mprj_io_vtrip_sel[31]
port 424 nsew
rlabel metal2 s 41713 540217 42193 540273 6 mprj_io_in[31]
port 425 nsew
rlabel metal5 s 6598 399840 19088 412360 6 mprj_io[32]
port 426 nsew
rlabel metal2 s 41713 407741 42193 407797 6 mprj_io_analog_en[32]
port 427 nsew
rlabel metal2 s 41713 406453 42193 406509 6 mprj_io_analog_pol[32]
port 428 nsew
rlabel metal2 s 41713 403417 42193 403473 6 mprj_io_analog_sel[32]
port 429 nsew
rlabel metal2 s 41713 407097 42193 407153 6 mprj_io_dm[96]
port 430 nsew
rlabel metal2 s 41713 408937 42193 408993 6 mprj_io_dm[97]
port 431 nsew
rlabel metal2 s 41713 402773 42193 402829 6 mprj_io_dm[98]
port 432 nsew
rlabel metal2 s 41713 404613 42193 404669 6 mprj_io_enh[32]
port 433 nsew
rlabel metal2 s 41713 403969 42193 404025 6 mprj_io_hldh_n[32]
port 434 nsew
rlabel metal2 s 41713 402129 42193 402185 6 mprj_io_holdover[32]
port 435 nsew
rlabel metal2 s 41713 399093 42193 399149 6 mprj_io_ib_mode_sel[32]
port 436 nsew
rlabel metal2 s 41713 405901 42193 405957 6 mprj_io_inp_dis[32]
port 437 nsew
rlabel metal2 s 41713 398449 42193 398505 6 mprj_io_oeb[32]
port 438 nsew
rlabel metal2 s 41713 401577 42193 401633 6 mprj_io_out[32]
port 439 nsew
rlabel metal2 s 41713 410777 42193 410833 6 mprj_io_slow_sel[32]
port 440 nsew
rlabel metal2 s 41713 399737 42193 399793 6 mprj_io_vtrip_sel[32]
port 441 nsew
rlabel metal2 s 41713 412617 42193 412673 6 mprj_io_in[32]
port 442 nsew
rlabel metal5 s 6598 356640 19088 369160 6 mprj_io[33]
port 443 nsew
rlabel metal2 s 41713 364541 42193 364597 6 mprj_io_analog_en[33]
port 444 nsew
rlabel metal2 s 41713 363253 42193 363309 6 mprj_io_analog_pol[33]
port 445 nsew
rlabel metal2 s 41713 360217 42193 360273 6 mprj_io_analog_sel[33]
port 446 nsew
rlabel metal2 s 41713 365737 42193 365793 6 mprj_io_dm[100]
port 447 nsew
rlabel metal2 s 41713 359573 42193 359629 6 mprj_io_dm[101]
port 448 nsew
rlabel metal2 s 41713 363897 42193 363953 6 mprj_io_dm[99]
port 449 nsew
rlabel metal2 s 41713 361413 42193 361469 6 mprj_io_enh[33]
port 450 nsew
rlabel metal2 s 41713 360769 42193 360825 6 mprj_io_hldh_n[33]
port 451 nsew
rlabel metal2 s 41713 358929 42193 358985 6 mprj_io_holdover[33]
port 452 nsew
rlabel metal2 s 41713 355893 42193 355949 6 mprj_io_ib_mode_sel[33]
port 453 nsew
rlabel metal2 s 41713 362701 42193 362757 6 mprj_io_inp_dis[33]
port 454 nsew
rlabel metal2 s 41713 355249 42193 355305 6 mprj_io_oeb[33]
port 455 nsew
rlabel metal2 s 41713 358377 42193 358433 6 mprj_io_out[33]
port 456 nsew
rlabel metal2 s 41713 367577 42193 367633 6 mprj_io_slow_sel[33]
port 457 nsew
rlabel metal2 s 41713 356537 42193 356593 6 mprj_io_vtrip_sel[33]
port 458 nsew
rlabel metal2 s 41713 369417 42193 369473 6 mprj_io_in[33]
port 459 nsew
rlabel metal5 s 6598 313440 19088 325960 6 mprj_io[34]
port 460 nsew
rlabel metal2 s 41713 321341 42193 321397 6 mprj_io_analog_en[34]
port 461 nsew
rlabel metal2 s 41713 320053 42193 320109 6 mprj_io_analog_pol[34]
port 462 nsew
rlabel metal2 s 41713 317017 42193 317073 6 mprj_io_analog_sel[34]
port 463 nsew
rlabel metal2 s 41713 320697 42193 320753 6 mprj_io_dm[102]
port 464 nsew
rlabel metal2 s 41713 322537 42193 322593 6 mprj_io_dm[103]
port 465 nsew
rlabel metal2 s 41713 316373 42193 316429 6 mprj_io_dm[104]
port 466 nsew
rlabel metal2 s 41713 318213 42193 318269 6 mprj_io_enh[34]
port 467 nsew
rlabel metal2 s 41713 317569 42193 317625 6 mprj_io_hldh_n[34]
port 468 nsew
rlabel metal2 s 41713 315729 42193 315785 6 mprj_io_holdover[34]
port 469 nsew
rlabel metal2 s 41713 312693 42193 312749 6 mprj_io_ib_mode_sel[34]
port 470 nsew
rlabel metal2 s 41713 319501 42193 319557 6 mprj_io_inp_dis[34]
port 471 nsew
rlabel metal2 s 41713 312049 42193 312105 6 mprj_io_oeb[34]
port 472 nsew
rlabel metal2 s 41713 315177 42193 315233 6 mprj_io_out[34]
port 473 nsew
rlabel metal2 s 41713 324377 42193 324433 6 mprj_io_slow_sel[34]
port 474 nsew
rlabel metal2 s 41713 313337 42193 313393 6 mprj_io_vtrip_sel[34]
port 475 nsew
rlabel metal2 s 41713 326217 42193 326273 6 mprj_io_in[34]
port 476 nsew
rlabel metal5 s 6598 270240 19088 282760 6 mprj_io[35]
port 477 nsew
rlabel metal2 s 41713 278141 42193 278197 6 mprj_io_analog_en[35]
port 478 nsew
rlabel metal2 s 41713 276853 42193 276909 6 mprj_io_analog_pol[35]
port 479 nsew
rlabel metal2 s 41713 273817 42193 273873 6 mprj_io_analog_sel[35]
port 480 nsew
rlabel metal2 s 41713 277497 42193 277553 6 mprj_io_dm[105]
port 481 nsew
rlabel metal2 s 41713 279337 42193 279393 6 mprj_io_dm[106]
port 482 nsew
rlabel metal2 s 41713 273173 42193 273229 6 mprj_io_dm[107]
port 483 nsew
rlabel metal2 s 41713 275013 42193 275069 6 mprj_io_enh[35]
port 484 nsew
rlabel metal2 s 41713 274369 42193 274425 6 mprj_io_hldh_n[35]
port 485 nsew
rlabel metal2 s 41713 272529 42193 272585 6 mprj_io_holdover[35]
port 486 nsew
rlabel metal2 s 41713 269493 42193 269549 6 mprj_io_ib_mode_sel[35]
port 487 nsew
rlabel metal2 s 41713 276301 42193 276357 6 mprj_io_inp_dis[35]
port 488 nsew
rlabel metal2 s 41713 268849 42193 268905 6 mprj_io_oeb[35]
port 489 nsew
rlabel metal2 s 41713 271977 42193 272033 6 mprj_io_out[35]
port 490 nsew
rlabel metal2 s 41713 281177 42193 281233 6 mprj_io_slow_sel[35]
port 491 nsew
rlabel metal2 s 41713 270137 42193 270193 6 mprj_io_vtrip_sel[35]
port 492 nsew
rlabel metal2 s 41713 283017 42193 283073 6 mprj_io_in[35]
port 493 nsew
rlabel metal5 s 6598 227040 19088 239560 6 mprj_io[36]
port 494 nsew
rlabel metal2 s 41713 234941 42193 234997 6 mprj_io_analog_en[36]
port 495 nsew
rlabel metal2 s 41713 233653 42193 233709 6 mprj_io_analog_pol[36]
port 496 nsew
rlabel metal2 s 41713 230617 42193 230673 6 mprj_io_analog_sel[36]
port 497 nsew
rlabel metal2 s 41713 234297 42193 234353 6 mprj_io_dm[108]
port 498 nsew
rlabel metal2 s 41713 236137 42193 236193 6 mprj_io_dm[109]
port 499 nsew
rlabel metal2 s 41713 229973 42193 230029 6 mprj_io_dm[110]
port 500 nsew
rlabel metal2 s 41713 231813 42193 231869 6 mprj_io_enh[36]
port 501 nsew
rlabel metal2 s 41713 231169 42193 231225 6 mprj_io_hldh_n[36]
port 502 nsew
rlabel metal2 s 41713 229329 42193 229385 6 mprj_io_holdover[36]
port 503 nsew
rlabel metal2 s 41713 226293 42193 226349 6 mprj_io_ib_mode_sel[36]
port 504 nsew
rlabel metal2 s 41713 233101 42193 233157 6 mprj_io_inp_dis[36]
port 505 nsew
rlabel metal2 s 41713 225649 42193 225705 6 mprj_io_oeb[36]
port 506 nsew
rlabel metal2 s 41713 228777 42193 228833 6 mprj_io_out[36]
port 507 nsew
rlabel metal2 s 41713 237977 42193 238033 6 mprj_io_slow_sel[36]
port 508 nsew
rlabel metal2 s 41713 226937 42193 226993 6 mprj_io_vtrip_sel[36]
port 509 nsew
rlabel metal2 s 41713 239817 42193 239873 6 mprj_io_in[36]
port 510 nsew
rlabel metal5 s 6598 183840 19088 196360 6 mprj_io[37]
port 511 nsew
rlabel metal2 s 41713 191741 42193 191797 6 mprj_io_analog_en[37]
port 512 nsew
rlabel metal2 s 41713 190453 42193 190509 6 mprj_io_analog_pol[37]
port 513 nsew
rlabel metal2 s 41713 187417 42193 187473 6 mprj_io_analog_sel[37]
port 514 nsew
rlabel metal2 s 41713 191097 42193 191153 6 mprj_io_dm[111]
port 515 nsew
rlabel metal2 s 41713 192937 42193 192993 6 mprj_io_dm[112]
port 516 nsew
rlabel metal2 s 41713 186773 42193 186829 6 mprj_io_dm[113]
port 517 nsew
rlabel metal2 s 41713 188613 42193 188669 6 mprj_io_enh[37]
port 518 nsew
rlabel metal2 s 41713 187969 42193 188025 6 mprj_io_hldh_n[37]
port 519 nsew
rlabel metal2 s 41713 186129 42193 186185 6 mprj_io_holdover[37]
port 520 nsew
rlabel metal2 s 41713 183093 42193 183149 6 mprj_io_ib_mode_sel[37]
port 521 nsew
rlabel metal2 s 41713 189901 42193 189957 6 mprj_io_inp_dis[37]
port 522 nsew
rlabel metal2 s 41713 182449 42193 182505 6 mprj_io_oeb[37]
port 523 nsew
rlabel metal2 s 41713 185577 42193 185633 6 mprj_io_out[37]
port 524 nsew
rlabel metal2 s 41713 194777 42193 194833 6 mprj_io_slow_sel[37]
port 525 nsew
rlabel metal2 s 41713 183737 42193 183793 6 mprj_io_vtrip_sel[37]
port 526 nsew
rlabel metal2 s 41713 196617 42193 196673 6 mprj_io_in[37]
port 527 nsew
rlabel metal5 s 284240 1018512 296760 1031002 6 mprj_io[19]
port 528 nsew
rlabel metal2 s 292141 995407 292197 995887 6 mprj_io_analog_en[19]
port 529 nsew
rlabel metal2 s 290853 995407 290909 995887 6 mprj_io_analog_pol[19]
port 530 nsew
rlabel metal2 s 287817 995407 287873 995887 6 mprj_io_analog_sel[19]
port 531 nsew
rlabel metal2 s 291497 995407 291553 995887 6 mprj_io_dm[57]
port 532 nsew
rlabel metal2 s 293337 995407 293393 995887 6 mprj_io_dm[58]
port 533 nsew
rlabel metal2 s 287173 995407 287229 995887 6 mprj_io_dm[59]
port 534 nsew
rlabel metal2 s 289013 995407 289069 995887 6 mprj_io_enh[19]
port 535 nsew
rlabel metal2 s 288369 995407 288425 995887 6 mprj_io_hldh_n[19]
port 536 nsew
rlabel metal2 s 286529 995407 286585 995887 6 mprj_io_holdover[19]
port 537 nsew
rlabel metal2 s 283493 995407 283549 995887 6 mprj_io_ib_mode_sel[19]
port 538 nsew
rlabel metal2 s 290301 995407 290357 995887 6 mprj_io_inp_dis[19]
port 539 nsew
rlabel metal2 s 282849 995407 282905 995887 6 mprj_io_oeb[19]
port 540 nsew
rlabel metal2 s 285977 995407 286033 995887 6 mprj_io_out[19]
port 541 nsew
rlabel metal2 s 295177 995407 295233 995887 6 mprj_io_slow_sel[19]
port 542 nsew
rlabel metal2 s 284137 995407 284193 995887 6 mprj_io_vtrip_sel[19]
port 543 nsew
rlabel metal2 s 297017 995407 297073 995887 6 mprj_io_in[19]
port 544 nsew
rlabel metal5 s 232640 1018512 245160 1031002 6 mprj_io[20]
port 545 nsew
rlabel metal2 s 240541 995407 240597 995887 6 mprj_io_analog_en[20]
port 546 nsew
rlabel metal2 s 239253 995407 239309 995887 6 mprj_io_analog_pol[20]
port 547 nsew
rlabel metal2 s 236217 995407 236273 995887 6 mprj_io_analog_sel[20]
port 548 nsew
rlabel metal2 s 239897 995407 239953 995887 6 mprj_io_dm[60]
port 549 nsew
rlabel metal2 s 241737 995407 241793 995887 6 mprj_io_dm[61]
port 550 nsew
rlabel metal2 s 235573 995407 235629 995887 6 mprj_io_dm[62]
port 551 nsew
rlabel metal2 s 237413 995407 237469 995887 6 mprj_io_enh[20]
port 552 nsew
rlabel metal2 s 236769 995407 236825 995887 6 mprj_io_hldh_n[20]
port 553 nsew
rlabel metal2 s 234929 995407 234985 995887 6 mprj_io_holdover[20]
port 554 nsew
rlabel metal2 s 231893 995407 231949 995887 6 mprj_io_ib_mode_sel[20]
port 555 nsew
rlabel metal2 s 238701 995407 238757 995887 6 mprj_io_inp_dis[20]
port 556 nsew
rlabel metal2 s 231249 995407 231305 995887 6 mprj_io_oeb[20]
port 557 nsew
rlabel metal2 s 234377 995407 234433 995887 6 mprj_io_out[20]
port 558 nsew
rlabel metal2 s 243577 995407 243633 995887 6 mprj_io_slow_sel[20]
port 559 nsew
rlabel metal2 s 232537 995407 232593 995887 6 mprj_io_vtrip_sel[20]
port 560 nsew
rlabel metal2 s 245417 995407 245473 995887 6 mprj_io_in[20]
port 561 nsew
rlabel metal5 s 181240 1018512 193760 1031002 6 mprj_io[21]
port 562 nsew
rlabel metal2 s 189141 995407 189197 995887 6 mprj_io_analog_en[21]
port 563 nsew
rlabel metal2 s 187853 995407 187909 995887 6 mprj_io_analog_pol[21]
port 564 nsew
rlabel metal2 s 184817 995407 184873 995887 6 mprj_io_analog_sel[21]
port 565 nsew
rlabel metal2 s 188497 995407 188553 995887 6 mprj_io_dm[63]
port 566 nsew
rlabel metal2 s 190337 995407 190393 995887 6 mprj_io_dm[64]
port 567 nsew
rlabel metal2 s 184173 995407 184229 995887 6 mprj_io_dm[65]
port 568 nsew
rlabel metal2 s 186013 995407 186069 995887 6 mprj_io_enh[21]
port 569 nsew
rlabel metal2 s 185369 995407 185425 995887 6 mprj_io_hldh_n[21]
port 570 nsew
rlabel metal2 s 183529 995407 183585 995887 6 mprj_io_holdover[21]
port 571 nsew
rlabel metal2 s 180493 995407 180549 995887 6 mprj_io_ib_mode_sel[21]
port 572 nsew
rlabel metal2 s 187301 995407 187357 995887 6 mprj_io_inp_dis[21]
port 573 nsew
rlabel metal2 s 179849 995407 179905 995887 6 mprj_io_oeb[21]
port 574 nsew
rlabel metal2 s 182977 995407 183033 995887 6 mprj_io_out[21]
port 575 nsew
rlabel metal2 s 192177 995407 192233 995887 6 mprj_io_slow_sel[21]
port 576 nsew
rlabel metal2 s 181137 995407 181193 995887 6 mprj_io_vtrip_sel[21]
port 577 nsew
rlabel metal2 s 194017 995407 194073 995887 6 mprj_io_in[21]
port 578 nsew
rlabel metal5 s 129840 1018512 142360 1031002 6 mprj_io[22]
port 579 nsew
rlabel metal2 s 137741 995407 137797 995887 6 mprj_io_analog_en[22]
port 580 nsew
rlabel metal2 s 136453 995407 136509 995887 6 mprj_io_analog_pol[22]
port 581 nsew
rlabel metal2 s 133417 995407 133473 995887 6 mprj_io_analog_sel[22]
port 582 nsew
rlabel metal2 s 137097 995407 137153 995887 6 mprj_io_dm[66]
port 583 nsew
rlabel metal2 s 138937 995407 138993 995887 6 mprj_io_dm[67]
port 584 nsew
rlabel metal2 s 132773 995407 132829 995887 6 mprj_io_dm[68]
port 585 nsew
rlabel metal2 s 134613 995407 134669 995887 6 mprj_io_enh[22]
port 586 nsew
rlabel metal2 s 133969 995407 134025 995887 6 mprj_io_hldh_n[22]
port 587 nsew
rlabel metal2 s 132129 995407 132185 995887 6 mprj_io_holdover[22]
port 588 nsew
rlabel metal2 s 129093 995407 129149 995887 6 mprj_io_ib_mode_sel[22]
port 589 nsew
rlabel metal2 s 135901 995407 135957 995887 6 mprj_io_inp_dis[22]
port 590 nsew
rlabel metal2 s 128449 995407 128505 995887 6 mprj_io_oeb[22]
port 591 nsew
rlabel metal2 s 131577 995407 131633 995887 6 mprj_io_out[22]
port 592 nsew
rlabel metal2 s 140777 995407 140833 995887 6 mprj_io_slow_sel[22]
port 593 nsew
rlabel metal2 s 129737 995407 129793 995887 6 mprj_io_vtrip_sel[22]
port 594 nsew
rlabel metal2 s 142617 995407 142673 995887 6 mprj_io_in[22]
port 595 nsew
rlabel metal5 s 78440 1018512 90960 1031002 6 mprj_io[23]
port 596 nsew
rlabel metal2 s 86341 995407 86397 995887 6 mprj_io_analog_en[23]
port 597 nsew
rlabel metal2 s 85053 995407 85109 995887 6 mprj_io_analog_pol[23]
port 598 nsew
rlabel metal2 s 82017 995407 82073 995887 6 mprj_io_analog_sel[23]
port 599 nsew
rlabel metal2 s 85697 995407 85753 995887 6 mprj_io_dm[69]
port 600 nsew
rlabel metal2 s 87537 995407 87593 995887 6 mprj_io_dm[70]
port 601 nsew
rlabel metal2 s 81373 995407 81429 995887 6 mprj_io_dm[71]
port 602 nsew
rlabel metal2 s 83213 995407 83269 995887 6 mprj_io_enh[23]
port 603 nsew
rlabel metal2 s 82569 995407 82625 995887 6 mprj_io_hldh_n[23]
port 604 nsew
rlabel metal2 s 80729 995407 80785 995887 6 mprj_io_holdover[23]
port 605 nsew
rlabel metal2 s 77693 995407 77749 995887 6 mprj_io_ib_mode_sel[23]
port 606 nsew
rlabel metal2 s 84501 995407 84557 995887 6 mprj_io_inp_dis[23]
port 607 nsew
rlabel metal2 s 77049 995407 77105 995887 6 mprj_io_oeb[23]
port 608 nsew
rlabel metal2 s 80177 995407 80233 995887 6 mprj_io_out[23]
port 609 nsew
rlabel metal2 s 89377 995407 89433 995887 6 mprj_io_slow_sel[23]
port 610 nsew
rlabel metal2 s 78337 995407 78393 995887 6 mprj_io_vtrip_sel[23]
port 611 nsew
rlabel metal2 s 91217 995407 91273 995887 6 mprj_io_in[23]
port 612 nsew
rlabel metal5 s 6598 956440 19088 968960 6 mprj_io[24]
port 613 nsew
rlabel metal2 s 41713 964341 42193 964397 6 mprj_io_analog_en[24]
port 614 nsew
rlabel metal2 s 41713 963053 42193 963109 6 mprj_io_analog_pol[24]
port 615 nsew
rlabel metal2 s 41713 960017 42193 960073 6 mprj_io_analog_sel[24]
port 616 nsew
rlabel metal2 s 41713 963697 42193 963753 6 mprj_io_dm[72]
port 617 nsew
rlabel metal2 s 41713 965537 42193 965593 6 mprj_io_dm[73]
port 618 nsew
rlabel metal2 s 41713 959373 42193 959429 6 mprj_io_dm[74]
port 619 nsew
rlabel metal2 s 41713 961213 42193 961269 6 mprj_io_enh[24]
port 620 nsew
rlabel metal2 s 41713 960569 42193 960625 6 mprj_io_hldh_n[24]
port 621 nsew
rlabel metal2 s 41713 958729 42193 958785 6 mprj_io_holdover[24]
port 622 nsew
rlabel metal2 s 41713 955693 42193 955749 6 mprj_io_ib_mode_sel[24]
port 623 nsew
rlabel metal2 s 41713 962501 42193 962557 6 mprj_io_inp_dis[24]
port 624 nsew
rlabel metal2 s 41713 955049 42193 955105 6 mprj_io_oeb[24]
port 625 nsew
rlabel metal2 s 41713 958177 42193 958233 6 mprj_io_out[24]
port 626 nsew
rlabel metal2 s 41713 967377 42193 967433 6 mprj_io_slow_sel[24]
port 627 nsew
rlabel metal2 s 41713 956337 42193 956393 6 mprj_io_vtrip_sel[24]
port 628 nsew
rlabel metal2 s 41713 969217 42193 969273 6 mprj_io_in[24]
port 629 nsew
rlabel metal5 s 6598 786640 19088 799160 6 mprj_io[25]
port 630 nsew
rlabel metal2 s 41713 794541 42193 794597 6 mprj_io_analog_en[25]
port 631 nsew
rlabel metal2 s 41713 793253 42193 793309 6 mprj_io_analog_pol[25]
port 632 nsew
rlabel metal2 s 41713 790217 42193 790273 6 mprj_io_analog_sel[25]
port 633 nsew
rlabel metal2 s 41713 793897 42193 793953 6 mprj_io_dm[75]
port 634 nsew
rlabel metal2 s 41713 795737 42193 795793 6 mprj_io_dm[76]
port 635 nsew
rlabel metal2 s 41713 789573 42193 789629 6 mprj_io_dm[77]
port 636 nsew
rlabel metal2 s 41713 791413 42193 791469 6 mprj_io_enh[25]
port 637 nsew
rlabel metal2 s 41713 790769 42193 790825 6 mprj_io_hldh_n[25]
port 638 nsew
rlabel metal2 s 41713 788929 42193 788985 6 mprj_io_holdover[25]
port 639 nsew
rlabel metal2 s 41713 785893 42193 785949 6 mprj_io_ib_mode_sel[25]
port 640 nsew
rlabel metal2 s 41713 792701 42193 792757 6 mprj_io_inp_dis[25]
port 641 nsew
rlabel metal2 s 41713 785249 42193 785305 6 mprj_io_oeb[25]
port 642 nsew
rlabel metal2 s 41713 788377 42193 788433 6 mprj_io_out[25]
port 643 nsew
rlabel metal2 s 41713 797577 42193 797633 6 mprj_io_slow_sel[25]
port 644 nsew
rlabel metal2 s 41713 786537 42193 786593 6 mprj_io_vtrip_sel[25]
port 645 nsew
rlabel metal2 s 41713 799417 42193 799473 6 mprj_io_in[25]
port 646 nsew
rlabel metal5 s 6598 743440 19088 755960 6 mprj_io[26]
port 647 nsew
rlabel metal2 s 41713 751341 42193 751397 6 mprj_io_analog_en[26]
port 648 nsew
rlabel metal2 s 41713 750053 42193 750109 6 mprj_io_analog_pol[26]
port 649 nsew
rlabel metal2 s 41713 747017 42193 747073 6 mprj_io_analog_sel[26]
port 650 nsew
rlabel metal2 s 41713 750697 42193 750753 6 mprj_io_dm[78]
port 651 nsew
rlabel metal2 s 41713 752537 42193 752593 6 mprj_io_dm[79]
port 652 nsew
rlabel metal2 s 41713 746373 42193 746429 6 mprj_io_dm[80]
port 653 nsew
rlabel metal2 s 41713 748213 42193 748269 6 mprj_io_enh[26]
port 654 nsew
rlabel metal2 s 41713 747569 42193 747625 6 mprj_io_hldh_n[26]
port 655 nsew
rlabel metal2 s 41713 745729 42193 745785 6 mprj_io_holdover[26]
port 656 nsew
rlabel metal2 s 41713 742693 42193 742749 6 mprj_io_ib_mode_sel[26]
port 657 nsew
rlabel metal2 s 41713 749501 42193 749557 6 mprj_io_inp_dis[26]
port 658 nsew
rlabel metal2 s 41713 742049 42193 742105 6 mprj_io_oeb[26]
port 659 nsew
rlabel metal2 s 41713 745177 42193 745233 6 mprj_io_out[26]
port 660 nsew
rlabel metal2 s 41713 754377 42193 754433 6 mprj_io_slow_sel[26]
port 661 nsew
rlabel metal2 s 41713 743337 42193 743393 6 mprj_io_vtrip_sel[26]
port 662 nsew
rlabel metal2 s 41713 756217 42193 756273 6 mprj_io_in[26]
port 663 nsew
rlabel metal5 s 6598 700240 19088 712760 6 mprj_io[27]
port 664 nsew
rlabel metal2 s 41713 708141 42193 708197 6 mprj_io_analog_en[27]
port 665 nsew
rlabel metal2 s 41713 706853 42193 706909 6 mprj_io_analog_pol[27]
port 666 nsew
rlabel metal2 s 41713 703817 42193 703873 6 mprj_io_analog_sel[27]
port 667 nsew
rlabel metal2 s 41713 707497 42193 707553 6 mprj_io_dm[81]
port 668 nsew
rlabel metal2 s 41713 709337 42193 709393 6 mprj_io_dm[82]
port 669 nsew
rlabel metal2 s 41713 703173 42193 703229 6 mprj_io_dm[83]
port 670 nsew
rlabel metal2 s 41713 705013 42193 705069 6 mprj_io_enh[27]
port 671 nsew
rlabel metal2 s 41713 704369 42193 704425 6 mprj_io_hldh_n[27]
port 672 nsew
rlabel metal2 s 41713 702529 42193 702585 6 mprj_io_holdover[27]
port 673 nsew
rlabel metal2 s 41713 699493 42193 699549 6 mprj_io_ib_mode_sel[27]
port 674 nsew
rlabel metal2 s 41713 706301 42193 706357 6 mprj_io_inp_dis[27]
port 675 nsew
rlabel metal2 s 41713 698849 42193 698905 6 mprj_io_oeb[27]
port 676 nsew
rlabel metal2 s 41713 701977 42193 702033 6 mprj_io_out[27]
port 677 nsew
rlabel metal2 s 41713 711177 42193 711233 6 mprj_io_slow_sel[27]
port 678 nsew
rlabel metal2 s 41713 700137 42193 700193 6 mprj_io_vtrip_sel[27]
port 679 nsew
rlabel metal2 s 41713 713017 42193 713073 6 mprj_io_in[27]
port 680 nsew
rlabel metal3 s 675385 338675 675451 338678 6 porb_h
port 681 nsew
rlabel metal3 s 673545 338675 673611 338678 6 porb_h
port 681 nsew
rlabel metal3 s 673545 338678 675451 338738 6 porb_h
port 681 nsew
rlabel metal3 s 675385 338738 675451 338741 6 porb_h
port 681 nsew
rlabel metal3 s 673545 338738 673611 338741 6 porb_h
port 681 nsew
rlabel metal3 s 675293 888659 675359 888662 6 porb_h
port 681 nsew
rlabel metal3 s 673453 888659 673519 888662 6 porb_h
port 681 nsew
rlabel metal3 s 673453 888662 675359 888722 6 porb_h
port 681 nsew
rlabel metal3 s 675293 888722 675359 888725 6 porb_h
port 681 nsew
rlabel metal3 s 673453 888722 673519 888725 6 porb_h
port 681 nsew
rlabel metal3 s 173801 990659 173867 990662 6 porb_h
port 681 nsew
rlabel metal3 s 160093 990659 160159 990662 6 porb_h
port 681 nsew
rlabel metal3 s 160093 990662 173867 990722 6 porb_h
port 681 nsew
rlabel metal3 s 173801 990722 173867 990725 6 porb_h
port 681 nsew
rlabel metal3 s 160093 990722 160159 990725 6 porb_h
port 681 nsew
rlabel via2 s 675390 338680 675446 338736 6 porb_h
port 681 nsew
rlabel via2 s 673550 338680 673606 338736 6 porb_h
port 681 nsew
rlabel via2 s 675298 888664 675354 888720 6 porb_h
port 681 nsew
rlabel via2 s 673458 888664 673514 888720 6 porb_h
port 681 nsew
rlabel via2 s 173806 990664 173862 990720 6 porb_h
port 681 nsew
rlabel via2 s 160098 990664 160154 990720 6 porb_h
port 681 nsew
rlabel metal2 s 145091 39706 145143 40000 6 porb_h
port 681 nsew
rlabel metal2 s 145103 40000 145131 40174 6 porb_h
port 681 nsew
rlabel metal2 s 145103 40174 145144 40202 6 porb_h
port 681 nsew
rlabel metal2 s 527455 41713 527511 41942 6 porb_h
port 681 nsew
rlabel metal2 s 523131 41713 523187 41806 6 porb_h
port 681 nsew
rlabel metal2 s 523131 41806 523264 41834 6 porb_h
port 681 nsew
rlabel metal2 s 523236 41834 523264 41890 6 porb_h
port 681 nsew
rlabel metal2 s 527364 41890 527416 41942 6 porb_h
port 681 nsew
rlabel metal2 s 527364 41942 527511 41954 6 porb_h
port 681 nsew
rlabel metal2 s 523224 41890 523276 41954 6 porb_h
port 681 nsew
rlabel metal2 s 527376 41954 527511 41970 6 porb_h
port 681 nsew
rlabel metal2 s 527455 41970 527511 42193 6 porb_h
port 681 nsew
rlabel metal2 s 523131 41834 523187 42193 6 porb_h
port 681 nsew
rlabel metal2 s 472655 41713 472711 41806 6 porb_h
port 681 nsew
rlabel metal2 s 468331 41713 468387 41806 6 porb_h
port 681 nsew
rlabel metal2 s 472544 41806 472711 41822 6 porb_h
port 681 nsew
rlabel metal2 s 468312 41806 468524 41822 6 porb_h
port 681 nsew
rlabel metal2 s 417855 41713 417911 41820 6 porb_h
port 681 nsew
rlabel metal2 s 413531 41713 413587 41820 6 porb_h
port 681 nsew
rlabel metal2 s 472532 41822 472711 41834 6 porb_h
port 681 nsew
rlabel metal2 s 472655 41834 472711 42193 6 porb_h
port 681 nsew
rlabel metal2 s 472532 41834 472584 41886 6 porb_h
port 681 nsew
rlabel metal2 s 468312 41822 468536 41834 6 porb_h
port 681 nsew
rlabel metal2 s 468484 41834 468536 41886 6 porb_h
port 681 nsew
rlabel metal2 s 468312 41834 468387 42193 6 porb_h
port 681 nsew
rlabel metal2 s 527468 42193 527496 47126 6 porb_h
port 681 nsew
rlabel metal2 s 468312 42193 468340 47126 6 porb_h
port 681 nsew
rlabel metal2 s 417855 41820 417924 42193 6 porb_h
port 681 nsew
rlabel metal2 s 413531 41820 413600 42193 6 porb_h
port 681 nsew
rlabel metal2 s 363055 41713 363111 42193 6 porb_h
port 681 nsew
rlabel metal2 s 358731 41713 358787 42193 6 porb_h
port 681 nsew
rlabel metal2 s 308255 41713 308311 41806 6 porb_h
port 681 nsew
rlabel metal2 s 303931 41713 303987 41806 6 porb_h
port 681 nsew
rlabel metal2 s 199655 41713 199711 41806 6 porb_h
port 681 nsew
rlabel metal2 s 195331 41713 195387 41806 6 porb_h
port 681 nsew
rlabel metal2 s 308232 41806 308311 42193 6 porb_h
port 681 nsew
rlabel metal2 s 303908 41806 303987 42193 6 porb_h
port 681 nsew
rlabel metal2 s 199580 41806 199711 41822 6 porb_h
port 681 nsew
rlabel metal2 s 195331 41806 195468 41822 6 porb_h
port 681 nsew
rlabel metal2 s 199568 41822 199711 41834 6 porb_h
port 681 nsew
rlabel metal2 s 199655 41834 199711 42193 6 porb_h
port 681 nsew
rlabel metal2 s 199568 41834 199620 41886 6 porb_h
port 681 nsew
rlabel metal2 s 195331 41822 195480 41834 6 porb_h
port 681 nsew
rlabel metal2 s 195428 41834 195480 41886 6 porb_h
port 681 nsew
rlabel metal2 s 195331 41834 195387 42193 6 porb_h
port 681 nsew
rlabel metal2 s 417896 42193 417924 47058 6 porb_h
port 681 nsew
rlabel metal2 s 413572 42193 413600 47058 6 porb_h
port 681 nsew
rlabel metal2 s 363064 42193 363092 47058 6 porb_h
port 681 nsew
rlabel metal2 s 358740 42193 358768 47058 6 porb_h
port 681 nsew
rlabel metal2 s 308232 42193 308260 47058 6 porb_h
port 681 nsew
rlabel metal2 s 303908 42193 303936 47058 6 porb_h
port 681 nsew
rlabel metal2 s 417884 47058 417936 47122 6 porb_h
port 681 nsew
rlabel metal2 s 413560 47058 413612 47122 6 porb_h
port 681 nsew
rlabel metal2 s 363052 47058 363104 47122 6 porb_h
port 681 nsew
rlabel metal2 s 358728 47058 358780 47122 6 porb_h
port 681 nsew
rlabel metal2 s 308220 47058 308272 47122 6 porb_h
port 681 nsew
rlabel metal2 s 303896 47058 303948 47122 6 porb_h
port 681 nsew
rlabel metal2 s 527456 47126 527508 47190 6 porb_h
port 681 nsew
rlabel metal2 s 468300 47126 468352 47190 6 porb_h
port 681 nsew
rlabel metal2 s 527468 47190 527496 47806 6 porb_h
port 681 nsew
rlabel metal2 s 199672 42193 199700 47262 6 porb_h
port 681 nsew
rlabel metal2 s 195348 42193 195376 44202 6 porb_h
port 681 nsew
rlabel metal2 s 145116 40202 145144 44202 6 porb_h
port 681 nsew
rlabel metal2 s 195336 44202 195388 44266 6 porb_h
port 681 nsew
rlabel metal2 s 145104 44202 145156 44266 6 porb_h
port 681 nsew
rlabel metal2 s 145116 44266 145144 45630 6 porb_h
port 681 nsew
rlabel metal2 s 145104 45630 145156 45694 6 porb_h
port 681 nsew
rlabel metal2 s 42248 45630 42300 45694 6 porb_h
port 681 nsew
rlabel metal2 s 199660 47262 199712 47326 6 porb_h
port 681 nsew
rlabel metal2 s 673552 47806 673604 47870 6 porb_h
port 681 nsew
rlabel metal2 s 527456 47806 527508 47870 6 porb_h
port 681 nsew
rlabel metal2 s 673564 47870 673592 112746 6 porb_h
port 681 nsew
rlabel metal2 s 675392 112746 675444 112810 6 porb_h
port 681 nsew
rlabel metal2 s 673552 112746 673604 112810 6 porb_h
port 681 nsew
rlabel metal2 s 675404 112810 675432 113255 6 porb_h
port 681 nsew
rlabel metal2 s 675404 113255 675887 113283 6 porb_h
port 681 nsew
rlabel metal2 s 675407 113283 675887 113311 6 porb_h
port 681 nsew
rlabel metal2 s 673564 112810 673592 158306 6 porb_h
port 681 nsew
rlabel metal2 s 675392 158306 675444 158370 6 porb_h
port 681 nsew
rlabel metal2 s 673552 158306 673604 158370 6 porb_h
port 681 nsew
rlabel metal2 s 675404 158370 675432 158455 6 porb_h
port 681 nsew
rlabel metal2 s 675404 158455 675887 158508 6 porb_h
port 681 nsew
rlabel metal2 s 675407 158508 675887 158511 6 porb_h
port 681 nsew
rlabel metal2 s 675407 203455 675887 203483 6 porb_h
port 681 nsew
rlabel metal2 s 675404 203483 675887 203511 6 porb_h
port 681 nsew
rlabel metal2 s 675404 203511 675432 203866 6 porb_h
port 681 nsew
rlabel metal2 s 673564 158370 673592 203866 6 porb_h
port 681 nsew
rlabel metal2 s 42260 45694 42288 184198 6 porb_h
port 681 nsew
rlabel metal2 s 41892 184198 42288 184214 6 porb_h
port 681 nsew
rlabel metal2 s 42432 184214 42484 184278 6 porb_h
port 681 nsew
rlabel metal2 s 41892 184214 42300 184226 6 porb_h
port 681 nsew
rlabel metal2 s 42248 184226 42300 184278 6 porb_h
port 681 nsew
rlabel metal2 s 675392 203866 675444 203930 6 porb_h
port 681 nsew
rlabel metal2 s 673828 203866 673880 203930 6 porb_h
port 681 nsew
rlabel metal2 s 673552 203866 673604 203930 6 porb_h
port 681 nsew
rlabel metal2 s 673840 203930 673868 248134 6 porb_h
port 681 nsew
rlabel metal2 s 42444 184278 42472 228006 6 porb_h
port 681 nsew
rlabel metal2 s 42260 184278 42288 184309 6 porb_h
port 681 nsew
rlabel metal2 s 41892 184226 41920 184289 6 porb_h
port 681 nsew
rlabel metal2 s 41713 184289 42193 184345 6 porb_h
port 681 nsew
rlabel metal2 s 41713 227489 42193 227545 6 porb_h
port 681 nsew
rlabel metal2 s 41800 227545 41828 228006 6 porb_h
port 681 nsew
rlabel metal2 s 42708 228006 42760 228070 6 porb_h
port 681 nsew
rlabel metal2 s 42432 228006 42484 228070 6 porb_h
port 681 nsew
rlabel metal2 s 41788 228006 41840 228070 6 porb_h
port 681 nsew
rlabel metal2 s 42720 228070 42748 246978 6 porb_h
port 681 nsew
rlabel metal2 s 42708 246978 42760 247042 6 porb_h
port 681 nsew
rlabel metal2 s 42340 246978 42392 247042 6 porb_h
port 681 nsew
rlabel metal2 s 675392 248134 675444 248198 6 porb_h
port 681 nsew
rlabel metal2 s 673828 248134 673880 248198 6 porb_h
port 681 nsew
rlabel metal2 s 675404 248198 675432 248655 6 porb_h
port 681 nsew
rlabel metal2 s 675404 248655 675887 248676 6 porb_h
port 681 nsew
rlabel metal2 s 675407 248676 675887 248711 6 porb_h
port 681 nsew
rlabel metal2 s 673840 248198 673868 293150 6 porb_h
port 681 nsew
rlabel metal2 s 42352 247042 42380 270234 6 porb_h
port 681 nsew
rlabel metal2 s 42708 270234 42760 270298 6 porb_h
port 681 nsew
rlabel metal2 s 42340 270234 42392 270298 6 porb_h
port 681 nsew
rlabel metal2 s 41788 270234 41840 270298 6 porb_h
port 681 nsew
rlabel metal2 s 42720 270298 42748 281998 6 porb_h
port 681 nsew
rlabel metal2 s 41800 270298 41828 270689 6 porb_h
port 681 nsew
rlabel metal2 s 41713 270689 42193 270745 6 porb_h
port 681 nsew
rlabel metal2 s 42708 281998 42760 282062 6 porb_h
port 681 nsew
rlabel metal2 s 42708 282202 42760 282266 6 porb_h
port 681 nsew
rlabel metal2 s 675392 293150 675444 293214 6 porb_h
port 681 nsew
rlabel metal2 s 673828 293150 673880 293214 6 porb_h
port 681 nsew
rlabel metal2 s 675404 293214 675432 293655 6 porb_h
port 681 nsew
rlabel metal2 s 673840 293214 673868 293270 6 porb_h
port 681 nsew
rlabel metal2 s 673564 293270 673868 293298 6 porb_h
port 681 nsew
rlabel metal2 s 675404 293655 675887 293692 6 porb_h
port 681 nsew
rlabel metal2 s 675407 293692 675887 293711 6 porb_h
port 681 nsew
rlabel metal2 s 675407 338655 675887 338671 6 porb_h
port 681 nsew
rlabel metal2 s 673564 293298 673592 338671 6 porb_h
port 681 nsew
rlabel metal2 s 42720 282266 42748 307906 6 porb_h
port 681 nsew
rlabel metal2 s 42708 307906 42760 307970 6 porb_h
port 681 nsew
rlabel metal2 s 42432 307906 42484 307970 6 porb_h
port 681 nsew
rlabel metal2 s 42444 307970 42472 313754 6 porb_h
port 681 nsew
rlabel metal2 s 42432 313754 42484 313818 6 porb_h
port 681 nsew
rlabel metal2 s 41788 313754 41840 313818 6 porb_h
port 681 nsew
rlabel metal2 s 675390 338671 675887 338711 6 porb_h
port 681 nsew
rlabel metal2 s 675390 338711 675446 338745 6 porb_h
port 681 nsew
rlabel metal2 s 673550 338671 673606 338745 6 porb_h
port 681 nsew
rlabel metal2 s 675407 383855 675887 383860 6 porb_h
port 681 nsew
rlabel metal2 s 675404 383860 675887 383911 6 porb_h
port 681 nsew
rlabel metal2 s 675404 383911 675432 383998 6 porb_h
port 681 nsew
rlabel metal2 s 673564 338745 673592 383998 6 porb_h
port 681 nsew
rlabel metal2 s 42444 313818 42472 356662 6 porb_h
port 681 nsew
rlabel metal2 s 41800 313818 41828 313889 6 porb_h
port 681 nsew
rlabel metal2 s 41713 313889 42193 313945 6 porb_h
port 681 nsew
rlabel metal2 s 42432 356662 42484 356726 6 porb_h
port 681 nsew
rlabel metal2 s 41788 356662 41840 356726 6 porb_h
port 681 nsew
rlabel metal2 s 675392 383998 675444 384062 6 porb_h
port 681 nsew
rlabel metal2 s 673552 383998 673604 384062 6 porb_h
port 681 nsew
rlabel metal2 s 42444 356726 42472 400114 6 porb_h
port 681 nsew
rlabel metal2 s 41800 356726 41828 357089 6 porb_h
port 681 nsew
rlabel metal2 s 41713 357089 42193 357145 6 porb_h
port 681 nsew
rlabel metal2 s 42432 400114 42484 400178 6 porb_h
port 681 nsew
rlabel metal2 s 41972 400114 42024 400178 6 porb_h
port 681 nsew
rlabel metal2 s 42444 400178 42472 528430 6 porb_h
port 681 nsew
rlabel metal2 s 41984 400178 42012 400289 6 porb_h
port 681 nsew
rlabel metal2 s 41713 400289 42193 400345 6 porb_h
port 681 nsew
rlabel metal2 s 41713 527889 42193 527945 6 porb_h
port 681 nsew
rlabel metal2 s 41800 527945 41828 528430 6 porb_h
port 681 nsew
rlabel metal2 s 42616 528430 42668 528494 6 porb_h
port 681 nsew
rlabel metal2 s 42432 528430 42484 528494 6 porb_h
port 681 nsew
rlabel metal2 s 41788 528430 41840 528494 6 porb_h
port 681 nsew
rlabel metal2 s 675407 561055 675887 561068 6 porb_h
port 681 nsew
rlabel metal2 s 675404 561068 675887 561111 6 porb_h
port 681 nsew
rlabel metal2 s 675404 561111 675432 561478 6 porb_h
port 681 nsew
rlabel metal2 s 675392 561478 675444 561542 6 porb_h
port 681 nsew
rlabel metal2 s 673644 561478 673696 561542 6 porb_h
port 681 nsew
rlabel metal2 s 675407 606255 675887 606283 6 porb_h
port 681 nsew
rlabel metal2 s 675404 606283 675887 606311 6 porb_h
port 681 nsew
rlabel metal2 s 675404 606311 675432 606698 6 porb_h
port 681 nsew
rlabel metal2 s 673656 561542 673684 606698 6 porb_h
port 681 nsew
rlabel metal2 s 42628 528494 42656 571610 6 porb_h
port 681 nsew
rlabel metal2 s 41713 571089 42193 571145 6 porb_h
port 681 nsew
rlabel metal2 s 41722 571145 41828 571146 6 porb_h
port 681 nsew
rlabel metal2 s 41800 571146 41828 571610 6 porb_h
port 681 nsew
rlabel metal2 s 42616 571610 42668 571674 6 porb_h
port 681 nsew
rlabel metal2 s 41788 571610 41840 571674 6 porb_h
port 681 nsew
rlabel metal2 s 42628 571674 42656 584190 6 porb_h
port 681 nsew
rlabel metal2 s 42616 584190 42668 584254 6 porb_h
port 681 nsew
rlabel metal2 s 42248 584190 42300 584254 6 porb_h
port 681 nsew
rlabel metal2 s 675392 606698 675444 606762 6 porb_h
port 681 nsew
rlabel metal2 s 673644 606698 673696 606762 6 porb_h
port 681 nsew
rlabel metal2 s 675407 651255 675887 651283 6 porb_h
port 681 nsew
rlabel metal2 s 675404 651283 675887 651311 6 porb_h
port 681 nsew
rlabel metal2 s 675404 651311 675432 651714 6 porb_h
port 681 nsew
rlabel metal2 s 673656 606762 673684 651714 6 porb_h
port 681 nsew
rlabel metal2 s 42260 584254 42288 614450 6 porb_h
port 681 nsew
rlabel metal2 s 41713 614289 42193 614345 6 porb_h
port 681 nsew
rlabel metal2 s 41892 614345 41920 614450 6 porb_h
port 681 nsew
rlabel metal2 s 42616 614450 42668 614514 6 porb_h
port 681 nsew
rlabel metal2 s 42248 614450 42300 614514 6 porb_h
port 681 nsew
rlabel metal2 s 41880 614450 41932 614514 6 porb_h
port 681 nsew
rlabel metal2 s 42628 614514 42656 633218 6 porb_h
port 681 nsew
rlabel metal2 s 42616 633218 42668 633282 6 porb_h
port 681 nsew
rlabel metal2 s 42340 633218 42392 633282 6 porb_h
port 681 nsew
rlabel metal2 s 675392 651714 675444 651778 6 porb_h
port 681 nsew
rlabel metal2 s 673644 651714 673696 651778 6 porb_h
port 681 nsew
rlabel metal2 s 673656 651778 673684 695914 6 porb_h
port 681 nsew
rlabel metal2 s 42352 633282 42380 657086 6 porb_h
port 681 nsew
rlabel metal2 s 42616 657086 42668 657150 6 porb_h
port 681 nsew
rlabel metal2 s 42340 657086 42392 657150 6 porb_h
port 681 nsew
rlabel metal2 s 41788 657086 41840 657150 6 porb_h
port 681 nsew
rlabel metal2 s 675392 695914 675444 695978 6 porb_h
port 681 nsew
rlabel metal2 s 673644 695914 673696 695978 6 porb_h
port 681 nsew
rlabel metal2 s 675404 695978 675432 696455 6 porb_h
port 681 nsew
rlabel metal2 s 675404 696455 675887 696469 6 porb_h
port 681 nsew
rlabel metal2 s 675312 696469 675887 696497 6 porb_h
port 681 nsew
rlabel metal2 s 675407 696497 675887 696511 6 porb_h
port 681 nsew
rlabel metal2 s 675312 696497 675340 710670 6 porb_h
port 681 nsew
rlabel metal2 s 42628 657150 42656 700810 6 porb_h
port 681 nsew
rlabel metal2 s 41800 657150 41828 657478 6 porb_h
port 681 nsew
rlabel metal2 s 41722 657478 41828 657489 6 porb_h
port 681 nsew
rlabel metal2 s 41713 657489 42193 657545 6 porb_h
port 681 nsew
rlabel metal2 s 41713 700689 42193 700745 6 porb_h
port 681 nsew
rlabel metal2 s 41722 700745 41828 700754 6 porb_h
port 681 nsew
rlabel metal2 s 41800 700754 41828 700810 6 porb_h
port 681 nsew
rlabel metal2 s 42616 700810 42668 700874 6 porb_h
port 681 nsew
rlabel metal2 s 41788 700810 41840 700874 6 porb_h
port 681 nsew
rlabel metal2 s 675300 710670 675352 710734 6 porb_h
port 681 nsew
rlabel metal2 s 674012 710670 674064 710734 6 porb_h
port 681 nsew
rlabel metal2 s 674024 710734 674052 720394 6 porb_h
port 681 nsew
rlabel metal2 s 674196 720394 674248 720458 6 porb_h
port 681 nsew
rlabel metal2 s 674012 720394 674064 720458 6 porb_h
port 681 nsew
rlabel metal2 s 675407 741455 675887 741483 6 porb_h
port 681 nsew
rlabel metal2 s 675404 741483 675887 741511 6 porb_h
port 681 nsew
rlabel metal2 s 675404 741511 675432 741882 6 porb_h
port 681 nsew
rlabel metal2 s 674208 720458 674236 741882 6 porb_h
port 681 nsew
rlabel metal2 s 675392 741882 675444 741946 6 porb_h
port 681 nsew
rlabel metal2 s 674196 741882 674248 741946 6 porb_h
port 681 nsew
rlabel metal2 s 673552 741882 673604 741946 6 porb_h
port 681 nsew
rlabel metal2 s 673564 741946 673592 768606 6 porb_h
port 681 nsew
rlabel metal2 s 42628 700874 42656 744398 6 porb_h
port 681 nsew
rlabel metal2 s 41713 743889 42193 743945 6 porb_h
port 681 nsew
rlabel metal2 s 41800 743945 41828 744398 6 porb_h
port 681 nsew
rlabel metal2 s 42616 744398 42668 744462 6 porb_h
port 681 nsew
rlabel metal2 s 41788 744398 41840 744462 6 porb_h
port 681 nsew
rlabel metal2 s 674012 768606 674064 768670 6 porb_h
port 681 nsew
rlabel metal2 s 673552 768606 673604 768670 6 porb_h
port 681 nsew
rlabel metal2 s 675312 786386 675340 786422 6 porb_h
port 681 nsew
rlabel metal2 s 674024 768670 674052 786422 6 porb_h
port 681 nsew
rlabel metal2 s 675407 786455 675887 786469 6 porb_h
port 681 nsew
rlabel metal2 s 675300 786422 675352 786469 6 porb_h
port 681 nsew
rlabel metal2 s 675300 786469 675887 786486 6 porb_h
port 681 nsew
rlabel metal2 s 674012 786422 674064 786486 6 porb_h
port 681 nsew
rlabel metal2 s 675312 786486 675887 786497 6 porb_h
port 681 nsew
rlabel metal2 s 675407 786497 675887 786511 6 porb_h
port 681 nsew
rlabel metal2 s 675312 786497 675340 797574 6 porb_h
port 681 nsew
rlabel metal2 s 42628 744462 42656 787170 6 porb_h
port 681 nsew
rlabel metal2 s 41722 787086 41828 787089 6 porb_h
port 681 nsew
rlabel metal2 s 42260 787139 42288 787170 6 porb_h
port 681 nsew
rlabel metal2 s 41713 787089 42193 787145 6 porb_h
port 681 nsew
rlabel metal2 s 42616 787170 42668 787234 6 porb_h
port 681 nsew
rlabel metal2 s 42248 787170 42300 787222 6 porb_h
port 681 nsew
rlabel metal2 s 41800 787145 41828 787222 6 porb_h
port 681 nsew
rlabel metal2 s 41800 787222 42300 787234 6 porb_h
port 681 nsew
rlabel metal2 s 41800 787234 42288 787250 6 porb_h
port 681 nsew
rlabel metal2 s 42260 787250 42288 788038 6 porb_h
port 681 nsew
rlabel metal2 s 42260 788038 42472 788066 6 porb_h
port 681 nsew
rlabel metal2 s 675300 797574 675352 797638 6 porb_h
port 681 nsew
rlabel metal2 s 674104 797574 674156 797638 6 porb_h
port 681 nsew
rlabel metal2 s 674116 797638 674144 821034 6 porb_h
port 681 nsew
rlabel metal2 s 674104 821034 674156 821098 6 porb_h
port 681 nsew
rlabel metal2 s 673552 821034 673604 821098 6 porb_h
port 681 nsew
rlabel metal2 s 673564 821098 673592 830758 6 porb_h
port 681 nsew
rlabel metal2 s 673644 830758 673696 830822 6 porb_h
port 681 nsew
rlabel metal2 s 673552 830758 673604 830822 6 porb_h
port 681 nsew
rlabel metal2 s 673656 830822 673684 836198 6 porb_h
port 681 nsew
rlabel metal2 s 673644 836198 673696 836262 6 porb_h
port 681 nsew
rlabel metal2 s 673552 836266 673604 836330 6 porb_h
port 681 nsew
rlabel metal2 s 673564 836330 673592 850054 6 porb_h
port 681 nsew
rlabel metal2 s 673564 850054 673684 850082 6 porb_h
port 681 nsew
rlabel metal2 s 673656 850082 673684 855494 6 porb_h
port 681 nsew
rlabel metal2 s 673656 855494 673776 855522 6 porb_h
port 681 nsew
rlabel metal2 s 673748 855522 673776 869382 6 porb_h
port 681 nsew
rlabel metal2 s 675208 869382 675260 869446 6 porb_h
port 681 nsew
rlabel metal2 s 673736 869382 673788 869446 6 porb_h
port 681 nsew
rlabel metal2 s 675407 875655 675887 875669 6 porb_h
port 681 nsew
rlabel metal2 s 675220 869446 675248 875669 6 porb_h
port 681 nsew
rlabel metal2 s 675220 875669 675887 875697 6 porb_h
port 681 nsew
rlabel metal2 s 675407 875697 675887 875711 6 porb_h
port 681 nsew
rlabel metal2 s 675312 875697 675340 888655 6 porb_h
port 681 nsew
rlabel metal2 s 675298 888655 675354 888729 6 porb_h
port 681 nsew
rlabel metal2 s 673458 888655 673514 888729 6 porb_h
port 681 nsew
rlabel metal2 s 673472 888729 673500 888762 6 porb_h
port 681 nsew
rlabel metal2 s 673460 888762 673512 888826 6 porb_h
port 681 nsew
rlabel metal2 s 673184 888762 673236 888826 6 porb_h
port 681 nsew
rlabel metal2 s 673196 888826 673224 908006 6 porb_h
port 681 nsew
rlabel metal2 s 673460 908006 673512 908070 6 porb_h
port 681 nsew
rlabel metal2 s 673184 908006 673236 908070 6 porb_h
port 681 nsew
rlabel metal2 s 675407 964855 675887 964883 6 porb_h
port 681 nsew
rlabel metal2 s 675404 964883 675887 964911 6 porb_h
port 681 nsew
rlabel metal2 s 675404 964911 675432 965262 6 porb_h
port 681 nsew
rlabel metal2 s 673472 908070 673500 965262 6 porb_h
port 681 nsew
rlabel metal2 s 42444 788066 42472 956422 6 porb_h
port 681 nsew
rlabel metal2 s 42432 956422 42484 956486 6 porb_h
port 681 nsew
rlabel metal2 s 41788 956422 41840 956486 6 porb_h
port 681 nsew
rlabel metal2 s 675392 965262 675444 965326 6 porb_h
port 681 nsew
rlabel metal2 s 673460 965262 673512 965326 6 porb_h
port 681 nsew
rlabel metal2 s 673472 965326 673500 990014 6 porb_h
port 681 nsew
rlabel metal2 s 673460 990014 673512 990078 6 porb_h
port 681 nsew
rlabel metal2 s 42444 956486 42472 990082 6 porb_h
port 681 nsew
rlabel metal2 s 41800 956486 41828 956889 6 porb_h
port 681 nsew
rlabel metal2 s 41713 956889 42193 956945 6 porb_h
port 681 nsew
rlabel metal2 s 628656 990082 628708 990146 6 porb_h
port 681 nsew
rlabel metal2 s 79048 990082 79100 990146 6 porb_h
port 681 nsew
rlabel metal2 s 42432 990082 42484 990146 6 porb_h
port 681 nsew
rlabel metal2 s 628668 990146 628696 990694 6 porb_h
port 681 nsew
rlabel metal2 s 246948 990422 247000 990486 6 porb_h
port 681 nsew
rlabel metal2 s 233056 990422 233108 990486 6 porb_h
port 681 nsew
rlabel metal2 s 202880 990422 202932 990486 6 porb_h
port 681 nsew
rlabel metal2 s 187700 990422 187752 990486 6 porb_h
port 681 nsew
rlabel metal2 s 187608 990422 187660 990486 6 porb_h
port 681 nsew
rlabel metal2 s 181720 990422 181772 990486 6 porb_h
port 681 nsew
rlabel metal2 s 160100 990422 160152 990486 6 porb_h
port 681 nsew
rlabel metal2 s 143264 990422 143316 990486 6 porb_h
port 681 nsew
rlabel metal2 s 438688 990542 438808 990558 6 porb_h
port 681 nsew
rlabel metal2 s 286968 990490 287020 990554 6 porb_h
port 681 nsew
rlabel metal2 s 450268 990558 450320 990622 6 porb_h
port 681 nsew
rlabel metal2 s 438688 990558 438820 990570 6 porb_h
port 681 nsew
rlabel metal2 s 438768 990570 438820 990622 6 porb_h
port 681 nsew
rlabel metal2 s 628656 990694 628708 990758 6 porb_h
port 681 nsew
rlabel metal2 s 526904 990694 526956 990758 6 porb_h
port 681 nsew
rlabel metal2 s 482928 990694 482980 990758 6 porb_h
port 681 nsew
rlabel metal2 s 628668 990758 628696 995407 6 porb_h
port 681 nsew
rlabel metal2 s 526916 990758 526944 995407 6 porb_h
port 681 nsew
rlabel metal2 s 482940 990758 482968 992258 6 porb_h
port 681 nsew
rlabel metal2 s 463620 990814 463832 990830 6 porb_h
port 681 nsew
rlabel metal2 s 450280 990622 450308 990830 6 porb_h
port 681 nsew
rlabel metal2 s 438688 990570 438716 990830 6 porb_h
port 681 nsew
rlabel metal2 s 419540 990558 419592 990622 6 porb_h
port 681 nsew
rlabel metal2 s 386512 990558 386564 990622 6 porb_h
port 681 nsew
rlabel metal2 s 419552 990622 419580 990830 6 porb_h
port 681 nsew
rlabel metal2 s 463608 990830 463832 990842 6 porb_h
port 681 nsew
rlabel metal2 s 463804 990842 463832 992258 6 porb_h
port 681 nsew
rlabel metal2 s 463608 990842 463660 990894 6 porb_h
port 681 nsew
rlabel metal2 s 450268 990830 450320 990894 6 porb_h
port 681 nsew
rlabel metal2 s 438676 990830 438728 990894 6 porb_h
port 681 nsew
rlabel metal2 s 419540 990830 419592 990894 6 porb_h
port 681 nsew
rlabel metal2 s 482928 992258 482980 992322 6 porb_h
port 681 nsew
rlabel metal2 s 475476 992258 475528 992322 6 porb_h
port 681 nsew
rlabel metal2 s 463792 992258 463844 992322 6 porb_h
port 681 nsew
rlabel metal2 s 475488 992322 475516 995407 6 porb_h
port 681 nsew
rlabel metal2 s 628668 995407 628745 995466 6 porb_h
port 681 nsew
rlabel metal2 s 628689 995466 628745 995887 6 porb_h
port 681 nsew
rlabel metal2 s 526889 995407 526945 995887 6 porb_h
port 681 nsew
rlabel metal2 s 475488 995407 475545 995452 6 porb_h
port 681 nsew
rlabel metal2 s 386524 990622 386552 995407 6 porb_h
port 681 nsew
rlabel metal2 s 286980 990554 287008 990762 6 porb_h
port 681 nsew
rlabel metal2 s 246960 990486 246988 990762 6 porb_h
port 681 nsew
rlabel metal2 s 233068 990486 233096 990694 6 porb_h
port 681 nsew
rlabel metal2 s 202892 990486 202920 990694 6 porb_h
port 681 nsew
rlabel metal2 s 187712 990486 187740 990694 6 porb_h
port 681 nsew
rlabel metal2 s 187620 990486 187648 990694 6 porb_h
port 681 nsew
rlabel metal2 s 181732 990486 181760 990558 6 porb_h
port 681 nsew
rlabel metal2 s 181720 990558 181772 990622 6 porb_h
port 681 nsew
rlabel metal2 s 179328 990558 179380 990622 6 porb_h
port 681 nsew
rlabel metal2 s 233056 990694 233108 990758 6 porb_h
port 681 nsew
rlabel metal2 s 202880 990694 202932 990758 6 porb_h
port 681 nsew
rlabel metal2 s 187700 990694 187752 990758 6 porb_h
port 681 nsew
rlabel metal2 s 187608 990694 187660 990758 6 porb_h
port 681 nsew
rlabel metal2 s 286968 990762 287020 990826 6 porb_h
port 681 nsew
rlabel metal2 s 284668 990762 284720 990826 6 porb_h
port 681 nsew
rlabel metal2 s 246948 990762 247000 990826 6 porb_h
port 681 nsew
rlabel metal2 s 284680 990826 284708 995407 6 porb_h
port 681 nsew
rlabel metal2 s 233068 990758 233096 995407 6 porb_h
port 681 nsew
rlabel metal2 s 386489 995407 386552 995452 6 porb_h
port 681 nsew
rlabel metal2 s 475489 995452 475545 995887 6 porb_h
port 681 nsew
rlabel metal2 s 386489 995452 386545 995887 6 porb_h
port 681 nsew
rlabel metal2 s 284680 995407 284745 995452 6 porb_h
port 681 nsew
rlabel metal2 s 284689 995452 284745 995887 6 porb_h
port 681 nsew
rlabel metal2 s 233068 995407 233145 995466 6 porb_h
port 681 nsew
rlabel metal2 s 181732 990622 181760 995407 6 porb_h
port 681 nsew
rlabel metal2 s 179340 990622 179368 990762 6 porb_h
port 681 nsew
rlabel metal2 s 160112 990486 160140 990655 6 porb_h
port 681 nsew
rlabel metal2 s 173806 990655 173862 990729 6 porb_h
port 681 nsew
rlabel metal2 s 160098 990655 160154 990729 6 porb_h
port 681 nsew
rlabel metal2 s 173820 990729 173848 990762 6 porb_h
port 681 nsew
rlabel metal2 s 143276 990486 143304 990762 6 porb_h
port 681 nsew
rlabel metal2 s 130108 990558 130160 990622 6 porb_h
port 681 nsew
rlabel metal2 s 110512 990558 110564 990622 6 porb_h
port 681 nsew
rlabel metal2 s 130120 990622 130148 990762 6 porb_h
port 681 nsew
rlabel metal2 s 110524 990622 110552 990678 6 porb_h
port 681 nsew
rlabel metal2 s 110432 990678 110552 990706 6 porb_h
port 681 nsew
rlabel metal2 s 110432 990706 110460 990762 6 porb_h
port 681 nsew
rlabel metal2 s 79060 990146 79088 990762 6 porb_h
port 681 nsew
rlabel metal2 s 179328 990762 179380 990826 6 porb_h
port 681 nsew
rlabel metal2 s 173808 990762 173860 990826 6 porb_h
port 681 nsew
rlabel metal2 s 143264 990762 143316 990826 6 porb_h
port 681 nsew
rlabel metal2 s 130108 990762 130160 990826 6 porb_h
port 681 nsew
rlabel metal2 s 110420 990762 110472 990826 6 porb_h
port 681 nsew
rlabel metal2 s 79048 990762 79100 990826 6 porb_h
port 681 nsew
rlabel metal2 s 130292 990830 130344 990894 6 porb_h
port 681 nsew
rlabel metal2 s 130304 990894 130332 995407 6 porb_h
port 681 nsew
rlabel metal2 s 79060 990826 79088 992174 6 porb_h
port 681 nsew
rlabel metal2 s 78876 992174 79088 992202 6 porb_h
port 681 nsew
rlabel metal2 s 78876 992202 78904 995407 6 porb_h
port 681 nsew
rlabel metal2 s 181689 995407 181760 995466 6 porb_h
port 681 nsew
rlabel metal2 s 233089 995466 233145 995887 6 porb_h
port 681 nsew
rlabel metal2 s 181689 995466 181745 995887 6 porb_h
port 681 nsew
rlabel metal2 s 130289 995407 130345 995887 6 porb_h
port 681 nsew
rlabel metal2 s 78876 995407 78945 995452 6 porb_h
port 681 nsew
rlabel metal2 s 78889 995452 78945 995887 6 porb_h
port 681 nsew
rlabel via1 s 472532 41828 472584 41880 6 porb_h
port 681 nsew
rlabel via1 s 468484 41828 468536 41880 6 porb_h
port 681 nsew
rlabel via1 s 199568 41828 199620 41880 6 porb_h
port 681 nsew
rlabel via1 s 195428 41828 195480 41880 6 porb_h
port 681 nsew
rlabel via1 s 527364 41896 527416 41948 6 porb_h
port 681 nsew
rlabel via1 s 523224 41896 523276 41948 6 porb_h
port 681 nsew
rlabel via1 s 195336 44208 195388 44260 6 porb_h
port 681 nsew
rlabel via1 s 145104 44208 145156 44260 6 porb_h
port 681 nsew
rlabel via1 s 145104 45636 145156 45688 6 porb_h
port 681 nsew
rlabel via1 s 42248 45636 42300 45688 6 porb_h
port 681 nsew
rlabel via1 s 417884 47064 417936 47116 6 porb_h
port 681 nsew
rlabel via1 s 413560 47064 413612 47116 6 porb_h
port 681 nsew
rlabel via1 s 363052 47064 363104 47116 6 porb_h
port 681 nsew
rlabel via1 s 358728 47064 358780 47116 6 porb_h
port 681 nsew
rlabel via1 s 308220 47064 308272 47116 6 porb_h
port 681 nsew
rlabel via1 s 303896 47064 303948 47116 6 porb_h
port 681 nsew
rlabel via1 s 527456 47132 527508 47184 6 porb_h
port 681 nsew
rlabel via1 s 468300 47132 468352 47184 6 porb_h
port 681 nsew
rlabel via1 s 199660 47268 199712 47320 6 porb_h
port 681 nsew
rlabel via1 s 673552 47812 673604 47864 6 porb_h
port 681 nsew
rlabel via1 s 527456 47812 527508 47864 6 porb_h
port 681 nsew
rlabel via1 s 675392 112752 675444 112804 6 porb_h
port 681 nsew
rlabel via1 s 673552 112752 673604 112804 6 porb_h
port 681 nsew
rlabel via1 s 675392 158312 675444 158364 6 porb_h
port 681 nsew
rlabel via1 s 673552 158312 673604 158364 6 porb_h
port 681 nsew
rlabel via1 s 42432 184220 42484 184272 6 porb_h
port 681 nsew
rlabel via1 s 42248 184220 42300 184272 6 porb_h
port 681 nsew
rlabel via1 s 675392 203872 675444 203924 6 porb_h
port 681 nsew
rlabel via1 s 673828 203872 673880 203924 6 porb_h
port 681 nsew
rlabel via1 s 673552 203872 673604 203924 6 porb_h
port 681 nsew
rlabel via1 s 42708 228012 42760 228064 6 porb_h
port 681 nsew
rlabel via1 s 42432 228012 42484 228064 6 porb_h
port 681 nsew
rlabel via1 s 41788 228012 41840 228064 6 porb_h
port 681 nsew
rlabel via1 s 42708 246984 42760 247036 6 porb_h
port 681 nsew
rlabel via1 s 42340 246984 42392 247036 6 porb_h
port 681 nsew
rlabel via1 s 675392 248140 675444 248192 6 porb_h
port 681 nsew
rlabel via1 s 673828 248140 673880 248192 6 porb_h
port 681 nsew
rlabel via1 s 42708 270240 42760 270292 6 porb_h
port 681 nsew
rlabel via1 s 42340 270240 42392 270292 6 porb_h
port 681 nsew
rlabel via1 s 41788 270240 41840 270292 6 porb_h
port 681 nsew
rlabel via1 s 42708 282004 42760 282056 6 porb_h
port 681 nsew
rlabel via1 s 42708 282208 42760 282260 6 porb_h
port 681 nsew
rlabel via1 s 675392 293156 675444 293208 6 porb_h
port 681 nsew
rlabel via1 s 673828 293156 673880 293208 6 porb_h
port 681 nsew
rlabel via1 s 42708 307912 42760 307964 6 porb_h
port 681 nsew
rlabel via1 s 42432 307912 42484 307964 6 porb_h
port 681 nsew
rlabel via1 s 42432 313760 42484 313812 6 porb_h
port 681 nsew
rlabel via1 s 41788 313760 41840 313812 6 porb_h
port 681 nsew
rlabel via1 s 42432 356668 42484 356720 6 porb_h
port 681 nsew
rlabel via1 s 41788 356668 41840 356720 6 porb_h
port 681 nsew
rlabel via1 s 675392 384004 675444 384056 6 porb_h
port 681 nsew
rlabel via1 s 673552 384004 673604 384056 6 porb_h
port 681 nsew
rlabel via1 s 42432 400120 42484 400172 6 porb_h
port 681 nsew
rlabel via1 s 41972 400120 42024 400172 6 porb_h
port 681 nsew
rlabel via1 s 42616 528436 42668 528488 6 porb_h
port 681 nsew
rlabel via1 s 42432 528436 42484 528488 6 porb_h
port 681 nsew
rlabel via1 s 41788 528436 41840 528488 6 porb_h
port 681 nsew
rlabel via1 s 675392 561484 675444 561536 6 porb_h
port 681 nsew
rlabel via1 s 673644 561484 673696 561536 6 porb_h
port 681 nsew
rlabel via1 s 42616 571616 42668 571668 6 porb_h
port 681 nsew
rlabel via1 s 41788 571616 41840 571668 6 porb_h
port 681 nsew
rlabel via1 s 42616 584196 42668 584248 6 porb_h
port 681 nsew
rlabel via1 s 42248 584196 42300 584248 6 porb_h
port 681 nsew
rlabel via1 s 675392 606704 675444 606756 6 porb_h
port 681 nsew
rlabel via1 s 673644 606704 673696 606756 6 porb_h
port 681 nsew
rlabel via1 s 42616 614456 42668 614508 6 porb_h
port 681 nsew
rlabel via1 s 42248 614456 42300 614508 6 porb_h
port 681 nsew
rlabel via1 s 41880 614456 41932 614508 6 porb_h
port 681 nsew
rlabel via1 s 42616 633224 42668 633276 6 porb_h
port 681 nsew
rlabel via1 s 42340 633224 42392 633276 6 porb_h
port 681 nsew
rlabel via1 s 675392 651720 675444 651772 6 porb_h
port 681 nsew
rlabel via1 s 673644 651720 673696 651772 6 porb_h
port 681 nsew
rlabel via1 s 42616 657092 42668 657144 6 porb_h
port 681 nsew
rlabel via1 s 42340 657092 42392 657144 6 porb_h
port 681 nsew
rlabel via1 s 41788 657092 41840 657144 6 porb_h
port 681 nsew
rlabel via1 s 675392 695920 675444 695972 6 porb_h
port 681 nsew
rlabel via1 s 673644 695920 673696 695972 6 porb_h
port 681 nsew
rlabel via1 s 42616 700816 42668 700868 6 porb_h
port 681 nsew
rlabel via1 s 41788 700816 41840 700868 6 porb_h
port 681 nsew
rlabel via1 s 675300 710676 675352 710728 6 porb_h
port 681 nsew
rlabel via1 s 674012 710676 674064 710728 6 porb_h
port 681 nsew
rlabel via1 s 674196 720400 674248 720452 6 porb_h
port 681 nsew
rlabel via1 s 674012 720400 674064 720452 6 porb_h
port 681 nsew
rlabel via1 s 675392 741888 675444 741940 6 porb_h
port 681 nsew
rlabel via1 s 674196 741888 674248 741940 6 porb_h
port 681 nsew
rlabel via1 s 673552 741888 673604 741940 6 porb_h
port 681 nsew
rlabel via1 s 42616 744404 42668 744456 6 porb_h
port 681 nsew
rlabel via1 s 41788 744404 41840 744456 6 porb_h
port 681 nsew
rlabel via1 s 674012 768612 674064 768664 6 porb_h
port 681 nsew
rlabel via1 s 673552 768612 673604 768664 6 porb_h
port 681 nsew
rlabel via1 s 675300 786428 675352 786480 6 porb_h
port 681 nsew
rlabel via1 s 674012 786428 674064 786480 6 porb_h
port 681 nsew
rlabel via1 s 42616 787176 42668 787228 6 porb_h
port 681 nsew
rlabel via1 s 42248 787176 42300 787228 6 porb_h
port 681 nsew
rlabel via1 s 675300 797580 675352 797632 6 porb_h
port 681 nsew
rlabel via1 s 674104 797580 674156 797632 6 porb_h
port 681 nsew
rlabel via1 s 674104 821040 674156 821092 6 porb_h
port 681 nsew
rlabel via1 s 673552 821040 673604 821092 6 porb_h
port 681 nsew
rlabel via1 s 673644 830764 673696 830816 6 porb_h
port 681 nsew
rlabel via1 s 673552 830764 673604 830816 6 porb_h
port 681 nsew
rlabel via1 s 673644 836204 673696 836256 6 porb_h
port 681 nsew
rlabel via1 s 673552 836272 673604 836324 6 porb_h
port 681 nsew
rlabel via1 s 675208 869388 675260 869440 6 porb_h
port 681 nsew
rlabel via1 s 673736 869388 673788 869440 6 porb_h
port 681 nsew
rlabel via1 s 673460 888768 673512 888820 6 porb_h
port 681 nsew
rlabel via1 s 673184 888768 673236 888820 6 porb_h
port 681 nsew
rlabel via1 s 673460 908012 673512 908064 6 porb_h
port 681 nsew
rlabel via1 s 673184 908012 673236 908064 6 porb_h
port 681 nsew
rlabel via1 s 42432 956428 42484 956480 6 porb_h
port 681 nsew
rlabel via1 s 41788 956428 41840 956480 6 porb_h
port 681 nsew
rlabel via1 s 675392 965268 675444 965320 6 porb_h
port 681 nsew
rlabel via1 s 673460 965268 673512 965320 6 porb_h
port 681 nsew
rlabel via1 s 673460 990020 673512 990072 6 porb_h
port 681 nsew
rlabel via1 s 628656 990088 628708 990140 6 porb_h
port 681 nsew
rlabel via1 s 79048 990088 79100 990140 6 porb_h
port 681 nsew
rlabel via1 s 42432 990088 42484 990140 6 porb_h
port 681 nsew
rlabel via1 s 246948 990428 247000 990480 6 porb_h
port 681 nsew
rlabel via1 s 233056 990428 233108 990480 6 porb_h
port 681 nsew
rlabel via1 s 202880 990428 202932 990480 6 porb_h
port 681 nsew
rlabel via1 s 187700 990428 187752 990480 6 porb_h
port 681 nsew
rlabel via1 s 187608 990428 187660 990480 6 porb_h
port 681 nsew
rlabel via1 s 181720 990428 181772 990480 6 porb_h
port 681 nsew
rlabel via1 s 160100 990428 160152 990480 6 porb_h
port 681 nsew
rlabel via1 s 143264 990428 143316 990480 6 porb_h
port 681 nsew
rlabel via1 s 450268 990564 450320 990616 6 porb_h
port 681 nsew
rlabel via1 s 438768 990564 438820 990616 6 porb_h
port 681 nsew
rlabel via1 s 419540 990564 419592 990616 6 porb_h
port 681 nsew
rlabel via1 s 286968 990496 287020 990548 6 porb_h
port 681 nsew
rlabel via1 s 386512 990564 386564 990616 6 porb_h
port 681 nsew
rlabel via1 s 181720 990564 181772 990616 6 porb_h
port 681 nsew
rlabel via1 s 179328 990564 179380 990616 6 porb_h
port 681 nsew
rlabel via1 s 130108 990564 130160 990616 6 porb_h
port 681 nsew
rlabel via1 s 110512 990564 110564 990616 6 porb_h
port 681 nsew
rlabel via1 s 628656 990700 628708 990752 6 porb_h
port 681 nsew
rlabel via1 s 526904 990700 526956 990752 6 porb_h
port 681 nsew
rlabel via1 s 482928 990700 482980 990752 6 porb_h
port 681 nsew
rlabel via1 s 233056 990700 233108 990752 6 porb_h
port 681 nsew
rlabel via1 s 202880 990700 202932 990752 6 porb_h
port 681 nsew
rlabel via1 s 187700 990700 187752 990752 6 porb_h
port 681 nsew
rlabel via1 s 187608 990700 187660 990752 6 porb_h
port 681 nsew
rlabel via1 s 286968 990768 287020 990820 6 porb_h
port 681 nsew
rlabel via1 s 284668 990768 284720 990820 6 porb_h
port 681 nsew
rlabel via1 s 246948 990768 247000 990820 6 porb_h
port 681 nsew
rlabel via1 s 179328 990768 179380 990820 6 porb_h
port 681 nsew
rlabel via1 s 173808 990768 173860 990820 6 porb_h
port 681 nsew
rlabel via1 s 143264 990768 143316 990820 6 porb_h
port 681 nsew
rlabel via1 s 463608 990836 463660 990888 6 porb_h
port 681 nsew
rlabel via1 s 450268 990836 450320 990888 6 porb_h
port 681 nsew
rlabel via1 s 438676 990836 438728 990888 6 porb_h
port 681 nsew
rlabel via1 s 419540 990836 419592 990888 6 porb_h
port 681 nsew
rlabel via1 s 130108 990768 130160 990820 6 porb_h
port 681 nsew
rlabel via1 s 110420 990768 110472 990820 6 porb_h
port 681 nsew
rlabel via1 s 79048 990768 79100 990820 6 porb_h
port 681 nsew
rlabel via1 s 130292 990836 130344 990888 6 porb_h
port 681 nsew
rlabel via1 s 482928 992264 482980 992316 6 porb_h
port 681 nsew
rlabel via1 s 475476 992264 475528 992316 6 porb_h
port 681 nsew
rlabel via1 s 463792 992264 463844 992316 6 porb_h
port 681 nsew
rlabel metal1 s 472526 41828 472590 41840 6 porb_h
port 681 nsew
rlabel metal1 s 468478 41828 468542 41840 6 porb_h
port 681 nsew
rlabel metal1 s 468478 41840 472590 41868 6 porb_h
port 681 nsew
rlabel metal1 s 472526 41868 472590 41880 6 porb_h
port 681 nsew
rlabel metal1 s 468478 41868 468542 41880 6 porb_h
port 681 nsew
rlabel metal1 s 199562 41828 199626 41840 6 porb_h
port 681 nsew
rlabel metal1 s 195422 41828 195486 41840 6 porb_h
port 681 nsew
rlabel metal1 s 195422 41840 199626 41868 6 porb_h
port 681 nsew
rlabel metal1 s 199562 41868 199626 41880 6 porb_h
port 681 nsew
rlabel metal1 s 195422 41868 195486 41880 6 porb_h
port 681 nsew
rlabel metal1 s 527358 41896 527422 41908 6 porb_h
port 681 nsew
rlabel metal1 s 523218 41896 523282 41908 6 porb_h
port 681 nsew
rlabel metal1 s 523218 41908 527422 41936 6 porb_h
port 681 nsew
rlabel metal1 s 527358 41936 527422 41948 6 porb_h
port 681 nsew
rlabel metal1 s 523218 41936 523282 41948 6 porb_h
port 681 nsew
rlabel metal1 s 195330 44208 195394 44220 6 porb_h
port 681 nsew
rlabel metal1 s 145098 44208 145162 44220 6 porb_h
port 681 nsew
rlabel metal1 s 145098 44220 195394 44248 6 porb_h
port 681 nsew
rlabel metal1 s 195330 44248 195394 44260 6 porb_h
port 681 nsew
rlabel metal1 s 145098 44248 145162 44260 6 porb_h
port 681 nsew
rlabel metal1 s 145098 45636 145162 45648 6 porb_h
port 681 nsew
rlabel metal1 s 42242 45636 42306 45648 6 porb_h
port 681 nsew
rlabel metal1 s 42242 45648 145162 45676 6 porb_h
port 681 nsew
rlabel metal1 s 145098 45676 145162 45688 6 porb_h
port 681 nsew
rlabel metal1 s 42242 45676 42306 45688 6 porb_h
port 681 nsew
rlabel metal1 s 417878 47064 417942 47076 6 porb_h
port 681 nsew
rlabel metal1 s 413554 47064 413618 47076 6 porb_h
port 681 nsew
rlabel metal1 s 363046 47064 363110 47076 6 porb_h
port 681 nsew
rlabel metal1 s 358722 47064 358786 47076 6 porb_h
port 681 nsew
rlabel metal1 s 308214 47064 308278 47076 6 porb_h
port 681 nsew
rlabel metal1 s 303890 47064 303954 47076 6 porb_h
port 681 nsew
rlabel metal1 s 285692 47076 417942 47104 6 porb_h
port 681 nsew
rlabel metal1 s 417878 47104 417942 47116 6 porb_h
port 681 nsew
rlabel metal1 s 413554 47104 413618 47116 6 porb_h
port 681 nsew
rlabel metal1 s 363046 47104 363110 47116 6 porb_h
port 681 nsew
rlabel metal1 s 358722 47104 358786 47116 6 porb_h
port 681 nsew
rlabel metal1 s 308214 47104 308278 47116 6 porb_h
port 681 nsew
rlabel metal1 s 303890 47104 303954 47116 6 porb_h
port 681 nsew
rlabel metal1 s 527450 47132 527514 47144 6 porb_h
port 681 nsew
rlabel metal1 s 468294 47132 468358 47144 6 porb_h
port 681 nsew
rlabel metal1 s 417896 47116 417924 47144 6 porb_h
port 681 nsew
rlabel metal1 s 417896 47144 527514 47172 6 porb_h
port 681 nsew
rlabel metal1 s 527450 47172 527514 47184 6 porb_h
port 681 nsew
rlabel metal1 s 468294 47172 468358 47184 6 porb_h
port 681 nsew
rlabel metal1 s 285692 47104 285720 47212 6 porb_h
port 681 nsew
rlabel metal1 s 276032 47212 285720 47240 6 porb_h
port 681 nsew
rlabel metal1 s 276032 47240 276060 47280 6 porb_h
port 681 nsew
rlabel metal1 s 199654 47268 199718 47280 6 porb_h
port 681 nsew
rlabel metal1 s 199654 47280 276060 47308 6 porb_h
port 681 nsew
rlabel metal1 s 199654 47308 199718 47320 6 porb_h
port 681 nsew
rlabel metal1 s 673546 47812 673610 47824 6 porb_h
port 681 nsew
rlabel metal1 s 527450 47812 527514 47824 6 porb_h
port 681 nsew
rlabel metal1 s 527450 47824 673610 47852 6 porb_h
port 681 nsew
rlabel metal1 s 673546 47852 673610 47864 6 porb_h
port 681 nsew
rlabel metal1 s 527450 47852 527514 47864 6 porb_h
port 681 nsew
rlabel metal1 s 675386 112752 675450 112764 6 porb_h
port 681 nsew
rlabel metal1 s 673546 112752 673610 112764 6 porb_h
port 681 nsew
rlabel metal1 s 673546 112764 675450 112792 6 porb_h
port 681 nsew
rlabel metal1 s 675386 112792 675450 112804 6 porb_h
port 681 nsew
rlabel metal1 s 673546 112792 673610 112804 6 porb_h
port 681 nsew
rlabel metal1 s 675386 158312 675450 158324 6 porb_h
port 681 nsew
rlabel metal1 s 673546 158312 673610 158324 6 porb_h
port 681 nsew
rlabel metal1 s 673546 158324 675450 158352 6 porb_h
port 681 nsew
rlabel metal1 s 675386 158352 675450 158364 6 porb_h
port 681 nsew
rlabel metal1 s 673546 158352 673610 158364 6 porb_h
port 681 nsew
rlabel metal1 s 42426 184220 42490 184232 6 porb_h
port 681 nsew
rlabel metal1 s 42242 184220 42306 184232 6 porb_h
port 681 nsew
rlabel metal1 s 42242 184232 42490 184260 6 porb_h
port 681 nsew
rlabel metal1 s 42426 184260 42490 184272 6 porb_h
port 681 nsew
rlabel metal1 s 42242 184260 42306 184272 6 porb_h
port 681 nsew
rlabel metal1 s 675386 203872 675450 203884 6 porb_h
port 681 nsew
rlabel metal1 s 673822 203872 673886 203884 6 porb_h
port 681 nsew
rlabel metal1 s 673546 203872 673610 203884 6 porb_h
port 681 nsew
rlabel metal1 s 673546 203884 675450 203912 6 porb_h
port 681 nsew
rlabel metal1 s 675386 203912 675450 203924 6 porb_h
port 681 nsew
rlabel metal1 s 673822 203912 673886 203924 6 porb_h
port 681 nsew
rlabel metal1 s 673546 203912 673610 203924 6 porb_h
port 681 nsew
rlabel metal1 s 42702 228012 42766 228024 6 porb_h
port 681 nsew
rlabel metal1 s 42426 228012 42490 228024 6 porb_h
port 681 nsew
rlabel metal1 s 41782 228012 41846 228024 6 porb_h
port 681 nsew
rlabel metal1 s 41782 228024 42766 228052 6 porb_h
port 681 nsew
rlabel metal1 s 42702 228052 42766 228064 6 porb_h
port 681 nsew
rlabel metal1 s 42426 228052 42490 228064 6 porb_h
port 681 nsew
rlabel metal1 s 41782 228052 41846 228064 6 porb_h
port 681 nsew
rlabel metal1 s 42702 246984 42766 246996 6 porb_h
port 681 nsew
rlabel metal1 s 42334 246984 42398 246996 6 porb_h
port 681 nsew
rlabel metal1 s 42334 246996 42766 247024 6 porb_h
port 681 nsew
rlabel metal1 s 42702 247024 42766 247036 6 porb_h
port 681 nsew
rlabel metal1 s 42334 247024 42398 247036 6 porb_h
port 681 nsew
rlabel metal1 s 675386 248140 675450 248152 6 porb_h
port 681 nsew
rlabel metal1 s 673822 248140 673886 248152 6 porb_h
port 681 nsew
rlabel metal1 s 673822 248152 675450 248180 6 porb_h
port 681 nsew
rlabel metal1 s 675386 248180 675450 248192 6 porb_h
port 681 nsew
rlabel metal1 s 673822 248180 673886 248192 6 porb_h
port 681 nsew
rlabel metal1 s 42702 270240 42766 270252 6 porb_h
port 681 nsew
rlabel metal1 s 42334 270240 42398 270252 6 porb_h
port 681 nsew
rlabel metal1 s 41782 270240 41846 270252 6 porb_h
port 681 nsew
rlabel metal1 s 41782 270252 42766 270280 6 porb_h
port 681 nsew
rlabel metal1 s 42702 270280 42766 270292 6 porb_h
port 681 nsew
rlabel metal1 s 42334 270280 42398 270292 6 porb_h
port 681 nsew
rlabel metal1 s 41782 270280 41846 270292 6 porb_h
port 681 nsew
rlabel metal1 s 42702 282004 42766 282056 6 porb_h
port 681 nsew
rlabel metal1 s 42720 282056 42748 282208 6 porb_h
port 681 nsew
rlabel metal1 s 42702 282208 42766 282260 6 porb_h
port 681 nsew
rlabel metal1 s 675386 293156 675450 293168 6 porb_h
port 681 nsew
rlabel metal1 s 673822 293156 673886 293168 6 porb_h
port 681 nsew
rlabel metal1 s 673822 293168 675450 293196 6 porb_h
port 681 nsew
rlabel metal1 s 675386 293196 675450 293208 6 porb_h
port 681 nsew
rlabel metal1 s 673822 293196 673886 293208 6 porb_h
port 681 nsew
rlabel metal1 s 42702 307912 42766 307924 6 porb_h
port 681 nsew
rlabel metal1 s 42426 307912 42490 307924 6 porb_h
port 681 nsew
rlabel metal1 s 42426 307924 42766 307952 6 porb_h
port 681 nsew
rlabel metal1 s 42702 307952 42766 307964 6 porb_h
port 681 nsew
rlabel metal1 s 42426 307952 42490 307964 6 porb_h
port 681 nsew
rlabel metal1 s 42426 313760 42490 313772 6 porb_h
port 681 nsew
rlabel metal1 s 41782 313760 41846 313772 6 porb_h
port 681 nsew
rlabel metal1 s 41782 313772 42490 313800 6 porb_h
port 681 nsew
rlabel metal1 s 42426 313800 42490 313812 6 porb_h
port 681 nsew
rlabel metal1 s 41782 313800 41846 313812 6 porb_h
port 681 nsew
rlabel metal1 s 42426 356668 42490 356680 6 porb_h
port 681 nsew
rlabel metal1 s 41782 356668 41846 356680 6 porb_h
port 681 nsew
rlabel metal1 s 41782 356680 42490 356708 6 porb_h
port 681 nsew
rlabel metal1 s 42426 356708 42490 356720 6 porb_h
port 681 nsew
rlabel metal1 s 41782 356708 41846 356720 6 porb_h
port 681 nsew
rlabel metal1 s 675386 384004 675450 384016 6 porb_h
port 681 nsew
rlabel metal1 s 673546 384004 673610 384016 6 porb_h
port 681 nsew
rlabel metal1 s 673546 384016 675450 384044 6 porb_h
port 681 nsew
rlabel metal1 s 675386 384044 675450 384056 6 porb_h
port 681 nsew
rlabel metal1 s 673546 384044 673610 384056 6 porb_h
port 681 nsew
rlabel metal1 s 42426 400120 42490 400132 6 porb_h
port 681 nsew
rlabel metal1 s 41966 400120 42030 400132 6 porb_h
port 681 nsew
rlabel metal1 s 41966 400132 42490 400160 6 porb_h
port 681 nsew
rlabel metal1 s 42426 400160 42490 400172 6 porb_h
port 681 nsew
rlabel metal1 s 41966 400160 42030 400172 6 porb_h
port 681 nsew
rlabel metal1 s 42610 528436 42674 528448 6 porb_h
port 681 nsew
rlabel metal1 s 42426 528436 42490 528448 6 porb_h
port 681 nsew
rlabel metal1 s 41782 528436 41846 528448 6 porb_h
port 681 nsew
rlabel metal1 s 41782 528448 42674 528476 6 porb_h
port 681 nsew
rlabel metal1 s 42610 528476 42674 528488 6 porb_h
port 681 nsew
rlabel metal1 s 42426 528476 42490 528488 6 porb_h
port 681 nsew
rlabel metal1 s 41782 528476 41846 528488 6 porb_h
port 681 nsew
rlabel metal1 s 675386 561484 675450 561496 6 porb_h
port 681 nsew
rlabel metal1 s 673638 561484 673702 561496 6 porb_h
port 681 nsew
rlabel metal1 s 673638 561496 675450 561524 6 porb_h
port 681 nsew
rlabel metal1 s 675386 561524 675450 561536 6 porb_h
port 681 nsew
rlabel metal1 s 673638 561524 673702 561536 6 porb_h
port 681 nsew
rlabel metal1 s 42610 571616 42674 571628 6 porb_h
port 681 nsew
rlabel metal1 s 41782 571616 41846 571628 6 porb_h
port 681 nsew
rlabel metal1 s 41782 571628 42674 571656 6 porb_h
port 681 nsew
rlabel metal1 s 42610 571656 42674 571668 6 porb_h
port 681 nsew
rlabel metal1 s 41782 571656 41846 571668 6 porb_h
port 681 nsew
rlabel metal1 s 42610 584196 42674 584208 6 porb_h
port 681 nsew
rlabel metal1 s 42242 584196 42306 584208 6 porb_h
port 681 nsew
rlabel metal1 s 42242 584208 42674 584236 6 porb_h
port 681 nsew
rlabel metal1 s 42610 584236 42674 584248 6 porb_h
port 681 nsew
rlabel metal1 s 42242 584236 42306 584248 6 porb_h
port 681 nsew
rlabel metal1 s 675386 606704 675450 606716 6 porb_h
port 681 nsew
rlabel metal1 s 673638 606704 673702 606716 6 porb_h
port 681 nsew
rlabel metal1 s 673638 606716 675450 606744 6 porb_h
port 681 nsew
rlabel metal1 s 675386 606744 675450 606756 6 porb_h
port 681 nsew
rlabel metal1 s 673638 606744 673702 606756 6 porb_h
port 681 nsew
rlabel metal1 s 42610 614456 42674 614468 6 porb_h
port 681 nsew
rlabel metal1 s 42242 614456 42306 614468 6 porb_h
port 681 nsew
rlabel metal1 s 41874 614456 41938 614468 6 porb_h
port 681 nsew
rlabel metal1 s 41874 614468 42674 614496 6 porb_h
port 681 nsew
rlabel metal1 s 42610 614496 42674 614508 6 porb_h
port 681 nsew
rlabel metal1 s 42242 614496 42306 614508 6 porb_h
port 681 nsew
rlabel metal1 s 41874 614496 41938 614508 6 porb_h
port 681 nsew
rlabel metal1 s 42610 633224 42674 633236 6 porb_h
port 681 nsew
rlabel metal1 s 42334 633224 42398 633236 6 porb_h
port 681 nsew
rlabel metal1 s 42334 633236 42674 633264 6 porb_h
port 681 nsew
rlabel metal1 s 42610 633264 42674 633276 6 porb_h
port 681 nsew
rlabel metal1 s 42334 633264 42398 633276 6 porb_h
port 681 nsew
rlabel metal1 s 675386 651720 675450 651732 6 porb_h
port 681 nsew
rlabel metal1 s 673638 651720 673702 651732 6 porb_h
port 681 nsew
rlabel metal1 s 673638 651732 675450 651760 6 porb_h
port 681 nsew
rlabel metal1 s 675386 651760 675450 651772 6 porb_h
port 681 nsew
rlabel metal1 s 673638 651760 673702 651772 6 porb_h
port 681 nsew
rlabel metal1 s 42610 657092 42674 657104 6 porb_h
port 681 nsew
rlabel metal1 s 42334 657092 42398 657104 6 porb_h
port 681 nsew
rlabel metal1 s 41782 657092 41846 657104 6 porb_h
port 681 nsew
rlabel metal1 s 41782 657104 42674 657132 6 porb_h
port 681 nsew
rlabel metal1 s 42610 657132 42674 657144 6 porb_h
port 681 nsew
rlabel metal1 s 42334 657132 42398 657144 6 porb_h
port 681 nsew
rlabel metal1 s 41782 657132 41846 657144 6 porb_h
port 681 nsew
rlabel metal1 s 675386 695920 675450 695932 6 porb_h
port 681 nsew
rlabel metal1 s 673638 695920 673702 695932 6 porb_h
port 681 nsew
rlabel metal1 s 673638 695932 675450 695960 6 porb_h
port 681 nsew
rlabel metal1 s 675386 695960 675450 695972 6 porb_h
port 681 nsew
rlabel metal1 s 673638 695960 673702 695972 6 porb_h
port 681 nsew
rlabel metal1 s 42610 700816 42674 700828 6 porb_h
port 681 nsew
rlabel metal1 s 41782 700816 41846 700828 6 porb_h
port 681 nsew
rlabel metal1 s 41782 700828 42674 700856 6 porb_h
port 681 nsew
rlabel metal1 s 42610 700856 42674 700868 6 porb_h
port 681 nsew
rlabel metal1 s 41782 700856 41846 700868 6 porb_h
port 681 nsew
rlabel metal1 s 675294 710676 675358 710688 6 porb_h
port 681 nsew
rlabel metal1 s 674006 710676 674070 710688 6 porb_h
port 681 nsew
rlabel metal1 s 674006 710688 675358 710716 6 porb_h
port 681 nsew
rlabel metal1 s 675294 710716 675358 710728 6 porb_h
port 681 nsew
rlabel metal1 s 674006 710716 674070 710728 6 porb_h
port 681 nsew
rlabel metal1 s 674190 720400 674254 720412 6 porb_h
port 681 nsew
rlabel metal1 s 674006 720400 674070 720412 6 porb_h
port 681 nsew
rlabel metal1 s 674006 720412 674254 720440 6 porb_h
port 681 nsew
rlabel metal1 s 674190 720440 674254 720452 6 porb_h
port 681 nsew
rlabel metal1 s 674006 720440 674070 720452 6 porb_h
port 681 nsew
rlabel metal1 s 675386 741888 675450 741900 6 porb_h
port 681 nsew
rlabel metal1 s 674190 741888 674254 741900 6 porb_h
port 681 nsew
rlabel metal1 s 673546 741888 673610 741900 6 porb_h
port 681 nsew
rlabel metal1 s 673546 741900 675450 741928 6 porb_h
port 681 nsew
rlabel metal1 s 675386 741928 675450 741940 6 porb_h
port 681 nsew
rlabel metal1 s 674190 741928 674254 741940 6 porb_h
port 681 nsew
rlabel metal1 s 673546 741928 673610 741940 6 porb_h
port 681 nsew
rlabel metal1 s 42610 744404 42674 744416 6 porb_h
port 681 nsew
rlabel metal1 s 41782 744404 41846 744416 6 porb_h
port 681 nsew
rlabel metal1 s 41782 744416 42674 744444 6 porb_h
port 681 nsew
rlabel metal1 s 42610 744444 42674 744456 6 porb_h
port 681 nsew
rlabel metal1 s 41782 744444 41846 744456 6 porb_h
port 681 nsew
rlabel metal1 s 674006 768612 674070 768624 6 porb_h
port 681 nsew
rlabel metal1 s 673546 768612 673610 768624 6 porb_h
port 681 nsew
rlabel metal1 s 673546 768624 674070 768652 6 porb_h
port 681 nsew
rlabel metal1 s 674006 768652 674070 768664 6 porb_h
port 681 nsew
rlabel metal1 s 673546 768652 673610 768664 6 porb_h
port 681 nsew
rlabel metal1 s 675294 786428 675358 786440 6 porb_h
port 681 nsew
rlabel metal1 s 674006 786428 674070 786440 6 porb_h
port 681 nsew
rlabel metal1 s 674006 786440 675358 786468 6 porb_h
port 681 nsew
rlabel metal1 s 675294 786468 675358 786480 6 porb_h
port 681 nsew
rlabel metal1 s 674006 786468 674070 786480 6 porb_h
port 681 nsew
rlabel metal1 s 42610 787176 42674 787188 6 porb_h
port 681 nsew
rlabel metal1 s 42242 787176 42306 787188 6 porb_h
port 681 nsew
rlabel metal1 s 42242 787188 42674 787216 6 porb_h
port 681 nsew
rlabel metal1 s 42610 787216 42674 787228 6 porb_h
port 681 nsew
rlabel metal1 s 42242 787216 42306 787228 6 porb_h
port 681 nsew
rlabel metal1 s 675294 797580 675358 797592 6 porb_h
port 681 nsew
rlabel metal1 s 674098 797580 674162 797592 6 porb_h
port 681 nsew
rlabel metal1 s 674098 797592 675358 797620 6 porb_h
port 681 nsew
rlabel metal1 s 675294 797620 675358 797632 6 porb_h
port 681 nsew
rlabel metal1 s 674098 797620 674162 797632 6 porb_h
port 681 nsew
rlabel metal1 s 674098 821040 674162 821052 6 porb_h
port 681 nsew
rlabel metal1 s 673546 821040 673610 821052 6 porb_h
port 681 nsew
rlabel metal1 s 673546 821052 674162 821080 6 porb_h
port 681 nsew
rlabel metal1 s 674098 821080 674162 821092 6 porb_h
port 681 nsew
rlabel metal1 s 673546 821080 673610 821092 6 porb_h
port 681 nsew
rlabel metal1 s 673638 830764 673702 830776 6 porb_h
port 681 nsew
rlabel metal1 s 673546 830764 673610 830776 6 porb_h
port 681 nsew
rlabel metal1 s 673546 830776 673702 830804 6 porb_h
port 681 nsew
rlabel metal1 s 673638 830804 673702 830816 6 porb_h
port 681 nsew
rlabel metal1 s 673546 830804 673610 830816 6 porb_h
port 681 nsew
rlabel metal1 s 673638 836204 673702 836256 6 porb_h
port 681 nsew
rlabel metal1 s 673656 836256 673684 836284 6 porb_h
port 681 nsew
rlabel metal1 s 673546 836272 673610 836284 6 porb_h
port 681 nsew
rlabel metal1 s 673546 836284 673684 836312 6 porb_h
port 681 nsew
rlabel metal1 s 673546 836312 673610 836324 6 porb_h
port 681 nsew
rlabel metal1 s 675202 869388 675266 869400 6 porb_h
port 681 nsew
rlabel metal1 s 673730 869388 673794 869400 6 porb_h
port 681 nsew
rlabel metal1 s 673730 869400 675266 869428 6 porb_h
port 681 nsew
rlabel metal1 s 675202 869428 675266 869440 6 porb_h
port 681 nsew
rlabel metal1 s 673730 869428 673794 869440 6 porb_h
port 681 nsew
rlabel metal1 s 673454 888768 673518 888780 6 porb_h
port 681 nsew
rlabel metal1 s 673178 888768 673242 888780 6 porb_h
port 681 nsew
rlabel metal1 s 673178 888780 673518 888808 6 porb_h
port 681 nsew
rlabel metal1 s 673454 888808 673518 888820 6 porb_h
port 681 nsew
rlabel metal1 s 673178 888808 673242 888820 6 porb_h
port 681 nsew
rlabel metal1 s 673454 908012 673518 908024 6 porb_h
port 681 nsew
rlabel metal1 s 673178 908012 673242 908024 6 porb_h
port 681 nsew
rlabel metal1 s 673178 908024 673518 908052 6 porb_h
port 681 nsew
rlabel metal1 s 673454 908052 673518 908064 6 porb_h
port 681 nsew
rlabel metal1 s 673178 908052 673242 908064 6 porb_h
port 681 nsew
rlabel metal1 s 42426 956428 42490 956440 6 porb_h
port 681 nsew
rlabel metal1 s 41782 956428 41846 956440 6 porb_h
port 681 nsew
rlabel metal1 s 41782 956440 42490 956468 6 porb_h
port 681 nsew
rlabel metal1 s 42426 956468 42490 956480 6 porb_h
port 681 nsew
rlabel metal1 s 41782 956468 41846 956480 6 porb_h
port 681 nsew
rlabel metal1 s 675386 965268 675450 965280 6 porb_h
port 681 nsew
rlabel metal1 s 673454 965268 673518 965280 6 porb_h
port 681 nsew
rlabel metal1 s 673454 965280 675450 965308 6 porb_h
port 681 nsew
rlabel metal1 s 675386 965308 675450 965320 6 porb_h
port 681 nsew
rlabel metal1 s 673454 965308 673518 965320 6 porb_h
port 681 nsew
rlabel metal1 s 673454 990020 673518 990032 6 porb_h
port 681 nsew
rlabel metal1 s 628668 990032 673518 990060 6 porb_h
port 681 nsew
rlabel metal1 s 673454 990060 673518 990072 6 porb_h
port 681 nsew
rlabel metal1 s 628668 990060 628696 990088 6 porb_h
port 681 nsew
rlabel metal1 s 628650 990088 628714 990140 6 porb_h
port 681 nsew
rlabel metal1 s 79042 990088 79106 990100 6 porb_h
port 681 nsew
rlabel metal1 s 42426 990088 42490 990100 6 porb_h
port 681 nsew
rlabel metal1 s 42426 990100 79106 990128 6 porb_h
port 681 nsew
rlabel metal1 s 79042 990128 79106 990140 6 porb_h
port 681 nsew
rlabel metal1 s 42426 990128 42490 990140 6 porb_h
port 681 nsew
rlabel metal1 s 246942 990428 247006 990440 6 porb_h
port 681 nsew
rlabel metal1 s 233050 990428 233114 990440 6 porb_h
port 681 nsew
rlabel metal1 s 233050 990440 247006 990468 6 porb_h
port 681 nsew
rlabel metal1 s 246942 990468 247006 990480 6 porb_h
port 681 nsew
rlabel metal1 s 233050 990468 233114 990480 6 porb_h
port 681 nsew
rlabel metal1 s 202874 990428 202938 990440 6 porb_h
port 681 nsew
rlabel metal1 s 187694 990428 187758 990440 6 porb_h
port 681 nsew
rlabel metal1 s 187694 990440 202938 990468 6 porb_h
port 681 nsew
rlabel metal1 s 202874 990468 202938 990480 6 porb_h
port 681 nsew
rlabel metal1 s 187694 990468 187758 990480 6 porb_h
port 681 nsew
rlabel metal1 s 187602 990428 187666 990440 6 porb_h
port 681 nsew
rlabel metal1 s 181714 990428 181778 990440 6 porb_h
port 681 nsew
rlabel metal1 s 181714 990440 187666 990468 6 porb_h
port 681 nsew
rlabel metal1 s 187602 990468 187666 990480 6 porb_h
port 681 nsew
rlabel metal1 s 181714 990468 181778 990480 6 porb_h
port 681 nsew
rlabel metal1 s 160094 990428 160158 990440 6 porb_h
port 681 nsew
rlabel metal1 s 143258 990428 143322 990440 6 porb_h
port 681 nsew
rlabel metal1 s 143258 990440 160158 990468 6 porb_h
port 681 nsew
rlabel metal1 s 160094 990468 160158 990480 6 porb_h
port 681 nsew
rlabel metal1 s 143258 990468 143322 990480 6 porb_h
port 681 nsew
rlabel metal1 s 286962 990496 287026 990508 6 porb_h
port 681 nsew
rlabel metal1 s 405568 990508 405780 990536 6 porb_h
port 681 nsew
rlabel metal1 s 450262 990564 450326 990576 6 porb_h
port 681 nsew
rlabel metal1 s 438762 990564 438826 990576 6 porb_h
port 681 nsew
rlabel metal1 s 438762 990576 450326 990604 6 porb_h
port 681 nsew
rlabel metal1 s 450262 990604 450326 990616 6 porb_h
port 681 nsew
rlabel metal1 s 438762 990604 438826 990616 6 porb_h
port 681 nsew
rlabel metal1 s 419534 990564 419598 990576 6 porb_h
port 681 nsew
rlabel metal1 s 405752 990536 405780 990576 6 porb_h
port 681 nsew
rlabel metal1 s 405752 990576 419598 990604 6 porb_h
port 681 nsew
rlabel metal1 s 419534 990604 419598 990616 6 porb_h
port 681 nsew
rlabel metal1 s 405568 990536 405596 990644 6 porb_h
port 681 nsew
rlabel metal1 s 286962 990508 386552 990536 6 porb_h
port 681 nsew
rlabel metal1 s 386524 990536 386552 990564 6 porb_h
port 681 nsew
rlabel metal1 s 286962 990536 287026 990548 6 porb_h
port 681 nsew
rlabel metal1 s 386506 990564 386570 990576 6 porb_h
port 681 nsew
rlabel metal1 s 181714 990564 181778 990576 6 porb_h
port 681 nsew
rlabel metal1 s 179322 990564 179386 990576 6 porb_h
port 681 nsew
rlabel metal1 s 386419 990576 391888 990604 6 porb_h
port 681 nsew
rlabel metal1 s 179322 990576 181778 990604 6 porb_h
port 681 nsew
rlabel metal1 s 391860 990604 391888 990644 6 porb_h
port 681 nsew
rlabel metal1 s 386506 990604 386570 990616 6 porb_h
port 681 nsew
rlabel metal1 s 181714 990604 181778 990616 6 porb_h
port 681 nsew
rlabel metal1 s 179322 990604 179386 990616 6 porb_h
port 681 nsew
rlabel metal1 s 130102 990564 130166 990576 6 porb_h
port 681 nsew
rlabel metal1 s 110506 990564 110570 990576 6 porb_h
port 681 nsew
rlabel metal1 s 110506 990576 130166 990604 6 porb_h
port 681 nsew
rlabel metal1 s 130102 990604 130166 990616 6 porb_h
port 681 nsew
rlabel metal1 s 110506 990604 110570 990616 6 porb_h
port 681 nsew
rlabel metal1 s 391860 990644 405596 990672 6 porb_h
port 681 nsew
rlabel metal1 s 628650 990700 628714 990712 6 porb_h
port 681 nsew
rlabel metal1 s 526898 990700 526962 990712 6 porb_h
port 681 nsew
rlabel metal1 s 482922 990700 482986 990712 6 porb_h
port 681 nsew
rlabel metal1 s 482922 990712 628714 990740 6 porb_h
port 681 nsew
rlabel metal1 s 628650 990740 628714 990752 6 porb_h
port 681 nsew
rlabel metal1 s 526898 990740 526962 990752 6 porb_h
port 681 nsew
rlabel metal1 s 482922 990740 482986 990752 6 porb_h
port 681 nsew
rlabel metal1 s 233050 990700 233114 990712 6 porb_h
port 681 nsew
rlabel metal1 s 202874 990700 202938 990712 6 porb_h
port 681 nsew
rlabel metal1 s 202874 990712 233114 990740 6 porb_h
port 681 nsew
rlabel metal1 s 233050 990740 233114 990752 6 porb_h
port 681 nsew
rlabel metal1 s 202874 990740 202938 990752 6 porb_h
port 681 nsew
rlabel metal1 s 187694 990700 187758 990712 6 porb_h
port 681 nsew
rlabel metal1 s 187602 990700 187666 990712 6 porb_h
port 681 nsew
rlabel metal1 s 187602 990712 187758 990740 6 porb_h
port 681 nsew
rlabel metal1 s 187694 990740 187758 990752 6 porb_h
port 681 nsew
rlabel metal1 s 187602 990740 187666 990752 6 porb_h
port 681 nsew
rlabel metal1 s 286962 990768 287026 990780 6 porb_h
port 681 nsew
rlabel metal1 s 284662 990768 284726 990780 6 porb_h
port 681 nsew
rlabel metal1 s 246942 990768 247006 990780 6 porb_h
port 681 nsew
rlabel metal1 s 246942 990780 287026 990808 6 porb_h
port 681 nsew
rlabel metal1 s 286962 990808 287026 990820 6 porb_h
port 681 nsew
rlabel metal1 s 284662 990808 284726 990820 6 porb_h
port 681 nsew
rlabel metal1 s 246942 990808 247006 990820 6 porb_h
port 681 nsew
rlabel metal1 s 179322 990768 179386 990780 6 porb_h
port 681 nsew
rlabel metal1 s 173802 990768 173866 990780 6 porb_h
port 681 nsew
rlabel metal1 s 173802 990780 179386 990808 6 porb_h
port 681 nsew
rlabel metal1 s 179322 990808 179386 990820 6 porb_h
port 681 nsew
rlabel metal1 s 173802 990808 173866 990820 6 porb_h
port 681 nsew
rlabel metal1 s 143258 990768 143322 990780 6 porb_h
port 681 nsew
rlabel metal1 s 130396 990780 143322 990808 6 porb_h
port 681 nsew
rlabel metal1 s 143258 990808 143322 990820 6 porb_h
port 681 nsew
rlabel metal1 s 463602 990836 463666 990848 6 porb_h
port 681 nsew
rlabel metal1 s 450262 990836 450326 990848 6 porb_h
port 681 nsew
rlabel metal1 s 450262 990848 463666 990876 6 porb_h
port 681 nsew
rlabel metal1 s 463602 990876 463666 990888 6 porb_h
port 681 nsew
rlabel metal1 s 450262 990876 450326 990888 6 porb_h
port 681 nsew
rlabel metal1 s 438670 990836 438734 990848 6 porb_h
port 681 nsew
rlabel metal1 s 419534 990836 419598 990848 6 porb_h
port 681 nsew
rlabel metal1 s 419534 990848 438734 990876 6 porb_h
port 681 nsew
rlabel metal1 s 130396 990808 130424 990848 6 porb_h
port 681 nsew
rlabel metal1 s 130102 990768 130166 990820 6 porb_h
port 681 nsew
rlabel metal1 s 110414 990768 110478 990780 6 porb_h
port 681 nsew
rlabel metal1 s 79042 990768 79106 990780 6 porb_h
port 681 nsew
rlabel metal1 s 79042 990780 110478 990808 6 porb_h
port 681 nsew
rlabel metal1 s 110414 990808 110478 990820 6 porb_h
port 681 nsew
rlabel metal1 s 79042 990808 79106 990820 6 porb_h
port 681 nsew
rlabel metal1 s 130286 990836 130350 990848 6 porb_h
port 681 nsew
rlabel metal1 s 130120 990820 130148 990848 6 porb_h
port 681 nsew
rlabel metal1 s 130120 990848 130424 990876 6 porb_h
port 681 nsew
rlabel metal1 s 438670 990876 438734 990888 6 porb_h
port 681 nsew
rlabel metal1 s 419534 990876 419598 990888 6 porb_h
port 681 nsew
rlabel metal1 s 130286 990876 130350 990888 6 porb_h
port 681 nsew
rlabel metal1 s 482922 992264 482986 992276 6 porb_h
port 681 nsew
rlabel metal1 s 475470 992264 475534 992276 6 porb_h
port 681 nsew
rlabel metal1 s 463786 992264 463850 992276 6 porb_h
port 681 nsew
rlabel metal1 s 463786 992276 482986 992304 6 porb_h
port 681 nsew
rlabel metal1 s 482922 992304 482986 992316 6 porb_h
port 681 nsew
rlabel metal1 s 475470 992304 475534 992316 6 porb_h
port 681 nsew
rlabel metal1 s 463786 992304 463850 992316 6 porb_h
port 681 nsew
rlabel metal5 s 133840 6675 146380 19198 6 resetb
port 682 nsew
rlabel metal3 s 141820 37046 141966 37818 6 resetb_core_h
port 683 nsew
rlabel metal3 s 141667 37818 141966 37911 6 resetb_core_h
port 683 nsew
rlabel metal3 s 141873 37911 141966 37971 6 resetb_core_h
port 683 nsew
rlabel metal3 s 141667 37911 141820 37971 6 resetb_core_h
port 683 nsew
rlabel metal3 s 141667 37971 141873 38031 6 resetb_core_h
port 683 nsew
rlabel metal3 s 141667 38031 141813 40000 6 resetb_core_h
port 683 nsew
rlabel metal5 s 698028 909409 711514 920737 6 vccd1
port 684 nsew
rlabel metal5 s 698402 819640 710925 832180 6 vdda1
port 685 nsew
rlabel metal5 s 576820 1018402 589360 1030925 6 vssa1
port 686 nsew
rlabel metal5 s 698028 461609 711514 472937 6 vssd1
port 687 nsew
rlabel metal5 s 6086 913863 19572 925191 6 vccd2
port 688 nsew
rlabel metal5 s 6675 484220 19198 496760 6 vdda2
port 689 nsew
rlabel metal5 s 6675 828820 19198 841360 6 vssa2
port 690 nsew
rlabel metal5 s 6086 442663 19572 453991 6 vssd2
port 691 nsew
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 717600 1037600
string LEFview TRUE
string GDS_FILE chip_io.gds
string GDS_END 35112252
string GDS_START 34578978
<< end >>

