magic
tech sky130A
magscale 1 2
timestamp 1624232573
<< obsli1 >>
rect 1104 2159 148856 102833
<< obsm1 >>
rect 1104 1028 149026 103012
<< metal2 >>
rect 2318 104200 2374 105000
rect 6918 104200 6974 105000
rect 11610 104200 11666 105000
rect 16302 104200 16358 105000
rect 20994 104200 21050 105000
rect 25686 104200 25742 105000
rect 30378 104200 30434 105000
rect 35070 104200 35126 105000
rect 39762 104200 39818 105000
rect 44454 104200 44510 105000
rect 49146 104200 49202 105000
rect 53838 104200 53894 105000
rect 58530 104200 58586 105000
rect 63222 104200 63278 105000
rect 67914 104200 67970 105000
rect 72606 104200 72662 105000
rect 77298 104200 77354 105000
rect 81898 104200 81954 105000
rect 86590 104200 86646 105000
rect 91282 104200 91338 105000
rect 95974 104200 96030 105000
rect 100666 104200 100722 105000
rect 105358 104200 105414 105000
rect 110050 104200 110106 105000
rect 114742 104200 114798 105000
rect 119434 104200 119490 105000
rect 124126 104200 124182 105000
rect 128818 104200 128874 105000
rect 133510 104200 133566 105000
rect 138202 104200 138258 105000
rect 142894 104200 142950 105000
rect 147586 104200 147642 105000
rect 2318 0 2374 800
rect 6918 0 6974 800
rect 11610 0 11666 800
rect 16302 0 16358 800
rect 20994 0 21050 800
rect 25686 0 25742 800
rect 30378 0 30434 800
rect 35070 0 35126 800
rect 39762 0 39818 800
rect 44454 0 44510 800
rect 49146 0 49202 800
rect 53838 0 53894 800
rect 58530 0 58586 800
rect 63222 0 63278 800
rect 67914 0 67970 800
rect 72606 0 72662 800
rect 77298 0 77354 800
rect 81898 0 81954 800
rect 86590 0 86646 800
rect 91282 0 91338 800
rect 95974 0 96030 800
rect 100666 0 100722 800
rect 105358 0 105414 800
rect 110050 0 110106 800
rect 114742 0 114798 800
rect 119434 0 119490 800
rect 124126 0 124182 800
rect 128818 0 128874 800
rect 133510 0 133566 800
rect 138202 0 138258 800
rect 142894 0 142950 800
rect 147586 0 147642 800
<< obsm2 >>
rect 1400 104144 2262 104200
rect 2430 104144 6862 104200
rect 7030 104144 11554 104200
rect 11722 104144 16246 104200
rect 16414 104144 20938 104200
rect 21106 104144 25630 104200
rect 25798 104144 30322 104200
rect 30490 104144 35014 104200
rect 35182 104144 39706 104200
rect 39874 104144 44398 104200
rect 44566 104144 49090 104200
rect 49258 104144 53782 104200
rect 53950 104144 58474 104200
rect 58642 104144 63166 104200
rect 63334 104144 67858 104200
rect 68026 104144 72550 104200
rect 72718 104144 77242 104200
rect 77410 104144 81842 104200
rect 82010 104144 86534 104200
rect 86702 104144 91226 104200
rect 91394 104144 95918 104200
rect 96086 104144 100610 104200
rect 100778 104144 105302 104200
rect 105470 104144 109994 104200
rect 110162 104144 114686 104200
rect 114854 104144 119378 104200
rect 119546 104144 124070 104200
rect 124238 104144 128762 104200
rect 128930 104144 133454 104200
rect 133622 104144 138146 104200
rect 138314 104144 142838 104200
rect 143006 104144 147530 104200
rect 147698 104144 149020 104200
rect 1400 856 149020 104144
rect 1400 800 2262 856
rect 2430 800 6862 856
rect 7030 800 11554 856
rect 11722 800 16246 856
rect 16414 800 20938 856
rect 21106 800 25630 856
rect 25798 800 30322 856
rect 30490 800 35014 856
rect 35182 800 39706 856
rect 39874 800 44398 856
rect 44566 800 49090 856
rect 49258 800 53782 856
rect 53950 800 58474 856
rect 58642 800 63166 856
rect 63334 800 67858 856
rect 68026 800 72550 856
rect 72718 800 77242 856
rect 77410 800 81842 856
rect 82010 800 86534 856
rect 86702 800 91226 856
rect 91394 800 95918 856
rect 96086 800 100610 856
rect 100778 800 105302 856
rect 105470 800 109994 856
rect 110162 800 114686 856
rect 114854 800 119378 856
rect 119546 800 124070 856
rect 124238 800 128762 856
rect 128930 800 133454 856
rect 133622 800 138146 856
rect 138314 800 142838 856
rect 143006 800 147530 856
rect 147698 800 149020 856
<< metal3 >>
rect 0 101056 800 101176
rect 0 93576 800 93696
rect 0 86096 800 86216
rect 0 78616 800 78736
rect 0 71136 800 71256
rect 0 63656 800 63776
rect 0 56176 800 56296
rect 0 48560 800 48680
rect 0 41080 800 41200
rect 0 33600 800 33720
rect 0 26120 800 26240
rect 0 18640 800 18760
rect 0 11160 800 11280
rect 0 3680 800 3800
<< obsm3 >>
rect 800 101256 147831 102849
rect 880 100976 147831 101256
rect 800 93776 147831 100976
rect 880 93496 147831 93776
rect 800 86296 147831 93496
rect 880 86016 147831 86296
rect 800 78816 147831 86016
rect 880 78536 147831 78816
rect 800 71336 147831 78536
rect 880 71056 147831 71336
rect 800 63856 147831 71056
rect 880 63576 147831 63856
rect 800 56376 147831 63576
rect 880 56096 147831 56376
rect 800 48760 147831 56096
rect 880 48480 147831 48760
rect 800 41280 147831 48480
rect 880 41000 147831 41280
rect 800 33800 147831 41000
rect 880 33520 147831 33800
rect 800 26320 147831 33520
rect 880 26040 147831 26320
rect 800 18840 147831 26040
rect 880 18560 147831 18840
rect 800 11360 147831 18560
rect 880 11080 147831 11360
rect 800 3880 147831 11080
rect 880 3600 147831 3880
rect 800 2143 147831 3600
<< metal4 >>
rect 4208 2128 4528 102864
rect 19568 2128 19888 102864
rect 34928 2128 35248 102864
rect 50288 2128 50608 102864
rect 65648 2128 65968 102864
rect 81008 2128 81328 102864
rect 96368 2128 96688 102864
rect 111728 2128 112048 102864
rect 127088 2128 127408 102864
rect 142448 2128 142768 102864
<< obsm4 >>
rect 8891 8331 19488 96525
rect 19968 8331 34848 96525
rect 35328 8331 50208 96525
rect 50688 8331 65568 96525
rect 66048 8331 80928 96525
rect 81408 8331 96288 96525
rect 96768 8331 111648 96525
rect 112128 8331 127008 96525
rect 127488 8331 142368 96525
rect 142848 8331 143461 96525
<< labels >>
rlabel metal3 s 0 3680 800 3800 6 A[0]
port 1 nsew signal input
rlabel metal3 s 0 11160 800 11280 6 A[1]
port 2 nsew signal input
rlabel metal3 s 0 18640 800 18760 6 A[2]
port 3 nsew signal input
rlabel metal3 s 0 26120 800 26240 6 A[3]
port 4 nsew signal input
rlabel metal3 s 0 33600 800 33720 6 A[4]
port 5 nsew signal input
rlabel metal3 s 0 41080 800 41200 6 A[5]
port 6 nsew signal input
rlabel metal3 s 0 48560 800 48680 6 A[6]
port 7 nsew signal input
rlabel metal3 s 0 56176 800 56296 6 A[7]
port 8 nsew signal input
rlabel metal3 s 0 63656 800 63776 6 CLK
port 9 nsew signal input
rlabel metal2 s 2318 104200 2374 105000 6 Di[0]
port 10 nsew signal input
rlabel metal2 s 49146 104200 49202 105000 6 Di[10]
port 11 nsew signal input
rlabel metal2 s 53838 104200 53894 105000 6 Di[11]
port 12 nsew signal input
rlabel metal2 s 58530 104200 58586 105000 6 Di[12]
port 13 nsew signal input
rlabel metal2 s 63222 104200 63278 105000 6 Di[13]
port 14 nsew signal input
rlabel metal2 s 67914 104200 67970 105000 6 Di[14]
port 15 nsew signal input
rlabel metal2 s 72606 104200 72662 105000 6 Di[15]
port 16 nsew signal input
rlabel metal2 s 77298 104200 77354 105000 6 Di[16]
port 17 nsew signal input
rlabel metal2 s 81898 104200 81954 105000 6 Di[17]
port 18 nsew signal input
rlabel metal2 s 86590 104200 86646 105000 6 Di[18]
port 19 nsew signal input
rlabel metal2 s 91282 104200 91338 105000 6 Di[19]
port 20 nsew signal input
rlabel metal2 s 6918 104200 6974 105000 6 Di[1]
port 21 nsew signal input
rlabel metal2 s 95974 104200 96030 105000 6 Di[20]
port 22 nsew signal input
rlabel metal2 s 100666 104200 100722 105000 6 Di[21]
port 23 nsew signal input
rlabel metal2 s 105358 104200 105414 105000 6 Di[22]
port 24 nsew signal input
rlabel metal2 s 110050 104200 110106 105000 6 Di[23]
port 25 nsew signal input
rlabel metal2 s 114742 104200 114798 105000 6 Di[24]
port 26 nsew signal input
rlabel metal2 s 119434 104200 119490 105000 6 Di[25]
port 27 nsew signal input
rlabel metal2 s 124126 104200 124182 105000 6 Di[26]
port 28 nsew signal input
rlabel metal2 s 128818 104200 128874 105000 6 Di[27]
port 29 nsew signal input
rlabel metal2 s 133510 104200 133566 105000 6 Di[28]
port 30 nsew signal input
rlabel metal2 s 138202 104200 138258 105000 6 Di[29]
port 31 nsew signal input
rlabel metal2 s 11610 104200 11666 105000 6 Di[2]
port 32 nsew signal input
rlabel metal2 s 142894 104200 142950 105000 6 Di[30]
port 33 nsew signal input
rlabel metal2 s 147586 104200 147642 105000 6 Di[31]
port 34 nsew signal input
rlabel metal2 s 16302 104200 16358 105000 6 Di[3]
port 35 nsew signal input
rlabel metal2 s 20994 104200 21050 105000 6 Di[4]
port 36 nsew signal input
rlabel metal2 s 25686 104200 25742 105000 6 Di[5]
port 37 nsew signal input
rlabel metal2 s 30378 104200 30434 105000 6 Di[6]
port 38 nsew signal input
rlabel metal2 s 35070 104200 35126 105000 6 Di[7]
port 39 nsew signal input
rlabel metal2 s 39762 104200 39818 105000 6 Di[8]
port 40 nsew signal input
rlabel metal2 s 44454 104200 44510 105000 6 Di[9]
port 41 nsew signal input
rlabel metal2 s 2318 0 2374 800 6 Do[0]
port 42 nsew signal output
rlabel metal2 s 49146 0 49202 800 6 Do[10]
port 43 nsew signal output
rlabel metal2 s 53838 0 53894 800 6 Do[11]
port 44 nsew signal output
rlabel metal2 s 58530 0 58586 800 6 Do[12]
port 45 nsew signal output
rlabel metal2 s 63222 0 63278 800 6 Do[13]
port 46 nsew signal output
rlabel metal2 s 67914 0 67970 800 6 Do[14]
port 47 nsew signal output
rlabel metal2 s 72606 0 72662 800 6 Do[15]
port 48 nsew signal output
rlabel metal2 s 77298 0 77354 800 6 Do[16]
port 49 nsew signal output
rlabel metal2 s 81898 0 81954 800 6 Do[17]
port 50 nsew signal output
rlabel metal2 s 86590 0 86646 800 6 Do[18]
port 51 nsew signal output
rlabel metal2 s 91282 0 91338 800 6 Do[19]
port 52 nsew signal output
rlabel metal2 s 6918 0 6974 800 6 Do[1]
port 53 nsew signal output
rlabel metal2 s 95974 0 96030 800 6 Do[20]
port 54 nsew signal output
rlabel metal2 s 100666 0 100722 800 6 Do[21]
port 55 nsew signal output
rlabel metal2 s 105358 0 105414 800 6 Do[22]
port 56 nsew signal output
rlabel metal2 s 110050 0 110106 800 6 Do[23]
port 57 nsew signal output
rlabel metal2 s 114742 0 114798 800 6 Do[24]
port 58 nsew signal output
rlabel metal2 s 119434 0 119490 800 6 Do[25]
port 59 nsew signal output
rlabel metal2 s 124126 0 124182 800 6 Do[26]
port 60 nsew signal output
rlabel metal2 s 128818 0 128874 800 6 Do[27]
port 61 nsew signal output
rlabel metal2 s 133510 0 133566 800 6 Do[28]
port 62 nsew signal output
rlabel metal2 s 138202 0 138258 800 6 Do[29]
port 63 nsew signal output
rlabel metal2 s 11610 0 11666 800 6 Do[2]
port 64 nsew signal output
rlabel metal2 s 142894 0 142950 800 6 Do[30]
port 65 nsew signal output
rlabel metal2 s 147586 0 147642 800 6 Do[31]
port 66 nsew signal output
rlabel metal2 s 16302 0 16358 800 6 Do[3]
port 67 nsew signal output
rlabel metal2 s 20994 0 21050 800 6 Do[4]
port 68 nsew signal output
rlabel metal2 s 25686 0 25742 800 6 Do[5]
port 69 nsew signal output
rlabel metal2 s 30378 0 30434 800 6 Do[6]
port 70 nsew signal output
rlabel metal2 s 35070 0 35126 800 6 Do[7]
port 71 nsew signal output
rlabel metal2 s 39762 0 39818 800 6 Do[8]
port 72 nsew signal output
rlabel metal2 s 44454 0 44510 800 6 Do[9]
port 73 nsew signal output
rlabel metal3 s 0 101056 800 101176 6 EN
port 74 nsew signal input
rlabel metal3 s 0 71136 800 71256 6 WE[0]
port 75 nsew signal input
rlabel metal3 s 0 78616 800 78736 6 WE[1]
port 76 nsew signal input
rlabel metal3 s 0 86096 800 86216 6 WE[2]
port 77 nsew signal input
rlabel metal3 s 0 93576 800 93696 6 WE[3]
port 78 nsew signal input
rlabel metal4 s 127088 2128 127408 102864 6 VPWR
port 79 nsew power bidirectional
rlabel metal4 s 96368 2128 96688 102864 6 VPWR
port 80 nsew power bidirectional
rlabel metal4 s 65648 2128 65968 102864 6 VPWR
port 81 nsew power bidirectional
rlabel metal4 s 34928 2128 35248 102864 6 VPWR
port 82 nsew power bidirectional
rlabel metal4 s 4208 2128 4528 102864 6 VPWR
port 83 nsew power bidirectional
rlabel metal4 s 142448 2128 142768 102864 6 VGND
port 84 nsew ground bidirectional
rlabel metal4 s 111728 2128 112048 102864 6 VGND
port 85 nsew ground bidirectional
rlabel metal4 s 81008 2128 81328 102864 6 VGND
port 86 nsew ground bidirectional
rlabel metal4 s 50288 2128 50608 102864 6 VGND
port 87 nsew ground bidirectional
rlabel metal4 s 19568 2128 19888 102864 6 VGND
port 88 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 150000 105000
string LEFview TRUE
string GDS_FILE ../gds/DFFRAM.gds
string GDS_END 61631538
string GDS_START 181858
<< end >>

