.subckt sky130_fd_pr__diode_pw2nd_11v0 A C a=1 p=1
D A C  sky130_fd_pr__diode_pw2nd_11v0 area={a}
.ends
