magic
tech sky130A
magscale 1 2
timestamp 1633363087
<< isosubstrate >>
rect 988 2232 3818 5400
<< locali >>
rect 7113 5151 7147 5321
<< viali >>
rect 7205 11169 7239 11203
rect 7573 11169 7607 11203
rect 8861 11169 8895 11203
rect 9045 11169 9079 11203
rect 8217 11101 8251 11135
rect 7297 11033 7331 11067
rect 8125 11033 8159 11067
rect 9229 11033 9263 11067
rect 9137 10693 9171 10727
rect 6837 10625 6871 10659
rect 6285 10557 6319 10591
rect 8762 10557 8796 10591
rect 8953 10557 8987 10591
rect 9321 10557 9355 10591
rect 8493 10489 8527 10523
rect 6469 10421 6503 10455
rect 7021 10421 7055 10455
rect 9505 10421 9539 10455
rect 6101 10217 6135 10251
rect 9505 10217 9539 10251
rect 5917 10081 5951 10115
rect 6377 10081 6411 10115
rect 6745 10081 6779 10115
rect 7757 10081 7791 10115
rect 9321 10081 9355 10115
rect 7395 10013 7429 10047
rect 6561 9877 6595 9911
rect 7297 9877 7331 9911
rect 9137 9877 9171 9911
rect 7205 9537 7239 9571
rect 5089 9469 5123 9503
rect 6929 9469 6963 9503
rect 9045 9469 9079 9503
rect 9505 9469 9539 9503
rect 9137 9401 9171 9435
rect 6377 9333 6411 9367
rect 8677 9333 8711 9367
rect 8033 9129 8067 9163
rect 8953 9061 8987 9095
rect 5273 8993 5307 9027
rect 5365 8993 5399 9027
rect 5641 8993 5675 9027
rect 5917 8993 5951 9027
rect 6285 8993 6319 9027
rect 8217 8993 8251 9027
rect 9045 8993 9079 9027
rect 6561 8925 6595 8959
rect 9229 8925 9263 8959
rect 5825 8857 5859 8891
rect 8401 8857 8435 8891
rect 5089 8789 5123 8823
rect 5549 8789 5583 8823
rect 6101 8789 6135 8823
rect 8585 8789 8619 8823
rect 7849 8585 7883 8619
rect 8769 8517 8803 8551
rect 9321 8517 9355 8551
rect 4445 8449 4479 8483
rect 8125 8449 8159 8483
rect 4169 8381 4203 8415
rect 6101 8381 6135 8415
rect 8953 8381 8987 8415
rect 6377 8313 6411 8347
rect 9137 8313 9171 8347
rect 5917 8245 5951 8279
rect 8493 8041 8527 8075
rect 8953 8041 8987 8075
rect 6292 7905 6326 7939
rect 4261 7837 4295 7871
rect 4537 7837 4571 7871
rect 6009 7837 6043 7871
rect 6561 7837 6595 7871
rect 8677 7837 8711 7871
rect 8861 7837 8895 7871
rect 8033 7769 8067 7803
rect 9321 7701 9355 7735
rect 4077 7497 4111 7531
rect 8677 7429 8711 7463
rect 4169 7361 4203 7395
rect 4445 7361 4479 7395
rect 6377 7361 6411 7395
rect 7849 7361 7883 7395
rect 3893 7293 3927 7327
rect 6101 7293 6135 7327
rect 9045 7293 9079 7327
rect 9321 7293 9355 7327
rect 9603 7289 9637 7323
rect 9811 7293 9845 7327
rect 8125 7225 8159 7259
rect 8217 7225 8251 7259
rect 9229 7225 9263 7259
rect 5917 7157 5951 7191
rect 7021 6953 7055 6987
rect 8953 6885 8987 6919
rect 2605 6817 2639 6851
rect 4077 6817 4111 6851
rect 4261 6817 4295 6851
rect 6285 6817 6319 6851
rect 6561 6817 6595 6851
rect 6837 6817 6871 6851
rect 7113 6817 7147 6851
rect 9137 6817 9171 6851
rect 9229 6817 9263 6851
rect 9413 6817 9447 6851
rect 9609 6825 9643 6859
rect 9793 6809 9827 6843
rect 4537 6749 4571 6783
rect 6009 6749 6043 6783
rect 7481 6749 7515 6783
rect 4077 6681 4111 6715
rect 6745 6681 6779 6715
rect 6469 6613 6503 6647
rect 3985 6409 4019 6443
rect 3341 6341 3375 6375
rect 9229 6341 9263 6375
rect 4353 6273 4387 6307
rect 4629 6273 4663 6307
rect 6745 6273 6779 6307
rect 8217 6273 8251 6307
rect 3525 6205 3559 6239
rect 3801 6205 3835 6239
rect 4077 6205 4111 6239
rect 6469 6205 6503 6239
rect 8401 6205 8435 6239
rect 8677 6205 8711 6239
rect 9045 6205 9079 6239
rect 9321 6205 9355 6239
rect 4261 6069 4295 6103
rect 6101 6069 6135 6103
rect 8585 6069 8619 6103
rect 8861 6069 8895 6103
rect 9505 6069 9539 6103
rect 4353 5729 4387 5763
rect 6285 5729 6319 5763
rect 6561 5729 6595 5763
rect 6837 5729 6871 5763
rect 7113 5729 7147 5763
rect 4629 5661 4663 5695
rect 7389 5661 7423 5695
rect 7757 5661 7791 5695
rect 6101 5593 6135 5627
rect 6469 5525 6503 5559
rect 6745 5525 6779 5559
rect 7021 5525 7055 5559
rect 7297 5525 7331 5559
rect 9137 5525 9171 5559
rect 4537 5321 4571 5355
rect 7113 5321 7147 5355
rect 9321 5321 9355 5355
rect 4629 5185 4663 5219
rect 4905 5185 4939 5219
rect 7573 5185 7607 5219
rect 4353 5117 4387 5151
rect 6837 5117 6871 5151
rect 7113 5117 7147 5151
rect 7205 5117 7239 5151
rect 9137 5117 9171 5151
rect 9045 5049 9079 5083
rect 6377 4981 6411 5015
rect 7021 4981 7055 5015
rect 6193 4777 6227 4811
rect 6929 4709 6963 4743
rect 4445 4641 4479 4675
rect 6377 4641 6411 4675
rect 8769 4641 8803 4675
rect 9229 4641 9263 4675
rect 4721 4573 4755 4607
rect 6653 4573 6687 4607
rect 8401 4505 8435 4539
rect 6561 4437 6595 4471
rect 9137 4437 9171 4471
rect 6561 4097 6595 4131
rect 9321 4097 9355 4131
rect 4537 4029 4571 4063
rect 4813 4029 4847 4063
rect 9137 4029 9171 4063
rect 5089 3961 5123 3995
rect 9229 3961 9263 3995
rect 4721 3893 4755 3927
rect 8585 3893 8619 3927
rect 8769 3893 8803 3927
rect 6469 3689 6503 3723
rect 9045 3689 9079 3723
rect 6929 3621 6963 3655
rect 4721 3553 4755 3587
rect 6653 3553 6687 3587
rect 8585 3553 8619 3587
rect 8861 3553 8895 3587
rect 4997 3485 5031 3519
rect 8401 3485 8435 3519
rect 8769 3349 8803 3383
rect 6561 3145 6595 3179
rect 6929 3145 6963 3179
rect 8769 3145 8803 3179
rect 4813 3009 4847 3043
rect 5089 3009 5123 3043
rect 9229 3009 9263 3043
rect 9413 3009 9447 3043
rect 6837 2941 6871 2975
rect 7113 2941 7147 2975
rect 7573 2941 7607 2975
rect 7389 2873 7423 2907
rect 7297 2805 7331 2839
rect 8677 2805 8711 2839
rect 9137 2805 9171 2839
rect 8585 2601 8619 2635
rect 5089 2533 5123 2567
rect 4813 2397 4847 2431
rect 6837 2397 6871 2431
rect 7113 2397 7147 2431
rect 6561 2261 6595 2295
<< metal1 >>
rect 9674 13200 9680 13252
rect 9732 13240 9738 13252
rect 14182 13240 14188 13252
rect 9732 13212 14188 13240
rect 9732 13200 9738 13212
rect 14182 13200 14188 13212
rect 14240 13200 14246 13252
rect 9490 12656 9496 12708
rect 9548 12696 9554 12708
rect 14182 12696 14188 12708
rect 9548 12668 14188 12696
rect 9548 12656 9554 12668
rect 14182 12656 14188 12668
rect 14240 12656 14246 12708
rect 13078 12452 13084 12504
rect 13136 12492 13142 12504
rect 14182 12492 14188 12504
rect 13136 12464 14188 12492
rect 13136 12452 13142 12464
rect 14182 12452 14188 12464
rect 14240 12452 14246 12504
rect 920 11450 9844 11472
rect 920 11398 2748 11450
rect 2800 11398 2812 11450
rect 2864 11398 2876 11450
rect 2928 11398 2940 11450
rect 2992 11398 5848 11450
rect 5900 11398 5912 11450
rect 5964 11398 5976 11450
rect 6028 11398 6040 11450
rect 6092 11398 8948 11450
rect 9000 11398 9012 11450
rect 9064 11398 9076 11450
rect 9128 11398 9140 11450
rect 9192 11398 9844 11450
rect 920 11376 9844 11398
rect 8662 11268 8668 11280
rect 7208 11240 8668 11268
rect 7208 11209 7236 11240
rect 8662 11228 8668 11240
rect 8720 11228 8726 11280
rect 7193 11203 7251 11209
rect 7193 11169 7205 11203
rect 7239 11169 7251 11203
rect 7193 11163 7251 11169
rect 7561 11203 7619 11209
rect 7561 11169 7573 11203
rect 7607 11200 7619 11203
rect 8849 11203 8907 11209
rect 8849 11200 8861 11203
rect 7607 11172 8861 11200
rect 7607 11169 7619 11172
rect 7561 11163 7619 11169
rect 8849 11169 8861 11172
rect 8895 11169 8907 11203
rect 8849 11163 8907 11169
rect 8938 11160 8944 11212
rect 8996 11200 9002 11212
rect 9033 11203 9091 11209
rect 9033 11200 9045 11203
rect 8996 11172 9045 11200
rect 8996 11160 9002 11172
rect 9033 11169 9045 11172
rect 9079 11200 9091 11203
rect 9582 11200 9588 11212
rect 9079 11172 9588 11200
rect 9079 11169 9091 11172
rect 9033 11163 9091 11169
rect 9582 11160 9588 11172
rect 9640 11160 9646 11212
rect 13170 11160 13176 11212
rect 13228 11200 13234 11212
rect 14182 11200 14188 11212
rect 13228 11172 14188 11200
rect 13228 11160 13234 11172
rect 14182 11160 14188 11172
rect 14240 11160 14246 11212
rect 8018 11092 8024 11144
rect 8076 11132 8082 11144
rect 8205 11135 8263 11141
rect 8205 11132 8217 11135
rect 8076 11104 8217 11132
rect 8076 11092 8082 11104
rect 8205 11101 8217 11104
rect 8251 11101 8263 11135
rect 8205 11095 8263 11101
rect 4614 11024 4620 11076
rect 4672 11064 4678 11076
rect 7285 11067 7343 11073
rect 7285 11064 7297 11067
rect 4672 11036 7297 11064
rect 4672 11024 4678 11036
rect 7285 11033 7297 11036
rect 7331 11033 7343 11067
rect 8110 11064 8116 11076
rect 8071 11036 8116 11064
rect 7285 11027 7343 11033
rect 8110 11024 8116 11036
rect 8168 11024 8174 11076
rect 9217 11067 9275 11073
rect 9217 11033 9229 11067
rect 9263 11064 9275 11067
rect 14182 11064 14188 11076
rect 9263 11036 14188 11064
rect 9263 11033 9275 11036
rect 9217 11027 9275 11033
rect 14182 11024 14188 11036
rect 14240 11024 14246 11076
rect 920 10906 9844 10928
rect 920 10854 1198 10906
rect 1250 10854 1262 10906
rect 1314 10854 1326 10906
rect 1378 10854 1390 10906
rect 1442 10854 4298 10906
rect 4350 10854 4362 10906
rect 4414 10854 4426 10906
rect 4478 10854 4490 10906
rect 4542 10854 7398 10906
rect 7450 10854 7462 10906
rect 7514 10854 7526 10906
rect 7578 10854 7590 10906
rect 7642 10854 9844 10906
rect 920 10832 9844 10854
rect 6472 10764 9076 10792
rect 6270 10588 6276 10600
rect 6183 10560 6276 10588
rect 6270 10548 6276 10560
rect 6328 10588 6334 10600
rect 6472 10588 6500 10764
rect 8938 10724 8944 10736
rect 8772 10696 8944 10724
rect 6825 10659 6883 10665
rect 6825 10625 6837 10659
rect 6871 10656 6883 10659
rect 8386 10656 8392 10668
rect 6871 10628 8392 10656
rect 6871 10625 6883 10628
rect 6825 10619 6883 10625
rect 8386 10616 8392 10628
rect 8444 10616 8450 10668
rect 8772 10597 8800 10696
rect 8938 10684 8944 10696
rect 8996 10684 9002 10736
rect 6328 10560 6500 10588
rect 8750 10591 8808 10597
rect 6328 10548 6334 10560
rect 8750 10557 8762 10591
rect 8796 10557 8808 10591
rect 8938 10588 8944 10600
rect 8899 10560 8944 10588
rect 8750 10551 8808 10557
rect 8938 10548 8944 10560
rect 8996 10548 9002 10600
rect 9048 10588 9076 10764
rect 9125 10727 9183 10733
rect 9125 10693 9137 10727
rect 9171 10724 9183 10727
rect 14182 10724 14188 10736
rect 9171 10696 14188 10724
rect 9171 10693 9183 10696
rect 9125 10687 9183 10693
rect 14182 10684 14188 10696
rect 14240 10684 14246 10736
rect 9309 10591 9367 10597
rect 9309 10588 9321 10591
rect 9048 10560 9321 10588
rect 9309 10557 9321 10560
rect 9355 10557 9367 10591
rect 9309 10551 9367 10557
rect 8386 10520 8392 10532
rect 8050 10492 8392 10520
rect 8386 10480 8392 10492
rect 8444 10480 8450 10532
rect 8481 10523 8539 10529
rect 8481 10489 8493 10523
rect 8527 10520 8539 10523
rect 8570 10520 8576 10532
rect 8527 10492 8576 10520
rect 8527 10489 8539 10492
rect 8481 10483 8539 10489
rect 8570 10480 8576 10492
rect 8628 10520 8634 10532
rect 14274 10520 14280 10532
rect 8628 10492 14280 10520
rect 8628 10480 8634 10492
rect 14274 10480 14280 10492
rect 14332 10480 14338 10532
rect 6454 10452 6460 10464
rect 6415 10424 6460 10452
rect 6454 10412 6460 10424
rect 6512 10412 6518 10464
rect 7009 10455 7067 10461
rect 7009 10421 7021 10455
rect 7055 10452 7067 10455
rect 7190 10452 7196 10464
rect 7055 10424 7196 10452
rect 7055 10421 7067 10424
rect 7009 10415 7067 10421
rect 7190 10412 7196 10424
rect 7248 10412 7254 10464
rect 8294 10412 8300 10464
rect 8352 10452 8358 10464
rect 9493 10455 9551 10461
rect 9493 10452 9505 10455
rect 8352 10424 9505 10452
rect 8352 10412 8358 10424
rect 9493 10421 9505 10424
rect 9539 10421 9551 10455
rect 9493 10415 9551 10421
rect 920 10362 9844 10384
rect 920 10310 2748 10362
rect 2800 10310 2812 10362
rect 2864 10310 2876 10362
rect 2928 10310 2940 10362
rect 2992 10310 5848 10362
rect 5900 10310 5912 10362
rect 5964 10310 5976 10362
rect 6028 10310 6040 10362
rect 6092 10310 8948 10362
rect 9000 10310 9012 10362
rect 9064 10310 9076 10362
rect 9128 10310 9140 10362
rect 9192 10310 9844 10362
rect 920 10288 9844 10310
rect 6089 10251 6147 10257
rect 6089 10217 6101 10251
rect 6135 10248 6147 10251
rect 6135 10220 8156 10248
rect 6135 10217 6147 10220
rect 6089 10211 6147 10217
rect 7466 10180 7472 10192
rect 6380 10152 7472 10180
rect 5905 10115 5963 10121
rect 5905 10081 5917 10115
rect 5951 10112 5963 10115
rect 6270 10112 6276 10124
rect 5951 10084 6276 10112
rect 5951 10081 5963 10084
rect 5905 10075 5963 10081
rect 6270 10072 6276 10084
rect 6328 10072 6334 10124
rect 6380 10121 6408 10152
rect 7466 10140 7472 10152
rect 7524 10140 7530 10192
rect 8128 10166 8156 10220
rect 8386 10208 8392 10260
rect 8444 10248 8450 10260
rect 9493 10251 9551 10257
rect 9493 10248 9505 10251
rect 8444 10220 9505 10248
rect 8444 10208 8450 10220
rect 9493 10217 9505 10220
rect 9539 10217 9551 10251
rect 9493 10211 9551 10217
rect 6365 10115 6423 10121
rect 6365 10081 6377 10115
rect 6411 10081 6423 10115
rect 6730 10112 6736 10124
rect 6691 10084 6736 10112
rect 6365 10075 6423 10081
rect 6730 10072 6736 10084
rect 6788 10072 6794 10124
rect 7190 10072 7196 10124
rect 7248 10112 7254 10124
rect 7745 10115 7803 10121
rect 7745 10112 7757 10115
rect 7248 10084 7757 10112
rect 7248 10072 7254 10084
rect 7745 10081 7757 10084
rect 7791 10081 7803 10115
rect 7745 10075 7803 10081
rect 8570 10072 8576 10124
rect 8628 10112 8634 10124
rect 9309 10115 9367 10121
rect 9309 10112 9321 10115
rect 8628 10084 9321 10112
rect 8628 10072 8634 10084
rect 9309 10081 9321 10084
rect 9355 10081 9367 10115
rect 9309 10075 9367 10081
rect 7098 10044 7104 10056
rect 6380 10016 7104 10044
rect 6380 9988 6408 10016
rect 7098 10004 7104 10016
rect 7156 10044 7162 10056
rect 7383 10047 7441 10053
rect 7383 10044 7395 10047
rect 7156 10016 7395 10044
rect 7156 10004 7162 10016
rect 7383 10013 7395 10016
rect 7429 10013 7441 10047
rect 7383 10007 7441 10013
rect 6362 9936 6368 9988
rect 6420 9936 6426 9988
rect 6546 9908 6552 9920
rect 6507 9880 6552 9908
rect 6546 9868 6552 9880
rect 6604 9868 6610 9920
rect 7285 9911 7343 9917
rect 7285 9877 7297 9911
rect 7331 9908 7343 9911
rect 8110 9908 8116 9920
rect 7331 9880 8116 9908
rect 7331 9877 7343 9880
rect 7285 9871 7343 9877
rect 8110 9868 8116 9880
rect 8168 9868 8174 9920
rect 9125 9911 9183 9917
rect 9125 9877 9137 9911
rect 9171 9908 9183 9911
rect 9306 9908 9312 9920
rect 9171 9880 9312 9908
rect 9171 9877 9183 9880
rect 9125 9871 9183 9877
rect 9306 9868 9312 9880
rect 9364 9868 9370 9920
rect 920 9818 9844 9840
rect 920 9766 1198 9818
rect 1250 9766 1262 9818
rect 1314 9766 1326 9818
rect 1378 9766 1390 9818
rect 1442 9766 4298 9818
rect 4350 9766 4362 9818
rect 4414 9766 4426 9818
rect 4478 9766 4490 9818
rect 4542 9766 7398 9818
rect 7450 9766 7462 9818
rect 7514 9766 7526 9818
rect 7578 9766 7590 9818
rect 7642 9766 9844 9818
rect 920 9744 9844 9766
rect 14366 9704 14372 9716
rect 7024 9676 14372 9704
rect 7024 9568 7052 9676
rect 14366 9664 14372 9676
rect 14424 9664 14430 9716
rect 8202 9596 8208 9648
rect 8260 9636 8266 9648
rect 8260 9608 8708 9636
rect 8260 9596 8266 9608
rect 7190 9568 7196 9580
rect 5092 9540 7052 9568
rect 7151 9540 7196 9568
rect 5092 9509 5120 9540
rect 7190 9528 7196 9540
rect 7248 9528 7254 9580
rect 7282 9528 7288 9580
rect 7340 9568 7346 9580
rect 8680 9568 8708 9608
rect 8846 9596 8852 9648
rect 8904 9636 8910 9648
rect 14182 9636 14188 9648
rect 8904 9608 14188 9636
rect 8904 9596 8910 9608
rect 14182 9596 14188 9608
rect 14240 9596 14246 9648
rect 7340 9540 8524 9568
rect 8680 9540 9076 9568
rect 7340 9528 7346 9540
rect 5077 9503 5135 9509
rect 5077 9469 5089 9503
rect 5123 9469 5135 9503
rect 5077 9463 5135 9469
rect 5350 9460 5356 9512
rect 5408 9500 5414 9512
rect 6917 9503 6975 9509
rect 6917 9500 6929 9503
rect 5408 9472 6929 9500
rect 5408 9460 5414 9472
rect 6917 9469 6929 9472
rect 6963 9469 6975 9503
rect 6917 9463 6975 9469
rect 6546 9392 6552 9444
rect 6604 9432 6610 9444
rect 8496 9432 8524 9540
rect 9048 9509 9076 9540
rect 9033 9503 9091 9509
rect 9033 9469 9045 9503
rect 9079 9469 9091 9503
rect 9033 9463 9091 9469
rect 9493 9503 9551 9509
rect 9493 9469 9505 9503
rect 9539 9500 9551 9503
rect 9582 9500 9588 9512
rect 9539 9472 9588 9500
rect 9539 9469 9551 9472
rect 9493 9463 9551 9469
rect 9582 9460 9588 9472
rect 9640 9460 9646 9512
rect 9125 9435 9183 9441
rect 9125 9432 9137 9435
rect 6604 9404 7682 9432
rect 8496 9404 9137 9432
rect 6604 9392 6610 9404
rect 9125 9401 9137 9404
rect 9171 9401 9183 9435
rect 9125 9395 9183 9401
rect 5258 9324 5264 9376
rect 5316 9364 5322 9376
rect 6365 9367 6423 9373
rect 6365 9364 6377 9367
rect 5316 9336 6377 9364
rect 5316 9324 5322 9336
rect 6365 9333 6377 9336
rect 6411 9333 6423 9367
rect 6365 9327 6423 9333
rect 7834 9324 7840 9376
rect 7892 9364 7898 9376
rect 8665 9367 8723 9373
rect 8665 9364 8677 9367
rect 7892 9336 8677 9364
rect 7892 9324 7898 9336
rect 8665 9333 8677 9336
rect 8711 9333 8723 9367
rect 8665 9327 8723 9333
rect 920 9274 9844 9296
rect 920 9222 2748 9274
rect 2800 9222 2812 9274
rect 2864 9222 2876 9274
rect 2928 9222 2940 9274
rect 2992 9222 5848 9274
rect 5900 9222 5912 9274
rect 5964 9222 5976 9274
rect 6028 9222 6040 9274
rect 6092 9222 8948 9274
rect 9000 9222 9012 9274
rect 9064 9222 9076 9274
rect 9128 9222 9140 9274
rect 9192 9222 9844 9274
rect 920 9200 9844 9222
rect 8021 9163 8079 9169
rect 5920 9132 7880 9160
rect 4706 8984 4712 9036
rect 4764 9024 4770 9036
rect 5258 9024 5264 9036
rect 4764 8996 5264 9024
rect 4764 8984 4770 8996
rect 5258 8984 5264 8996
rect 5316 8984 5322 9036
rect 5920 9033 5948 9132
rect 6454 9052 6460 9104
rect 6512 9092 6518 9104
rect 6512 9064 7038 9092
rect 6512 9052 6518 9064
rect 5353 9027 5411 9033
rect 5353 8993 5365 9027
rect 5399 9024 5411 9027
rect 5629 9027 5687 9033
rect 5629 9024 5641 9027
rect 5399 8996 5641 9024
rect 5399 8993 5411 8996
rect 5353 8987 5411 8993
rect 5629 8993 5641 8996
rect 5675 8993 5687 9027
rect 5629 8987 5687 8993
rect 5905 9027 5963 9033
rect 5905 8993 5917 9027
rect 5951 8993 5963 9027
rect 6270 9024 6276 9036
rect 6231 8996 6276 9024
rect 5905 8987 5963 8993
rect 4154 8780 4160 8832
rect 4212 8820 4218 8832
rect 5077 8823 5135 8829
rect 5077 8820 5089 8823
rect 4212 8792 5089 8820
rect 4212 8780 4218 8792
rect 5077 8789 5089 8792
rect 5123 8820 5135 8823
rect 5350 8820 5356 8832
rect 5123 8792 5356 8820
rect 5123 8789 5135 8792
rect 5077 8783 5135 8789
rect 5350 8780 5356 8792
rect 5408 8780 5414 8832
rect 5534 8820 5540 8832
rect 5495 8792 5540 8820
rect 5534 8780 5540 8792
rect 5592 8780 5598 8832
rect 5644 8820 5672 8987
rect 6270 8984 6276 8996
rect 6328 8984 6334 9036
rect 7852 9024 7880 9132
rect 8021 9129 8033 9163
rect 8067 9160 8079 9163
rect 14182 9160 14188 9172
rect 8067 9132 14188 9160
rect 8067 9129 8079 9132
rect 8021 9123 8079 9129
rect 14182 9120 14188 9132
rect 14240 9120 14246 9172
rect 8941 9095 8999 9101
rect 8941 9061 8953 9095
rect 8987 9092 8999 9095
rect 9490 9092 9496 9104
rect 8987 9064 9496 9092
rect 8987 9061 8999 9064
rect 8941 9055 8999 9061
rect 9490 9052 9496 9064
rect 9548 9052 9554 9104
rect 8205 9027 8263 9033
rect 8205 9024 8217 9027
rect 7852 8996 8217 9024
rect 8205 8993 8217 8996
rect 8251 9024 8263 9027
rect 8846 9024 8852 9036
rect 8251 8996 8852 9024
rect 8251 8993 8263 8996
rect 8205 8987 8263 8993
rect 8846 8984 8852 8996
rect 8904 8984 8910 9036
rect 9033 9027 9091 9033
rect 9033 8993 9045 9027
rect 9079 9024 9091 9027
rect 9398 9024 9404 9036
rect 9079 8996 9404 9024
rect 9079 8993 9091 8996
rect 9033 8987 9091 8993
rect 9398 8984 9404 8996
rect 9456 8984 9462 9036
rect 6546 8956 6552 8968
rect 6507 8928 6552 8956
rect 6546 8916 6552 8928
rect 6604 8916 6610 8968
rect 8570 8956 8576 8968
rect 8404 8928 8576 8956
rect 8404 8897 8432 8928
rect 8570 8916 8576 8928
rect 8628 8916 8634 8968
rect 9217 8959 9275 8965
rect 9217 8925 9229 8959
rect 9263 8956 9275 8959
rect 9306 8956 9312 8968
rect 9263 8928 9312 8956
rect 9263 8925 9275 8928
rect 9217 8919 9275 8925
rect 9306 8916 9312 8928
rect 9364 8916 9370 8968
rect 5813 8891 5871 8897
rect 5813 8857 5825 8891
rect 5859 8888 5871 8891
rect 8389 8891 8447 8897
rect 5859 8860 6316 8888
rect 5859 8857 5871 8860
rect 5813 8851 5871 8857
rect 6089 8823 6147 8829
rect 6089 8820 6101 8823
rect 5644 8792 6101 8820
rect 6089 8789 6101 8792
rect 6135 8820 6147 8823
rect 6178 8820 6184 8832
rect 6135 8792 6184 8820
rect 6135 8789 6147 8792
rect 6089 8783 6147 8789
rect 6178 8780 6184 8792
rect 6236 8780 6242 8832
rect 6288 8820 6316 8860
rect 8389 8857 8401 8891
rect 8435 8857 8447 8891
rect 8389 8851 8447 8857
rect 6638 8820 6644 8832
rect 6288 8792 6644 8820
rect 6638 8780 6644 8792
rect 6696 8780 6702 8832
rect 8573 8823 8631 8829
rect 8573 8789 8585 8823
rect 8619 8820 8631 8823
rect 10502 8820 10508 8832
rect 8619 8792 10508 8820
rect 8619 8789 8631 8792
rect 8573 8783 8631 8789
rect 10502 8780 10508 8792
rect 10560 8780 10566 8832
rect 920 8730 9844 8752
rect 920 8678 1198 8730
rect 1250 8678 1262 8730
rect 1314 8678 1326 8730
rect 1378 8678 1390 8730
rect 1442 8678 4298 8730
rect 4350 8678 4362 8730
rect 4414 8678 4426 8730
rect 4478 8678 4490 8730
rect 4542 8678 7398 8730
rect 7450 8678 7462 8730
rect 7514 8678 7526 8730
rect 7578 8678 7590 8730
rect 7642 8678 9844 8730
rect 920 8656 9844 8678
rect 7837 8619 7895 8625
rect 7837 8585 7849 8619
rect 7883 8616 7895 8619
rect 14182 8616 14188 8628
rect 7883 8588 14188 8616
rect 7883 8585 7895 8588
rect 7837 8579 7895 8585
rect 14182 8576 14188 8588
rect 14240 8576 14246 8628
rect 8018 8508 8024 8560
rect 8076 8548 8082 8560
rect 8757 8551 8815 8557
rect 8757 8548 8769 8551
rect 8076 8520 8769 8548
rect 8076 8508 8082 8520
rect 8757 8517 8769 8520
rect 8803 8517 8815 8551
rect 8757 8511 8815 8517
rect 8846 8508 8852 8560
rect 8904 8548 8910 8560
rect 9309 8551 9367 8557
rect 9309 8548 9321 8551
rect 8904 8520 9321 8548
rect 8904 8508 8910 8520
rect 9309 8517 9321 8520
rect 9355 8517 9367 8551
rect 9309 8511 9367 8517
rect 4433 8483 4491 8489
rect 4433 8449 4445 8483
rect 4479 8480 4491 8483
rect 5166 8480 5172 8492
rect 4479 8452 5172 8480
rect 4479 8449 4491 8452
rect 4433 8443 4491 8449
rect 5166 8440 5172 8452
rect 5224 8440 5230 8492
rect 5442 8440 5448 8492
rect 5500 8480 5506 8492
rect 8110 8480 8116 8492
rect 5500 8452 7972 8480
rect 8071 8452 8116 8480
rect 5500 8440 5506 8452
rect 4154 8412 4160 8424
rect 4115 8384 4160 8412
rect 4154 8372 4160 8384
rect 4212 8372 4218 8424
rect 6086 8412 6092 8424
rect 6047 8384 6092 8412
rect 6086 8372 6092 8384
rect 6144 8372 6150 8424
rect 4890 8304 4896 8356
rect 4948 8304 4954 8356
rect 6362 8344 6368 8356
rect 6323 8316 6368 8344
rect 6362 8304 6368 8316
rect 6420 8304 6426 8356
rect 6638 8304 6644 8356
rect 6696 8344 6702 8356
rect 7944 8344 7972 8452
rect 8110 8440 8116 8452
rect 8168 8440 8174 8492
rect 8754 8372 8760 8424
rect 8812 8412 8818 8424
rect 8941 8415 8999 8421
rect 8941 8412 8953 8415
rect 8812 8384 8953 8412
rect 8812 8372 8818 8384
rect 8941 8381 8953 8384
rect 8987 8381 8999 8415
rect 8941 8375 8999 8381
rect 9125 8347 9183 8353
rect 9125 8344 9137 8347
rect 6696 8316 6854 8344
rect 7944 8316 9137 8344
rect 6696 8304 6702 8316
rect 9125 8313 9137 8316
rect 9171 8344 9183 8347
rect 9490 8344 9496 8356
rect 9171 8316 9496 8344
rect 9171 8313 9183 8316
rect 9125 8307 9183 8313
rect 9490 8304 9496 8316
rect 9548 8304 9554 8356
rect 5718 8236 5724 8288
rect 5776 8276 5782 8288
rect 5905 8279 5963 8285
rect 5905 8276 5917 8279
rect 5776 8248 5917 8276
rect 5776 8236 5782 8248
rect 5905 8245 5917 8248
rect 5951 8245 5963 8279
rect 5905 8239 5963 8245
rect 10502 8236 10508 8288
rect 10560 8276 10566 8288
rect 14182 8276 14188 8288
rect 10560 8248 14188 8276
rect 10560 8236 10566 8248
rect 14182 8236 14188 8248
rect 14240 8236 14246 8288
rect 920 8186 9844 8208
rect 920 8134 2748 8186
rect 2800 8134 2812 8186
rect 2864 8134 2876 8186
rect 2928 8134 2940 8186
rect 2992 8134 5848 8186
rect 5900 8134 5912 8186
rect 5964 8134 5976 8186
rect 6028 8134 6040 8186
rect 6092 8134 8948 8186
rect 9000 8134 9012 8186
rect 9064 8134 9076 8186
rect 9128 8134 9140 8186
rect 9192 8134 9844 8186
rect 920 8112 9844 8134
rect 5534 8032 5540 8084
rect 5592 8072 5598 8084
rect 8481 8075 8539 8081
rect 5592 8044 7052 8072
rect 5592 8032 5598 8044
rect 6822 8004 6828 8016
rect 5750 7976 6828 8004
rect 6822 7964 6828 7976
rect 6880 7964 6886 8016
rect 7024 7990 7052 8044
rect 8481 8041 8493 8075
rect 8527 8072 8539 8075
rect 8941 8075 8999 8081
rect 8941 8072 8953 8075
rect 8527 8044 8953 8072
rect 8527 8041 8539 8044
rect 8481 8035 8539 8041
rect 8941 8041 8953 8044
rect 8987 8072 8999 8075
rect 9582 8072 9588 8084
rect 8987 8044 9588 8072
rect 8987 8041 8999 8044
rect 8941 8035 8999 8041
rect 9582 8032 9588 8044
rect 9640 8032 9646 8084
rect 9306 8004 9312 8016
rect 8864 7976 9312 8004
rect 6178 7896 6184 7948
rect 6236 7936 6242 7948
rect 6280 7939 6338 7945
rect 6280 7936 6292 7939
rect 6236 7908 6292 7936
rect 6236 7896 6242 7908
rect 6280 7905 6292 7908
rect 6326 7905 6338 7939
rect 8864 7936 8892 7976
rect 9306 7964 9312 7976
rect 9364 7964 9370 8016
rect 6280 7899 6338 7905
rect 8680 7908 8892 7936
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 4249 7871 4307 7877
rect 4249 7868 4261 7871
rect 4212 7840 4261 7868
rect 4212 7828 4218 7840
rect 4249 7837 4261 7840
rect 4295 7837 4307 7871
rect 4249 7831 4307 7837
rect 4525 7871 4583 7877
rect 4525 7837 4537 7871
rect 4571 7868 4583 7871
rect 4982 7868 4988 7880
rect 4571 7840 4988 7868
rect 4571 7837 4583 7840
rect 4525 7831 4583 7837
rect 4982 7828 4988 7840
rect 5040 7828 5046 7880
rect 5166 7828 5172 7880
rect 5224 7868 5230 7880
rect 8680 7877 8708 7908
rect 5997 7871 6055 7877
rect 5997 7868 6009 7871
rect 5224 7840 6009 7868
rect 5224 7828 5230 7840
rect 5997 7837 6009 7840
rect 6043 7868 6055 7871
rect 6549 7871 6607 7877
rect 6549 7868 6561 7871
rect 6043 7840 6561 7868
rect 6043 7837 6055 7840
rect 5997 7831 6055 7837
rect 6549 7837 6561 7840
rect 6595 7837 6607 7871
rect 6549 7831 6607 7837
rect 8665 7871 8723 7877
rect 8665 7837 8677 7871
rect 8711 7837 8723 7871
rect 8846 7868 8852 7880
rect 8807 7840 8852 7868
rect 8665 7831 8723 7837
rect 8846 7828 8852 7840
rect 8904 7828 8910 7880
rect 8021 7803 8079 7809
rect 8021 7769 8033 7803
rect 8067 7800 8079 7803
rect 9582 7800 9588 7812
rect 8067 7772 9588 7800
rect 8067 7769 8079 7772
rect 8021 7763 8079 7769
rect 9582 7760 9588 7772
rect 9640 7760 9646 7812
rect 9309 7735 9367 7741
rect 9309 7701 9321 7735
rect 9355 7732 9367 7735
rect 14182 7732 14188 7744
rect 9355 7704 14188 7732
rect 9355 7701 9367 7704
rect 9309 7695 9367 7701
rect 14182 7692 14188 7704
rect 14240 7692 14246 7744
rect 920 7642 9844 7664
rect 920 7590 1198 7642
rect 1250 7590 1262 7642
rect 1314 7590 1326 7642
rect 1378 7590 1390 7642
rect 1442 7590 4298 7642
rect 4350 7590 4362 7642
rect 4414 7590 4426 7642
rect 4478 7590 4490 7642
rect 4542 7590 7398 7642
rect 7450 7590 7462 7642
rect 7514 7590 7526 7642
rect 7578 7590 7590 7642
rect 7642 7590 9844 7642
rect 920 7568 9844 7590
rect 4065 7531 4123 7537
rect 4065 7497 4077 7531
rect 4111 7528 4123 7531
rect 4890 7528 4896 7540
rect 4111 7500 4896 7528
rect 4111 7497 4123 7500
rect 4065 7491 4123 7497
rect 4890 7488 4896 7500
rect 4948 7488 4954 7540
rect 4982 7488 4988 7540
rect 5040 7528 5046 7540
rect 7834 7528 7840 7540
rect 5040 7500 7840 7528
rect 5040 7488 5046 7500
rect 7834 7488 7840 7500
rect 7892 7488 7898 7540
rect 8478 7488 8484 7540
rect 8536 7528 8542 7540
rect 14274 7528 14280 7540
rect 8536 7500 14280 7528
rect 8536 7488 8542 7500
rect 14274 7488 14280 7500
rect 14332 7488 14338 7540
rect 8294 7460 8300 7472
rect 7484 7432 8300 7460
rect 4062 7352 4068 7404
rect 4120 7392 4126 7404
rect 4157 7395 4215 7401
rect 4157 7392 4169 7395
rect 4120 7364 4169 7392
rect 4120 7352 4126 7364
rect 4157 7361 4169 7364
rect 4203 7361 4215 7395
rect 4157 7355 4215 7361
rect 4433 7395 4491 7401
rect 4433 7361 4445 7395
rect 4479 7392 4491 7395
rect 5718 7392 5724 7404
rect 4479 7364 5724 7392
rect 4479 7361 4491 7364
rect 4433 7355 4491 7361
rect 5718 7352 5724 7364
rect 5776 7392 5782 7404
rect 6365 7395 6423 7401
rect 6365 7392 6377 7395
rect 5776 7364 6377 7392
rect 5776 7352 5782 7364
rect 6365 7361 6377 7364
rect 6411 7361 6423 7395
rect 6365 7355 6423 7361
rect 3878 7324 3884 7336
rect 3839 7296 3884 7324
rect 3878 7284 3884 7296
rect 3936 7284 3942 7336
rect 6086 7324 6092 7336
rect 6047 7296 6092 7324
rect 6086 7284 6092 7296
rect 6144 7284 6150 7336
rect 7484 7310 7512 7432
rect 8294 7420 8300 7432
rect 8352 7420 8358 7472
rect 8662 7460 8668 7472
rect 8623 7432 8668 7460
rect 8662 7420 8668 7432
rect 8720 7420 8726 7472
rect 7837 7395 7895 7401
rect 7837 7361 7849 7395
rect 7883 7392 7895 7395
rect 14182 7392 14188 7404
rect 7883 7364 14188 7392
rect 7883 7361 7895 7364
rect 7837 7355 7895 7361
rect 9048 7333 9076 7364
rect 14182 7352 14188 7364
rect 14240 7352 14246 7404
rect 9033 7327 9091 7333
rect 9033 7293 9045 7327
rect 9079 7293 9091 7327
rect 9306 7324 9312 7336
rect 9267 7296 9312 7324
rect 9033 7287 9091 7293
rect 9306 7284 9312 7296
rect 9364 7284 9370 7336
rect 9597 7323 9643 7335
rect 9597 7289 9603 7323
rect 9637 7289 9643 7323
rect 9597 7277 9643 7289
rect 9799 7327 9857 7333
rect 9799 7293 9811 7327
rect 9845 7324 9857 7327
rect 9845 7296 10070 7324
rect 9845 7293 9857 7296
rect 9799 7287 9857 7293
rect 5442 7216 5448 7268
rect 5500 7216 5506 7268
rect 8110 7256 8116 7268
rect 8071 7228 8116 7256
rect 8110 7216 8116 7228
rect 8168 7216 8174 7268
rect 8205 7259 8263 7265
rect 8205 7225 8217 7259
rect 8251 7225 8263 7259
rect 8205 7219 8263 7225
rect 9217 7259 9275 7265
rect 9217 7225 9229 7259
rect 9263 7225 9275 7259
rect 9217 7219 9275 7225
rect 5718 7148 5724 7200
rect 5776 7188 5782 7200
rect 5905 7191 5963 7197
rect 5905 7188 5917 7191
rect 5776 7160 5917 7188
rect 5776 7148 5782 7160
rect 5905 7157 5917 7160
rect 5951 7157 5963 7191
rect 8220 7188 8248 7219
rect 9232 7188 9260 7219
rect 8220 7160 9260 7188
rect 9606 7212 9634 7277
rect 9606 7184 9998 7212
rect 5905 7151 5963 7157
rect 920 7098 9844 7120
rect 920 7046 2748 7098
rect 2800 7046 2812 7098
rect 2864 7046 2876 7098
rect 2928 7046 2940 7098
rect 2992 7046 5848 7098
rect 5900 7046 5912 7098
rect 5964 7046 5976 7098
rect 6028 7046 6040 7098
rect 6092 7046 8948 7098
rect 9000 7046 9012 7098
rect 9064 7046 9076 7098
rect 9128 7046 9140 7098
rect 9192 7046 9844 7098
rect 920 7024 9844 7046
rect 4614 6984 4620 6996
rect 4080 6956 4620 6984
rect 4080 6857 4108 6956
rect 4614 6944 4620 6956
rect 4672 6944 4678 6996
rect 6178 6944 6184 6996
rect 6236 6944 6242 6996
rect 6914 6944 6920 6996
rect 6972 6984 6978 6996
rect 7009 6987 7067 6993
rect 7009 6984 7021 6987
rect 6972 6956 7021 6984
rect 6972 6944 6978 6956
rect 7009 6953 7021 6956
rect 7055 6953 7067 6987
rect 7009 6947 7067 6953
rect 4154 6876 4160 6928
rect 4212 6916 4218 6928
rect 4212 6888 4292 6916
rect 4212 6876 4218 6888
rect 4264 6857 4292 6888
rect 4982 6876 4988 6928
rect 5040 6876 5046 6928
rect 6196 6916 6224 6944
rect 6638 6916 6644 6928
rect 6196 6888 6644 6916
rect 6638 6876 6644 6888
rect 6696 6916 6702 6928
rect 6696 6888 6960 6916
rect 6696 6876 6702 6888
rect 2593 6851 2651 6857
rect 2593 6817 2605 6851
rect 2639 6848 2651 6851
rect 4065 6851 4123 6857
rect 2639 6820 2774 6848
rect 2639 6817 2651 6820
rect 2593 6811 2651 6817
rect 2746 6780 2774 6820
rect 4065 6817 4077 6851
rect 4111 6817 4123 6851
rect 4065 6811 4123 6817
rect 4249 6851 4307 6857
rect 4249 6817 4261 6851
rect 4295 6817 4307 6851
rect 6178 6848 6184 6860
rect 4249 6811 4307 6817
rect 5920 6820 6184 6848
rect 4154 6780 4160 6792
rect 2746 6752 4160 6780
rect 4154 6740 4160 6752
rect 4212 6740 4218 6792
rect 4525 6783 4583 6789
rect 4525 6749 4537 6783
rect 4571 6780 4583 6783
rect 5920 6780 5948 6820
rect 6178 6808 6184 6820
rect 6236 6808 6242 6860
rect 6270 6808 6276 6860
rect 6328 6848 6334 6860
rect 6328 6820 6373 6848
rect 6328 6808 6334 6820
rect 6454 6808 6460 6860
rect 6512 6848 6518 6860
rect 6549 6851 6607 6857
rect 6549 6848 6561 6851
rect 6512 6820 6561 6848
rect 6512 6808 6518 6820
rect 6549 6817 6561 6820
rect 6595 6848 6607 6851
rect 6825 6851 6883 6857
rect 6825 6848 6837 6851
rect 6595 6820 6837 6848
rect 6595 6817 6607 6820
rect 6549 6811 6607 6817
rect 6825 6817 6837 6820
rect 6871 6817 6883 6851
rect 6932 6848 6960 6888
rect 8018 6876 8024 6928
rect 8076 6876 8082 6928
rect 8941 6919 8999 6925
rect 8941 6885 8953 6919
rect 8987 6916 8999 6919
rect 9306 6916 9312 6928
rect 8987 6888 9312 6916
rect 8987 6885 8999 6888
rect 8941 6879 8999 6885
rect 9140 6857 9168 6888
rect 9306 6876 9312 6888
rect 9364 6876 9370 6928
rect 7101 6851 7159 6857
rect 7101 6848 7113 6851
rect 6932 6820 7113 6848
rect 6825 6811 6883 6817
rect 7101 6817 7113 6820
rect 7147 6817 7159 6851
rect 7101 6811 7159 6817
rect 9125 6851 9183 6857
rect 9125 6817 9137 6851
rect 9171 6817 9183 6851
rect 9125 6811 9183 6817
rect 9217 6851 9275 6857
rect 9217 6817 9229 6851
rect 9263 6817 9275 6851
rect 9398 6848 9404 6860
rect 9359 6820 9404 6848
rect 9217 6811 9275 6817
rect 4571 6752 5948 6780
rect 5997 6783 6055 6789
rect 4571 6749 4583 6752
rect 4525 6743 4583 6749
rect 5997 6749 6009 6783
rect 6043 6780 6055 6783
rect 7469 6783 7527 6789
rect 6043 6752 7052 6780
rect 6043 6749 6055 6752
rect 5997 6743 6055 6749
rect 4065 6715 4123 6721
rect 4065 6681 4077 6715
rect 4111 6681 4123 6715
rect 4065 6675 4123 6681
rect 4080 6644 4108 6675
rect 5534 6672 5540 6724
rect 5592 6712 5598 6724
rect 6733 6715 6791 6721
rect 6733 6712 6745 6715
rect 5592 6684 6745 6712
rect 5592 6672 5598 6684
rect 6733 6681 6745 6684
rect 6779 6681 6791 6715
rect 7024 6712 7052 6752
rect 7469 6749 7481 6783
rect 7515 6780 7527 6783
rect 7834 6780 7840 6792
rect 7515 6752 7840 6780
rect 7515 6749 7527 6752
rect 7469 6743 7527 6749
rect 7834 6740 7840 6752
rect 7892 6740 7898 6792
rect 7024 6684 7144 6712
rect 6733 6675 6791 6681
rect 5902 6644 5908 6656
rect 4080 6616 5908 6644
rect 5902 6604 5908 6616
rect 5960 6604 5966 6656
rect 6454 6644 6460 6656
rect 6415 6616 6460 6644
rect 6454 6604 6460 6616
rect 6512 6604 6518 6656
rect 7116 6644 7144 6684
rect 8478 6672 8484 6724
rect 8536 6712 8542 6724
rect 8754 6712 8760 6724
rect 8536 6684 8760 6712
rect 8536 6672 8542 6684
rect 8754 6672 8760 6684
rect 8812 6672 8818 6724
rect 9232 6712 9260 6811
rect 9398 6808 9404 6820
rect 9456 6808 9462 6860
rect 9597 6859 9655 6865
rect 9597 6856 9609 6859
rect 9550 6825 9609 6856
rect 9643 6825 9655 6859
rect 9550 6819 9655 6825
rect 9781 6843 9839 6849
rect 9398 6712 9404 6724
rect 9232 6684 9404 6712
rect 9398 6672 9404 6684
rect 9456 6672 9462 6724
rect 7742 6644 7748 6656
rect 7116 6616 7748 6644
rect 7742 6604 7748 6616
rect 7800 6644 7806 6656
rect 9550 6644 9578 6819
rect 9781 6809 9793 6843
rect 9827 6840 9839 6843
rect 9970 6840 9998 7184
rect 9827 6812 9998 6840
rect 9827 6809 9839 6812
rect 9781 6803 9839 6809
rect 7800 6616 9578 6644
rect 10042 6644 10070 7296
rect 13170 6644 13176 6656
rect 10042 6616 13176 6644
rect 7800 6604 7806 6616
rect 13170 6604 13176 6616
rect 13228 6604 13234 6656
rect 920 6554 9844 6576
rect 920 6502 1198 6554
rect 1250 6502 1262 6554
rect 1314 6502 1326 6554
rect 1378 6502 1390 6554
rect 1442 6502 4298 6554
rect 4350 6502 4362 6554
rect 4414 6502 4426 6554
rect 4478 6502 4490 6554
rect 4542 6502 7398 6554
rect 7450 6502 7462 6554
rect 7514 6502 7526 6554
rect 7578 6502 7590 6554
rect 7642 6502 9844 6554
rect 920 6480 9844 6502
rect 3973 6443 4031 6449
rect 3973 6409 3985 6443
rect 4019 6440 4031 6443
rect 4982 6440 4988 6452
rect 4019 6412 4988 6440
rect 4019 6409 4031 6412
rect 3973 6403 4031 6409
rect 4982 6400 4988 6412
rect 5040 6400 5046 6452
rect 5902 6400 5908 6452
rect 5960 6440 5966 6452
rect 5960 6412 12434 6440
rect 5960 6400 5966 6412
rect 3329 6375 3387 6381
rect 3329 6341 3341 6375
rect 3375 6372 3387 6375
rect 4062 6372 4068 6384
rect 3375 6344 4068 6372
rect 3375 6341 3387 6344
rect 3329 6335 3387 6341
rect 4062 6332 4068 6344
rect 4120 6372 4126 6384
rect 4120 6344 4384 6372
rect 4120 6332 4126 6344
rect 4356 6316 4384 6344
rect 5718 6332 5724 6384
rect 5776 6332 5782 6384
rect 8018 6332 8024 6384
rect 8076 6372 8082 6384
rect 9217 6375 9275 6381
rect 9217 6372 9229 6375
rect 8076 6344 9229 6372
rect 8076 6332 8082 6344
rect 9217 6341 9229 6344
rect 9263 6341 9275 6375
rect 12406 6372 12434 6412
rect 13078 6372 13084 6384
rect 12406 6344 13084 6372
rect 9217 6335 9275 6341
rect 13078 6332 13084 6344
rect 13136 6332 13142 6384
rect 4338 6304 4344 6316
rect 4251 6276 4344 6304
rect 4338 6264 4344 6276
rect 4396 6264 4402 6316
rect 4617 6307 4675 6313
rect 4617 6273 4629 6307
rect 4663 6304 4675 6307
rect 5736 6304 5764 6332
rect 6733 6307 6791 6313
rect 6733 6304 6745 6307
rect 4663 6276 6745 6304
rect 4663 6273 4675 6276
rect 4617 6267 4675 6273
rect 6733 6273 6745 6276
rect 6779 6273 6791 6307
rect 6733 6267 6791 6273
rect 8205 6307 8263 6313
rect 8205 6273 8217 6307
rect 8251 6304 8263 6307
rect 14182 6304 14188 6316
rect 8251 6276 14188 6304
rect 8251 6273 8263 6276
rect 8205 6267 8263 6273
rect 14182 6264 14188 6276
rect 14240 6264 14246 6316
rect 3513 6239 3571 6245
rect 3513 6205 3525 6239
rect 3559 6205 3571 6239
rect 3786 6236 3792 6248
rect 3747 6208 3792 6236
rect 3513 6199 3571 6205
rect 3528 6168 3556 6199
rect 3786 6196 3792 6208
rect 3844 6196 3850 6248
rect 3878 6196 3884 6248
rect 3936 6236 3942 6248
rect 4065 6239 4123 6245
rect 4065 6236 4077 6239
rect 3936 6208 4077 6236
rect 3936 6196 3942 6208
rect 4065 6205 4077 6208
rect 4111 6205 4123 6239
rect 4065 6199 4123 6205
rect 6457 6239 6515 6245
rect 6457 6205 6469 6239
rect 6503 6205 6515 6239
rect 6457 6199 6515 6205
rect 8389 6239 8447 6245
rect 8389 6205 8401 6239
rect 8435 6236 8447 6239
rect 8570 6236 8576 6248
rect 8435 6208 8576 6236
rect 8435 6205 8447 6208
rect 8389 6199 8447 6205
rect 4706 6168 4712 6180
rect 3528 6140 4712 6168
rect 4706 6128 4712 6140
rect 4764 6128 4770 6180
rect 6472 6168 6500 6199
rect 8570 6196 8576 6208
rect 8628 6236 8634 6248
rect 8665 6239 8723 6245
rect 8665 6236 8677 6239
rect 8628 6208 8677 6236
rect 8628 6196 8634 6208
rect 8665 6205 8677 6208
rect 8711 6205 8723 6239
rect 8665 6199 8723 6205
rect 8754 6196 8760 6248
rect 8812 6236 8818 6248
rect 9033 6239 9091 6245
rect 9033 6236 9045 6239
rect 8812 6208 9045 6236
rect 8812 6196 8818 6208
rect 9033 6205 9045 6208
rect 9079 6236 9091 6239
rect 9309 6239 9367 6245
rect 9309 6236 9321 6239
rect 9079 6208 9321 6236
rect 9079 6205 9091 6208
rect 9033 6199 9091 6205
rect 9309 6205 9321 6208
rect 9355 6205 9367 6239
rect 9309 6199 9367 6205
rect 6638 6168 6644 6180
rect 4249 6103 4307 6109
rect 4249 6069 4261 6103
rect 4295 6100 4307 6103
rect 5092 6100 5120 6154
rect 6472 6140 6644 6168
rect 6638 6128 6644 6140
rect 6696 6128 6702 6180
rect 7958 6140 9536 6168
rect 4295 6072 5120 6100
rect 4295 6069 4307 6072
rect 4249 6063 4307 6069
rect 5534 6060 5540 6112
rect 5592 6100 5598 6112
rect 6089 6103 6147 6109
rect 6089 6100 6101 6103
rect 5592 6072 6101 6100
rect 5592 6060 5598 6072
rect 6089 6069 6101 6072
rect 6135 6069 6147 6103
rect 6089 6063 6147 6069
rect 8478 6060 8484 6112
rect 8536 6100 8542 6112
rect 8573 6103 8631 6109
rect 8573 6100 8585 6103
rect 8536 6072 8585 6100
rect 8536 6060 8542 6072
rect 8573 6069 8585 6072
rect 8619 6069 8631 6103
rect 8573 6063 8631 6069
rect 8754 6060 8760 6112
rect 8812 6100 8818 6112
rect 9508 6109 9536 6140
rect 8849 6103 8907 6109
rect 8849 6100 8861 6103
rect 8812 6072 8861 6100
rect 8812 6060 8818 6072
rect 8849 6069 8861 6072
rect 8895 6069 8907 6103
rect 8849 6063 8907 6069
rect 9493 6103 9551 6109
rect 9493 6069 9505 6103
rect 9539 6069 9551 6103
rect 9493 6063 9551 6069
rect 9582 6060 9588 6112
rect 9640 6100 9646 6112
rect 14182 6100 14188 6112
rect 9640 6072 14188 6100
rect 9640 6060 9646 6072
rect 14182 6060 14188 6072
rect 14240 6060 14246 6112
rect 920 6010 9844 6032
rect 920 5958 2748 6010
rect 2800 5958 2812 6010
rect 2864 5958 2876 6010
rect 2928 5958 2940 6010
rect 2992 5958 5848 6010
rect 5900 5958 5912 6010
rect 5964 5958 5976 6010
rect 6028 5958 6040 6010
rect 6092 5958 8948 6010
rect 9000 5958 9012 6010
rect 9064 5958 9076 6010
rect 9128 5958 9140 6010
rect 9192 5958 9844 6010
rect 920 5936 9844 5958
rect 3786 5856 3792 5908
rect 3844 5896 3850 5908
rect 8570 5896 8576 5908
rect 3844 5868 5948 5896
rect 3844 5856 3850 5868
rect 5074 5788 5080 5840
rect 5132 5788 5138 5840
rect 4338 5760 4344 5772
rect 4299 5732 4344 5760
rect 4338 5720 4344 5732
rect 4396 5720 4402 5772
rect 5920 5760 5948 5868
rect 6656 5868 8576 5896
rect 6656 5828 6684 5868
rect 8570 5856 8576 5868
rect 8628 5856 8634 5908
rect 9306 5828 9312 5840
rect 6380 5800 6684 5828
rect 8786 5800 9312 5828
rect 6270 5760 6276 5772
rect 5920 5732 6276 5760
rect 6270 5720 6276 5732
rect 6328 5760 6334 5772
rect 6380 5760 6408 5800
rect 9306 5788 9312 5800
rect 9364 5788 9370 5840
rect 6328 5732 6408 5760
rect 6328 5720 6334 5732
rect 6454 5720 6460 5772
rect 6512 5760 6518 5772
rect 6549 5763 6607 5769
rect 6549 5760 6561 5763
rect 6512 5732 6561 5760
rect 6512 5720 6518 5732
rect 6549 5729 6561 5732
rect 6595 5729 6607 5763
rect 6549 5723 6607 5729
rect 6825 5763 6883 5769
rect 6825 5729 6837 5763
rect 6871 5760 6883 5763
rect 7101 5763 7159 5769
rect 7101 5760 7113 5763
rect 6871 5732 7113 5760
rect 6871 5729 6883 5732
rect 6825 5723 6883 5729
rect 7101 5729 7113 5732
rect 7147 5760 7159 5763
rect 7147 5732 7880 5760
rect 7147 5729 7159 5732
rect 7101 5723 7159 5729
rect 4617 5695 4675 5701
rect 4617 5661 4629 5695
rect 4663 5692 4675 5695
rect 6362 5692 6368 5704
rect 4663 5664 6368 5692
rect 4663 5661 4675 5664
rect 4617 5655 4675 5661
rect 6362 5652 6368 5664
rect 6420 5652 6426 5704
rect 6086 5624 6092 5636
rect 6047 5596 6092 5624
rect 6086 5584 6092 5596
rect 6144 5584 6150 5636
rect 6564 5624 6592 5723
rect 6638 5652 6644 5704
rect 6696 5692 6702 5704
rect 7377 5695 7435 5701
rect 7377 5692 7389 5695
rect 6696 5664 7389 5692
rect 6696 5652 6702 5664
rect 7377 5661 7389 5664
rect 7423 5661 7435 5695
rect 7742 5692 7748 5704
rect 7703 5664 7748 5692
rect 7377 5655 7435 5661
rect 7742 5652 7748 5664
rect 7800 5652 7806 5704
rect 7852 5692 7880 5732
rect 8754 5692 8760 5704
rect 7852 5664 8760 5692
rect 8754 5652 8760 5664
rect 8812 5692 8818 5704
rect 9122 5692 9128 5704
rect 8812 5664 9128 5692
rect 8812 5652 8818 5664
rect 9122 5652 9128 5664
rect 9180 5652 9186 5704
rect 6288 5596 6592 5624
rect 3878 5516 3884 5568
rect 3936 5556 3942 5568
rect 6288 5556 6316 5596
rect 6454 5556 6460 5568
rect 3936 5528 6316 5556
rect 6415 5528 6460 5556
rect 3936 5516 3942 5528
rect 6454 5516 6460 5528
rect 6512 5516 6518 5568
rect 6546 5516 6552 5568
rect 6604 5556 6610 5568
rect 6733 5559 6791 5565
rect 6733 5556 6745 5559
rect 6604 5528 6745 5556
rect 6604 5516 6610 5528
rect 6733 5525 6745 5528
rect 6779 5525 6791 5559
rect 7006 5556 7012 5568
rect 6967 5528 7012 5556
rect 6733 5519 6791 5525
rect 7006 5516 7012 5528
rect 7064 5516 7070 5568
rect 7285 5559 7343 5565
rect 7285 5525 7297 5559
rect 7331 5556 7343 5559
rect 7926 5556 7932 5568
rect 7331 5528 7932 5556
rect 7331 5525 7343 5528
rect 7285 5519 7343 5525
rect 7926 5516 7932 5528
rect 7984 5516 7990 5568
rect 8754 5516 8760 5568
rect 8812 5556 8818 5568
rect 9125 5559 9183 5565
rect 9125 5556 9137 5559
rect 8812 5528 9137 5556
rect 8812 5516 8818 5528
rect 9125 5525 9137 5528
rect 9171 5556 9183 5559
rect 9171 5528 9904 5556
rect 9171 5525 9183 5528
rect 9125 5519 9183 5525
rect 9876 5488 9904 5528
rect 14182 5488 14188 5500
rect 4048 5466 9844 5488
rect 4048 5414 4298 5466
rect 4350 5414 4362 5466
rect 4414 5414 4426 5466
rect 4478 5414 4490 5466
rect 4542 5414 7398 5466
rect 7450 5414 7462 5466
rect 7514 5414 7526 5466
rect 7578 5414 7590 5466
rect 7642 5414 9844 5466
rect 9876 5460 14188 5488
rect 14182 5448 14188 5460
rect 14240 5448 14246 5500
rect 4048 5392 9844 5414
rect 4525 5355 4583 5361
rect 4525 5321 4537 5355
rect 4571 5352 4583 5355
rect 5074 5352 5080 5364
rect 4571 5324 5080 5352
rect 4571 5321 4583 5324
rect 4525 5315 4583 5321
rect 5074 5312 5080 5324
rect 5132 5312 5138 5364
rect 6638 5312 6644 5364
rect 6696 5352 6702 5364
rect 6822 5352 6828 5364
rect 6696 5324 6828 5352
rect 6696 5312 6702 5324
rect 6822 5312 6828 5324
rect 6880 5352 6886 5364
rect 7101 5355 7159 5361
rect 7101 5352 7113 5355
rect 6880 5324 7113 5352
rect 6880 5312 6886 5324
rect 7101 5321 7113 5324
rect 7147 5321 7159 5355
rect 9306 5352 9312 5364
rect 9267 5324 9312 5352
rect 7101 5315 7159 5321
rect 9306 5312 9312 5324
rect 9364 5312 9370 5364
rect 4614 5216 4620 5228
rect 4575 5188 4620 5216
rect 4614 5176 4620 5188
rect 4672 5176 4678 5228
rect 4893 5219 4951 5225
rect 4893 5185 4905 5219
rect 4939 5216 4951 5219
rect 6086 5216 6092 5228
rect 4939 5188 6092 5216
rect 4939 5185 4951 5188
rect 4893 5179 4951 5185
rect 6086 5176 6092 5188
rect 6144 5176 6150 5228
rect 6178 5176 6184 5228
rect 6236 5216 6242 5228
rect 6730 5216 6736 5228
rect 6236 5188 6736 5216
rect 6236 5176 6242 5188
rect 6730 5176 6736 5188
rect 6788 5216 6794 5228
rect 7561 5219 7619 5225
rect 7561 5216 7573 5219
rect 6788 5188 7573 5216
rect 6788 5176 6794 5188
rect 7561 5185 7573 5188
rect 7607 5185 7619 5219
rect 7561 5179 7619 5185
rect 4341 5151 4399 5157
rect 4341 5117 4353 5151
rect 4387 5117 4399 5151
rect 4341 5111 4399 5117
rect 4356 5080 4384 5111
rect 6454 5108 6460 5160
rect 6512 5148 6518 5160
rect 6825 5151 6883 5157
rect 6825 5148 6837 5151
rect 6512 5120 6837 5148
rect 6512 5108 6518 5120
rect 6825 5117 6837 5120
rect 6871 5117 6883 5151
rect 6825 5111 6883 5117
rect 7101 5151 7159 5157
rect 7101 5117 7113 5151
rect 7147 5148 7159 5151
rect 7193 5151 7251 5157
rect 7193 5148 7205 5151
rect 7147 5120 7205 5148
rect 7147 5117 7159 5120
rect 7101 5111 7159 5117
rect 7193 5117 7205 5120
rect 7239 5117 7251 5151
rect 9122 5148 9128 5160
rect 9083 5120 9128 5148
rect 7193 5111 7251 5117
rect 9122 5108 9128 5120
rect 9180 5108 9186 5160
rect 4798 5080 4804 5092
rect 4356 5052 4804 5080
rect 4798 5040 4804 5052
rect 4856 5040 4862 5092
rect 6118 5052 7052 5080
rect 6365 5015 6423 5021
rect 6365 4981 6377 5015
rect 6411 5012 6423 5015
rect 6638 5012 6644 5024
rect 6411 4984 6644 5012
rect 6411 4981 6423 4984
rect 6365 4975 6423 4981
rect 6638 4972 6644 4984
rect 6696 4972 6702 5024
rect 7024 5021 7052 5052
rect 7926 5040 7932 5092
rect 7984 5040 7990 5092
rect 9033 5083 9091 5089
rect 9033 5049 9045 5083
rect 9079 5080 9091 5083
rect 9079 5052 9904 5080
rect 9079 5049 9091 5052
rect 9033 5043 9091 5049
rect 7009 5015 7067 5021
rect 7009 4981 7021 5015
rect 7055 4981 7067 5015
rect 7009 4975 7067 4981
rect 4048 4922 9844 4944
rect 4048 4870 5848 4922
rect 5900 4870 5912 4922
rect 5964 4870 5976 4922
rect 6028 4870 6040 4922
rect 6092 4870 8948 4922
rect 9000 4870 9012 4922
rect 9064 4870 9076 4922
rect 9128 4870 9140 4922
rect 9192 4870 9844 4922
rect 4048 4848 9844 4870
rect 6181 4811 6239 4817
rect 6181 4777 6193 4811
rect 6227 4808 6239 4811
rect 6362 4808 6368 4820
rect 6227 4780 6368 4808
rect 6227 4777 6239 4780
rect 6181 4771 6239 4777
rect 6362 4768 6368 4780
rect 6420 4768 6426 4820
rect 4614 4740 4620 4752
rect 4448 4712 4620 4740
rect 4448 4681 4476 4712
rect 4614 4700 4620 4712
rect 4672 4700 4678 4752
rect 5718 4700 5724 4752
rect 5776 4700 5782 4752
rect 6638 4700 6644 4752
rect 6696 4740 6702 4752
rect 6917 4743 6975 4749
rect 6917 4740 6929 4743
rect 6696 4712 6929 4740
rect 6696 4700 6702 4712
rect 6917 4709 6929 4712
rect 6963 4709 6975 4743
rect 6917 4703 6975 4709
rect 7006 4700 7012 4752
rect 7064 4740 7070 4752
rect 7064 4712 7406 4740
rect 7064 4700 7070 4712
rect 4433 4675 4491 4681
rect 4433 4641 4445 4675
rect 4479 4641 4491 4675
rect 4433 4635 4491 4641
rect 6365 4675 6423 4681
rect 6365 4641 6377 4675
rect 6411 4672 6423 4675
rect 6454 4672 6460 4684
rect 6411 4644 6460 4672
rect 6411 4641 6423 4644
rect 6365 4635 6423 4641
rect 4706 4604 4712 4616
rect 4667 4576 4712 4604
rect 4706 4564 4712 4576
rect 4764 4564 4770 4616
rect 5350 4564 5356 4616
rect 5408 4604 5414 4616
rect 6380 4604 6408 4635
rect 6454 4632 6460 4644
rect 6512 4632 6518 4684
rect 8754 4672 8760 4684
rect 8715 4644 8760 4672
rect 8754 4632 8760 4644
rect 8812 4632 8818 4684
rect 9217 4675 9275 4681
rect 9217 4641 9229 4675
rect 9263 4672 9275 4675
rect 9876 4672 9904 5052
rect 14182 4672 14188 4684
rect 9263 4644 14188 4672
rect 9263 4641 9275 4644
rect 9217 4635 9275 4641
rect 14182 4632 14188 4644
rect 14240 4632 14246 4684
rect 5408 4576 6408 4604
rect 6641 4607 6699 4613
rect 5408 4564 5414 4576
rect 6641 4573 6653 4607
rect 6687 4604 6699 4607
rect 6914 4604 6920 4616
rect 6687 4576 6920 4604
rect 6687 4573 6699 4576
rect 6641 4567 6699 4573
rect 6914 4564 6920 4576
rect 6972 4564 6978 4616
rect 8389 4539 8447 4545
rect 8389 4505 8401 4539
rect 8435 4536 8447 4539
rect 14182 4536 14188 4548
rect 8435 4508 14188 4536
rect 8435 4505 8447 4508
rect 8389 4499 8447 4505
rect 6362 4428 6368 4480
rect 6420 4468 6426 4480
rect 6549 4471 6607 4477
rect 6549 4468 6561 4471
rect 6420 4440 6561 4468
rect 6420 4428 6426 4440
rect 6549 4437 6561 4440
rect 6595 4437 6607 4471
rect 6549 4431 6607 4437
rect 7006 4428 7012 4480
rect 7064 4468 7070 4480
rect 8404 4468 8432 4499
rect 14182 4496 14188 4508
rect 14240 4496 14246 4548
rect 9122 4468 9128 4480
rect 7064 4440 8432 4468
rect 9083 4440 9128 4468
rect 7064 4428 7070 4440
rect 9122 4428 9128 4440
rect 9180 4428 9186 4480
rect 4048 4378 9844 4400
rect 4048 4326 4298 4378
rect 4350 4326 4362 4378
rect 4414 4326 4426 4378
rect 4478 4326 4490 4378
rect 4542 4326 7398 4378
rect 7450 4326 7462 4378
rect 7514 4326 7526 4378
rect 7578 4326 7590 4378
rect 7642 4326 9844 4378
rect 4048 4304 9844 4326
rect 4798 4264 4804 4276
rect 4632 4236 4804 4264
rect 4632 4128 4660 4236
rect 4798 4224 4804 4236
rect 4856 4264 4862 4276
rect 5258 4264 5264 4276
rect 4856 4236 5264 4264
rect 4856 4224 4862 4236
rect 5258 4224 5264 4236
rect 5316 4224 5322 4276
rect 9122 4156 9128 4208
rect 9180 4196 9186 4208
rect 9180 4168 9352 4196
rect 9180 4156 9186 4168
rect 4540 4100 4660 4128
rect 4540 4069 4568 4100
rect 4706 4088 4712 4140
rect 4764 4128 4770 4140
rect 9324 4137 9352 4168
rect 9398 4156 9404 4208
rect 9456 4196 9462 4208
rect 12526 4196 12532 4208
rect 9456 4168 12532 4196
rect 9456 4156 9462 4168
rect 12526 4156 12532 4168
rect 12584 4156 12590 4208
rect 6549 4131 6607 4137
rect 6549 4128 6561 4131
rect 4764 4100 6561 4128
rect 4764 4088 4770 4100
rect 6549 4097 6561 4100
rect 6595 4097 6607 4131
rect 6549 4091 6607 4097
rect 9309 4131 9367 4137
rect 9309 4097 9321 4131
rect 9355 4097 9367 4131
rect 9309 4091 9367 4097
rect 4525 4063 4583 4069
rect 4525 4029 4537 4063
rect 4571 4029 4583 4063
rect 4525 4023 4583 4029
rect 4614 4020 4620 4072
rect 4672 4060 4678 4072
rect 4801 4063 4859 4069
rect 4801 4060 4813 4063
rect 4672 4032 4813 4060
rect 4672 4020 4678 4032
rect 4801 4029 4813 4032
rect 4847 4029 4859 4063
rect 4801 4023 4859 4029
rect 6914 4020 6920 4072
rect 6972 4060 6978 4072
rect 9125 4063 9183 4069
rect 9125 4060 9137 4063
rect 6972 4032 9137 4060
rect 6972 4020 6978 4032
rect 9125 4029 9137 4032
rect 9171 4029 9183 4063
rect 9125 4023 9183 4029
rect 5074 3992 5080 4004
rect 5035 3964 5080 3992
rect 5074 3952 5080 3964
rect 5132 3952 5138 4004
rect 6362 3992 6368 4004
rect 6302 3964 6368 3992
rect 6362 3952 6368 3964
rect 6420 3952 6426 4004
rect 9217 3995 9275 4001
rect 9217 3992 9229 3995
rect 8588 3964 9229 3992
rect 8588 3936 8616 3964
rect 9217 3961 9229 3964
rect 9263 3961 9275 3995
rect 9217 3955 9275 3961
rect 4709 3927 4767 3933
rect 4709 3893 4721 3927
rect 4755 3924 4767 3927
rect 5718 3924 5724 3936
rect 4755 3896 5724 3924
rect 4755 3893 4767 3896
rect 4709 3887 4767 3893
rect 5718 3884 5724 3896
rect 5776 3884 5782 3936
rect 8570 3924 8576 3936
rect 8531 3896 8576 3924
rect 8570 3884 8576 3896
rect 8628 3884 8634 3936
rect 8754 3924 8760 3936
rect 8715 3896 8760 3924
rect 8754 3884 8760 3896
rect 8812 3884 8818 3936
rect 4048 3834 9844 3856
rect 4048 3782 5848 3834
rect 5900 3782 5912 3834
rect 5964 3782 5976 3834
rect 6028 3782 6040 3834
rect 6092 3782 8948 3834
rect 9000 3782 9012 3834
rect 9064 3782 9076 3834
rect 9128 3782 9140 3834
rect 9192 3782 9844 3834
rect 4048 3760 9844 3782
rect 5074 3680 5080 3732
rect 5132 3720 5138 3732
rect 6457 3723 6515 3729
rect 6457 3720 6469 3723
rect 5132 3692 6469 3720
rect 5132 3680 5138 3692
rect 6457 3689 6469 3692
rect 6503 3720 6515 3723
rect 9033 3723 9091 3729
rect 6503 3692 6960 3720
rect 6503 3689 6515 3692
rect 6457 3683 6515 3689
rect 6546 3652 6552 3664
rect 6210 3624 6552 3652
rect 6546 3612 6552 3624
rect 6604 3612 6610 3664
rect 6822 3652 6828 3664
rect 6656 3624 6828 3652
rect 4614 3544 4620 3596
rect 4672 3584 4678 3596
rect 6656 3593 6684 3624
rect 6822 3612 6828 3624
rect 6880 3612 6886 3664
rect 6932 3661 6960 3692
rect 9033 3689 9045 3723
rect 9079 3689 9091 3723
rect 9033 3683 9091 3689
rect 6917 3655 6975 3661
rect 6917 3621 6929 3655
rect 6963 3621 6975 3655
rect 9048 3652 9076 3683
rect 8142 3624 9076 3652
rect 6917 3615 6975 3621
rect 4709 3587 4767 3593
rect 4709 3584 4721 3587
rect 4672 3556 4721 3584
rect 4672 3544 4678 3556
rect 4709 3553 4721 3556
rect 4755 3553 4767 3587
rect 6641 3587 6699 3593
rect 6641 3584 6653 3587
rect 4709 3547 4767 3553
rect 6564 3556 6653 3584
rect 6564 3528 6592 3556
rect 6641 3553 6653 3556
rect 6687 3553 6699 3587
rect 6641 3547 6699 3553
rect 8478 3544 8484 3596
rect 8536 3584 8542 3596
rect 8573 3587 8631 3593
rect 8573 3584 8585 3587
rect 8536 3556 8585 3584
rect 8536 3544 8542 3556
rect 8573 3553 8585 3556
rect 8619 3584 8631 3587
rect 8849 3587 8907 3593
rect 8849 3584 8861 3587
rect 8619 3556 8861 3584
rect 8619 3553 8631 3556
rect 8573 3547 8631 3553
rect 8849 3553 8861 3556
rect 8895 3553 8907 3587
rect 8849 3547 8907 3553
rect 4985 3519 5043 3525
rect 4985 3485 4997 3519
rect 5031 3516 5043 3519
rect 5534 3516 5540 3528
rect 5031 3488 5540 3516
rect 5031 3485 5043 3488
rect 4985 3479 5043 3485
rect 5534 3476 5540 3488
rect 5592 3516 5598 3528
rect 6178 3516 6184 3528
rect 5592 3488 6184 3516
rect 5592 3476 5598 3488
rect 6178 3476 6184 3488
rect 6236 3476 6242 3528
rect 6546 3476 6552 3528
rect 6604 3476 6610 3528
rect 8389 3519 8447 3525
rect 8389 3485 8401 3519
rect 8435 3516 8447 3519
rect 14182 3516 14188 3528
rect 8435 3488 14188 3516
rect 8435 3485 8447 3488
rect 8389 3479 8447 3485
rect 14182 3476 14188 3488
rect 14240 3476 14246 3528
rect 7098 3340 7104 3392
rect 7156 3380 7162 3392
rect 8757 3383 8815 3389
rect 8757 3380 8769 3383
rect 7156 3352 8769 3380
rect 7156 3340 7162 3352
rect 8757 3349 8769 3352
rect 8803 3349 8815 3383
rect 8757 3343 8815 3349
rect 4048 3290 9844 3312
rect 4048 3238 4298 3290
rect 4350 3238 4362 3290
rect 4414 3238 4426 3290
rect 4478 3238 4490 3290
rect 4542 3238 7398 3290
rect 7450 3238 7462 3290
rect 7514 3238 7526 3290
rect 7578 3238 7590 3290
rect 7642 3238 9844 3290
rect 4048 3216 9844 3238
rect 6549 3179 6607 3185
rect 6549 3145 6561 3179
rect 6595 3176 6607 3179
rect 6730 3176 6736 3188
rect 6595 3148 6736 3176
rect 6595 3145 6607 3148
rect 6549 3139 6607 3145
rect 6730 3136 6736 3148
rect 6788 3136 6794 3188
rect 6914 3176 6920 3188
rect 6875 3148 6920 3176
rect 6914 3136 6920 3148
rect 6972 3136 6978 3188
rect 8757 3179 8815 3185
rect 8757 3145 8769 3179
rect 8803 3176 8815 3179
rect 8846 3176 8852 3188
rect 8803 3148 8852 3176
rect 8803 3145 8815 3148
rect 8757 3139 8815 3145
rect 8846 3136 8852 3148
rect 8904 3136 8910 3188
rect 8478 3108 8484 3120
rect 7116 3080 8484 3108
rect 4614 3000 4620 3052
rect 4672 3040 4678 3052
rect 4801 3043 4859 3049
rect 4801 3040 4813 3043
rect 4672 3012 4813 3040
rect 4672 3000 4678 3012
rect 4801 3009 4813 3012
rect 4847 3009 4859 3043
rect 4801 3003 4859 3009
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3040 5135 3043
rect 6638 3040 6644 3052
rect 5123 3012 6644 3040
rect 5123 3009 5135 3012
rect 5077 3003 5135 3009
rect 6638 3000 6644 3012
rect 6696 3000 6702 3052
rect 6825 2975 6883 2981
rect 6825 2941 6837 2975
rect 6871 2972 6883 2975
rect 7006 2972 7012 2984
rect 6871 2944 7012 2972
rect 6871 2941 6883 2944
rect 6825 2935 6883 2941
rect 7006 2932 7012 2944
rect 7064 2932 7070 2984
rect 7116 2981 7144 3080
rect 8478 3068 8484 3080
rect 8536 3068 8542 3120
rect 8754 3000 8760 3052
rect 8812 3040 8818 3052
rect 9217 3043 9275 3049
rect 9217 3040 9229 3043
rect 8812 3012 9229 3040
rect 8812 3000 8818 3012
rect 9217 3009 9229 3012
rect 9263 3009 9275 3043
rect 9398 3040 9404 3052
rect 9359 3012 9404 3040
rect 9217 3003 9275 3009
rect 9398 3000 9404 3012
rect 9456 3000 9462 3052
rect 7101 2975 7159 2981
rect 7101 2941 7113 2975
rect 7147 2941 7159 2975
rect 7558 2972 7564 2984
rect 7519 2944 7564 2972
rect 7101 2935 7159 2941
rect 7558 2932 7564 2944
rect 7616 2932 7622 2984
rect 12434 2932 12440 2984
rect 12492 2972 12498 2984
rect 14182 2972 14188 2984
rect 12492 2944 14188 2972
rect 12492 2932 12498 2944
rect 14182 2932 14188 2944
rect 14240 2932 14246 2984
rect 5350 2864 5356 2916
rect 5408 2904 5414 2916
rect 7377 2907 7435 2913
rect 5408 2876 5566 2904
rect 5408 2864 5414 2876
rect 7377 2873 7389 2907
rect 7423 2904 7435 2907
rect 12618 2904 12624 2916
rect 7423 2876 12624 2904
rect 7423 2873 7435 2876
rect 7377 2867 7435 2873
rect 12618 2864 12624 2876
rect 12676 2864 12682 2916
rect 7282 2836 7288 2848
rect 7243 2808 7288 2836
rect 7282 2796 7288 2808
rect 7340 2796 7346 2848
rect 8570 2796 8576 2848
rect 8628 2836 8634 2848
rect 8665 2839 8723 2845
rect 8665 2836 8677 2839
rect 8628 2808 8677 2836
rect 8628 2796 8634 2808
rect 8665 2805 8677 2808
rect 8711 2836 8723 2839
rect 9125 2839 9183 2845
rect 9125 2836 9137 2839
rect 8711 2808 9137 2836
rect 8711 2805 8723 2808
rect 8665 2799 8723 2805
rect 9125 2805 9137 2808
rect 9171 2836 9183 2839
rect 14274 2836 14280 2848
rect 9171 2808 14280 2836
rect 9171 2805 9183 2808
rect 9125 2799 9183 2805
rect 14274 2796 14280 2808
rect 14332 2796 14338 2848
rect 4048 2746 9844 2768
rect 4048 2694 5848 2746
rect 5900 2694 5912 2746
rect 5964 2694 5976 2746
rect 6028 2694 6040 2746
rect 6092 2694 8948 2746
rect 9000 2694 9012 2746
rect 9064 2694 9076 2746
rect 9128 2694 9140 2746
rect 9192 2694 9844 2746
rect 4048 2672 9844 2694
rect 7282 2592 7288 2644
rect 7340 2632 7346 2644
rect 8573 2635 8631 2641
rect 7340 2604 7604 2632
rect 7340 2592 7346 2604
rect 4706 2524 4712 2576
rect 4764 2564 4770 2576
rect 5077 2567 5135 2573
rect 5077 2564 5089 2567
rect 4764 2536 5089 2564
rect 4764 2524 4770 2536
rect 5077 2533 5089 2536
rect 5123 2533 5135 2567
rect 7098 2564 7104 2576
rect 6302 2536 7104 2564
rect 5077 2527 5135 2533
rect 7098 2524 7104 2536
rect 7156 2524 7162 2576
rect 7576 2550 7604 2604
rect 8573 2601 8585 2635
rect 8619 2632 8631 2635
rect 14182 2632 14188 2644
rect 8619 2604 14188 2632
rect 8619 2601 8631 2604
rect 8573 2595 8631 2601
rect 14182 2592 14188 2604
rect 14240 2592 14246 2644
rect 4801 2431 4859 2437
rect 4801 2397 4813 2431
rect 4847 2428 4859 2431
rect 6546 2428 6552 2440
rect 4847 2400 6552 2428
rect 4847 2397 4859 2400
rect 4801 2391 4859 2397
rect 6546 2388 6552 2400
rect 6604 2428 6610 2440
rect 6825 2431 6883 2437
rect 6825 2428 6837 2431
rect 6604 2400 6837 2428
rect 6604 2388 6610 2400
rect 6825 2397 6837 2400
rect 6871 2397 6883 2431
rect 7101 2431 7159 2437
rect 7101 2428 7113 2431
rect 6825 2391 6883 2397
rect 6932 2400 7113 2428
rect 6178 2320 6184 2372
rect 6236 2360 6242 2372
rect 6932 2360 6960 2400
rect 7101 2397 7113 2400
rect 7147 2397 7159 2431
rect 7101 2391 7159 2397
rect 7558 2388 7564 2440
rect 7616 2428 7622 2440
rect 14182 2428 14188 2440
rect 7616 2400 14188 2428
rect 7616 2388 7622 2400
rect 14182 2388 14188 2400
rect 14240 2388 14246 2440
rect 6236 2332 6960 2360
rect 6236 2320 6242 2332
rect 6549 2295 6607 2301
rect 6549 2261 6561 2295
rect 6595 2292 6607 2295
rect 12434 2292 12440 2304
rect 6595 2264 12440 2292
rect 6595 2261 6607 2264
rect 6549 2255 6607 2261
rect 12434 2252 12440 2264
rect 12492 2252 12498 2304
rect 4048 2202 9844 2224
rect 4048 2150 4298 2202
rect 4350 2150 4362 2202
rect 4414 2150 4426 2202
rect 4478 2150 4490 2202
rect 4542 2150 7398 2202
rect 7450 2150 7462 2202
rect 7514 2150 7526 2202
rect 7578 2150 7590 2202
rect 7642 2150 9844 2202
rect 4048 2128 9844 2150
rect 12526 1980 12532 2032
rect 12584 2020 12590 2032
rect 14274 2020 14280 2032
rect 12584 1992 14280 2020
rect 12584 1980 12590 1992
rect 14274 1980 14280 1992
rect 14332 1980 14338 2032
rect 8662 1300 8668 1352
rect 8720 1340 8726 1352
rect 14274 1340 14280 1352
rect 8720 1312 14280 1340
rect 8720 1300 8726 1312
rect 14274 1300 14280 1312
rect 14332 1300 14338 1352
rect 12618 1028 12624 1080
rect 12676 1068 12682 1080
rect 14274 1068 14280 1080
rect 12676 1040 14280 1068
rect 12676 1028 12682 1040
rect 14274 1028 14280 1040
rect 14332 1028 14338 1080
<< via1 >>
rect 9680 13200 9732 13252
rect 14188 13200 14240 13252
rect 9496 12656 9548 12708
rect 14188 12656 14240 12708
rect 13084 12452 13136 12504
rect 14188 12452 14240 12504
rect 2748 11398 2800 11450
rect 2812 11398 2864 11450
rect 2876 11398 2928 11450
rect 2940 11398 2992 11450
rect 5848 11398 5900 11450
rect 5912 11398 5964 11450
rect 5976 11398 6028 11450
rect 6040 11398 6092 11450
rect 8948 11398 9000 11450
rect 9012 11398 9064 11450
rect 9076 11398 9128 11450
rect 9140 11398 9192 11450
rect 8668 11228 8720 11280
rect 8944 11160 8996 11212
rect 9588 11160 9640 11212
rect 13176 11160 13228 11212
rect 14188 11160 14240 11212
rect 8024 11092 8076 11144
rect 4620 11024 4672 11076
rect 8116 11067 8168 11076
rect 8116 11033 8125 11067
rect 8125 11033 8159 11067
rect 8159 11033 8168 11067
rect 8116 11024 8168 11033
rect 14188 11024 14240 11076
rect 1198 10854 1250 10906
rect 1262 10854 1314 10906
rect 1326 10854 1378 10906
rect 1390 10854 1442 10906
rect 4298 10854 4350 10906
rect 4362 10854 4414 10906
rect 4426 10854 4478 10906
rect 4490 10854 4542 10906
rect 7398 10854 7450 10906
rect 7462 10854 7514 10906
rect 7526 10854 7578 10906
rect 7590 10854 7642 10906
rect 6276 10591 6328 10600
rect 6276 10557 6285 10591
rect 6285 10557 6319 10591
rect 6319 10557 6328 10591
rect 8392 10616 8444 10668
rect 8944 10684 8996 10736
rect 6276 10548 6328 10557
rect 8944 10591 8996 10600
rect 8944 10557 8953 10591
rect 8953 10557 8987 10591
rect 8987 10557 8996 10591
rect 8944 10548 8996 10557
rect 14188 10684 14240 10736
rect 8392 10480 8444 10532
rect 8576 10480 8628 10532
rect 14280 10480 14332 10532
rect 6460 10455 6512 10464
rect 6460 10421 6469 10455
rect 6469 10421 6503 10455
rect 6503 10421 6512 10455
rect 6460 10412 6512 10421
rect 7196 10412 7248 10464
rect 8300 10412 8352 10464
rect 2748 10310 2800 10362
rect 2812 10310 2864 10362
rect 2876 10310 2928 10362
rect 2940 10310 2992 10362
rect 5848 10310 5900 10362
rect 5912 10310 5964 10362
rect 5976 10310 6028 10362
rect 6040 10310 6092 10362
rect 8948 10310 9000 10362
rect 9012 10310 9064 10362
rect 9076 10310 9128 10362
rect 9140 10310 9192 10362
rect 6276 10072 6328 10124
rect 7472 10140 7524 10192
rect 8392 10208 8444 10260
rect 6736 10115 6788 10124
rect 6736 10081 6745 10115
rect 6745 10081 6779 10115
rect 6779 10081 6788 10115
rect 6736 10072 6788 10081
rect 7196 10072 7248 10124
rect 8576 10072 8628 10124
rect 7104 10004 7156 10056
rect 6368 9936 6420 9988
rect 6552 9911 6604 9920
rect 6552 9877 6561 9911
rect 6561 9877 6595 9911
rect 6595 9877 6604 9911
rect 6552 9868 6604 9877
rect 8116 9868 8168 9920
rect 9312 9868 9364 9920
rect 1198 9766 1250 9818
rect 1262 9766 1314 9818
rect 1326 9766 1378 9818
rect 1390 9766 1442 9818
rect 4298 9766 4350 9818
rect 4362 9766 4414 9818
rect 4426 9766 4478 9818
rect 4490 9766 4542 9818
rect 7398 9766 7450 9818
rect 7462 9766 7514 9818
rect 7526 9766 7578 9818
rect 7590 9766 7642 9818
rect 14372 9664 14424 9716
rect 8208 9596 8260 9648
rect 7196 9571 7248 9580
rect 7196 9537 7205 9571
rect 7205 9537 7239 9571
rect 7239 9537 7248 9571
rect 7196 9528 7248 9537
rect 7288 9528 7340 9580
rect 8852 9596 8904 9648
rect 14188 9596 14240 9648
rect 5356 9460 5408 9512
rect 6552 9392 6604 9444
rect 9588 9460 9640 9512
rect 5264 9324 5316 9376
rect 7840 9324 7892 9376
rect 2748 9222 2800 9274
rect 2812 9222 2864 9274
rect 2876 9222 2928 9274
rect 2940 9222 2992 9274
rect 5848 9222 5900 9274
rect 5912 9222 5964 9274
rect 5976 9222 6028 9274
rect 6040 9222 6092 9274
rect 8948 9222 9000 9274
rect 9012 9222 9064 9274
rect 9076 9222 9128 9274
rect 9140 9222 9192 9274
rect 4712 8984 4764 9036
rect 5264 9027 5316 9036
rect 5264 8993 5273 9027
rect 5273 8993 5307 9027
rect 5307 8993 5316 9027
rect 5264 8984 5316 8993
rect 6460 9052 6512 9104
rect 6276 9027 6328 9036
rect 4160 8780 4212 8832
rect 5356 8780 5408 8832
rect 5540 8823 5592 8832
rect 5540 8789 5549 8823
rect 5549 8789 5583 8823
rect 5583 8789 5592 8823
rect 5540 8780 5592 8789
rect 6276 8993 6285 9027
rect 6285 8993 6319 9027
rect 6319 8993 6328 9027
rect 6276 8984 6328 8993
rect 14188 9120 14240 9172
rect 9496 9052 9548 9104
rect 8852 8984 8904 9036
rect 9404 8984 9456 9036
rect 6552 8959 6604 8968
rect 6552 8925 6561 8959
rect 6561 8925 6595 8959
rect 6595 8925 6604 8959
rect 6552 8916 6604 8925
rect 8576 8916 8628 8968
rect 9312 8916 9364 8968
rect 6184 8780 6236 8832
rect 6644 8780 6696 8832
rect 10508 8780 10560 8832
rect 1198 8678 1250 8730
rect 1262 8678 1314 8730
rect 1326 8678 1378 8730
rect 1390 8678 1442 8730
rect 4298 8678 4350 8730
rect 4362 8678 4414 8730
rect 4426 8678 4478 8730
rect 4490 8678 4542 8730
rect 7398 8678 7450 8730
rect 7462 8678 7514 8730
rect 7526 8678 7578 8730
rect 7590 8678 7642 8730
rect 14188 8576 14240 8628
rect 8024 8508 8076 8560
rect 8852 8508 8904 8560
rect 5172 8440 5224 8492
rect 5448 8440 5500 8492
rect 8116 8483 8168 8492
rect 4160 8415 4212 8424
rect 4160 8381 4169 8415
rect 4169 8381 4203 8415
rect 4203 8381 4212 8415
rect 4160 8372 4212 8381
rect 6092 8415 6144 8424
rect 6092 8381 6101 8415
rect 6101 8381 6135 8415
rect 6135 8381 6144 8415
rect 6092 8372 6144 8381
rect 4896 8304 4948 8356
rect 6368 8347 6420 8356
rect 6368 8313 6377 8347
rect 6377 8313 6411 8347
rect 6411 8313 6420 8347
rect 6368 8304 6420 8313
rect 6644 8304 6696 8356
rect 8116 8449 8125 8483
rect 8125 8449 8159 8483
rect 8159 8449 8168 8483
rect 8116 8440 8168 8449
rect 8760 8372 8812 8424
rect 9496 8304 9548 8356
rect 5724 8236 5776 8288
rect 10508 8236 10560 8288
rect 14188 8236 14240 8288
rect 2748 8134 2800 8186
rect 2812 8134 2864 8186
rect 2876 8134 2928 8186
rect 2940 8134 2992 8186
rect 5848 8134 5900 8186
rect 5912 8134 5964 8186
rect 5976 8134 6028 8186
rect 6040 8134 6092 8186
rect 8948 8134 9000 8186
rect 9012 8134 9064 8186
rect 9076 8134 9128 8186
rect 9140 8134 9192 8186
rect 5540 8032 5592 8084
rect 6828 7964 6880 8016
rect 9588 8032 9640 8084
rect 6184 7896 6236 7948
rect 9312 7964 9364 8016
rect 4160 7828 4212 7880
rect 4988 7828 5040 7880
rect 5172 7828 5224 7880
rect 8852 7871 8904 7880
rect 8852 7837 8861 7871
rect 8861 7837 8895 7871
rect 8895 7837 8904 7871
rect 8852 7828 8904 7837
rect 9588 7760 9640 7812
rect 14188 7692 14240 7744
rect 1198 7590 1250 7642
rect 1262 7590 1314 7642
rect 1326 7590 1378 7642
rect 1390 7590 1442 7642
rect 4298 7590 4350 7642
rect 4362 7590 4414 7642
rect 4426 7590 4478 7642
rect 4490 7590 4542 7642
rect 7398 7590 7450 7642
rect 7462 7590 7514 7642
rect 7526 7590 7578 7642
rect 7590 7590 7642 7642
rect 4896 7488 4948 7540
rect 4988 7488 5040 7540
rect 7840 7488 7892 7540
rect 8484 7488 8536 7540
rect 14280 7488 14332 7540
rect 4068 7352 4120 7404
rect 5724 7352 5776 7404
rect 3884 7327 3936 7336
rect 3884 7293 3893 7327
rect 3893 7293 3927 7327
rect 3927 7293 3936 7327
rect 3884 7284 3936 7293
rect 6092 7327 6144 7336
rect 6092 7293 6101 7327
rect 6101 7293 6135 7327
rect 6135 7293 6144 7327
rect 6092 7284 6144 7293
rect 8300 7420 8352 7472
rect 8668 7463 8720 7472
rect 8668 7429 8677 7463
rect 8677 7429 8711 7463
rect 8711 7429 8720 7463
rect 8668 7420 8720 7429
rect 14188 7352 14240 7404
rect 9312 7327 9364 7336
rect 9312 7293 9321 7327
rect 9321 7293 9355 7327
rect 9355 7293 9364 7327
rect 9312 7284 9364 7293
rect 5448 7216 5500 7268
rect 8116 7259 8168 7268
rect 8116 7225 8125 7259
rect 8125 7225 8159 7259
rect 8159 7225 8168 7259
rect 8116 7216 8168 7225
rect 5724 7148 5776 7200
rect 2748 7046 2800 7098
rect 2812 7046 2864 7098
rect 2876 7046 2928 7098
rect 2940 7046 2992 7098
rect 5848 7046 5900 7098
rect 5912 7046 5964 7098
rect 5976 7046 6028 7098
rect 6040 7046 6092 7098
rect 8948 7046 9000 7098
rect 9012 7046 9064 7098
rect 9076 7046 9128 7098
rect 9140 7046 9192 7098
rect 4620 6944 4672 6996
rect 6184 6944 6236 6996
rect 6920 6944 6972 6996
rect 4160 6876 4212 6928
rect 4988 6876 5040 6928
rect 6644 6876 6696 6928
rect 4160 6740 4212 6792
rect 6184 6808 6236 6860
rect 6276 6851 6328 6860
rect 6276 6817 6285 6851
rect 6285 6817 6319 6851
rect 6319 6817 6328 6851
rect 6276 6808 6328 6817
rect 6460 6808 6512 6860
rect 8024 6876 8076 6928
rect 9312 6876 9364 6928
rect 9404 6851 9456 6860
rect 5540 6672 5592 6724
rect 7840 6740 7892 6792
rect 5908 6604 5960 6656
rect 6460 6647 6512 6656
rect 6460 6613 6469 6647
rect 6469 6613 6503 6647
rect 6503 6613 6512 6647
rect 6460 6604 6512 6613
rect 8484 6672 8536 6724
rect 8760 6672 8812 6724
rect 9404 6817 9413 6851
rect 9413 6817 9447 6851
rect 9447 6817 9456 6851
rect 9404 6808 9456 6817
rect 9404 6672 9456 6724
rect 7748 6604 7800 6656
rect 13176 6604 13228 6656
rect 1198 6502 1250 6554
rect 1262 6502 1314 6554
rect 1326 6502 1378 6554
rect 1390 6502 1442 6554
rect 4298 6502 4350 6554
rect 4362 6502 4414 6554
rect 4426 6502 4478 6554
rect 4490 6502 4542 6554
rect 7398 6502 7450 6554
rect 7462 6502 7514 6554
rect 7526 6502 7578 6554
rect 7590 6502 7642 6554
rect 4988 6400 5040 6452
rect 5908 6400 5960 6452
rect 4068 6332 4120 6384
rect 5724 6332 5776 6384
rect 8024 6332 8076 6384
rect 13084 6332 13136 6384
rect 4344 6307 4396 6316
rect 4344 6273 4353 6307
rect 4353 6273 4387 6307
rect 4387 6273 4396 6307
rect 4344 6264 4396 6273
rect 14188 6264 14240 6316
rect 3792 6239 3844 6248
rect 3792 6205 3801 6239
rect 3801 6205 3835 6239
rect 3835 6205 3844 6239
rect 3792 6196 3844 6205
rect 3884 6196 3936 6248
rect 4712 6128 4764 6180
rect 8576 6196 8628 6248
rect 8760 6196 8812 6248
rect 6644 6128 6696 6180
rect 5540 6060 5592 6112
rect 8484 6060 8536 6112
rect 8760 6060 8812 6112
rect 9588 6060 9640 6112
rect 14188 6060 14240 6112
rect 2748 5958 2800 6010
rect 2812 5958 2864 6010
rect 2876 5958 2928 6010
rect 2940 5958 2992 6010
rect 5848 5958 5900 6010
rect 5912 5958 5964 6010
rect 5976 5958 6028 6010
rect 6040 5958 6092 6010
rect 8948 5958 9000 6010
rect 9012 5958 9064 6010
rect 9076 5958 9128 6010
rect 9140 5958 9192 6010
rect 3792 5856 3844 5908
rect 5080 5788 5132 5840
rect 4344 5763 4396 5772
rect 4344 5729 4353 5763
rect 4353 5729 4387 5763
rect 4387 5729 4396 5763
rect 4344 5720 4396 5729
rect 8576 5856 8628 5908
rect 6276 5763 6328 5772
rect 6276 5729 6285 5763
rect 6285 5729 6319 5763
rect 6319 5729 6328 5763
rect 9312 5788 9364 5840
rect 6276 5720 6328 5729
rect 6460 5720 6512 5772
rect 6368 5652 6420 5704
rect 6092 5627 6144 5636
rect 6092 5593 6101 5627
rect 6101 5593 6135 5627
rect 6135 5593 6144 5627
rect 6092 5584 6144 5593
rect 6644 5652 6696 5704
rect 7748 5695 7800 5704
rect 7748 5661 7757 5695
rect 7757 5661 7791 5695
rect 7791 5661 7800 5695
rect 7748 5652 7800 5661
rect 8760 5652 8812 5704
rect 9128 5652 9180 5704
rect 3884 5516 3936 5568
rect 6460 5559 6512 5568
rect 6460 5525 6469 5559
rect 6469 5525 6503 5559
rect 6503 5525 6512 5559
rect 6460 5516 6512 5525
rect 6552 5516 6604 5568
rect 7012 5559 7064 5568
rect 7012 5525 7021 5559
rect 7021 5525 7055 5559
rect 7055 5525 7064 5559
rect 7012 5516 7064 5525
rect 7932 5516 7984 5568
rect 8760 5516 8812 5568
rect 4298 5414 4350 5466
rect 4362 5414 4414 5466
rect 4426 5414 4478 5466
rect 4490 5414 4542 5466
rect 7398 5414 7450 5466
rect 7462 5414 7514 5466
rect 7526 5414 7578 5466
rect 7590 5414 7642 5466
rect 14188 5448 14240 5500
rect 5080 5312 5132 5364
rect 6644 5312 6696 5364
rect 6828 5312 6880 5364
rect 9312 5355 9364 5364
rect 9312 5321 9321 5355
rect 9321 5321 9355 5355
rect 9355 5321 9364 5355
rect 9312 5312 9364 5321
rect 4620 5219 4672 5228
rect 4620 5185 4629 5219
rect 4629 5185 4663 5219
rect 4663 5185 4672 5219
rect 4620 5176 4672 5185
rect 6092 5176 6144 5228
rect 6184 5176 6236 5228
rect 6736 5176 6788 5228
rect 6460 5108 6512 5160
rect 9128 5151 9180 5160
rect 9128 5117 9137 5151
rect 9137 5117 9171 5151
rect 9171 5117 9180 5151
rect 9128 5108 9180 5117
rect 4804 5040 4856 5092
rect 6644 4972 6696 5024
rect 7932 5040 7984 5092
rect 5848 4870 5900 4922
rect 5912 4870 5964 4922
rect 5976 4870 6028 4922
rect 6040 4870 6092 4922
rect 8948 4870 9000 4922
rect 9012 4870 9064 4922
rect 9076 4870 9128 4922
rect 9140 4870 9192 4922
rect 6368 4768 6420 4820
rect 4620 4700 4672 4752
rect 5724 4700 5776 4752
rect 6644 4700 6696 4752
rect 7012 4700 7064 4752
rect 4712 4607 4764 4616
rect 4712 4573 4721 4607
rect 4721 4573 4755 4607
rect 4755 4573 4764 4607
rect 4712 4564 4764 4573
rect 5356 4564 5408 4616
rect 6460 4632 6512 4684
rect 8760 4675 8812 4684
rect 8760 4641 8769 4675
rect 8769 4641 8803 4675
rect 8803 4641 8812 4675
rect 8760 4632 8812 4641
rect 14188 4632 14240 4684
rect 6920 4564 6972 4616
rect 6368 4428 6420 4480
rect 7012 4428 7064 4480
rect 14188 4496 14240 4548
rect 9128 4471 9180 4480
rect 9128 4437 9137 4471
rect 9137 4437 9171 4471
rect 9171 4437 9180 4471
rect 9128 4428 9180 4437
rect 4298 4326 4350 4378
rect 4362 4326 4414 4378
rect 4426 4326 4478 4378
rect 4490 4326 4542 4378
rect 7398 4326 7450 4378
rect 7462 4326 7514 4378
rect 7526 4326 7578 4378
rect 7590 4326 7642 4378
rect 4804 4224 4856 4276
rect 5264 4224 5316 4276
rect 9128 4156 9180 4208
rect 4712 4088 4764 4140
rect 9404 4156 9456 4208
rect 12532 4156 12584 4208
rect 4620 4020 4672 4072
rect 6920 4020 6972 4072
rect 5080 3995 5132 4004
rect 5080 3961 5089 3995
rect 5089 3961 5123 3995
rect 5123 3961 5132 3995
rect 5080 3952 5132 3961
rect 6368 3952 6420 4004
rect 5724 3884 5776 3936
rect 8576 3927 8628 3936
rect 8576 3893 8585 3927
rect 8585 3893 8619 3927
rect 8619 3893 8628 3927
rect 8576 3884 8628 3893
rect 8760 3927 8812 3936
rect 8760 3893 8769 3927
rect 8769 3893 8803 3927
rect 8803 3893 8812 3927
rect 8760 3884 8812 3893
rect 5848 3782 5900 3834
rect 5912 3782 5964 3834
rect 5976 3782 6028 3834
rect 6040 3782 6092 3834
rect 8948 3782 9000 3834
rect 9012 3782 9064 3834
rect 9076 3782 9128 3834
rect 9140 3782 9192 3834
rect 5080 3680 5132 3732
rect 6552 3612 6604 3664
rect 4620 3544 4672 3596
rect 6828 3612 6880 3664
rect 8484 3544 8536 3596
rect 5540 3476 5592 3528
rect 6184 3476 6236 3528
rect 6552 3476 6604 3528
rect 14188 3476 14240 3528
rect 7104 3340 7156 3392
rect 4298 3238 4350 3290
rect 4362 3238 4414 3290
rect 4426 3238 4478 3290
rect 4490 3238 4542 3290
rect 7398 3238 7450 3290
rect 7462 3238 7514 3290
rect 7526 3238 7578 3290
rect 7590 3238 7642 3290
rect 6736 3136 6788 3188
rect 6920 3179 6972 3188
rect 6920 3145 6929 3179
rect 6929 3145 6963 3179
rect 6963 3145 6972 3179
rect 6920 3136 6972 3145
rect 8852 3136 8904 3188
rect 4620 3000 4672 3052
rect 6644 3000 6696 3052
rect 7012 2932 7064 2984
rect 8484 3068 8536 3120
rect 8760 3000 8812 3052
rect 9404 3043 9456 3052
rect 9404 3009 9413 3043
rect 9413 3009 9447 3043
rect 9447 3009 9456 3043
rect 9404 3000 9456 3009
rect 7564 2975 7616 2984
rect 7564 2941 7573 2975
rect 7573 2941 7607 2975
rect 7607 2941 7616 2975
rect 7564 2932 7616 2941
rect 12440 2932 12492 2984
rect 14188 2932 14240 2984
rect 5356 2864 5408 2916
rect 12624 2864 12676 2916
rect 7288 2839 7340 2848
rect 7288 2805 7297 2839
rect 7297 2805 7331 2839
rect 7331 2805 7340 2839
rect 7288 2796 7340 2805
rect 8576 2796 8628 2848
rect 14280 2796 14332 2848
rect 5848 2694 5900 2746
rect 5912 2694 5964 2746
rect 5976 2694 6028 2746
rect 6040 2694 6092 2746
rect 8948 2694 9000 2746
rect 9012 2694 9064 2746
rect 9076 2694 9128 2746
rect 9140 2694 9192 2746
rect 7288 2592 7340 2644
rect 4712 2524 4764 2576
rect 7104 2524 7156 2576
rect 14188 2592 14240 2644
rect 6552 2388 6604 2440
rect 6184 2320 6236 2372
rect 7564 2388 7616 2440
rect 14188 2388 14240 2440
rect 12440 2252 12492 2304
rect 4298 2150 4350 2202
rect 4362 2150 4414 2202
rect 4426 2150 4478 2202
rect 4490 2150 4542 2202
rect 7398 2150 7450 2202
rect 7462 2150 7514 2202
rect 7526 2150 7578 2202
rect 7590 2150 7642 2202
rect 12532 1980 12584 2032
rect 14280 1980 14332 2032
rect 8668 1300 8720 1352
rect 14280 1300 14332 1352
rect 12624 1028 12676 1080
rect 14280 1028 14332 1080
<< metal2 >>
rect 14186 13696 14242 13705
rect 14186 13631 14242 13640
rect 14200 13258 14228 13631
rect 9680 13252 9732 13258
rect 9680 13194 9732 13200
rect 14188 13252 14240 13258
rect 14188 13194 14240 13200
rect 9496 12708 9548 12714
rect 9496 12650 9548 12656
rect 2722 11452 3018 11472
rect 2778 11450 2802 11452
rect 2858 11450 2882 11452
rect 2938 11450 2962 11452
rect 2800 11398 2802 11450
rect 2864 11398 2876 11450
rect 2938 11398 2940 11450
rect 2778 11396 2802 11398
rect 2858 11396 2882 11398
rect 2938 11396 2962 11398
rect 2722 11376 3018 11396
rect 5822 11452 6118 11472
rect 5878 11450 5902 11452
rect 5958 11450 5982 11452
rect 6038 11450 6062 11452
rect 5900 11398 5902 11450
rect 5964 11398 5976 11450
rect 6038 11398 6040 11450
rect 5878 11396 5902 11398
rect 5958 11396 5982 11398
rect 6038 11396 6062 11398
rect 5822 11376 6118 11396
rect 8922 11452 9218 11472
rect 8978 11450 9002 11452
rect 9058 11450 9082 11452
rect 9138 11450 9162 11452
rect 9000 11398 9002 11450
rect 9064 11398 9076 11450
rect 9138 11398 9140 11450
rect 8978 11396 9002 11398
rect 9058 11396 9082 11398
rect 9138 11396 9162 11398
rect 8922 11376 9218 11396
rect 8668 11280 8720 11286
rect 8668 11222 8720 11228
rect 8024 11144 8076 11150
rect 8024 11086 8076 11092
rect 4620 11076 4672 11082
rect 4620 11018 4672 11024
rect 1172 10908 1468 10928
rect 1228 10906 1252 10908
rect 1308 10906 1332 10908
rect 1388 10906 1412 10908
rect 1250 10854 1252 10906
rect 1314 10854 1326 10906
rect 1388 10854 1390 10906
rect 1228 10852 1252 10854
rect 1308 10852 1332 10854
rect 1388 10852 1412 10854
rect 1172 10832 1468 10852
rect 4272 10908 4568 10928
rect 4328 10906 4352 10908
rect 4408 10906 4432 10908
rect 4488 10906 4512 10908
rect 4350 10854 4352 10906
rect 4414 10854 4426 10906
rect 4488 10854 4490 10906
rect 4328 10852 4352 10854
rect 4408 10852 4432 10854
rect 4488 10852 4512 10854
rect 4272 10832 4568 10852
rect 2722 10364 3018 10384
rect 2778 10362 2802 10364
rect 2858 10362 2882 10364
rect 2938 10362 2962 10364
rect 2800 10310 2802 10362
rect 2864 10310 2876 10362
rect 2938 10310 2940 10362
rect 2778 10308 2802 10310
rect 2858 10308 2882 10310
rect 2938 10308 2962 10310
rect 2722 10288 3018 10308
rect 1172 9820 1468 9840
rect 1228 9818 1252 9820
rect 1308 9818 1332 9820
rect 1388 9818 1412 9820
rect 1250 9766 1252 9818
rect 1314 9766 1326 9818
rect 1388 9766 1390 9818
rect 1228 9764 1252 9766
rect 1308 9764 1332 9766
rect 1388 9764 1412 9766
rect 1172 9744 1468 9764
rect 4272 9820 4568 9840
rect 4328 9818 4352 9820
rect 4408 9818 4432 9820
rect 4488 9818 4512 9820
rect 4350 9766 4352 9818
rect 4414 9766 4426 9818
rect 4488 9766 4490 9818
rect 4328 9764 4352 9766
rect 4408 9764 4432 9766
rect 4488 9764 4512 9766
rect 4272 9744 4568 9764
rect 2722 9276 3018 9296
rect 2778 9274 2802 9276
rect 2858 9274 2882 9276
rect 2938 9274 2962 9276
rect 2800 9222 2802 9274
rect 2864 9222 2876 9274
rect 2938 9222 2940 9274
rect 2778 9220 2802 9222
rect 2858 9220 2882 9222
rect 2938 9220 2962 9222
rect 2722 9200 3018 9220
rect 4160 8832 4212 8838
rect 4160 8774 4212 8780
rect 1172 8732 1468 8752
rect 1228 8730 1252 8732
rect 1308 8730 1332 8732
rect 1388 8730 1412 8732
rect 1250 8678 1252 8730
rect 1314 8678 1326 8730
rect 1388 8678 1390 8730
rect 1228 8676 1252 8678
rect 1308 8676 1332 8678
rect 1388 8676 1412 8678
rect 1172 8656 1468 8676
rect 4172 8430 4200 8774
rect 4272 8732 4568 8752
rect 4328 8730 4352 8732
rect 4408 8730 4432 8732
rect 4488 8730 4512 8732
rect 4350 8678 4352 8730
rect 4414 8678 4426 8730
rect 4488 8678 4490 8730
rect 4328 8676 4352 8678
rect 4408 8676 4432 8678
rect 4488 8676 4512 8678
rect 4272 8656 4568 8676
rect 4160 8424 4212 8430
rect 4160 8366 4212 8372
rect 2722 8188 3018 8208
rect 2778 8186 2802 8188
rect 2858 8186 2882 8188
rect 2938 8186 2962 8188
rect 2800 8134 2802 8186
rect 2864 8134 2876 8186
rect 2938 8134 2940 8186
rect 2778 8132 2802 8134
rect 2858 8132 2882 8134
rect 2938 8132 2962 8134
rect 2722 8112 3018 8132
rect 4172 7970 4200 8366
rect 4080 7942 4200 7970
rect 1172 7644 1468 7664
rect 1228 7642 1252 7644
rect 1308 7642 1332 7644
rect 1388 7642 1412 7644
rect 1250 7590 1252 7642
rect 1314 7590 1326 7642
rect 1388 7590 1390 7642
rect 1228 7588 1252 7590
rect 1308 7588 1332 7590
rect 1388 7588 1412 7590
rect 1172 7568 1468 7588
rect 4080 7410 4108 7942
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 4068 7404 4120 7410
rect 4068 7346 4120 7352
rect 3884 7336 3936 7342
rect 3884 7278 3936 7284
rect 2722 7100 3018 7120
rect 2778 7098 2802 7100
rect 2858 7098 2882 7100
rect 2938 7098 2962 7100
rect 2800 7046 2802 7098
rect 2864 7046 2876 7098
rect 2938 7046 2940 7098
rect 2778 7044 2802 7046
rect 2858 7044 2882 7046
rect 2938 7044 2962 7046
rect 2722 7024 3018 7044
rect 1172 6556 1468 6576
rect 1228 6554 1252 6556
rect 1308 6554 1332 6556
rect 1388 6554 1412 6556
rect 1250 6502 1252 6554
rect 1314 6502 1326 6554
rect 1388 6502 1390 6554
rect 1228 6500 1252 6502
rect 1308 6500 1332 6502
rect 1388 6500 1412 6502
rect 1172 6480 1468 6500
rect 3896 6254 3924 7278
rect 4172 6934 4200 7822
rect 4272 7644 4568 7664
rect 4328 7642 4352 7644
rect 4408 7642 4432 7644
rect 4488 7642 4512 7644
rect 4350 7590 4352 7642
rect 4414 7590 4426 7642
rect 4488 7590 4490 7642
rect 4328 7588 4352 7590
rect 4408 7588 4432 7590
rect 4488 7588 4512 7590
rect 4272 7568 4568 7588
rect 4632 7002 4660 11018
rect 7372 10908 7668 10928
rect 7428 10906 7452 10908
rect 7508 10906 7532 10908
rect 7588 10906 7612 10908
rect 7450 10854 7452 10906
rect 7514 10854 7526 10906
rect 7588 10854 7590 10906
rect 7428 10852 7452 10854
rect 7508 10852 7532 10854
rect 7588 10852 7612 10854
rect 7372 10832 7668 10852
rect 6276 10600 6328 10606
rect 6276 10542 6328 10548
rect 6734 10568 6790 10577
rect 5822 10364 6118 10384
rect 5878 10362 5902 10364
rect 5958 10362 5982 10364
rect 6038 10362 6062 10364
rect 5900 10310 5902 10362
rect 5964 10310 5976 10362
rect 6038 10310 6040 10362
rect 5878 10308 5902 10310
rect 5958 10308 5982 10310
rect 6038 10308 6062 10310
rect 5822 10288 6118 10308
rect 6288 10130 6316 10542
rect 6734 10503 6790 10512
rect 6460 10464 6512 10470
rect 6460 10406 6512 10412
rect 6276 10124 6328 10130
rect 6276 10066 6328 10072
rect 5356 9512 5408 9518
rect 5356 9454 5408 9460
rect 5264 9376 5316 9382
rect 5264 9318 5316 9324
rect 5276 9042 5304 9318
rect 4712 9036 4764 9042
rect 4712 8978 4764 8984
rect 5264 9036 5316 9042
rect 5264 8978 5316 8984
rect 4620 6996 4672 7002
rect 4620 6938 4672 6944
rect 4160 6928 4212 6934
rect 4080 6876 4160 6882
rect 4080 6870 4212 6876
rect 4080 6854 4200 6870
rect 4080 6390 4108 6854
rect 4160 6792 4212 6798
rect 4160 6734 4212 6740
rect 4068 6384 4120 6390
rect 4068 6326 4120 6332
rect 3792 6248 3844 6254
rect 3792 6190 3844 6196
rect 3884 6248 3936 6254
rect 3884 6190 3936 6196
rect 2722 6012 3018 6032
rect 2778 6010 2802 6012
rect 2858 6010 2882 6012
rect 2938 6010 2962 6012
rect 2800 5958 2802 6010
rect 2864 5958 2876 6010
rect 2938 5958 2940 6010
rect 2778 5956 2802 5958
rect 2858 5956 2882 5958
rect 2938 5956 2962 5958
rect 2722 5936 3018 5956
rect 3804 5914 3832 6190
rect 3792 5908 3844 5914
rect 3792 5850 3844 5856
rect 3896 5574 3924 6190
rect 3884 5568 3936 5574
rect 3884 5510 3936 5516
rect 4172 4049 4200 6734
rect 4272 6556 4568 6576
rect 4328 6554 4352 6556
rect 4408 6554 4432 6556
rect 4488 6554 4512 6556
rect 4350 6502 4352 6554
rect 4414 6502 4426 6554
rect 4488 6502 4490 6554
rect 4328 6500 4352 6502
rect 4408 6500 4432 6502
rect 4488 6500 4512 6502
rect 4272 6480 4568 6500
rect 4344 6316 4396 6322
rect 4344 6258 4396 6264
rect 4356 5778 4384 6258
rect 4724 6186 4752 8978
rect 5368 8838 5396 9454
rect 5822 9276 6118 9296
rect 5878 9274 5902 9276
rect 5958 9274 5982 9276
rect 6038 9274 6062 9276
rect 5900 9222 5902 9274
rect 5964 9222 5976 9274
rect 6038 9222 6040 9274
rect 5878 9220 5902 9222
rect 5958 9220 5982 9222
rect 6038 9220 6062 9222
rect 5822 9200 6118 9220
rect 6288 9194 6316 10066
rect 6368 9988 6420 9994
rect 6368 9930 6420 9936
rect 6196 9166 6316 9194
rect 6196 8838 6224 9166
rect 6380 9058 6408 9930
rect 6472 9110 6500 10406
rect 6748 10130 6776 10503
rect 7196 10464 7248 10470
rect 7196 10406 7248 10412
rect 7208 10130 7236 10406
rect 7472 10192 7524 10198
rect 7470 10160 7472 10169
rect 7524 10160 7526 10169
rect 6736 10124 6788 10130
rect 6736 10066 6788 10072
rect 7196 10124 7248 10130
rect 7470 10095 7526 10104
rect 7196 10066 7248 10072
rect 7104 10056 7156 10062
rect 7104 9998 7156 10004
rect 6552 9920 6604 9926
rect 6552 9862 6604 9868
rect 6564 9450 6592 9862
rect 7116 9466 7144 9998
rect 7208 9586 7236 10066
rect 7372 9820 7668 9840
rect 7428 9818 7452 9820
rect 7508 9818 7532 9820
rect 7588 9818 7612 9820
rect 7450 9766 7452 9818
rect 7514 9766 7526 9818
rect 7588 9766 7590 9818
rect 7428 9764 7452 9766
rect 7508 9764 7532 9766
rect 7588 9764 7612 9766
rect 7372 9744 7668 9764
rect 7196 9580 7248 9586
rect 7196 9522 7248 9528
rect 7288 9580 7340 9586
rect 7288 9522 7340 9528
rect 7300 9466 7328 9522
rect 6552 9444 6604 9450
rect 7116 9438 7328 9466
rect 6552 9386 6604 9392
rect 7840 9376 7892 9382
rect 7840 9318 7892 9324
rect 6288 9042 6408 9058
rect 6460 9104 6512 9110
rect 6460 9046 6512 9052
rect 6276 9036 6408 9042
rect 6328 9030 6408 9036
rect 6276 8978 6328 8984
rect 5356 8832 5408 8838
rect 5356 8774 5408 8780
rect 5540 8832 5592 8838
rect 5540 8774 5592 8780
rect 6184 8832 6236 8838
rect 6184 8774 6236 8780
rect 5368 8514 5396 8774
rect 5368 8498 5488 8514
rect 5172 8492 5224 8498
rect 5368 8492 5500 8498
rect 5368 8486 5448 8492
rect 5172 8434 5224 8440
rect 5448 8434 5500 8440
rect 4896 8356 4948 8362
rect 4896 8298 4948 8304
rect 4908 7546 4936 8298
rect 5184 7886 5212 8434
rect 5552 8090 5580 8774
rect 6288 8514 6316 8978
rect 6552 8968 6604 8974
rect 6552 8910 6604 8916
rect 6104 8486 6316 8514
rect 6104 8430 6132 8486
rect 6092 8424 6144 8430
rect 6092 8366 6144 8372
rect 5724 8288 5776 8294
rect 5724 8230 5776 8236
rect 5540 8084 5592 8090
rect 5540 8026 5592 8032
rect 4988 7880 5040 7886
rect 4988 7822 5040 7828
rect 5172 7880 5224 7886
rect 5172 7822 5224 7828
rect 5000 7546 5028 7822
rect 4896 7540 4948 7546
rect 4896 7482 4948 7488
rect 4988 7540 5040 7546
rect 4988 7482 5040 7488
rect 5736 7410 5764 8230
rect 5822 8188 6118 8208
rect 5878 8186 5902 8188
rect 5958 8186 5982 8188
rect 6038 8186 6062 8188
rect 5900 8134 5902 8186
rect 5964 8134 5976 8186
rect 6038 8134 6040 8186
rect 5878 8132 5902 8134
rect 5958 8132 5982 8134
rect 6038 8132 6062 8134
rect 5822 8112 6118 8132
rect 6196 7954 6224 8486
rect 6368 8356 6420 8362
rect 6368 8298 6420 8304
rect 6184 7948 6236 7954
rect 6184 7890 6236 7896
rect 6196 7426 6224 7890
rect 5724 7404 5776 7410
rect 5724 7346 5776 7352
rect 6104 7398 6224 7426
rect 6104 7342 6132 7398
rect 6092 7336 6144 7342
rect 6092 7278 6144 7284
rect 5448 7268 5500 7274
rect 5448 7210 5500 7216
rect 4988 6928 5040 6934
rect 4988 6870 5040 6876
rect 5000 6458 5028 6870
rect 5460 6746 5488 7210
rect 5724 7200 5776 7206
rect 5724 7142 5776 7148
rect 5460 6730 5580 6746
rect 5460 6724 5592 6730
rect 5460 6718 5540 6724
rect 5540 6666 5592 6672
rect 4988 6452 5040 6458
rect 4988 6394 5040 6400
rect 5736 6390 5764 7142
rect 5822 7100 6118 7120
rect 5878 7098 5902 7100
rect 5958 7098 5982 7100
rect 6038 7098 6062 7100
rect 5900 7046 5902 7098
rect 5964 7046 5976 7098
rect 6038 7046 6040 7098
rect 5878 7044 5902 7046
rect 5958 7044 5982 7046
rect 6038 7044 6062 7046
rect 5822 7024 6118 7044
rect 6196 7002 6224 7398
rect 6184 6996 6236 7002
rect 6184 6938 6236 6944
rect 6184 6860 6236 6866
rect 6184 6802 6236 6808
rect 6276 6860 6328 6866
rect 6276 6802 6328 6808
rect 5908 6656 5960 6662
rect 5908 6598 5960 6604
rect 5920 6458 5948 6598
rect 5908 6452 5960 6458
rect 5908 6394 5960 6400
rect 5724 6384 5776 6390
rect 5724 6326 5776 6332
rect 4712 6180 4764 6186
rect 4712 6122 4764 6128
rect 5540 6112 5592 6118
rect 5540 6054 5592 6060
rect 5080 5840 5132 5846
rect 5080 5782 5132 5788
rect 4344 5772 4396 5778
rect 4344 5714 4396 5720
rect 4356 5658 4384 5714
rect 4356 5630 4660 5658
rect 4272 5468 4568 5488
rect 4328 5466 4352 5468
rect 4408 5466 4432 5468
rect 4488 5466 4512 5468
rect 4350 5414 4352 5466
rect 4414 5414 4426 5466
rect 4488 5414 4490 5466
rect 4328 5412 4352 5414
rect 4408 5412 4432 5414
rect 4488 5412 4512 5414
rect 4272 5392 4568 5412
rect 4632 5234 4660 5630
rect 5092 5370 5120 5782
rect 5080 5364 5132 5370
rect 5080 5306 5132 5312
rect 4620 5228 4672 5234
rect 4620 5170 4672 5176
rect 4632 4758 4660 5170
rect 4804 5092 4856 5098
rect 4804 5034 4856 5040
rect 4620 4752 4672 4758
rect 4620 4694 4672 4700
rect 4272 4380 4568 4400
rect 4328 4378 4352 4380
rect 4408 4378 4432 4380
rect 4488 4378 4512 4380
rect 4350 4326 4352 4378
rect 4414 4326 4426 4378
rect 4488 4326 4490 4378
rect 4328 4324 4352 4326
rect 4408 4324 4432 4326
rect 4488 4324 4512 4326
rect 4272 4304 4568 4324
rect 4632 4078 4660 4694
rect 4712 4616 4764 4622
rect 4712 4558 4764 4564
rect 4724 4146 4752 4558
rect 4816 4282 4844 5034
rect 5356 4616 5408 4622
rect 5356 4558 5408 4564
rect 5368 4298 5396 4558
rect 5276 4282 5396 4298
rect 4804 4276 4856 4282
rect 4804 4218 4856 4224
rect 5264 4276 5396 4282
rect 5316 4270 5396 4276
rect 5264 4218 5316 4224
rect 4712 4140 4764 4146
rect 4712 4082 4764 4088
rect 4620 4072 4672 4078
rect 4158 4040 4214 4049
rect 4620 4014 4672 4020
rect 4158 3975 4214 3984
rect 4632 3602 4660 4014
rect 4620 3596 4672 3602
rect 4620 3538 4672 3544
rect 4272 3292 4568 3312
rect 4328 3290 4352 3292
rect 4408 3290 4432 3292
rect 4488 3290 4512 3292
rect 4350 3238 4352 3290
rect 4414 3238 4426 3290
rect 4488 3238 4490 3290
rect 4328 3236 4352 3238
rect 4408 3236 4432 3238
rect 4488 3236 4512 3238
rect 4272 3216 4568 3236
rect 4632 3058 4660 3538
rect 4620 3052 4672 3058
rect 4620 2994 4672 3000
rect 4724 2582 4752 4082
rect 5080 4004 5132 4010
rect 5080 3946 5132 3952
rect 5092 3738 5120 3946
rect 5080 3732 5132 3738
rect 5080 3674 5132 3680
rect 5368 2922 5396 4270
rect 5552 3534 5580 6054
rect 5822 6012 6118 6032
rect 5878 6010 5902 6012
rect 5958 6010 5982 6012
rect 6038 6010 6062 6012
rect 5900 5958 5902 6010
rect 5964 5958 5976 6010
rect 6038 5958 6040 6010
rect 5878 5956 5902 5958
rect 5958 5956 5982 5958
rect 6038 5956 6062 5958
rect 5822 5936 6118 5956
rect 6090 5672 6146 5681
rect 6090 5607 6092 5616
rect 6144 5607 6146 5616
rect 6092 5578 6144 5584
rect 6104 5234 6132 5578
rect 6196 5234 6224 6802
rect 6288 5778 6316 6802
rect 6276 5772 6328 5778
rect 6276 5714 6328 5720
rect 6380 5710 6408 8298
rect 6460 6860 6512 6866
rect 6460 6802 6512 6808
rect 6472 6662 6500 6802
rect 6460 6656 6512 6662
rect 6460 6598 6512 6604
rect 6472 5778 6500 6598
rect 6460 5772 6512 5778
rect 6460 5714 6512 5720
rect 6368 5704 6420 5710
rect 6564 5681 6592 8910
rect 6644 8832 6696 8838
rect 6644 8774 6696 8780
rect 6656 8362 6684 8774
rect 7372 8732 7668 8752
rect 7428 8730 7452 8732
rect 7508 8730 7532 8732
rect 7588 8730 7612 8732
rect 7450 8678 7452 8730
rect 7514 8678 7526 8730
rect 7588 8678 7590 8730
rect 7428 8676 7452 8678
rect 7508 8676 7532 8678
rect 7588 8676 7612 8678
rect 7372 8656 7668 8676
rect 6644 8356 6696 8362
rect 6644 8298 6696 8304
rect 6828 8016 6880 8022
rect 6880 7964 6960 7970
rect 6828 7958 6960 7964
rect 6840 7942 6960 7958
rect 6932 7002 6960 7942
rect 7372 7644 7668 7664
rect 7428 7642 7452 7644
rect 7508 7642 7532 7644
rect 7588 7642 7612 7644
rect 7450 7590 7452 7642
rect 7514 7590 7526 7642
rect 7588 7590 7590 7642
rect 7428 7588 7452 7590
rect 7508 7588 7532 7590
rect 7588 7588 7612 7590
rect 7372 7568 7668 7588
rect 7852 7546 7880 9318
rect 8036 8566 8064 11086
rect 8116 11076 8168 11082
rect 8116 11018 8168 11024
rect 8128 10010 8156 11018
rect 8404 10674 8616 10690
rect 8392 10668 8616 10674
rect 8444 10662 8616 10668
rect 8392 10610 8444 10616
rect 8588 10538 8616 10662
rect 8392 10532 8444 10538
rect 8392 10474 8444 10480
rect 8576 10532 8628 10538
rect 8576 10474 8628 10480
rect 8300 10464 8352 10470
rect 8300 10406 8352 10412
rect 8128 9982 8248 10010
rect 8116 9920 8168 9926
rect 8116 9862 8168 9868
rect 8024 8560 8076 8566
rect 8024 8502 8076 8508
rect 8128 8498 8156 9862
rect 8220 9654 8248 9982
rect 8208 9648 8260 9654
rect 8208 9590 8260 9596
rect 8116 8492 8168 8498
rect 8116 8434 8168 8440
rect 7840 7540 7892 7546
rect 7840 7482 7892 7488
rect 6920 6996 6972 7002
rect 6920 6938 6972 6944
rect 6644 6928 6696 6934
rect 6644 6870 6696 6876
rect 6656 6186 6684 6870
rect 7852 6798 7880 7482
rect 8312 7478 8340 10406
rect 8404 10266 8432 10474
rect 8680 10282 8708 11222
rect 8944 11212 8996 11218
rect 8944 11154 8996 11160
rect 8956 10742 8984 11154
rect 8944 10736 8996 10742
rect 8944 10678 8996 10684
rect 8944 10600 8996 10606
rect 8942 10568 8944 10577
rect 8996 10568 8998 10577
rect 8392 10260 8444 10266
rect 8392 10202 8444 10208
rect 8496 10254 8708 10282
rect 8864 10526 8942 10554
rect 8496 7546 8524 10254
rect 8574 10160 8630 10169
rect 8574 10095 8576 10104
rect 8628 10095 8630 10104
rect 8576 10066 8628 10072
rect 8588 9058 8616 10066
rect 8864 9654 8892 10526
rect 8942 10503 8998 10512
rect 8922 10364 9218 10384
rect 8978 10362 9002 10364
rect 9058 10362 9082 10364
rect 9138 10362 9162 10364
rect 9000 10310 9002 10362
rect 9064 10310 9076 10362
rect 9138 10310 9140 10362
rect 8978 10308 9002 10310
rect 9058 10308 9082 10310
rect 9138 10308 9162 10310
rect 8922 10288 9218 10308
rect 9312 9920 9364 9926
rect 9312 9862 9364 9868
rect 8852 9648 8904 9654
rect 8852 9590 8904 9596
rect 8864 9194 8892 9590
rect 8922 9276 9218 9296
rect 8978 9274 9002 9276
rect 9058 9274 9082 9276
rect 9138 9274 9162 9276
rect 9000 9222 9002 9274
rect 9064 9222 9076 9274
rect 9138 9222 9140 9274
rect 8978 9220 9002 9222
rect 9058 9220 9082 9222
rect 9138 9220 9162 9222
rect 8922 9200 9218 9220
rect 8772 9166 8892 9194
rect 8588 9030 8708 9058
rect 8576 8968 8628 8974
rect 8576 8910 8628 8916
rect 8484 7540 8536 7546
rect 8484 7482 8536 7488
rect 8300 7472 8352 7478
rect 8300 7414 8352 7420
rect 8496 7290 8524 7482
rect 8128 7274 8524 7290
rect 8116 7268 8524 7274
rect 8168 7262 8524 7268
rect 8116 7210 8168 7216
rect 8024 6928 8076 6934
rect 8024 6870 8076 6876
rect 7840 6792 7892 6798
rect 7840 6734 7892 6740
rect 7748 6656 7800 6662
rect 7748 6598 7800 6604
rect 7372 6556 7668 6576
rect 7428 6554 7452 6556
rect 7508 6554 7532 6556
rect 7588 6554 7612 6556
rect 7450 6502 7452 6554
rect 7514 6502 7526 6554
rect 7588 6502 7590 6554
rect 7428 6500 7452 6502
rect 7508 6500 7532 6502
rect 7588 6500 7612 6502
rect 7372 6480 7668 6500
rect 6644 6180 6696 6186
rect 6644 6122 6696 6128
rect 6656 5710 6684 6122
rect 7760 5710 7788 6598
rect 8036 6390 8064 6870
rect 8484 6724 8536 6730
rect 8484 6666 8536 6672
rect 8024 6384 8076 6390
rect 8024 6326 8076 6332
rect 8496 6118 8524 6666
rect 8588 6254 8616 8910
rect 8680 7562 8708 9030
rect 8772 8430 8800 9166
rect 8852 9036 8904 9042
rect 8852 8978 8904 8984
rect 8864 8566 8892 8978
rect 9324 8974 9352 9862
rect 9508 9110 9536 12650
rect 9588 11212 9640 11218
rect 9588 11154 9640 11160
rect 9600 9518 9628 11154
rect 9588 9512 9640 9518
rect 9588 9454 9640 9460
rect 9496 9104 9548 9110
rect 9496 9046 9548 9052
rect 9404 9036 9456 9042
rect 9404 8978 9456 8984
rect 9312 8968 9364 8974
rect 9312 8910 9364 8916
rect 8852 8560 8904 8566
rect 8852 8502 8904 8508
rect 8760 8424 8812 8430
rect 8760 8366 8812 8372
rect 8922 8188 9218 8208
rect 8978 8186 9002 8188
rect 9058 8186 9082 8188
rect 9138 8186 9162 8188
rect 9000 8134 9002 8186
rect 9064 8134 9076 8186
rect 9138 8134 9140 8186
rect 8978 8132 9002 8134
rect 9058 8132 9082 8134
rect 9138 8132 9162 8134
rect 8922 8112 9218 8132
rect 9324 8022 9352 8910
rect 9312 8016 9364 8022
rect 9312 7958 9364 7964
rect 8852 7880 8904 7886
rect 8852 7822 8904 7828
rect 8680 7534 8800 7562
rect 8668 7472 8720 7478
rect 8668 7414 8720 7420
rect 8576 6248 8628 6254
rect 8576 6190 8628 6196
rect 8484 6112 8536 6118
rect 8484 6054 8536 6060
rect 6644 5704 6696 5710
rect 6368 5646 6420 5652
rect 6550 5672 6606 5681
rect 6092 5228 6144 5234
rect 6092 5170 6144 5176
rect 6184 5228 6236 5234
rect 6184 5170 6236 5176
rect 5822 4924 6118 4944
rect 5878 4922 5902 4924
rect 5958 4922 5982 4924
rect 6038 4922 6062 4924
rect 5900 4870 5902 4922
rect 5964 4870 5976 4922
rect 6038 4870 6040 4922
rect 5878 4868 5902 4870
rect 5958 4868 5982 4870
rect 6038 4868 6062 4870
rect 5822 4848 6118 4868
rect 6380 4826 6408 5646
rect 6644 5646 6696 5652
rect 7748 5704 7800 5710
rect 7748 5646 7800 5652
rect 6550 5607 6606 5616
rect 6460 5568 6512 5574
rect 6460 5510 6512 5516
rect 6552 5568 6604 5574
rect 6552 5510 6604 5516
rect 6472 5166 6500 5510
rect 6460 5160 6512 5166
rect 6460 5102 6512 5108
rect 6368 4820 6420 4826
rect 6368 4762 6420 4768
rect 5724 4752 5776 4758
rect 5724 4694 5776 4700
rect 5736 3942 5764 4694
rect 6472 4690 6500 5102
rect 6460 4684 6512 4690
rect 6460 4626 6512 4632
rect 6368 4480 6420 4486
rect 6368 4422 6420 4428
rect 6380 4010 6408 4422
rect 6368 4004 6420 4010
rect 6368 3946 6420 3952
rect 5724 3936 5776 3942
rect 5724 3878 5776 3884
rect 5822 3836 6118 3856
rect 5878 3834 5902 3836
rect 5958 3834 5982 3836
rect 6038 3834 6062 3836
rect 5900 3782 5902 3834
rect 5964 3782 5976 3834
rect 6038 3782 6040 3834
rect 5878 3780 5902 3782
rect 5958 3780 5982 3782
rect 6038 3780 6062 3782
rect 5822 3760 6118 3780
rect 6564 3670 6592 5510
rect 6656 5370 6684 5646
rect 7012 5568 7064 5574
rect 7012 5510 7064 5516
rect 7932 5568 7984 5574
rect 7932 5510 7984 5516
rect 6644 5364 6696 5370
rect 6644 5306 6696 5312
rect 6828 5364 6880 5370
rect 6828 5306 6880 5312
rect 6736 5228 6788 5234
rect 6736 5170 6788 5176
rect 6644 5024 6696 5030
rect 6644 4966 6696 4972
rect 6656 4758 6684 4966
rect 6644 4752 6696 4758
rect 6644 4694 6696 4700
rect 6552 3664 6604 3670
rect 6552 3606 6604 3612
rect 5540 3528 5592 3534
rect 5540 3470 5592 3476
rect 6184 3528 6236 3534
rect 6184 3470 6236 3476
rect 6552 3528 6604 3534
rect 6552 3470 6604 3476
rect 5356 2916 5408 2922
rect 5356 2858 5408 2864
rect 5822 2748 6118 2768
rect 5878 2746 5902 2748
rect 5958 2746 5982 2748
rect 6038 2746 6062 2748
rect 5900 2694 5902 2746
rect 5964 2694 5976 2746
rect 6038 2694 6040 2746
rect 5878 2692 5902 2694
rect 5958 2692 5982 2694
rect 6038 2692 6062 2694
rect 5822 2672 6118 2692
rect 4712 2576 4764 2582
rect 4712 2518 4764 2524
rect 6196 2378 6224 3470
rect 6564 2446 6592 3470
rect 6656 3058 6684 4694
rect 6748 3194 6776 5170
rect 6840 4570 6868 5306
rect 7024 4758 7052 5510
rect 7372 5468 7668 5488
rect 7428 5466 7452 5468
rect 7508 5466 7532 5468
rect 7588 5466 7612 5468
rect 7450 5414 7452 5466
rect 7514 5414 7526 5466
rect 7588 5414 7590 5466
rect 7428 5412 7452 5414
rect 7508 5412 7532 5414
rect 7588 5412 7612 5414
rect 7372 5392 7668 5412
rect 7944 5098 7972 5510
rect 7932 5092 7984 5098
rect 7932 5034 7984 5040
rect 7012 4752 7064 4758
rect 7012 4694 7064 4700
rect 6920 4616 6972 4622
rect 6840 4564 6920 4570
rect 6840 4558 6972 4564
rect 6840 4542 6960 4558
rect 6840 3670 6868 4542
rect 7012 4480 7064 4486
rect 7012 4422 7064 4428
rect 6920 4072 6972 4078
rect 6920 4014 6972 4020
rect 6828 3664 6880 3670
rect 6828 3606 6880 3612
rect 6932 3194 6960 4014
rect 6736 3188 6788 3194
rect 6736 3130 6788 3136
rect 6920 3188 6972 3194
rect 6920 3130 6972 3136
rect 6644 3052 6696 3058
rect 6644 2994 6696 3000
rect 7024 2990 7052 4422
rect 7372 4380 7668 4400
rect 7428 4378 7452 4380
rect 7508 4378 7532 4380
rect 7588 4378 7612 4380
rect 7450 4326 7452 4378
rect 7514 4326 7526 4378
rect 7588 4326 7590 4378
rect 7428 4324 7452 4326
rect 7508 4324 7532 4326
rect 7588 4324 7612 4326
rect 7372 4304 7668 4324
rect 8496 3602 8524 6054
rect 8588 5914 8616 6190
rect 8576 5908 8628 5914
rect 8576 5850 8628 5856
rect 8576 3936 8628 3942
rect 8576 3878 8628 3884
rect 8484 3596 8536 3602
rect 8484 3538 8536 3544
rect 7104 3392 7156 3398
rect 7104 3334 7156 3340
rect 7012 2984 7064 2990
rect 7012 2926 7064 2932
rect 7116 2582 7144 3334
rect 7372 3292 7668 3312
rect 7428 3290 7452 3292
rect 7508 3290 7532 3292
rect 7588 3290 7612 3292
rect 7450 3238 7452 3290
rect 7514 3238 7526 3290
rect 7588 3238 7590 3290
rect 7428 3236 7452 3238
rect 7508 3236 7532 3238
rect 7588 3236 7612 3238
rect 7372 3216 7668 3236
rect 8496 3126 8524 3538
rect 8484 3120 8536 3126
rect 8484 3062 8536 3068
rect 7564 2984 7616 2990
rect 7564 2926 7616 2932
rect 7288 2848 7340 2854
rect 7288 2790 7340 2796
rect 7300 2650 7328 2790
rect 7288 2644 7340 2650
rect 7288 2586 7340 2592
rect 7104 2576 7156 2582
rect 7104 2518 7156 2524
rect 7576 2446 7604 2926
rect 8588 2854 8616 3878
rect 8576 2848 8628 2854
rect 8576 2790 8628 2796
rect 6552 2440 6604 2446
rect 6552 2382 6604 2388
rect 7564 2440 7616 2446
rect 7564 2382 7616 2388
rect 6184 2372 6236 2378
rect 6184 2314 6236 2320
rect 4272 2204 4568 2224
rect 4328 2202 4352 2204
rect 4408 2202 4432 2204
rect 4488 2202 4512 2204
rect 4350 2150 4352 2202
rect 4414 2150 4426 2202
rect 4488 2150 4490 2202
rect 4328 2148 4352 2150
rect 4408 2148 4432 2150
rect 4488 2148 4512 2150
rect 4272 2128 4568 2148
rect 7372 2204 7668 2224
rect 7428 2202 7452 2204
rect 7508 2202 7532 2204
rect 7588 2202 7612 2204
rect 7450 2150 7452 2202
rect 7514 2150 7526 2202
rect 7588 2150 7590 2202
rect 7428 2148 7452 2150
rect 7508 2148 7532 2150
rect 7588 2148 7612 2150
rect 7372 2128 7668 2148
rect 8680 1358 8708 7414
rect 8772 6730 8800 7534
rect 8760 6724 8812 6730
rect 8760 6666 8812 6672
rect 8760 6248 8812 6254
rect 8760 6190 8812 6196
rect 8772 6118 8800 6190
rect 8760 6112 8812 6118
rect 8760 6054 8812 6060
rect 8772 5710 8800 6054
rect 8760 5704 8812 5710
rect 8760 5646 8812 5652
rect 8760 5568 8812 5574
rect 8760 5510 8812 5516
rect 8772 4690 8800 5510
rect 8760 4684 8812 4690
rect 8760 4626 8812 4632
rect 8760 3936 8812 3942
rect 8760 3878 8812 3884
rect 8772 3058 8800 3878
rect 8864 3194 8892 7822
rect 9312 7336 9364 7342
rect 9312 7278 9364 7284
rect 8922 7100 9218 7120
rect 8978 7098 9002 7100
rect 9058 7098 9082 7100
rect 9138 7098 9162 7100
rect 9000 7046 9002 7098
rect 9064 7046 9076 7098
rect 9138 7046 9140 7098
rect 8978 7044 9002 7046
rect 9058 7044 9082 7046
rect 9138 7044 9162 7046
rect 8922 7024 9218 7044
rect 9324 6934 9352 7278
rect 9312 6928 9364 6934
rect 9312 6870 9364 6876
rect 9416 6866 9444 8978
rect 9600 8922 9628 9454
rect 9508 8894 9628 8922
rect 9508 8362 9536 8894
rect 9692 8514 9720 13194
rect 14186 13152 14242 13161
rect 14186 13087 14242 13096
rect 14200 12714 14228 13087
rect 14188 12708 14240 12714
rect 14188 12650 14240 12656
rect 14186 12608 14242 12617
rect 14186 12543 14242 12552
rect 14200 12510 14228 12543
rect 13084 12504 13136 12510
rect 13084 12446 13136 12452
rect 14188 12504 14240 12510
rect 14188 12446 14240 12452
rect 10508 8832 10560 8838
rect 10508 8774 10560 8780
rect 9600 8486 9720 8514
rect 9496 8356 9548 8362
rect 9496 8298 9548 8304
rect 9600 8090 9628 8486
rect 10520 8294 10548 8774
rect 10508 8288 10560 8294
rect 10508 8230 10560 8236
rect 9588 8084 9640 8090
rect 9588 8026 9640 8032
rect 9588 7812 9640 7818
rect 9588 7754 9640 7760
rect 9404 6860 9456 6866
rect 9404 6802 9456 6808
rect 9404 6724 9456 6730
rect 9404 6666 9456 6672
rect 8922 6012 9218 6032
rect 8978 6010 9002 6012
rect 9058 6010 9082 6012
rect 9138 6010 9162 6012
rect 9000 5958 9002 6010
rect 9064 5958 9076 6010
rect 9138 5958 9140 6010
rect 8978 5956 9002 5958
rect 9058 5956 9082 5958
rect 9138 5956 9162 5958
rect 8922 5936 9218 5956
rect 9312 5840 9364 5846
rect 9312 5782 9364 5788
rect 9128 5704 9180 5710
rect 9128 5646 9180 5652
rect 9140 5166 9168 5646
rect 9324 5370 9352 5782
rect 9312 5364 9364 5370
rect 9312 5306 9364 5312
rect 9128 5160 9180 5166
rect 9128 5102 9180 5108
rect 8922 4924 9218 4944
rect 8978 4922 9002 4924
rect 9058 4922 9082 4924
rect 9138 4922 9162 4924
rect 9000 4870 9002 4922
rect 9064 4870 9076 4922
rect 9138 4870 9140 4922
rect 8978 4868 9002 4870
rect 9058 4868 9082 4870
rect 9138 4868 9162 4870
rect 8922 4848 9218 4868
rect 9128 4480 9180 4486
rect 9128 4422 9180 4428
rect 9140 4214 9168 4422
rect 9416 4214 9444 6666
rect 9600 6118 9628 7754
rect 13096 6390 13124 12446
rect 14186 12200 14242 12209
rect 14186 12135 14242 12144
rect 14200 11218 14228 12135
rect 14278 11656 14334 11665
rect 14278 11591 14334 11600
rect 13176 11212 13228 11218
rect 13176 11154 13228 11160
rect 14188 11212 14240 11218
rect 14188 11154 14240 11160
rect 13188 6662 13216 11154
rect 14186 11112 14242 11121
rect 14186 11047 14188 11056
rect 14240 11047 14242 11056
rect 14188 11018 14240 11024
rect 14188 10736 14240 10742
rect 14188 10678 14240 10684
rect 14200 10169 14228 10678
rect 14292 10538 14320 11591
rect 14370 10704 14426 10713
rect 14370 10639 14426 10648
rect 14280 10532 14332 10538
rect 14280 10474 14332 10480
rect 14186 10160 14242 10169
rect 14186 10095 14242 10104
rect 14384 9722 14412 10639
rect 14372 9716 14424 9722
rect 14372 9658 14424 9664
rect 14188 9648 14240 9654
rect 14186 9616 14188 9625
rect 14240 9616 14242 9625
rect 14186 9551 14242 9560
rect 14186 9208 14242 9217
rect 14186 9143 14188 9152
rect 14240 9143 14242 9152
rect 14188 9114 14240 9120
rect 14186 8664 14242 8673
rect 14186 8599 14188 8608
rect 14240 8599 14242 8608
rect 14188 8570 14240 8576
rect 14188 8288 14240 8294
rect 14188 8230 14240 8236
rect 14200 8129 14228 8230
rect 14186 8120 14242 8129
rect 14186 8055 14242 8064
rect 14188 7744 14240 7750
rect 14186 7712 14188 7721
rect 14240 7712 14242 7721
rect 14186 7647 14242 7656
rect 14280 7540 14332 7546
rect 14280 7482 14332 7488
rect 14188 7404 14240 7410
rect 14188 7346 14240 7352
rect 14200 7177 14228 7346
rect 14186 7168 14242 7177
rect 14186 7103 14242 7112
rect 13176 6656 13228 6662
rect 14292 6633 14320 7482
rect 13176 6598 13228 6604
rect 14278 6624 14334 6633
rect 14278 6559 14334 6568
rect 13084 6384 13136 6390
rect 13084 6326 13136 6332
rect 14188 6316 14240 6322
rect 14188 6258 14240 6264
rect 14200 6225 14228 6258
rect 14186 6216 14242 6225
rect 14186 6151 14242 6160
rect 9588 6112 9640 6118
rect 9588 6054 9640 6060
rect 14188 6112 14240 6118
rect 14188 6054 14240 6060
rect 14200 5681 14228 6054
rect 14186 5672 14242 5681
rect 14186 5607 14242 5616
rect 14188 5500 14240 5506
rect 14188 5442 14240 5448
rect 14200 5137 14228 5442
rect 14186 5128 14242 5137
rect 14186 5063 14242 5072
rect 14186 4720 14242 4729
rect 14186 4655 14188 4664
rect 14240 4655 14242 4664
rect 14188 4626 14240 4632
rect 14188 4548 14240 4554
rect 14188 4490 14240 4496
rect 9128 4208 9180 4214
rect 9128 4150 9180 4156
rect 9404 4208 9456 4214
rect 9404 4150 9456 4156
rect 12532 4208 12584 4214
rect 14200 4185 14228 4490
rect 12532 4150 12584 4156
rect 14186 4176 14242 4185
rect 8922 3836 9218 3856
rect 8978 3834 9002 3836
rect 9058 3834 9082 3836
rect 9138 3834 9162 3836
rect 9000 3782 9002 3834
rect 9064 3782 9076 3834
rect 9138 3782 9140 3834
rect 8978 3780 9002 3782
rect 9058 3780 9082 3782
rect 9138 3780 9162 3782
rect 8922 3760 9218 3780
rect 8852 3188 8904 3194
rect 8852 3130 8904 3136
rect 9416 3058 9444 4150
rect 8760 3052 8812 3058
rect 8760 2994 8812 3000
rect 9404 3052 9456 3058
rect 9404 2994 9456 3000
rect 12440 2984 12492 2990
rect 12440 2926 12492 2932
rect 8922 2748 9218 2768
rect 8978 2746 9002 2748
rect 9058 2746 9082 2748
rect 9138 2746 9162 2748
rect 9000 2694 9002 2746
rect 9064 2694 9076 2746
rect 9138 2694 9140 2746
rect 8978 2692 9002 2694
rect 9058 2692 9082 2694
rect 9138 2692 9162 2694
rect 8922 2672 9218 2692
rect 12452 2310 12480 2926
rect 12440 2304 12492 2310
rect 12440 2246 12492 2252
rect 12544 2038 12572 4150
rect 14186 4111 14242 4120
rect 14186 3632 14242 3641
rect 14186 3567 14242 3576
rect 14200 3534 14228 3567
rect 14188 3528 14240 3534
rect 14188 3470 14240 3476
rect 14186 3224 14242 3233
rect 14186 3159 14242 3168
rect 14200 2990 14228 3159
rect 14188 2984 14240 2990
rect 14188 2926 14240 2932
rect 12624 2916 12676 2922
rect 12624 2858 12676 2864
rect 12532 2032 12584 2038
rect 12532 1974 12584 1980
rect 8668 1352 8720 1358
rect 8668 1294 8720 1300
rect 12636 1086 12664 2858
rect 14280 2848 14332 2854
rect 14280 2790 14332 2796
rect 14186 2680 14242 2689
rect 14186 2615 14188 2624
rect 14240 2615 14242 2624
rect 14188 2586 14240 2592
rect 14188 2440 14240 2446
rect 14188 2382 14240 2388
rect 12624 1080 12676 1086
rect 12624 1022 12676 1028
rect 14200 241 14228 2382
rect 14292 2145 14320 2790
rect 14278 2136 14334 2145
rect 14278 2071 14334 2080
rect 14280 2032 14332 2038
rect 14280 1974 14332 1980
rect 14292 1737 14320 1974
rect 14278 1728 14334 1737
rect 14278 1663 14334 1672
rect 14280 1352 14332 1358
rect 14280 1294 14332 1300
rect 14292 1193 14320 1294
rect 14278 1184 14334 1193
rect 14278 1119 14334 1128
rect 14280 1080 14332 1086
rect 14280 1022 14332 1028
rect 14292 649 14320 1022
rect 14278 640 14334 649
rect 14278 575 14334 584
rect 14186 232 14242 241
rect 14186 167 14242 176
<< via2 >>
rect 14186 13640 14242 13696
rect 2722 11450 2778 11452
rect 2802 11450 2858 11452
rect 2882 11450 2938 11452
rect 2962 11450 3018 11452
rect 2722 11398 2748 11450
rect 2748 11398 2778 11450
rect 2802 11398 2812 11450
rect 2812 11398 2858 11450
rect 2882 11398 2928 11450
rect 2928 11398 2938 11450
rect 2962 11398 2992 11450
rect 2992 11398 3018 11450
rect 2722 11396 2778 11398
rect 2802 11396 2858 11398
rect 2882 11396 2938 11398
rect 2962 11396 3018 11398
rect 5822 11450 5878 11452
rect 5902 11450 5958 11452
rect 5982 11450 6038 11452
rect 6062 11450 6118 11452
rect 5822 11398 5848 11450
rect 5848 11398 5878 11450
rect 5902 11398 5912 11450
rect 5912 11398 5958 11450
rect 5982 11398 6028 11450
rect 6028 11398 6038 11450
rect 6062 11398 6092 11450
rect 6092 11398 6118 11450
rect 5822 11396 5878 11398
rect 5902 11396 5958 11398
rect 5982 11396 6038 11398
rect 6062 11396 6118 11398
rect 8922 11450 8978 11452
rect 9002 11450 9058 11452
rect 9082 11450 9138 11452
rect 9162 11450 9218 11452
rect 8922 11398 8948 11450
rect 8948 11398 8978 11450
rect 9002 11398 9012 11450
rect 9012 11398 9058 11450
rect 9082 11398 9128 11450
rect 9128 11398 9138 11450
rect 9162 11398 9192 11450
rect 9192 11398 9218 11450
rect 8922 11396 8978 11398
rect 9002 11396 9058 11398
rect 9082 11396 9138 11398
rect 9162 11396 9218 11398
rect 1172 10906 1228 10908
rect 1252 10906 1308 10908
rect 1332 10906 1388 10908
rect 1412 10906 1468 10908
rect 1172 10854 1198 10906
rect 1198 10854 1228 10906
rect 1252 10854 1262 10906
rect 1262 10854 1308 10906
rect 1332 10854 1378 10906
rect 1378 10854 1388 10906
rect 1412 10854 1442 10906
rect 1442 10854 1468 10906
rect 1172 10852 1228 10854
rect 1252 10852 1308 10854
rect 1332 10852 1388 10854
rect 1412 10852 1468 10854
rect 4272 10906 4328 10908
rect 4352 10906 4408 10908
rect 4432 10906 4488 10908
rect 4512 10906 4568 10908
rect 4272 10854 4298 10906
rect 4298 10854 4328 10906
rect 4352 10854 4362 10906
rect 4362 10854 4408 10906
rect 4432 10854 4478 10906
rect 4478 10854 4488 10906
rect 4512 10854 4542 10906
rect 4542 10854 4568 10906
rect 4272 10852 4328 10854
rect 4352 10852 4408 10854
rect 4432 10852 4488 10854
rect 4512 10852 4568 10854
rect 2722 10362 2778 10364
rect 2802 10362 2858 10364
rect 2882 10362 2938 10364
rect 2962 10362 3018 10364
rect 2722 10310 2748 10362
rect 2748 10310 2778 10362
rect 2802 10310 2812 10362
rect 2812 10310 2858 10362
rect 2882 10310 2928 10362
rect 2928 10310 2938 10362
rect 2962 10310 2992 10362
rect 2992 10310 3018 10362
rect 2722 10308 2778 10310
rect 2802 10308 2858 10310
rect 2882 10308 2938 10310
rect 2962 10308 3018 10310
rect 1172 9818 1228 9820
rect 1252 9818 1308 9820
rect 1332 9818 1388 9820
rect 1412 9818 1468 9820
rect 1172 9766 1198 9818
rect 1198 9766 1228 9818
rect 1252 9766 1262 9818
rect 1262 9766 1308 9818
rect 1332 9766 1378 9818
rect 1378 9766 1388 9818
rect 1412 9766 1442 9818
rect 1442 9766 1468 9818
rect 1172 9764 1228 9766
rect 1252 9764 1308 9766
rect 1332 9764 1388 9766
rect 1412 9764 1468 9766
rect 4272 9818 4328 9820
rect 4352 9818 4408 9820
rect 4432 9818 4488 9820
rect 4512 9818 4568 9820
rect 4272 9766 4298 9818
rect 4298 9766 4328 9818
rect 4352 9766 4362 9818
rect 4362 9766 4408 9818
rect 4432 9766 4478 9818
rect 4478 9766 4488 9818
rect 4512 9766 4542 9818
rect 4542 9766 4568 9818
rect 4272 9764 4328 9766
rect 4352 9764 4408 9766
rect 4432 9764 4488 9766
rect 4512 9764 4568 9766
rect 2722 9274 2778 9276
rect 2802 9274 2858 9276
rect 2882 9274 2938 9276
rect 2962 9274 3018 9276
rect 2722 9222 2748 9274
rect 2748 9222 2778 9274
rect 2802 9222 2812 9274
rect 2812 9222 2858 9274
rect 2882 9222 2928 9274
rect 2928 9222 2938 9274
rect 2962 9222 2992 9274
rect 2992 9222 3018 9274
rect 2722 9220 2778 9222
rect 2802 9220 2858 9222
rect 2882 9220 2938 9222
rect 2962 9220 3018 9222
rect 1172 8730 1228 8732
rect 1252 8730 1308 8732
rect 1332 8730 1388 8732
rect 1412 8730 1468 8732
rect 1172 8678 1198 8730
rect 1198 8678 1228 8730
rect 1252 8678 1262 8730
rect 1262 8678 1308 8730
rect 1332 8678 1378 8730
rect 1378 8678 1388 8730
rect 1412 8678 1442 8730
rect 1442 8678 1468 8730
rect 1172 8676 1228 8678
rect 1252 8676 1308 8678
rect 1332 8676 1388 8678
rect 1412 8676 1468 8678
rect 4272 8730 4328 8732
rect 4352 8730 4408 8732
rect 4432 8730 4488 8732
rect 4512 8730 4568 8732
rect 4272 8678 4298 8730
rect 4298 8678 4328 8730
rect 4352 8678 4362 8730
rect 4362 8678 4408 8730
rect 4432 8678 4478 8730
rect 4478 8678 4488 8730
rect 4512 8678 4542 8730
rect 4542 8678 4568 8730
rect 4272 8676 4328 8678
rect 4352 8676 4408 8678
rect 4432 8676 4488 8678
rect 4512 8676 4568 8678
rect 2722 8186 2778 8188
rect 2802 8186 2858 8188
rect 2882 8186 2938 8188
rect 2962 8186 3018 8188
rect 2722 8134 2748 8186
rect 2748 8134 2778 8186
rect 2802 8134 2812 8186
rect 2812 8134 2858 8186
rect 2882 8134 2928 8186
rect 2928 8134 2938 8186
rect 2962 8134 2992 8186
rect 2992 8134 3018 8186
rect 2722 8132 2778 8134
rect 2802 8132 2858 8134
rect 2882 8132 2938 8134
rect 2962 8132 3018 8134
rect 1172 7642 1228 7644
rect 1252 7642 1308 7644
rect 1332 7642 1388 7644
rect 1412 7642 1468 7644
rect 1172 7590 1198 7642
rect 1198 7590 1228 7642
rect 1252 7590 1262 7642
rect 1262 7590 1308 7642
rect 1332 7590 1378 7642
rect 1378 7590 1388 7642
rect 1412 7590 1442 7642
rect 1442 7590 1468 7642
rect 1172 7588 1228 7590
rect 1252 7588 1308 7590
rect 1332 7588 1388 7590
rect 1412 7588 1468 7590
rect 2722 7098 2778 7100
rect 2802 7098 2858 7100
rect 2882 7098 2938 7100
rect 2962 7098 3018 7100
rect 2722 7046 2748 7098
rect 2748 7046 2778 7098
rect 2802 7046 2812 7098
rect 2812 7046 2858 7098
rect 2882 7046 2928 7098
rect 2928 7046 2938 7098
rect 2962 7046 2992 7098
rect 2992 7046 3018 7098
rect 2722 7044 2778 7046
rect 2802 7044 2858 7046
rect 2882 7044 2938 7046
rect 2962 7044 3018 7046
rect 1172 6554 1228 6556
rect 1252 6554 1308 6556
rect 1332 6554 1388 6556
rect 1412 6554 1468 6556
rect 1172 6502 1198 6554
rect 1198 6502 1228 6554
rect 1252 6502 1262 6554
rect 1262 6502 1308 6554
rect 1332 6502 1378 6554
rect 1378 6502 1388 6554
rect 1412 6502 1442 6554
rect 1442 6502 1468 6554
rect 1172 6500 1228 6502
rect 1252 6500 1308 6502
rect 1332 6500 1388 6502
rect 1412 6500 1468 6502
rect 4272 7642 4328 7644
rect 4352 7642 4408 7644
rect 4432 7642 4488 7644
rect 4512 7642 4568 7644
rect 4272 7590 4298 7642
rect 4298 7590 4328 7642
rect 4352 7590 4362 7642
rect 4362 7590 4408 7642
rect 4432 7590 4478 7642
rect 4478 7590 4488 7642
rect 4512 7590 4542 7642
rect 4542 7590 4568 7642
rect 4272 7588 4328 7590
rect 4352 7588 4408 7590
rect 4432 7588 4488 7590
rect 4512 7588 4568 7590
rect 7372 10906 7428 10908
rect 7452 10906 7508 10908
rect 7532 10906 7588 10908
rect 7612 10906 7668 10908
rect 7372 10854 7398 10906
rect 7398 10854 7428 10906
rect 7452 10854 7462 10906
rect 7462 10854 7508 10906
rect 7532 10854 7578 10906
rect 7578 10854 7588 10906
rect 7612 10854 7642 10906
rect 7642 10854 7668 10906
rect 7372 10852 7428 10854
rect 7452 10852 7508 10854
rect 7532 10852 7588 10854
rect 7612 10852 7668 10854
rect 5822 10362 5878 10364
rect 5902 10362 5958 10364
rect 5982 10362 6038 10364
rect 6062 10362 6118 10364
rect 5822 10310 5848 10362
rect 5848 10310 5878 10362
rect 5902 10310 5912 10362
rect 5912 10310 5958 10362
rect 5982 10310 6028 10362
rect 6028 10310 6038 10362
rect 6062 10310 6092 10362
rect 6092 10310 6118 10362
rect 5822 10308 5878 10310
rect 5902 10308 5958 10310
rect 5982 10308 6038 10310
rect 6062 10308 6118 10310
rect 6734 10512 6790 10568
rect 2722 6010 2778 6012
rect 2802 6010 2858 6012
rect 2882 6010 2938 6012
rect 2962 6010 3018 6012
rect 2722 5958 2748 6010
rect 2748 5958 2778 6010
rect 2802 5958 2812 6010
rect 2812 5958 2858 6010
rect 2882 5958 2928 6010
rect 2928 5958 2938 6010
rect 2962 5958 2992 6010
rect 2992 5958 3018 6010
rect 2722 5956 2778 5958
rect 2802 5956 2858 5958
rect 2882 5956 2938 5958
rect 2962 5956 3018 5958
rect 4272 6554 4328 6556
rect 4352 6554 4408 6556
rect 4432 6554 4488 6556
rect 4512 6554 4568 6556
rect 4272 6502 4298 6554
rect 4298 6502 4328 6554
rect 4352 6502 4362 6554
rect 4362 6502 4408 6554
rect 4432 6502 4478 6554
rect 4478 6502 4488 6554
rect 4512 6502 4542 6554
rect 4542 6502 4568 6554
rect 4272 6500 4328 6502
rect 4352 6500 4408 6502
rect 4432 6500 4488 6502
rect 4512 6500 4568 6502
rect 5822 9274 5878 9276
rect 5902 9274 5958 9276
rect 5982 9274 6038 9276
rect 6062 9274 6118 9276
rect 5822 9222 5848 9274
rect 5848 9222 5878 9274
rect 5902 9222 5912 9274
rect 5912 9222 5958 9274
rect 5982 9222 6028 9274
rect 6028 9222 6038 9274
rect 6062 9222 6092 9274
rect 6092 9222 6118 9274
rect 5822 9220 5878 9222
rect 5902 9220 5958 9222
rect 5982 9220 6038 9222
rect 6062 9220 6118 9222
rect 7470 10140 7472 10160
rect 7472 10140 7524 10160
rect 7524 10140 7526 10160
rect 7470 10104 7526 10140
rect 7372 9818 7428 9820
rect 7452 9818 7508 9820
rect 7532 9818 7588 9820
rect 7612 9818 7668 9820
rect 7372 9766 7398 9818
rect 7398 9766 7428 9818
rect 7452 9766 7462 9818
rect 7462 9766 7508 9818
rect 7532 9766 7578 9818
rect 7578 9766 7588 9818
rect 7612 9766 7642 9818
rect 7642 9766 7668 9818
rect 7372 9764 7428 9766
rect 7452 9764 7508 9766
rect 7532 9764 7588 9766
rect 7612 9764 7668 9766
rect 5822 8186 5878 8188
rect 5902 8186 5958 8188
rect 5982 8186 6038 8188
rect 6062 8186 6118 8188
rect 5822 8134 5848 8186
rect 5848 8134 5878 8186
rect 5902 8134 5912 8186
rect 5912 8134 5958 8186
rect 5982 8134 6028 8186
rect 6028 8134 6038 8186
rect 6062 8134 6092 8186
rect 6092 8134 6118 8186
rect 5822 8132 5878 8134
rect 5902 8132 5958 8134
rect 5982 8132 6038 8134
rect 6062 8132 6118 8134
rect 5822 7098 5878 7100
rect 5902 7098 5958 7100
rect 5982 7098 6038 7100
rect 6062 7098 6118 7100
rect 5822 7046 5848 7098
rect 5848 7046 5878 7098
rect 5902 7046 5912 7098
rect 5912 7046 5958 7098
rect 5982 7046 6028 7098
rect 6028 7046 6038 7098
rect 6062 7046 6092 7098
rect 6092 7046 6118 7098
rect 5822 7044 5878 7046
rect 5902 7044 5958 7046
rect 5982 7044 6038 7046
rect 6062 7044 6118 7046
rect 4272 5466 4328 5468
rect 4352 5466 4408 5468
rect 4432 5466 4488 5468
rect 4512 5466 4568 5468
rect 4272 5414 4298 5466
rect 4298 5414 4328 5466
rect 4352 5414 4362 5466
rect 4362 5414 4408 5466
rect 4432 5414 4478 5466
rect 4478 5414 4488 5466
rect 4512 5414 4542 5466
rect 4542 5414 4568 5466
rect 4272 5412 4328 5414
rect 4352 5412 4408 5414
rect 4432 5412 4488 5414
rect 4512 5412 4568 5414
rect 4272 4378 4328 4380
rect 4352 4378 4408 4380
rect 4432 4378 4488 4380
rect 4512 4378 4568 4380
rect 4272 4326 4298 4378
rect 4298 4326 4328 4378
rect 4352 4326 4362 4378
rect 4362 4326 4408 4378
rect 4432 4326 4478 4378
rect 4478 4326 4488 4378
rect 4512 4326 4542 4378
rect 4542 4326 4568 4378
rect 4272 4324 4328 4326
rect 4352 4324 4408 4326
rect 4432 4324 4488 4326
rect 4512 4324 4568 4326
rect 4158 3984 4214 4040
rect 4272 3290 4328 3292
rect 4352 3290 4408 3292
rect 4432 3290 4488 3292
rect 4512 3290 4568 3292
rect 4272 3238 4298 3290
rect 4298 3238 4328 3290
rect 4352 3238 4362 3290
rect 4362 3238 4408 3290
rect 4432 3238 4478 3290
rect 4478 3238 4488 3290
rect 4512 3238 4542 3290
rect 4542 3238 4568 3290
rect 4272 3236 4328 3238
rect 4352 3236 4408 3238
rect 4432 3236 4488 3238
rect 4512 3236 4568 3238
rect 5822 6010 5878 6012
rect 5902 6010 5958 6012
rect 5982 6010 6038 6012
rect 6062 6010 6118 6012
rect 5822 5958 5848 6010
rect 5848 5958 5878 6010
rect 5902 5958 5912 6010
rect 5912 5958 5958 6010
rect 5982 5958 6028 6010
rect 6028 5958 6038 6010
rect 6062 5958 6092 6010
rect 6092 5958 6118 6010
rect 5822 5956 5878 5958
rect 5902 5956 5958 5958
rect 5982 5956 6038 5958
rect 6062 5956 6118 5958
rect 6090 5636 6146 5672
rect 6090 5616 6092 5636
rect 6092 5616 6144 5636
rect 6144 5616 6146 5636
rect 7372 8730 7428 8732
rect 7452 8730 7508 8732
rect 7532 8730 7588 8732
rect 7612 8730 7668 8732
rect 7372 8678 7398 8730
rect 7398 8678 7428 8730
rect 7452 8678 7462 8730
rect 7462 8678 7508 8730
rect 7532 8678 7578 8730
rect 7578 8678 7588 8730
rect 7612 8678 7642 8730
rect 7642 8678 7668 8730
rect 7372 8676 7428 8678
rect 7452 8676 7508 8678
rect 7532 8676 7588 8678
rect 7612 8676 7668 8678
rect 7372 7642 7428 7644
rect 7452 7642 7508 7644
rect 7532 7642 7588 7644
rect 7612 7642 7668 7644
rect 7372 7590 7398 7642
rect 7398 7590 7428 7642
rect 7452 7590 7462 7642
rect 7462 7590 7508 7642
rect 7532 7590 7578 7642
rect 7578 7590 7588 7642
rect 7612 7590 7642 7642
rect 7642 7590 7668 7642
rect 7372 7588 7428 7590
rect 7452 7588 7508 7590
rect 7532 7588 7588 7590
rect 7612 7588 7668 7590
rect 8942 10548 8944 10568
rect 8944 10548 8996 10568
rect 8996 10548 8998 10568
rect 8574 10124 8630 10160
rect 8574 10104 8576 10124
rect 8576 10104 8628 10124
rect 8628 10104 8630 10124
rect 8942 10512 8998 10548
rect 8922 10362 8978 10364
rect 9002 10362 9058 10364
rect 9082 10362 9138 10364
rect 9162 10362 9218 10364
rect 8922 10310 8948 10362
rect 8948 10310 8978 10362
rect 9002 10310 9012 10362
rect 9012 10310 9058 10362
rect 9082 10310 9128 10362
rect 9128 10310 9138 10362
rect 9162 10310 9192 10362
rect 9192 10310 9218 10362
rect 8922 10308 8978 10310
rect 9002 10308 9058 10310
rect 9082 10308 9138 10310
rect 9162 10308 9218 10310
rect 8922 9274 8978 9276
rect 9002 9274 9058 9276
rect 9082 9274 9138 9276
rect 9162 9274 9218 9276
rect 8922 9222 8948 9274
rect 8948 9222 8978 9274
rect 9002 9222 9012 9274
rect 9012 9222 9058 9274
rect 9082 9222 9128 9274
rect 9128 9222 9138 9274
rect 9162 9222 9192 9274
rect 9192 9222 9218 9274
rect 8922 9220 8978 9222
rect 9002 9220 9058 9222
rect 9082 9220 9138 9222
rect 9162 9220 9218 9222
rect 7372 6554 7428 6556
rect 7452 6554 7508 6556
rect 7532 6554 7588 6556
rect 7612 6554 7668 6556
rect 7372 6502 7398 6554
rect 7398 6502 7428 6554
rect 7452 6502 7462 6554
rect 7462 6502 7508 6554
rect 7532 6502 7578 6554
rect 7578 6502 7588 6554
rect 7612 6502 7642 6554
rect 7642 6502 7668 6554
rect 7372 6500 7428 6502
rect 7452 6500 7508 6502
rect 7532 6500 7588 6502
rect 7612 6500 7668 6502
rect 8922 8186 8978 8188
rect 9002 8186 9058 8188
rect 9082 8186 9138 8188
rect 9162 8186 9218 8188
rect 8922 8134 8948 8186
rect 8948 8134 8978 8186
rect 9002 8134 9012 8186
rect 9012 8134 9058 8186
rect 9082 8134 9128 8186
rect 9128 8134 9138 8186
rect 9162 8134 9192 8186
rect 9192 8134 9218 8186
rect 8922 8132 8978 8134
rect 9002 8132 9058 8134
rect 9082 8132 9138 8134
rect 9162 8132 9218 8134
rect 5822 4922 5878 4924
rect 5902 4922 5958 4924
rect 5982 4922 6038 4924
rect 6062 4922 6118 4924
rect 5822 4870 5848 4922
rect 5848 4870 5878 4922
rect 5902 4870 5912 4922
rect 5912 4870 5958 4922
rect 5982 4870 6028 4922
rect 6028 4870 6038 4922
rect 6062 4870 6092 4922
rect 6092 4870 6118 4922
rect 5822 4868 5878 4870
rect 5902 4868 5958 4870
rect 5982 4868 6038 4870
rect 6062 4868 6118 4870
rect 6550 5616 6606 5672
rect 5822 3834 5878 3836
rect 5902 3834 5958 3836
rect 5982 3834 6038 3836
rect 6062 3834 6118 3836
rect 5822 3782 5848 3834
rect 5848 3782 5878 3834
rect 5902 3782 5912 3834
rect 5912 3782 5958 3834
rect 5982 3782 6028 3834
rect 6028 3782 6038 3834
rect 6062 3782 6092 3834
rect 6092 3782 6118 3834
rect 5822 3780 5878 3782
rect 5902 3780 5958 3782
rect 5982 3780 6038 3782
rect 6062 3780 6118 3782
rect 5822 2746 5878 2748
rect 5902 2746 5958 2748
rect 5982 2746 6038 2748
rect 6062 2746 6118 2748
rect 5822 2694 5848 2746
rect 5848 2694 5878 2746
rect 5902 2694 5912 2746
rect 5912 2694 5958 2746
rect 5982 2694 6028 2746
rect 6028 2694 6038 2746
rect 6062 2694 6092 2746
rect 6092 2694 6118 2746
rect 5822 2692 5878 2694
rect 5902 2692 5958 2694
rect 5982 2692 6038 2694
rect 6062 2692 6118 2694
rect 7372 5466 7428 5468
rect 7452 5466 7508 5468
rect 7532 5466 7588 5468
rect 7612 5466 7668 5468
rect 7372 5414 7398 5466
rect 7398 5414 7428 5466
rect 7452 5414 7462 5466
rect 7462 5414 7508 5466
rect 7532 5414 7578 5466
rect 7578 5414 7588 5466
rect 7612 5414 7642 5466
rect 7642 5414 7668 5466
rect 7372 5412 7428 5414
rect 7452 5412 7508 5414
rect 7532 5412 7588 5414
rect 7612 5412 7668 5414
rect 7372 4378 7428 4380
rect 7452 4378 7508 4380
rect 7532 4378 7588 4380
rect 7612 4378 7668 4380
rect 7372 4326 7398 4378
rect 7398 4326 7428 4378
rect 7452 4326 7462 4378
rect 7462 4326 7508 4378
rect 7532 4326 7578 4378
rect 7578 4326 7588 4378
rect 7612 4326 7642 4378
rect 7642 4326 7668 4378
rect 7372 4324 7428 4326
rect 7452 4324 7508 4326
rect 7532 4324 7588 4326
rect 7612 4324 7668 4326
rect 7372 3290 7428 3292
rect 7452 3290 7508 3292
rect 7532 3290 7588 3292
rect 7612 3290 7668 3292
rect 7372 3238 7398 3290
rect 7398 3238 7428 3290
rect 7452 3238 7462 3290
rect 7462 3238 7508 3290
rect 7532 3238 7578 3290
rect 7578 3238 7588 3290
rect 7612 3238 7642 3290
rect 7642 3238 7668 3290
rect 7372 3236 7428 3238
rect 7452 3236 7508 3238
rect 7532 3236 7588 3238
rect 7612 3236 7668 3238
rect 4272 2202 4328 2204
rect 4352 2202 4408 2204
rect 4432 2202 4488 2204
rect 4512 2202 4568 2204
rect 4272 2150 4298 2202
rect 4298 2150 4328 2202
rect 4352 2150 4362 2202
rect 4362 2150 4408 2202
rect 4432 2150 4478 2202
rect 4478 2150 4488 2202
rect 4512 2150 4542 2202
rect 4542 2150 4568 2202
rect 4272 2148 4328 2150
rect 4352 2148 4408 2150
rect 4432 2148 4488 2150
rect 4512 2148 4568 2150
rect 7372 2202 7428 2204
rect 7452 2202 7508 2204
rect 7532 2202 7588 2204
rect 7612 2202 7668 2204
rect 7372 2150 7398 2202
rect 7398 2150 7428 2202
rect 7452 2150 7462 2202
rect 7462 2150 7508 2202
rect 7532 2150 7578 2202
rect 7578 2150 7588 2202
rect 7612 2150 7642 2202
rect 7642 2150 7668 2202
rect 7372 2148 7428 2150
rect 7452 2148 7508 2150
rect 7532 2148 7588 2150
rect 7612 2148 7668 2150
rect 8922 7098 8978 7100
rect 9002 7098 9058 7100
rect 9082 7098 9138 7100
rect 9162 7098 9218 7100
rect 8922 7046 8948 7098
rect 8948 7046 8978 7098
rect 9002 7046 9012 7098
rect 9012 7046 9058 7098
rect 9082 7046 9128 7098
rect 9128 7046 9138 7098
rect 9162 7046 9192 7098
rect 9192 7046 9218 7098
rect 8922 7044 8978 7046
rect 9002 7044 9058 7046
rect 9082 7044 9138 7046
rect 9162 7044 9218 7046
rect 14186 13096 14242 13152
rect 14186 12552 14242 12608
rect 8922 6010 8978 6012
rect 9002 6010 9058 6012
rect 9082 6010 9138 6012
rect 9162 6010 9218 6012
rect 8922 5958 8948 6010
rect 8948 5958 8978 6010
rect 9002 5958 9012 6010
rect 9012 5958 9058 6010
rect 9082 5958 9128 6010
rect 9128 5958 9138 6010
rect 9162 5958 9192 6010
rect 9192 5958 9218 6010
rect 8922 5956 8978 5958
rect 9002 5956 9058 5958
rect 9082 5956 9138 5958
rect 9162 5956 9218 5958
rect 8922 4922 8978 4924
rect 9002 4922 9058 4924
rect 9082 4922 9138 4924
rect 9162 4922 9218 4924
rect 8922 4870 8948 4922
rect 8948 4870 8978 4922
rect 9002 4870 9012 4922
rect 9012 4870 9058 4922
rect 9082 4870 9128 4922
rect 9128 4870 9138 4922
rect 9162 4870 9192 4922
rect 9192 4870 9218 4922
rect 8922 4868 8978 4870
rect 9002 4868 9058 4870
rect 9082 4868 9138 4870
rect 9162 4868 9218 4870
rect 14186 12144 14242 12200
rect 14278 11600 14334 11656
rect 14186 11076 14242 11112
rect 14186 11056 14188 11076
rect 14188 11056 14240 11076
rect 14240 11056 14242 11076
rect 14370 10648 14426 10704
rect 14186 10104 14242 10160
rect 14186 9596 14188 9616
rect 14188 9596 14240 9616
rect 14240 9596 14242 9616
rect 14186 9560 14242 9596
rect 14186 9172 14242 9208
rect 14186 9152 14188 9172
rect 14188 9152 14240 9172
rect 14240 9152 14242 9172
rect 14186 8628 14242 8664
rect 14186 8608 14188 8628
rect 14188 8608 14240 8628
rect 14240 8608 14242 8628
rect 14186 8064 14242 8120
rect 14186 7692 14188 7712
rect 14188 7692 14240 7712
rect 14240 7692 14242 7712
rect 14186 7656 14242 7692
rect 14186 7112 14242 7168
rect 14278 6568 14334 6624
rect 14186 6160 14242 6216
rect 14186 5616 14242 5672
rect 14186 5072 14242 5128
rect 14186 4684 14242 4720
rect 14186 4664 14188 4684
rect 14188 4664 14240 4684
rect 14240 4664 14242 4684
rect 8922 3834 8978 3836
rect 9002 3834 9058 3836
rect 9082 3834 9138 3836
rect 9162 3834 9218 3836
rect 8922 3782 8948 3834
rect 8948 3782 8978 3834
rect 9002 3782 9012 3834
rect 9012 3782 9058 3834
rect 9082 3782 9128 3834
rect 9128 3782 9138 3834
rect 9162 3782 9192 3834
rect 9192 3782 9218 3834
rect 8922 3780 8978 3782
rect 9002 3780 9058 3782
rect 9082 3780 9138 3782
rect 9162 3780 9218 3782
rect 8922 2746 8978 2748
rect 9002 2746 9058 2748
rect 9082 2746 9138 2748
rect 9162 2746 9218 2748
rect 8922 2694 8948 2746
rect 8948 2694 8978 2746
rect 9002 2694 9012 2746
rect 9012 2694 9058 2746
rect 9082 2694 9128 2746
rect 9128 2694 9138 2746
rect 9162 2694 9192 2746
rect 9192 2694 9218 2746
rect 8922 2692 8978 2694
rect 9002 2692 9058 2694
rect 9082 2692 9138 2694
rect 9162 2692 9218 2694
rect 14186 4120 14242 4176
rect 14186 3576 14242 3632
rect 14186 3168 14242 3224
rect 14186 2644 14242 2680
rect 14186 2624 14188 2644
rect 14188 2624 14240 2644
rect 14240 2624 14242 2644
rect 14278 2080 14334 2136
rect 14278 1672 14334 1728
rect 14278 1128 14334 1184
rect 14278 584 14334 640
rect 14186 176 14242 232
<< metal3 >>
rect 14000 13696 34000 13728
rect 14000 13640 14186 13696
rect 14242 13640 34000 13696
rect 14000 13608 34000 13640
rect 14000 13152 34000 13184
rect 14000 13096 14186 13152
rect 14242 13096 34000 13152
rect 14000 13064 34000 13096
rect 14000 12608 34000 12640
rect 14000 12552 14186 12608
rect 14242 12552 34000 12608
rect 14000 12520 34000 12552
rect 14000 12200 34000 12232
rect 14000 12144 14186 12200
rect 14242 12144 34000 12200
rect 14000 12112 34000 12144
rect 14000 11656 34000 11688
rect 14000 11600 14278 11656
rect 14334 11600 34000 11656
rect 14000 11568 34000 11600
rect 2710 11456 3030 11457
rect 2710 11392 2718 11456
rect 2782 11392 2798 11456
rect 2862 11392 2878 11456
rect 2942 11392 2958 11456
rect 3022 11392 3030 11456
rect 2710 11391 3030 11392
rect 5810 11456 6130 11457
rect 5810 11392 5818 11456
rect 5882 11392 5898 11456
rect 5962 11392 5978 11456
rect 6042 11392 6058 11456
rect 6122 11392 6130 11456
rect 5810 11391 6130 11392
rect 8910 11456 9230 11457
rect 8910 11392 8918 11456
rect 8982 11392 8998 11456
rect 9062 11392 9078 11456
rect 9142 11392 9158 11456
rect 9222 11392 9230 11456
rect 8910 11391 9230 11392
rect 14000 11112 34000 11144
rect 14000 11056 14186 11112
rect 14242 11056 34000 11112
rect 14000 11024 34000 11056
rect 1160 10912 1480 10913
rect 1160 10848 1168 10912
rect 1232 10848 1248 10912
rect 1312 10848 1328 10912
rect 1392 10848 1408 10912
rect 1472 10848 1480 10912
rect 1160 10847 1480 10848
rect 4260 10912 4580 10913
rect 4260 10848 4268 10912
rect 4332 10848 4348 10912
rect 4412 10848 4428 10912
rect 4492 10848 4508 10912
rect 4572 10848 4580 10912
rect 4260 10847 4580 10848
rect 7360 10912 7680 10913
rect 7360 10848 7368 10912
rect 7432 10848 7448 10912
rect 7512 10848 7528 10912
rect 7592 10848 7608 10912
rect 7672 10848 7680 10912
rect 7360 10847 7680 10848
rect 14000 10704 34000 10736
rect 14000 10648 14370 10704
rect 14426 10648 34000 10704
rect 14000 10616 34000 10648
rect 6729 10570 6795 10573
rect 8937 10570 9003 10573
rect 6729 10568 9003 10570
rect 6729 10512 6734 10568
rect 6790 10512 8942 10568
rect 8998 10512 9003 10568
rect 6729 10510 9003 10512
rect 6729 10507 6795 10510
rect 8937 10507 9003 10510
rect 2710 10368 3030 10369
rect 2710 10304 2718 10368
rect 2782 10304 2798 10368
rect 2862 10304 2878 10368
rect 2942 10304 2958 10368
rect 3022 10304 3030 10368
rect 2710 10303 3030 10304
rect 5810 10368 6130 10369
rect 5810 10304 5818 10368
rect 5882 10304 5898 10368
rect 5962 10304 5978 10368
rect 6042 10304 6058 10368
rect 6122 10304 6130 10368
rect 5810 10303 6130 10304
rect 8910 10368 9230 10369
rect 8910 10304 8918 10368
rect 8982 10304 8998 10368
rect 9062 10304 9078 10368
rect 9142 10304 9158 10368
rect 9222 10304 9230 10368
rect 8910 10303 9230 10304
rect 7465 10162 7531 10165
rect 8569 10162 8635 10165
rect 7465 10160 8635 10162
rect 7465 10104 7470 10160
rect 7526 10104 8574 10160
rect 8630 10104 8635 10160
rect 7465 10102 8635 10104
rect 7465 10099 7531 10102
rect 8569 10099 8635 10102
rect 14000 10160 34000 10192
rect 14000 10104 14186 10160
rect 14242 10104 34000 10160
rect 14000 10072 34000 10104
rect 1160 9824 1480 9825
rect 1160 9760 1168 9824
rect 1232 9760 1248 9824
rect 1312 9760 1328 9824
rect 1392 9760 1408 9824
rect 1472 9760 1480 9824
rect 1160 9759 1480 9760
rect 4260 9824 4580 9825
rect 4260 9760 4268 9824
rect 4332 9760 4348 9824
rect 4412 9760 4428 9824
rect 4492 9760 4508 9824
rect 4572 9760 4580 9824
rect 4260 9759 4580 9760
rect 7360 9824 7680 9825
rect 7360 9760 7368 9824
rect 7432 9760 7448 9824
rect 7512 9760 7528 9824
rect 7592 9760 7608 9824
rect 7672 9760 7680 9824
rect 7360 9759 7680 9760
rect 14000 9616 34000 9648
rect 14000 9560 14186 9616
rect 14242 9560 34000 9616
rect 14000 9528 34000 9560
rect 2710 9280 3030 9281
rect 2710 9216 2718 9280
rect 2782 9216 2798 9280
rect 2862 9216 2878 9280
rect 2942 9216 2958 9280
rect 3022 9216 3030 9280
rect 2710 9215 3030 9216
rect 5810 9280 6130 9281
rect 5810 9216 5818 9280
rect 5882 9216 5898 9280
rect 5962 9216 5978 9280
rect 6042 9216 6058 9280
rect 6122 9216 6130 9280
rect 5810 9215 6130 9216
rect 8910 9280 9230 9281
rect 8910 9216 8918 9280
rect 8982 9216 8998 9280
rect 9062 9216 9078 9280
rect 9142 9216 9158 9280
rect 9222 9216 9230 9280
rect 8910 9215 9230 9216
rect 14000 9208 34000 9240
rect 14000 9152 14186 9208
rect 14242 9152 34000 9208
rect 14000 9120 34000 9152
rect 1160 8736 1480 8737
rect 1160 8672 1168 8736
rect 1232 8672 1248 8736
rect 1312 8672 1328 8736
rect 1392 8672 1408 8736
rect 1472 8672 1480 8736
rect 1160 8671 1480 8672
rect 4260 8736 4580 8737
rect 4260 8672 4268 8736
rect 4332 8672 4348 8736
rect 4412 8672 4428 8736
rect 4492 8672 4508 8736
rect 4572 8672 4580 8736
rect 4260 8671 4580 8672
rect 7360 8736 7680 8737
rect 7360 8672 7368 8736
rect 7432 8672 7448 8736
rect 7512 8672 7528 8736
rect 7592 8672 7608 8736
rect 7672 8672 7680 8736
rect 7360 8671 7680 8672
rect 14000 8664 34000 8696
rect 14000 8608 14186 8664
rect 14242 8608 34000 8664
rect 14000 8576 34000 8608
rect 2710 8192 3030 8193
rect 2710 8128 2718 8192
rect 2782 8128 2798 8192
rect 2862 8128 2878 8192
rect 2942 8128 2958 8192
rect 3022 8128 3030 8192
rect 2710 8127 3030 8128
rect 5810 8192 6130 8193
rect 5810 8128 5818 8192
rect 5882 8128 5898 8192
rect 5962 8128 5978 8192
rect 6042 8128 6058 8192
rect 6122 8128 6130 8192
rect 5810 8127 6130 8128
rect 8910 8192 9230 8193
rect 8910 8128 8918 8192
rect 8982 8128 8998 8192
rect 9062 8128 9078 8192
rect 9142 8128 9158 8192
rect 9222 8128 9230 8192
rect 8910 8127 9230 8128
rect 14000 8120 34000 8152
rect 14000 8064 14186 8120
rect 14242 8064 34000 8120
rect 14000 8032 34000 8064
rect 14000 7712 34000 7744
rect 14000 7656 14186 7712
rect 14242 7656 34000 7712
rect 1160 7648 1480 7649
rect 1160 7584 1168 7648
rect 1232 7584 1248 7648
rect 1312 7584 1328 7648
rect 1392 7584 1408 7648
rect 1472 7584 1480 7648
rect 1160 7583 1480 7584
rect 4260 7648 4580 7649
rect 4260 7584 4268 7648
rect 4332 7584 4348 7648
rect 4412 7584 4428 7648
rect 4492 7584 4508 7648
rect 4572 7584 4580 7648
rect 4260 7583 4580 7584
rect 7360 7648 7680 7649
rect 7360 7584 7368 7648
rect 7432 7584 7448 7648
rect 7512 7584 7528 7648
rect 7592 7584 7608 7648
rect 7672 7584 7680 7648
rect 14000 7624 34000 7656
rect 7360 7583 7680 7584
rect 14000 7168 34000 7200
rect 14000 7112 14186 7168
rect 14242 7112 34000 7168
rect 2710 7104 3030 7105
rect 2710 7040 2718 7104
rect 2782 7040 2798 7104
rect 2862 7040 2878 7104
rect 2942 7040 2958 7104
rect 3022 7040 3030 7104
rect 2710 7039 3030 7040
rect 5810 7104 6130 7105
rect 5810 7040 5818 7104
rect 5882 7040 5898 7104
rect 5962 7040 5978 7104
rect 6042 7040 6058 7104
rect 6122 7040 6130 7104
rect 5810 7039 6130 7040
rect 8910 7104 9230 7105
rect 8910 7040 8918 7104
rect 8982 7040 8998 7104
rect 9062 7040 9078 7104
rect 9142 7040 9158 7104
rect 9222 7040 9230 7104
rect 14000 7080 34000 7112
rect 8910 7039 9230 7040
rect 14000 6624 34000 6656
rect 14000 6568 14278 6624
rect 14334 6568 34000 6624
rect 1160 6560 1480 6561
rect 1160 6496 1168 6560
rect 1232 6496 1248 6560
rect 1312 6496 1328 6560
rect 1392 6496 1408 6560
rect 1472 6496 1480 6560
rect 1160 6495 1480 6496
rect 4260 6560 4580 6561
rect 4260 6496 4268 6560
rect 4332 6496 4348 6560
rect 4412 6496 4428 6560
rect 4492 6496 4508 6560
rect 4572 6496 4580 6560
rect 4260 6495 4580 6496
rect 7360 6560 7680 6561
rect 7360 6496 7368 6560
rect 7432 6496 7448 6560
rect 7512 6496 7528 6560
rect 7592 6496 7608 6560
rect 7672 6496 7680 6560
rect 14000 6536 34000 6568
rect 7360 6495 7680 6496
rect 14000 6216 34000 6248
rect 14000 6160 14186 6216
rect 14242 6160 34000 6216
rect 14000 6128 34000 6160
rect 2710 6016 3030 6017
rect 2710 5952 2718 6016
rect 2782 5952 2798 6016
rect 2862 5952 2878 6016
rect 2942 5952 2958 6016
rect 3022 5952 3030 6016
rect 2710 5951 3030 5952
rect 5810 6016 6130 6017
rect 5810 5952 5818 6016
rect 5882 5952 5898 6016
rect 5962 5952 5978 6016
rect 6042 5952 6058 6016
rect 6122 5952 6130 6016
rect 5810 5951 6130 5952
rect 8910 6016 9230 6017
rect 8910 5952 8918 6016
rect 8982 5952 8998 6016
rect 9062 5952 9078 6016
rect 9142 5952 9158 6016
rect 9222 5952 9230 6016
rect 8910 5951 9230 5952
rect 6085 5674 6151 5677
rect 6545 5674 6611 5677
rect 6085 5672 6611 5674
rect 6085 5616 6090 5672
rect 6146 5616 6550 5672
rect 6606 5616 6611 5672
rect 6085 5614 6611 5616
rect 6085 5611 6151 5614
rect 6545 5611 6611 5614
rect 14000 5672 34000 5704
rect 14000 5616 14186 5672
rect 14242 5616 34000 5672
rect 14000 5584 34000 5616
rect 4260 5472 4580 5473
rect 4260 5408 4268 5472
rect 4332 5408 4348 5472
rect 4412 5408 4428 5472
rect 4492 5408 4508 5472
rect 4572 5408 4580 5472
rect 4260 5407 4580 5408
rect 7360 5472 7680 5473
rect 7360 5408 7368 5472
rect 7432 5408 7448 5472
rect 7512 5408 7528 5472
rect 7592 5408 7608 5472
rect 7672 5408 7680 5472
rect 7360 5407 7680 5408
rect 14000 5128 34000 5160
rect 14000 5072 14186 5128
rect 14242 5072 34000 5128
rect 14000 5040 34000 5072
rect 5810 4928 6130 4929
rect 5810 4864 5818 4928
rect 5882 4864 5898 4928
rect 5962 4864 5978 4928
rect 6042 4864 6058 4928
rect 6122 4864 6130 4928
rect 5810 4863 6130 4864
rect 8910 4928 9230 4929
rect 8910 4864 8918 4928
rect 8982 4864 8998 4928
rect 9062 4864 9078 4928
rect 9142 4864 9158 4928
rect 9222 4864 9230 4928
rect 8910 4863 9230 4864
rect 14000 4720 34000 4752
rect 14000 4664 14186 4720
rect 14242 4664 34000 4720
rect 14000 4632 34000 4664
rect 4260 4384 4580 4385
rect 4260 4320 4268 4384
rect 4332 4320 4348 4384
rect 4412 4320 4428 4384
rect 4492 4320 4508 4384
rect 4572 4320 4580 4384
rect 4260 4319 4580 4320
rect 7360 4384 7680 4385
rect 7360 4320 7368 4384
rect 7432 4320 7448 4384
rect 7512 4320 7528 4384
rect 7592 4320 7608 4384
rect 7672 4320 7680 4384
rect 7360 4319 7680 4320
rect 14000 4176 34000 4208
rect 14000 4120 14186 4176
rect 14242 4120 34000 4176
rect 14000 4088 34000 4120
rect 4153 4042 4219 4045
rect 3558 4040 4219 4042
rect 3558 3984 4158 4040
rect 4214 3984 4219 4040
rect 3558 3982 4219 3984
rect 3558 3876 3618 3982
rect 4153 3979 4219 3982
rect 5810 3840 6130 3841
rect 5810 3776 5818 3840
rect 5882 3776 5898 3840
rect 5962 3776 5978 3840
rect 6042 3776 6058 3840
rect 6122 3776 6130 3840
rect 5810 3775 6130 3776
rect 8910 3840 9230 3841
rect 8910 3776 8918 3840
rect 8982 3776 8998 3840
rect 9062 3776 9078 3840
rect 9142 3776 9158 3840
rect 9222 3776 9230 3840
rect 8910 3775 9230 3776
rect 14000 3632 34000 3664
rect 14000 3576 14186 3632
rect 14242 3576 34000 3632
rect 14000 3544 34000 3576
rect 4260 3296 4580 3297
rect 4260 3232 4268 3296
rect 4332 3232 4348 3296
rect 4412 3232 4428 3296
rect 4492 3232 4508 3296
rect 4572 3232 4580 3296
rect 4260 3231 4580 3232
rect 7360 3296 7680 3297
rect 7360 3232 7368 3296
rect 7432 3232 7448 3296
rect 7512 3232 7528 3296
rect 7592 3232 7608 3296
rect 7672 3232 7680 3296
rect 7360 3231 7680 3232
rect 14000 3224 34000 3256
rect 14000 3168 14186 3224
rect 14242 3168 34000 3224
rect 14000 3136 34000 3168
rect 5810 2752 6130 2753
rect 5810 2688 5818 2752
rect 5882 2688 5898 2752
rect 5962 2688 5978 2752
rect 6042 2688 6058 2752
rect 6122 2688 6130 2752
rect 5810 2687 6130 2688
rect 8910 2752 9230 2753
rect 8910 2688 8918 2752
rect 8982 2688 8998 2752
rect 9062 2688 9078 2752
rect 9142 2688 9158 2752
rect 9222 2688 9230 2752
rect 8910 2687 9230 2688
rect 14000 2680 34000 2712
rect 14000 2624 14186 2680
rect 14242 2624 34000 2680
rect 14000 2592 34000 2624
rect 4260 2208 4580 2209
rect 4260 2144 4268 2208
rect 4332 2144 4348 2208
rect 4412 2144 4428 2208
rect 4492 2144 4508 2208
rect 4572 2144 4580 2208
rect 4260 2143 4580 2144
rect 7360 2208 7680 2209
rect 7360 2144 7368 2208
rect 7432 2144 7448 2208
rect 7512 2144 7528 2208
rect 7592 2144 7608 2208
rect 7672 2144 7680 2208
rect 7360 2143 7680 2144
rect 14000 2136 34000 2168
rect 14000 2080 14278 2136
rect 14334 2080 34000 2136
rect 14000 2048 34000 2080
rect 14000 1728 34000 1760
rect 14000 1672 14278 1728
rect 14334 1672 34000 1728
rect 14000 1640 34000 1672
rect 14000 1184 34000 1216
rect 14000 1128 14278 1184
rect 14334 1128 34000 1184
rect 14000 1096 34000 1128
rect 14000 640 34000 672
rect 14000 584 14278 640
rect 14334 584 34000 640
rect 14000 552 34000 584
rect 14000 232 34000 264
rect 14000 176 14186 232
rect 14242 176 34000 232
rect 14000 144 34000 176
<< via3 >>
rect 2718 11452 2782 11456
rect 2718 11396 2722 11452
rect 2722 11396 2778 11452
rect 2778 11396 2782 11452
rect 2718 11392 2782 11396
rect 2798 11452 2862 11456
rect 2798 11396 2802 11452
rect 2802 11396 2858 11452
rect 2858 11396 2862 11452
rect 2798 11392 2862 11396
rect 2878 11452 2942 11456
rect 2878 11396 2882 11452
rect 2882 11396 2938 11452
rect 2938 11396 2942 11452
rect 2878 11392 2942 11396
rect 2958 11452 3022 11456
rect 2958 11396 2962 11452
rect 2962 11396 3018 11452
rect 3018 11396 3022 11452
rect 2958 11392 3022 11396
rect 5818 11452 5882 11456
rect 5818 11396 5822 11452
rect 5822 11396 5878 11452
rect 5878 11396 5882 11452
rect 5818 11392 5882 11396
rect 5898 11452 5962 11456
rect 5898 11396 5902 11452
rect 5902 11396 5958 11452
rect 5958 11396 5962 11452
rect 5898 11392 5962 11396
rect 5978 11452 6042 11456
rect 5978 11396 5982 11452
rect 5982 11396 6038 11452
rect 6038 11396 6042 11452
rect 5978 11392 6042 11396
rect 6058 11452 6122 11456
rect 6058 11396 6062 11452
rect 6062 11396 6118 11452
rect 6118 11396 6122 11452
rect 6058 11392 6122 11396
rect 8918 11452 8982 11456
rect 8918 11396 8922 11452
rect 8922 11396 8978 11452
rect 8978 11396 8982 11452
rect 8918 11392 8982 11396
rect 8998 11452 9062 11456
rect 8998 11396 9002 11452
rect 9002 11396 9058 11452
rect 9058 11396 9062 11452
rect 8998 11392 9062 11396
rect 9078 11452 9142 11456
rect 9078 11396 9082 11452
rect 9082 11396 9138 11452
rect 9138 11396 9142 11452
rect 9078 11392 9142 11396
rect 9158 11452 9222 11456
rect 9158 11396 9162 11452
rect 9162 11396 9218 11452
rect 9218 11396 9222 11452
rect 9158 11392 9222 11396
rect 1168 10908 1232 10912
rect 1168 10852 1172 10908
rect 1172 10852 1228 10908
rect 1228 10852 1232 10908
rect 1168 10848 1232 10852
rect 1248 10908 1312 10912
rect 1248 10852 1252 10908
rect 1252 10852 1308 10908
rect 1308 10852 1312 10908
rect 1248 10848 1312 10852
rect 1328 10908 1392 10912
rect 1328 10852 1332 10908
rect 1332 10852 1388 10908
rect 1388 10852 1392 10908
rect 1328 10848 1392 10852
rect 1408 10908 1472 10912
rect 1408 10852 1412 10908
rect 1412 10852 1468 10908
rect 1468 10852 1472 10908
rect 1408 10848 1472 10852
rect 4268 10908 4332 10912
rect 4268 10852 4272 10908
rect 4272 10852 4328 10908
rect 4328 10852 4332 10908
rect 4268 10848 4332 10852
rect 4348 10908 4412 10912
rect 4348 10852 4352 10908
rect 4352 10852 4408 10908
rect 4408 10852 4412 10908
rect 4348 10848 4412 10852
rect 4428 10908 4492 10912
rect 4428 10852 4432 10908
rect 4432 10852 4488 10908
rect 4488 10852 4492 10908
rect 4428 10848 4492 10852
rect 4508 10908 4572 10912
rect 4508 10852 4512 10908
rect 4512 10852 4568 10908
rect 4568 10852 4572 10908
rect 4508 10848 4572 10852
rect 7368 10908 7432 10912
rect 7368 10852 7372 10908
rect 7372 10852 7428 10908
rect 7428 10852 7432 10908
rect 7368 10848 7432 10852
rect 7448 10908 7512 10912
rect 7448 10852 7452 10908
rect 7452 10852 7508 10908
rect 7508 10852 7512 10908
rect 7448 10848 7512 10852
rect 7528 10908 7592 10912
rect 7528 10852 7532 10908
rect 7532 10852 7588 10908
rect 7588 10852 7592 10908
rect 7528 10848 7592 10852
rect 7608 10908 7672 10912
rect 7608 10852 7612 10908
rect 7612 10852 7668 10908
rect 7668 10852 7672 10908
rect 7608 10848 7672 10852
rect 2718 10364 2782 10368
rect 2718 10308 2722 10364
rect 2722 10308 2778 10364
rect 2778 10308 2782 10364
rect 2718 10304 2782 10308
rect 2798 10364 2862 10368
rect 2798 10308 2802 10364
rect 2802 10308 2858 10364
rect 2858 10308 2862 10364
rect 2798 10304 2862 10308
rect 2878 10364 2942 10368
rect 2878 10308 2882 10364
rect 2882 10308 2938 10364
rect 2938 10308 2942 10364
rect 2878 10304 2942 10308
rect 2958 10364 3022 10368
rect 2958 10308 2962 10364
rect 2962 10308 3018 10364
rect 3018 10308 3022 10364
rect 2958 10304 3022 10308
rect 5818 10364 5882 10368
rect 5818 10308 5822 10364
rect 5822 10308 5878 10364
rect 5878 10308 5882 10364
rect 5818 10304 5882 10308
rect 5898 10364 5962 10368
rect 5898 10308 5902 10364
rect 5902 10308 5958 10364
rect 5958 10308 5962 10364
rect 5898 10304 5962 10308
rect 5978 10364 6042 10368
rect 5978 10308 5982 10364
rect 5982 10308 6038 10364
rect 6038 10308 6042 10364
rect 5978 10304 6042 10308
rect 6058 10364 6122 10368
rect 6058 10308 6062 10364
rect 6062 10308 6118 10364
rect 6118 10308 6122 10364
rect 6058 10304 6122 10308
rect 8918 10364 8982 10368
rect 8918 10308 8922 10364
rect 8922 10308 8978 10364
rect 8978 10308 8982 10364
rect 8918 10304 8982 10308
rect 8998 10364 9062 10368
rect 8998 10308 9002 10364
rect 9002 10308 9058 10364
rect 9058 10308 9062 10364
rect 8998 10304 9062 10308
rect 9078 10364 9142 10368
rect 9078 10308 9082 10364
rect 9082 10308 9138 10364
rect 9138 10308 9142 10364
rect 9078 10304 9142 10308
rect 9158 10364 9222 10368
rect 9158 10308 9162 10364
rect 9162 10308 9218 10364
rect 9218 10308 9222 10364
rect 9158 10304 9222 10308
rect 1168 9820 1232 9824
rect 1168 9764 1172 9820
rect 1172 9764 1228 9820
rect 1228 9764 1232 9820
rect 1168 9760 1232 9764
rect 1248 9820 1312 9824
rect 1248 9764 1252 9820
rect 1252 9764 1308 9820
rect 1308 9764 1312 9820
rect 1248 9760 1312 9764
rect 1328 9820 1392 9824
rect 1328 9764 1332 9820
rect 1332 9764 1388 9820
rect 1388 9764 1392 9820
rect 1328 9760 1392 9764
rect 1408 9820 1472 9824
rect 1408 9764 1412 9820
rect 1412 9764 1468 9820
rect 1468 9764 1472 9820
rect 1408 9760 1472 9764
rect 4268 9820 4332 9824
rect 4268 9764 4272 9820
rect 4272 9764 4328 9820
rect 4328 9764 4332 9820
rect 4268 9760 4332 9764
rect 4348 9820 4412 9824
rect 4348 9764 4352 9820
rect 4352 9764 4408 9820
rect 4408 9764 4412 9820
rect 4348 9760 4412 9764
rect 4428 9820 4492 9824
rect 4428 9764 4432 9820
rect 4432 9764 4488 9820
rect 4488 9764 4492 9820
rect 4428 9760 4492 9764
rect 4508 9820 4572 9824
rect 4508 9764 4512 9820
rect 4512 9764 4568 9820
rect 4568 9764 4572 9820
rect 4508 9760 4572 9764
rect 7368 9820 7432 9824
rect 7368 9764 7372 9820
rect 7372 9764 7428 9820
rect 7428 9764 7432 9820
rect 7368 9760 7432 9764
rect 7448 9820 7512 9824
rect 7448 9764 7452 9820
rect 7452 9764 7508 9820
rect 7508 9764 7512 9820
rect 7448 9760 7512 9764
rect 7528 9820 7592 9824
rect 7528 9764 7532 9820
rect 7532 9764 7588 9820
rect 7588 9764 7592 9820
rect 7528 9760 7592 9764
rect 7608 9820 7672 9824
rect 7608 9764 7612 9820
rect 7612 9764 7668 9820
rect 7668 9764 7672 9820
rect 7608 9760 7672 9764
rect 2718 9276 2782 9280
rect 2718 9220 2722 9276
rect 2722 9220 2778 9276
rect 2778 9220 2782 9276
rect 2718 9216 2782 9220
rect 2798 9276 2862 9280
rect 2798 9220 2802 9276
rect 2802 9220 2858 9276
rect 2858 9220 2862 9276
rect 2798 9216 2862 9220
rect 2878 9276 2942 9280
rect 2878 9220 2882 9276
rect 2882 9220 2938 9276
rect 2938 9220 2942 9276
rect 2878 9216 2942 9220
rect 2958 9276 3022 9280
rect 2958 9220 2962 9276
rect 2962 9220 3018 9276
rect 3018 9220 3022 9276
rect 2958 9216 3022 9220
rect 5818 9276 5882 9280
rect 5818 9220 5822 9276
rect 5822 9220 5878 9276
rect 5878 9220 5882 9276
rect 5818 9216 5882 9220
rect 5898 9276 5962 9280
rect 5898 9220 5902 9276
rect 5902 9220 5958 9276
rect 5958 9220 5962 9276
rect 5898 9216 5962 9220
rect 5978 9276 6042 9280
rect 5978 9220 5982 9276
rect 5982 9220 6038 9276
rect 6038 9220 6042 9276
rect 5978 9216 6042 9220
rect 6058 9276 6122 9280
rect 6058 9220 6062 9276
rect 6062 9220 6118 9276
rect 6118 9220 6122 9276
rect 6058 9216 6122 9220
rect 8918 9276 8982 9280
rect 8918 9220 8922 9276
rect 8922 9220 8978 9276
rect 8978 9220 8982 9276
rect 8918 9216 8982 9220
rect 8998 9276 9062 9280
rect 8998 9220 9002 9276
rect 9002 9220 9058 9276
rect 9058 9220 9062 9276
rect 8998 9216 9062 9220
rect 9078 9276 9142 9280
rect 9078 9220 9082 9276
rect 9082 9220 9138 9276
rect 9138 9220 9142 9276
rect 9078 9216 9142 9220
rect 9158 9276 9222 9280
rect 9158 9220 9162 9276
rect 9162 9220 9218 9276
rect 9218 9220 9222 9276
rect 9158 9216 9222 9220
rect 1168 8732 1232 8736
rect 1168 8676 1172 8732
rect 1172 8676 1228 8732
rect 1228 8676 1232 8732
rect 1168 8672 1232 8676
rect 1248 8732 1312 8736
rect 1248 8676 1252 8732
rect 1252 8676 1308 8732
rect 1308 8676 1312 8732
rect 1248 8672 1312 8676
rect 1328 8732 1392 8736
rect 1328 8676 1332 8732
rect 1332 8676 1388 8732
rect 1388 8676 1392 8732
rect 1328 8672 1392 8676
rect 1408 8732 1472 8736
rect 1408 8676 1412 8732
rect 1412 8676 1468 8732
rect 1468 8676 1472 8732
rect 1408 8672 1472 8676
rect 4268 8732 4332 8736
rect 4268 8676 4272 8732
rect 4272 8676 4328 8732
rect 4328 8676 4332 8732
rect 4268 8672 4332 8676
rect 4348 8732 4412 8736
rect 4348 8676 4352 8732
rect 4352 8676 4408 8732
rect 4408 8676 4412 8732
rect 4348 8672 4412 8676
rect 4428 8732 4492 8736
rect 4428 8676 4432 8732
rect 4432 8676 4488 8732
rect 4488 8676 4492 8732
rect 4428 8672 4492 8676
rect 4508 8732 4572 8736
rect 4508 8676 4512 8732
rect 4512 8676 4568 8732
rect 4568 8676 4572 8732
rect 4508 8672 4572 8676
rect 7368 8732 7432 8736
rect 7368 8676 7372 8732
rect 7372 8676 7428 8732
rect 7428 8676 7432 8732
rect 7368 8672 7432 8676
rect 7448 8732 7512 8736
rect 7448 8676 7452 8732
rect 7452 8676 7508 8732
rect 7508 8676 7512 8732
rect 7448 8672 7512 8676
rect 7528 8732 7592 8736
rect 7528 8676 7532 8732
rect 7532 8676 7588 8732
rect 7588 8676 7592 8732
rect 7528 8672 7592 8676
rect 7608 8732 7672 8736
rect 7608 8676 7612 8732
rect 7612 8676 7668 8732
rect 7668 8676 7672 8732
rect 7608 8672 7672 8676
rect 2718 8188 2782 8192
rect 2718 8132 2722 8188
rect 2722 8132 2778 8188
rect 2778 8132 2782 8188
rect 2718 8128 2782 8132
rect 2798 8188 2862 8192
rect 2798 8132 2802 8188
rect 2802 8132 2858 8188
rect 2858 8132 2862 8188
rect 2798 8128 2862 8132
rect 2878 8188 2942 8192
rect 2878 8132 2882 8188
rect 2882 8132 2938 8188
rect 2938 8132 2942 8188
rect 2878 8128 2942 8132
rect 2958 8188 3022 8192
rect 2958 8132 2962 8188
rect 2962 8132 3018 8188
rect 3018 8132 3022 8188
rect 2958 8128 3022 8132
rect 5818 8188 5882 8192
rect 5818 8132 5822 8188
rect 5822 8132 5878 8188
rect 5878 8132 5882 8188
rect 5818 8128 5882 8132
rect 5898 8188 5962 8192
rect 5898 8132 5902 8188
rect 5902 8132 5958 8188
rect 5958 8132 5962 8188
rect 5898 8128 5962 8132
rect 5978 8188 6042 8192
rect 5978 8132 5982 8188
rect 5982 8132 6038 8188
rect 6038 8132 6042 8188
rect 5978 8128 6042 8132
rect 6058 8188 6122 8192
rect 6058 8132 6062 8188
rect 6062 8132 6118 8188
rect 6118 8132 6122 8188
rect 6058 8128 6122 8132
rect 8918 8188 8982 8192
rect 8918 8132 8922 8188
rect 8922 8132 8978 8188
rect 8978 8132 8982 8188
rect 8918 8128 8982 8132
rect 8998 8188 9062 8192
rect 8998 8132 9002 8188
rect 9002 8132 9058 8188
rect 9058 8132 9062 8188
rect 8998 8128 9062 8132
rect 9078 8188 9142 8192
rect 9078 8132 9082 8188
rect 9082 8132 9138 8188
rect 9138 8132 9142 8188
rect 9078 8128 9142 8132
rect 9158 8188 9222 8192
rect 9158 8132 9162 8188
rect 9162 8132 9218 8188
rect 9218 8132 9222 8188
rect 9158 8128 9222 8132
rect 1168 7644 1232 7648
rect 1168 7588 1172 7644
rect 1172 7588 1228 7644
rect 1228 7588 1232 7644
rect 1168 7584 1232 7588
rect 1248 7644 1312 7648
rect 1248 7588 1252 7644
rect 1252 7588 1308 7644
rect 1308 7588 1312 7644
rect 1248 7584 1312 7588
rect 1328 7644 1392 7648
rect 1328 7588 1332 7644
rect 1332 7588 1388 7644
rect 1388 7588 1392 7644
rect 1328 7584 1392 7588
rect 1408 7644 1472 7648
rect 1408 7588 1412 7644
rect 1412 7588 1468 7644
rect 1468 7588 1472 7644
rect 1408 7584 1472 7588
rect 4268 7644 4332 7648
rect 4268 7588 4272 7644
rect 4272 7588 4328 7644
rect 4328 7588 4332 7644
rect 4268 7584 4332 7588
rect 4348 7644 4412 7648
rect 4348 7588 4352 7644
rect 4352 7588 4408 7644
rect 4408 7588 4412 7644
rect 4348 7584 4412 7588
rect 4428 7644 4492 7648
rect 4428 7588 4432 7644
rect 4432 7588 4488 7644
rect 4488 7588 4492 7644
rect 4428 7584 4492 7588
rect 4508 7644 4572 7648
rect 4508 7588 4512 7644
rect 4512 7588 4568 7644
rect 4568 7588 4572 7644
rect 4508 7584 4572 7588
rect 7368 7644 7432 7648
rect 7368 7588 7372 7644
rect 7372 7588 7428 7644
rect 7428 7588 7432 7644
rect 7368 7584 7432 7588
rect 7448 7644 7512 7648
rect 7448 7588 7452 7644
rect 7452 7588 7508 7644
rect 7508 7588 7512 7644
rect 7448 7584 7512 7588
rect 7528 7644 7592 7648
rect 7528 7588 7532 7644
rect 7532 7588 7588 7644
rect 7588 7588 7592 7644
rect 7528 7584 7592 7588
rect 7608 7644 7672 7648
rect 7608 7588 7612 7644
rect 7612 7588 7668 7644
rect 7668 7588 7672 7644
rect 7608 7584 7672 7588
rect 2718 7100 2782 7104
rect 2718 7044 2722 7100
rect 2722 7044 2778 7100
rect 2778 7044 2782 7100
rect 2718 7040 2782 7044
rect 2798 7100 2862 7104
rect 2798 7044 2802 7100
rect 2802 7044 2858 7100
rect 2858 7044 2862 7100
rect 2798 7040 2862 7044
rect 2878 7100 2942 7104
rect 2878 7044 2882 7100
rect 2882 7044 2938 7100
rect 2938 7044 2942 7100
rect 2878 7040 2942 7044
rect 2958 7100 3022 7104
rect 2958 7044 2962 7100
rect 2962 7044 3018 7100
rect 3018 7044 3022 7100
rect 2958 7040 3022 7044
rect 5818 7100 5882 7104
rect 5818 7044 5822 7100
rect 5822 7044 5878 7100
rect 5878 7044 5882 7100
rect 5818 7040 5882 7044
rect 5898 7100 5962 7104
rect 5898 7044 5902 7100
rect 5902 7044 5958 7100
rect 5958 7044 5962 7100
rect 5898 7040 5962 7044
rect 5978 7100 6042 7104
rect 5978 7044 5982 7100
rect 5982 7044 6038 7100
rect 6038 7044 6042 7100
rect 5978 7040 6042 7044
rect 6058 7100 6122 7104
rect 6058 7044 6062 7100
rect 6062 7044 6118 7100
rect 6118 7044 6122 7100
rect 6058 7040 6122 7044
rect 8918 7100 8982 7104
rect 8918 7044 8922 7100
rect 8922 7044 8978 7100
rect 8978 7044 8982 7100
rect 8918 7040 8982 7044
rect 8998 7100 9062 7104
rect 8998 7044 9002 7100
rect 9002 7044 9058 7100
rect 9058 7044 9062 7100
rect 8998 7040 9062 7044
rect 9078 7100 9142 7104
rect 9078 7044 9082 7100
rect 9082 7044 9138 7100
rect 9138 7044 9142 7100
rect 9078 7040 9142 7044
rect 9158 7100 9222 7104
rect 9158 7044 9162 7100
rect 9162 7044 9218 7100
rect 9218 7044 9222 7100
rect 9158 7040 9222 7044
rect 1168 6556 1232 6560
rect 1168 6500 1172 6556
rect 1172 6500 1228 6556
rect 1228 6500 1232 6556
rect 1168 6496 1232 6500
rect 1248 6556 1312 6560
rect 1248 6500 1252 6556
rect 1252 6500 1308 6556
rect 1308 6500 1312 6556
rect 1248 6496 1312 6500
rect 1328 6556 1392 6560
rect 1328 6500 1332 6556
rect 1332 6500 1388 6556
rect 1388 6500 1392 6556
rect 1328 6496 1392 6500
rect 1408 6556 1472 6560
rect 1408 6500 1412 6556
rect 1412 6500 1468 6556
rect 1468 6500 1472 6556
rect 1408 6496 1472 6500
rect 4268 6556 4332 6560
rect 4268 6500 4272 6556
rect 4272 6500 4328 6556
rect 4328 6500 4332 6556
rect 4268 6496 4332 6500
rect 4348 6556 4412 6560
rect 4348 6500 4352 6556
rect 4352 6500 4408 6556
rect 4408 6500 4412 6556
rect 4348 6496 4412 6500
rect 4428 6556 4492 6560
rect 4428 6500 4432 6556
rect 4432 6500 4488 6556
rect 4488 6500 4492 6556
rect 4428 6496 4492 6500
rect 4508 6556 4572 6560
rect 4508 6500 4512 6556
rect 4512 6500 4568 6556
rect 4568 6500 4572 6556
rect 4508 6496 4572 6500
rect 7368 6556 7432 6560
rect 7368 6500 7372 6556
rect 7372 6500 7428 6556
rect 7428 6500 7432 6556
rect 7368 6496 7432 6500
rect 7448 6556 7512 6560
rect 7448 6500 7452 6556
rect 7452 6500 7508 6556
rect 7508 6500 7512 6556
rect 7448 6496 7512 6500
rect 7528 6556 7592 6560
rect 7528 6500 7532 6556
rect 7532 6500 7588 6556
rect 7588 6500 7592 6556
rect 7528 6496 7592 6500
rect 7608 6556 7672 6560
rect 7608 6500 7612 6556
rect 7612 6500 7668 6556
rect 7668 6500 7672 6556
rect 7608 6496 7672 6500
rect 2718 6012 2782 6016
rect 2718 5956 2722 6012
rect 2722 5956 2778 6012
rect 2778 5956 2782 6012
rect 2718 5952 2782 5956
rect 2798 6012 2862 6016
rect 2798 5956 2802 6012
rect 2802 5956 2858 6012
rect 2858 5956 2862 6012
rect 2798 5952 2862 5956
rect 2878 6012 2942 6016
rect 2878 5956 2882 6012
rect 2882 5956 2938 6012
rect 2938 5956 2942 6012
rect 2878 5952 2942 5956
rect 2958 6012 3022 6016
rect 2958 5956 2962 6012
rect 2962 5956 3018 6012
rect 3018 5956 3022 6012
rect 2958 5952 3022 5956
rect 5818 6012 5882 6016
rect 5818 5956 5822 6012
rect 5822 5956 5878 6012
rect 5878 5956 5882 6012
rect 5818 5952 5882 5956
rect 5898 6012 5962 6016
rect 5898 5956 5902 6012
rect 5902 5956 5958 6012
rect 5958 5956 5962 6012
rect 5898 5952 5962 5956
rect 5978 6012 6042 6016
rect 5978 5956 5982 6012
rect 5982 5956 6038 6012
rect 6038 5956 6042 6012
rect 5978 5952 6042 5956
rect 6058 6012 6122 6016
rect 6058 5956 6062 6012
rect 6062 5956 6118 6012
rect 6118 5956 6122 6012
rect 6058 5952 6122 5956
rect 8918 6012 8982 6016
rect 8918 5956 8922 6012
rect 8922 5956 8978 6012
rect 8978 5956 8982 6012
rect 8918 5952 8982 5956
rect 8998 6012 9062 6016
rect 8998 5956 9002 6012
rect 9002 5956 9058 6012
rect 9058 5956 9062 6012
rect 8998 5952 9062 5956
rect 9078 6012 9142 6016
rect 9078 5956 9082 6012
rect 9082 5956 9138 6012
rect 9138 5956 9142 6012
rect 9078 5952 9142 5956
rect 9158 6012 9222 6016
rect 9158 5956 9162 6012
rect 9162 5956 9218 6012
rect 9218 5956 9222 6012
rect 9158 5952 9222 5956
rect 4268 5468 4332 5472
rect 4268 5412 4272 5468
rect 4272 5412 4328 5468
rect 4328 5412 4332 5468
rect 4268 5408 4332 5412
rect 4348 5468 4412 5472
rect 4348 5412 4352 5468
rect 4352 5412 4408 5468
rect 4408 5412 4412 5468
rect 4348 5408 4412 5412
rect 4428 5468 4492 5472
rect 4428 5412 4432 5468
rect 4432 5412 4488 5468
rect 4488 5412 4492 5468
rect 4428 5408 4492 5412
rect 4508 5468 4572 5472
rect 4508 5412 4512 5468
rect 4512 5412 4568 5468
rect 4568 5412 4572 5468
rect 4508 5408 4572 5412
rect 7368 5468 7432 5472
rect 7368 5412 7372 5468
rect 7372 5412 7428 5468
rect 7428 5412 7432 5468
rect 7368 5408 7432 5412
rect 7448 5468 7512 5472
rect 7448 5412 7452 5468
rect 7452 5412 7508 5468
rect 7508 5412 7512 5468
rect 7448 5408 7512 5412
rect 7528 5468 7592 5472
rect 7528 5412 7532 5468
rect 7532 5412 7588 5468
rect 7588 5412 7592 5468
rect 7528 5408 7592 5412
rect 7608 5468 7672 5472
rect 7608 5412 7612 5468
rect 7612 5412 7668 5468
rect 7668 5412 7672 5468
rect 7608 5408 7672 5412
rect 5818 4924 5882 4928
rect 5818 4868 5822 4924
rect 5822 4868 5878 4924
rect 5878 4868 5882 4924
rect 5818 4864 5882 4868
rect 5898 4924 5962 4928
rect 5898 4868 5902 4924
rect 5902 4868 5958 4924
rect 5958 4868 5962 4924
rect 5898 4864 5962 4868
rect 5978 4924 6042 4928
rect 5978 4868 5982 4924
rect 5982 4868 6038 4924
rect 6038 4868 6042 4924
rect 5978 4864 6042 4868
rect 6058 4924 6122 4928
rect 6058 4868 6062 4924
rect 6062 4868 6118 4924
rect 6118 4868 6122 4924
rect 6058 4864 6122 4868
rect 8918 4924 8982 4928
rect 8918 4868 8922 4924
rect 8922 4868 8978 4924
rect 8978 4868 8982 4924
rect 8918 4864 8982 4868
rect 8998 4924 9062 4928
rect 8998 4868 9002 4924
rect 9002 4868 9058 4924
rect 9058 4868 9062 4924
rect 8998 4864 9062 4868
rect 9078 4924 9142 4928
rect 9078 4868 9082 4924
rect 9082 4868 9138 4924
rect 9138 4868 9142 4924
rect 9078 4864 9142 4868
rect 9158 4924 9222 4928
rect 9158 4868 9162 4924
rect 9162 4868 9218 4924
rect 9218 4868 9222 4924
rect 9158 4864 9222 4868
rect 4268 4380 4332 4384
rect 4268 4324 4272 4380
rect 4272 4324 4328 4380
rect 4328 4324 4332 4380
rect 4268 4320 4332 4324
rect 4348 4380 4412 4384
rect 4348 4324 4352 4380
rect 4352 4324 4408 4380
rect 4408 4324 4412 4380
rect 4348 4320 4412 4324
rect 4428 4380 4492 4384
rect 4428 4324 4432 4380
rect 4432 4324 4488 4380
rect 4488 4324 4492 4380
rect 4428 4320 4492 4324
rect 4508 4380 4572 4384
rect 4508 4324 4512 4380
rect 4512 4324 4568 4380
rect 4568 4324 4572 4380
rect 4508 4320 4572 4324
rect 7368 4380 7432 4384
rect 7368 4324 7372 4380
rect 7372 4324 7428 4380
rect 7428 4324 7432 4380
rect 7368 4320 7432 4324
rect 7448 4380 7512 4384
rect 7448 4324 7452 4380
rect 7452 4324 7508 4380
rect 7508 4324 7512 4380
rect 7448 4320 7512 4324
rect 7528 4380 7592 4384
rect 7528 4324 7532 4380
rect 7532 4324 7588 4380
rect 7588 4324 7592 4380
rect 7528 4320 7592 4324
rect 7608 4380 7672 4384
rect 7608 4324 7612 4380
rect 7612 4324 7668 4380
rect 7668 4324 7672 4380
rect 7608 4320 7672 4324
rect 5818 3836 5882 3840
rect 5818 3780 5822 3836
rect 5822 3780 5878 3836
rect 5878 3780 5882 3836
rect 5818 3776 5882 3780
rect 5898 3836 5962 3840
rect 5898 3780 5902 3836
rect 5902 3780 5958 3836
rect 5958 3780 5962 3836
rect 5898 3776 5962 3780
rect 5978 3836 6042 3840
rect 5978 3780 5982 3836
rect 5982 3780 6038 3836
rect 6038 3780 6042 3836
rect 5978 3776 6042 3780
rect 6058 3836 6122 3840
rect 6058 3780 6062 3836
rect 6062 3780 6118 3836
rect 6118 3780 6122 3836
rect 6058 3776 6122 3780
rect 8918 3836 8982 3840
rect 8918 3780 8922 3836
rect 8922 3780 8978 3836
rect 8978 3780 8982 3836
rect 8918 3776 8982 3780
rect 8998 3836 9062 3840
rect 8998 3780 9002 3836
rect 9002 3780 9058 3836
rect 9058 3780 9062 3836
rect 8998 3776 9062 3780
rect 9078 3836 9142 3840
rect 9078 3780 9082 3836
rect 9082 3780 9138 3836
rect 9138 3780 9142 3836
rect 9078 3776 9142 3780
rect 9158 3836 9222 3840
rect 9158 3780 9162 3836
rect 9162 3780 9218 3836
rect 9218 3780 9222 3836
rect 9158 3776 9222 3780
rect 4268 3292 4332 3296
rect 4268 3236 4272 3292
rect 4272 3236 4328 3292
rect 4328 3236 4332 3292
rect 4268 3232 4332 3236
rect 4348 3292 4412 3296
rect 4348 3236 4352 3292
rect 4352 3236 4408 3292
rect 4408 3236 4412 3292
rect 4348 3232 4412 3236
rect 4428 3292 4492 3296
rect 4428 3236 4432 3292
rect 4432 3236 4488 3292
rect 4488 3236 4492 3292
rect 4428 3232 4492 3236
rect 4508 3292 4572 3296
rect 4508 3236 4512 3292
rect 4512 3236 4568 3292
rect 4568 3236 4572 3292
rect 4508 3232 4572 3236
rect 7368 3292 7432 3296
rect 7368 3236 7372 3292
rect 7372 3236 7428 3292
rect 7428 3236 7432 3292
rect 7368 3232 7432 3236
rect 7448 3292 7512 3296
rect 7448 3236 7452 3292
rect 7452 3236 7508 3292
rect 7508 3236 7512 3292
rect 7448 3232 7512 3236
rect 7528 3292 7592 3296
rect 7528 3236 7532 3292
rect 7532 3236 7588 3292
rect 7588 3236 7592 3292
rect 7528 3232 7592 3236
rect 7608 3292 7672 3296
rect 7608 3236 7612 3292
rect 7612 3236 7668 3292
rect 7668 3236 7672 3292
rect 7608 3232 7672 3236
rect 5818 2748 5882 2752
rect 5818 2692 5822 2748
rect 5822 2692 5878 2748
rect 5878 2692 5882 2748
rect 5818 2688 5882 2692
rect 5898 2748 5962 2752
rect 5898 2692 5902 2748
rect 5902 2692 5958 2748
rect 5958 2692 5962 2748
rect 5898 2688 5962 2692
rect 5978 2748 6042 2752
rect 5978 2692 5982 2748
rect 5982 2692 6038 2748
rect 6038 2692 6042 2748
rect 5978 2688 6042 2692
rect 6058 2748 6122 2752
rect 6058 2692 6062 2748
rect 6062 2692 6118 2748
rect 6118 2692 6122 2748
rect 6058 2688 6122 2692
rect 8918 2748 8982 2752
rect 8918 2692 8922 2748
rect 8922 2692 8978 2748
rect 8978 2692 8982 2748
rect 8918 2688 8982 2692
rect 8998 2748 9062 2752
rect 8998 2692 9002 2748
rect 9002 2692 9058 2748
rect 9058 2692 9062 2748
rect 8998 2688 9062 2692
rect 9078 2748 9142 2752
rect 9078 2692 9082 2748
rect 9082 2692 9138 2748
rect 9138 2692 9142 2748
rect 9078 2688 9142 2692
rect 9158 2748 9222 2752
rect 9158 2692 9162 2748
rect 9162 2692 9218 2748
rect 9218 2692 9222 2748
rect 9158 2688 9222 2692
rect 4268 2204 4332 2208
rect 4268 2148 4272 2204
rect 4272 2148 4328 2204
rect 4328 2148 4332 2204
rect 4268 2144 4332 2148
rect 4348 2204 4412 2208
rect 4348 2148 4352 2204
rect 4352 2148 4408 2204
rect 4408 2148 4412 2204
rect 4348 2144 4412 2148
rect 4428 2204 4492 2208
rect 4428 2148 4432 2204
rect 4432 2148 4488 2204
rect 4488 2148 4492 2204
rect 4428 2144 4492 2148
rect 4508 2204 4572 2208
rect 4508 2148 4512 2204
rect 4512 2148 4568 2204
rect 4568 2148 4572 2204
rect 4508 2144 4572 2148
rect 7368 2204 7432 2208
rect 7368 2148 7372 2204
rect 7372 2148 7428 2204
rect 7428 2148 7432 2204
rect 7368 2144 7432 2148
rect 7448 2204 7512 2208
rect 7448 2148 7452 2204
rect 7452 2148 7508 2204
rect 7508 2148 7512 2204
rect 7448 2144 7512 2148
rect 7528 2204 7592 2208
rect 7528 2148 7532 2204
rect 7532 2148 7588 2204
rect 7588 2148 7592 2204
rect 7528 2144 7592 2148
rect 7608 2204 7672 2208
rect 7608 2148 7612 2204
rect 7612 2148 7668 2204
rect 7668 2148 7672 2204
rect 7608 2144 7672 2148
<< metal4 >>
rect -1620 13922 -1300 13964
rect -1620 13686 -1578 13922
rect -1342 13686 -1300 13922
rect -1620 8244 -1300 13686
rect -1620 8008 -1578 8244
rect -1342 8008 -1300 8244
rect -1620 5144 -1300 8008
rect -1620 4908 -1578 5144
rect -1342 4908 -1300 5144
rect -1620 -86 -1300 4908
rect -960 13262 -640 13304
rect -960 13026 -918 13262
rect -682 13026 -640 13262
rect -960 9794 -640 13026
rect 2060 13262 2380 13964
rect 2060 13026 2102 13262
rect 2338 13026 2380 13262
rect -960 9558 -918 9794
rect -682 9558 -640 9794
rect -960 6694 -640 9558
rect -960 6458 -918 6694
rect -682 6458 -640 6694
rect -960 3594 -640 6458
rect -960 3358 -918 3594
rect -682 3358 -640 3594
rect -960 574 -640 3358
rect -300 12602 20 12644
rect -300 12366 -258 12602
rect -22 12366 20 12602
rect -300 10444 20 12366
rect -300 10208 -258 10444
rect -22 10208 20 10444
rect -300 7344 20 10208
rect -300 7108 -258 7344
rect -22 7108 20 7344
rect -300 4244 20 7108
rect -300 4008 -258 4244
rect -22 4008 20 4244
rect -300 1234 20 4008
rect 360 11942 680 11984
rect 360 11706 402 11942
rect 638 11706 680 11942
rect 360 8894 680 11706
rect 360 8658 402 8894
rect 638 8658 680 8894
rect 360 5794 680 8658
rect 360 5558 402 5794
rect 638 5558 680 5794
rect 1160 11942 1480 12644
rect 1160 11706 1202 11942
rect 1438 11706 1480 11942
rect 1160 10912 1480 11706
rect 1160 10848 1168 10912
rect 1232 10848 1248 10912
rect 1312 10848 1328 10912
rect 1392 10848 1408 10912
rect 1472 10848 1480 10912
rect 1160 9824 1480 10848
rect 1160 9760 1168 9824
rect 1232 9760 1248 9824
rect 1312 9760 1328 9824
rect 1392 9760 1408 9824
rect 1472 9760 1480 9824
rect 1160 8894 1480 9760
rect 1160 8736 1202 8894
rect 1438 8736 1480 8894
rect 1160 8672 1168 8736
rect 1472 8672 1480 8736
rect 1160 8658 1202 8672
rect 1438 8658 1480 8672
rect 1160 7648 1480 8658
rect 1160 7584 1168 7648
rect 1232 7584 1248 7648
rect 1312 7584 1328 7648
rect 1392 7584 1408 7648
rect 1472 7584 1480 7648
rect 1160 6560 1480 7584
rect 1160 6496 1168 6560
rect 1232 6496 1248 6560
rect 1312 6496 1328 6560
rect 1392 6496 1408 6560
rect 1472 6496 1480 6560
rect 1160 5632 1480 6496
rect 2060 9794 2380 13026
rect 3610 13922 3930 13964
rect 3610 13686 3652 13922
rect 3888 13686 3930 13922
rect 2060 9558 2102 9794
rect 2338 9558 2380 9794
rect 2060 6694 2380 9558
rect 2060 6458 2102 6694
rect 2338 6458 2380 6694
rect 2060 5680 2380 6458
rect 2710 12602 3030 12644
rect 2710 12366 2752 12602
rect 2988 12366 3030 12602
rect 2710 11456 3030 12366
rect 2710 11392 2718 11456
rect 2782 11392 2798 11456
rect 2862 11392 2878 11456
rect 2942 11392 2958 11456
rect 3022 11392 3030 11456
rect 2710 10444 3030 11392
rect 2710 10368 2752 10444
rect 2988 10368 3030 10444
rect 2710 10304 2718 10368
rect 3022 10304 3030 10368
rect 2710 10208 2752 10304
rect 2988 10208 3030 10304
rect 2710 9280 3030 10208
rect 2710 9216 2718 9280
rect 2782 9216 2798 9280
rect 2862 9216 2878 9280
rect 2942 9216 2958 9280
rect 3022 9216 3030 9280
rect 2710 8192 3030 9216
rect 2710 8128 2718 8192
rect 2782 8128 2798 8192
rect 2862 8128 2878 8192
rect 2942 8128 2958 8192
rect 3022 8128 3030 8192
rect 2710 7344 3030 8128
rect 2710 7108 2752 7344
rect 2988 7108 3030 7344
rect 2710 7104 3030 7108
rect 2710 7040 2718 7104
rect 2782 7040 2798 7104
rect 2862 7040 2878 7104
rect 2942 7040 2958 7104
rect 3022 7040 3030 7104
rect 2710 6016 3030 7040
rect 2710 5952 2718 6016
rect 2782 5952 2798 6016
rect 2862 5952 2878 6016
rect 2942 5952 2958 6016
rect 3022 5952 3030 6016
rect 2710 5632 3030 5952
rect 3610 8244 3930 13686
rect 5160 13262 5480 13964
rect 5160 13026 5202 13262
rect 5438 13026 5480 13262
rect 3610 8008 3652 8244
rect 3888 8008 3930 8244
rect 3610 5680 3930 8008
rect 4260 11942 4580 12644
rect 4260 11706 4302 11942
rect 4538 11706 4580 11942
rect 4260 10912 4580 11706
rect 4260 10848 4268 10912
rect 4332 10848 4348 10912
rect 4412 10848 4428 10912
rect 4492 10848 4508 10912
rect 4572 10848 4580 10912
rect 4260 9824 4580 10848
rect 4260 9760 4268 9824
rect 4332 9760 4348 9824
rect 4412 9760 4428 9824
rect 4492 9760 4508 9824
rect 4572 9760 4580 9824
rect 4260 8894 4580 9760
rect 4260 8736 4302 8894
rect 4538 8736 4580 8894
rect 4260 8672 4268 8736
rect 4572 8672 4580 8736
rect 4260 8658 4302 8672
rect 4538 8658 4580 8672
rect 4260 7648 4580 8658
rect 4260 7584 4268 7648
rect 4332 7584 4348 7648
rect 4412 7584 4428 7648
rect 4492 7584 4508 7648
rect 4572 7584 4580 7648
rect 4260 6560 4580 7584
rect 4260 6496 4268 6560
rect 4332 6496 4348 6560
rect 4412 6496 4428 6560
rect 4492 6496 4508 6560
rect 4572 6496 4580 6560
rect 4260 5794 4580 6496
rect 360 2694 680 5558
rect 4260 5558 4302 5794
rect 4538 5558 4580 5794
rect 4260 5472 4580 5558
rect 4260 5408 4268 5472
rect 4332 5408 4348 5472
rect 4412 5408 4428 5472
rect 4492 5408 4508 5472
rect 4572 5408 4580 5472
rect 1878 5144 2114 5186
rect 1878 4866 2114 4908
rect 2678 5144 2914 5186
rect 2678 4866 2914 4908
rect 4260 4384 4580 5408
rect 4260 4320 4268 4384
rect 4332 4320 4348 4384
rect 4412 4320 4428 4384
rect 4492 4320 4508 4384
rect 4572 4320 4580 4384
rect 1478 3594 1714 3636
rect 1478 3316 1714 3358
rect 2278 3594 2514 3636
rect 2278 3316 2514 3358
rect 3078 3594 3314 3636
rect 3078 3316 3314 3358
rect 360 2458 402 2694
rect 638 2458 680 2694
rect 360 1894 680 2458
rect 4260 3296 4580 4320
rect 4260 3232 4268 3296
rect 4332 3232 4348 3296
rect 4412 3232 4428 3296
rect 4492 3232 4508 3296
rect 4572 3232 4580 3296
rect 4260 2694 4580 3232
rect 4260 2458 4302 2694
rect 4538 2458 4580 2694
rect 4260 2208 4580 2458
rect 4260 2144 4268 2208
rect 4332 2144 4348 2208
rect 4412 2144 4428 2208
rect 4492 2144 4508 2208
rect 4572 2144 4580 2208
rect 360 1658 402 1894
rect 638 1658 680 1894
rect 360 1616 680 1658
rect 1160 1894 1480 2128
rect 1160 1658 1202 1894
rect 1438 1658 1480 1894
rect -300 998 -258 1234
rect -22 998 20 1234
rect -300 956 20 998
rect 1160 956 1480 1658
rect -960 338 -918 574
rect -682 338 -640 574
rect -960 296 -640 338
rect 2060 574 2380 2080
rect 2710 1234 3030 2128
rect 2710 998 2752 1234
rect 2988 998 3030 1234
rect 2710 956 3030 998
rect 2060 338 2102 574
rect 2338 338 2380 574
rect -1620 -322 -1578 -86
rect -1342 -322 -1300 -86
rect -1620 -364 -1300 -322
rect 2060 -364 2380 338
rect 3610 -86 3930 2080
rect 4260 1894 4580 2144
rect 4260 1658 4302 1894
rect 4538 1658 4580 1894
rect 4260 956 4580 1658
rect 5160 9794 5480 13026
rect 6710 13922 7030 13964
rect 6710 13686 6752 13922
rect 6988 13686 7030 13922
rect 5160 9558 5202 9794
rect 5438 9558 5480 9794
rect 5160 6694 5480 9558
rect 5160 6458 5202 6694
rect 5438 6458 5480 6694
rect 5160 3594 5480 6458
rect 5160 3358 5202 3594
rect 5438 3358 5480 3594
rect 3610 -322 3652 -86
rect 3888 -322 3930 -86
rect 3610 -364 3930 -322
rect 5160 574 5480 3358
rect 5810 12602 6130 12644
rect 5810 12366 5852 12602
rect 6088 12366 6130 12602
rect 5810 11456 6130 12366
rect 5810 11392 5818 11456
rect 5882 11392 5898 11456
rect 5962 11392 5978 11456
rect 6042 11392 6058 11456
rect 6122 11392 6130 11456
rect 5810 10444 6130 11392
rect 5810 10368 5852 10444
rect 6088 10368 6130 10444
rect 5810 10304 5818 10368
rect 6122 10304 6130 10368
rect 5810 10208 5852 10304
rect 6088 10208 6130 10304
rect 5810 9280 6130 10208
rect 5810 9216 5818 9280
rect 5882 9216 5898 9280
rect 5962 9216 5978 9280
rect 6042 9216 6058 9280
rect 6122 9216 6130 9280
rect 5810 8192 6130 9216
rect 5810 8128 5818 8192
rect 5882 8128 5898 8192
rect 5962 8128 5978 8192
rect 6042 8128 6058 8192
rect 6122 8128 6130 8192
rect 5810 7344 6130 8128
rect 5810 7108 5852 7344
rect 6088 7108 6130 7344
rect 5810 7104 6130 7108
rect 5810 7040 5818 7104
rect 5882 7040 5898 7104
rect 5962 7040 5978 7104
rect 6042 7040 6058 7104
rect 6122 7040 6130 7104
rect 5810 6016 6130 7040
rect 5810 5952 5818 6016
rect 5882 5952 5898 6016
rect 5962 5952 5978 6016
rect 6042 5952 6058 6016
rect 6122 5952 6130 6016
rect 5810 4928 6130 5952
rect 5810 4864 5818 4928
rect 5882 4864 5898 4928
rect 5962 4864 5978 4928
rect 6042 4864 6058 4928
rect 6122 4864 6130 4928
rect 5810 4244 6130 4864
rect 5810 4008 5852 4244
rect 6088 4008 6130 4244
rect 5810 3840 6130 4008
rect 5810 3776 5818 3840
rect 5882 3776 5898 3840
rect 5962 3776 5978 3840
rect 6042 3776 6058 3840
rect 6122 3776 6130 3840
rect 5810 2752 6130 3776
rect 5810 2688 5818 2752
rect 5882 2688 5898 2752
rect 5962 2688 5978 2752
rect 6042 2688 6058 2752
rect 6122 2688 6130 2752
rect 5810 1234 6130 2688
rect 5810 998 5852 1234
rect 6088 998 6130 1234
rect 5810 956 6130 998
rect 6710 8244 7030 13686
rect 8260 13262 8580 13964
rect 12064 13922 12384 13964
rect 12064 13686 12106 13922
rect 12342 13686 12384 13922
rect 8260 13026 8302 13262
rect 8538 13026 8580 13262
rect 6710 8008 6752 8244
rect 6988 8008 7030 8244
rect 6710 5144 7030 8008
rect 6710 4908 6752 5144
rect 6988 4908 7030 5144
rect 5160 338 5202 574
rect 5438 338 5480 574
rect 5160 -364 5480 338
rect 6710 -86 7030 4908
rect 7360 11942 7680 12644
rect 7360 11706 7402 11942
rect 7638 11706 7680 11942
rect 7360 10912 7680 11706
rect 7360 10848 7368 10912
rect 7432 10848 7448 10912
rect 7512 10848 7528 10912
rect 7592 10848 7608 10912
rect 7672 10848 7680 10912
rect 7360 9824 7680 10848
rect 7360 9760 7368 9824
rect 7432 9760 7448 9824
rect 7512 9760 7528 9824
rect 7592 9760 7608 9824
rect 7672 9760 7680 9824
rect 7360 8894 7680 9760
rect 7360 8736 7402 8894
rect 7638 8736 7680 8894
rect 7360 8672 7368 8736
rect 7672 8672 7680 8736
rect 7360 8658 7402 8672
rect 7638 8658 7680 8672
rect 7360 7648 7680 8658
rect 7360 7584 7368 7648
rect 7432 7584 7448 7648
rect 7512 7584 7528 7648
rect 7592 7584 7608 7648
rect 7672 7584 7680 7648
rect 7360 6560 7680 7584
rect 7360 6496 7368 6560
rect 7432 6496 7448 6560
rect 7512 6496 7528 6560
rect 7592 6496 7608 6560
rect 7672 6496 7680 6560
rect 7360 5794 7680 6496
rect 7360 5558 7402 5794
rect 7638 5558 7680 5794
rect 7360 5472 7680 5558
rect 7360 5408 7368 5472
rect 7432 5408 7448 5472
rect 7512 5408 7528 5472
rect 7592 5408 7608 5472
rect 7672 5408 7680 5472
rect 7360 4384 7680 5408
rect 7360 4320 7368 4384
rect 7432 4320 7448 4384
rect 7512 4320 7528 4384
rect 7592 4320 7608 4384
rect 7672 4320 7680 4384
rect 7360 3296 7680 4320
rect 7360 3232 7368 3296
rect 7432 3232 7448 3296
rect 7512 3232 7528 3296
rect 7592 3232 7608 3296
rect 7672 3232 7680 3296
rect 7360 2694 7680 3232
rect 7360 2458 7402 2694
rect 7638 2458 7680 2694
rect 7360 2208 7680 2458
rect 7360 2144 7368 2208
rect 7432 2144 7448 2208
rect 7512 2144 7528 2208
rect 7592 2144 7608 2208
rect 7672 2144 7680 2208
rect 7360 1894 7680 2144
rect 7360 1658 7402 1894
rect 7638 1658 7680 1894
rect 7360 956 7680 1658
rect 8260 9794 8580 13026
rect 11404 13262 11724 13304
rect 11404 13026 11446 13262
rect 11682 13026 11724 13262
rect 8260 9558 8302 9794
rect 8538 9558 8580 9794
rect 8260 6694 8580 9558
rect 8260 6458 8302 6694
rect 8538 6458 8580 6694
rect 8260 3594 8580 6458
rect 8260 3358 8302 3594
rect 8538 3358 8580 3594
rect 6710 -322 6752 -86
rect 6988 -322 7030 -86
rect 6710 -364 7030 -322
rect 8260 574 8580 3358
rect 8910 12602 9230 12644
rect 8910 12366 8952 12602
rect 9188 12366 9230 12602
rect 8910 11456 9230 12366
rect 10744 12602 11064 12644
rect 10744 12366 10786 12602
rect 11022 12366 11064 12602
rect 8910 11392 8918 11456
rect 8982 11392 8998 11456
rect 9062 11392 9078 11456
rect 9142 11392 9158 11456
rect 9222 11392 9230 11456
rect 8910 10444 9230 11392
rect 8910 10368 8952 10444
rect 9188 10368 9230 10444
rect 8910 10304 8918 10368
rect 9222 10304 9230 10368
rect 8910 10208 8952 10304
rect 9188 10208 9230 10304
rect 8910 9280 9230 10208
rect 8910 9216 8918 9280
rect 8982 9216 8998 9280
rect 9062 9216 9078 9280
rect 9142 9216 9158 9280
rect 9222 9216 9230 9280
rect 8910 8192 9230 9216
rect 8910 8128 8918 8192
rect 8982 8128 8998 8192
rect 9062 8128 9078 8192
rect 9142 8128 9158 8192
rect 9222 8128 9230 8192
rect 8910 7344 9230 8128
rect 8910 7108 8952 7344
rect 9188 7108 9230 7344
rect 8910 7104 9230 7108
rect 8910 7040 8918 7104
rect 8982 7040 8998 7104
rect 9062 7040 9078 7104
rect 9142 7040 9158 7104
rect 9222 7040 9230 7104
rect 8910 6016 9230 7040
rect 8910 5952 8918 6016
rect 8982 5952 8998 6016
rect 9062 5952 9078 6016
rect 9142 5952 9158 6016
rect 9222 5952 9230 6016
rect 8910 4928 9230 5952
rect 8910 4864 8918 4928
rect 8982 4864 8998 4928
rect 9062 4864 9078 4928
rect 9142 4864 9158 4928
rect 9222 4864 9230 4928
rect 8910 4244 9230 4864
rect 8910 4008 8952 4244
rect 9188 4008 9230 4244
rect 8910 3840 9230 4008
rect 8910 3776 8918 3840
rect 8982 3776 8998 3840
rect 9062 3776 9078 3840
rect 9142 3776 9158 3840
rect 9222 3776 9230 3840
rect 8910 2752 9230 3776
rect 8910 2688 8918 2752
rect 8982 2688 8998 2752
rect 9062 2688 9078 2752
rect 9142 2688 9158 2752
rect 9222 2688 9230 2752
rect 8910 1234 9230 2688
rect 10084 11942 10404 11984
rect 10084 11706 10126 11942
rect 10362 11706 10404 11942
rect 10084 8894 10404 11706
rect 10084 8658 10126 8894
rect 10362 8658 10404 8894
rect 10084 5794 10404 8658
rect 10084 5558 10126 5794
rect 10362 5558 10404 5794
rect 10084 2694 10404 5558
rect 10084 2458 10126 2694
rect 10362 2458 10404 2694
rect 10084 1894 10404 2458
rect 10084 1658 10126 1894
rect 10362 1658 10404 1894
rect 10084 1616 10404 1658
rect 10744 10444 11064 12366
rect 10744 10208 10786 10444
rect 11022 10208 11064 10444
rect 10744 7344 11064 10208
rect 10744 7108 10786 7344
rect 11022 7108 11064 7344
rect 10744 4244 11064 7108
rect 10744 4008 10786 4244
rect 11022 4008 11064 4244
rect 8910 998 8952 1234
rect 9188 998 9230 1234
rect 8910 956 9230 998
rect 10744 1234 11064 4008
rect 10744 998 10786 1234
rect 11022 998 11064 1234
rect 10744 956 11064 998
rect 11404 9794 11724 13026
rect 11404 9558 11446 9794
rect 11682 9558 11724 9794
rect 11404 6694 11724 9558
rect 11404 6458 11446 6694
rect 11682 6458 11724 6694
rect 11404 3594 11724 6458
rect 11404 3358 11446 3594
rect 11682 3358 11724 3594
rect 8260 338 8302 574
rect 8538 338 8580 574
rect 8260 -364 8580 338
rect 11404 574 11724 3358
rect 11404 338 11446 574
rect 11682 338 11724 574
rect 11404 296 11724 338
rect 12064 8244 12384 13686
rect 12064 8008 12106 8244
rect 12342 8008 12384 8244
rect 12064 5144 12384 8008
rect 12064 4908 12106 5144
rect 12342 4908 12384 5144
rect 12064 -86 12384 4908
rect 12064 -322 12106 -86
rect 12342 -322 12384 -86
rect 12064 -364 12384 -322
<< via4 >>
rect -1578 13686 -1342 13922
rect -1578 8008 -1342 8244
rect -1578 4908 -1342 5144
rect -918 13026 -682 13262
rect 2102 13026 2338 13262
rect -918 9558 -682 9794
rect -918 6458 -682 6694
rect -918 3358 -682 3594
rect -258 12366 -22 12602
rect -258 10208 -22 10444
rect -258 7108 -22 7344
rect -258 4008 -22 4244
rect 402 11706 638 11942
rect 402 8658 638 8894
rect 402 5558 638 5794
rect 1202 11706 1438 11942
rect 1202 8736 1438 8894
rect 1202 8672 1232 8736
rect 1232 8672 1248 8736
rect 1248 8672 1312 8736
rect 1312 8672 1328 8736
rect 1328 8672 1392 8736
rect 1392 8672 1408 8736
rect 1408 8672 1438 8736
rect 1202 8658 1438 8672
rect 3652 13686 3888 13922
rect 2102 9558 2338 9794
rect 2102 6458 2338 6694
rect 2752 12366 2988 12602
rect 2752 10368 2988 10444
rect 2752 10304 2782 10368
rect 2782 10304 2798 10368
rect 2798 10304 2862 10368
rect 2862 10304 2878 10368
rect 2878 10304 2942 10368
rect 2942 10304 2958 10368
rect 2958 10304 2988 10368
rect 2752 10208 2988 10304
rect 2752 7108 2988 7344
rect 5202 13026 5438 13262
rect 3652 8008 3888 8244
rect 4302 11706 4538 11942
rect 4302 8736 4538 8894
rect 4302 8672 4332 8736
rect 4332 8672 4348 8736
rect 4348 8672 4412 8736
rect 4412 8672 4428 8736
rect 4428 8672 4492 8736
rect 4492 8672 4508 8736
rect 4508 8672 4538 8736
rect 4302 8658 4538 8672
rect 4302 5558 4538 5794
rect 1878 4908 2114 5144
rect 2678 4908 2914 5144
rect 1478 3358 1714 3594
rect 2278 3358 2514 3594
rect 3078 3358 3314 3594
rect 402 2458 638 2694
rect 4302 2458 4538 2694
rect 402 1658 638 1894
rect 1202 1658 1438 1894
rect -258 998 -22 1234
rect -918 338 -682 574
rect 2752 998 2988 1234
rect 2102 338 2338 574
rect -1578 -322 -1342 -86
rect 4302 1658 4538 1894
rect 6752 13686 6988 13922
rect 5202 9558 5438 9794
rect 5202 6458 5438 6694
rect 5202 3358 5438 3594
rect 3652 -322 3888 -86
rect 5852 12366 6088 12602
rect 5852 10368 6088 10444
rect 5852 10304 5882 10368
rect 5882 10304 5898 10368
rect 5898 10304 5962 10368
rect 5962 10304 5978 10368
rect 5978 10304 6042 10368
rect 6042 10304 6058 10368
rect 6058 10304 6088 10368
rect 5852 10208 6088 10304
rect 5852 7108 6088 7344
rect 5852 4008 6088 4244
rect 5852 998 6088 1234
rect 12106 13686 12342 13922
rect 8302 13026 8538 13262
rect 6752 8008 6988 8244
rect 6752 4908 6988 5144
rect 5202 338 5438 574
rect 7402 11706 7638 11942
rect 7402 8736 7638 8894
rect 7402 8672 7432 8736
rect 7432 8672 7448 8736
rect 7448 8672 7512 8736
rect 7512 8672 7528 8736
rect 7528 8672 7592 8736
rect 7592 8672 7608 8736
rect 7608 8672 7638 8736
rect 7402 8658 7638 8672
rect 7402 5558 7638 5794
rect 7402 2458 7638 2694
rect 7402 1658 7638 1894
rect 11446 13026 11682 13262
rect 8302 9558 8538 9794
rect 8302 6458 8538 6694
rect 8302 3358 8538 3594
rect 6752 -322 6988 -86
rect 8952 12366 9188 12602
rect 10786 12366 11022 12602
rect 8952 10368 9188 10444
rect 8952 10304 8982 10368
rect 8982 10304 8998 10368
rect 8998 10304 9062 10368
rect 9062 10304 9078 10368
rect 9078 10304 9142 10368
rect 9142 10304 9158 10368
rect 9158 10304 9188 10368
rect 8952 10208 9188 10304
rect 8952 7108 9188 7344
rect 8952 4008 9188 4244
rect 10126 11706 10362 11942
rect 10126 8658 10362 8894
rect 10126 5558 10362 5794
rect 10126 2458 10362 2694
rect 10126 1658 10362 1894
rect 10786 10208 11022 10444
rect 10786 7108 11022 7344
rect 10786 4008 11022 4244
rect 8952 998 9188 1234
rect 10786 998 11022 1234
rect 11446 9558 11682 9794
rect 11446 6458 11682 6694
rect 11446 3358 11682 3594
rect 8302 338 8538 574
rect 11446 338 11682 574
rect 12106 8008 12342 8244
rect 12106 4908 12342 5144
rect 12106 -322 12342 -86
<< metal5 >>
rect -1620 13922 12384 13964
rect -1620 13686 -1578 13922
rect -1342 13686 3652 13922
rect 3888 13686 6752 13922
rect 6988 13686 12106 13922
rect 12342 13686 12384 13922
rect -1620 13644 12384 13686
rect -960 13262 11724 13304
rect -960 13026 -918 13262
rect -682 13026 2102 13262
rect 2338 13026 5202 13262
rect 5438 13026 8302 13262
rect 8538 13026 11446 13262
rect 11682 13026 11724 13262
rect -960 12984 11724 13026
rect -300 12602 11064 12644
rect -300 12366 -258 12602
rect -22 12366 2752 12602
rect 2988 12366 5852 12602
rect 6088 12366 8952 12602
rect 9188 12366 10786 12602
rect 11022 12366 11064 12602
rect -300 12324 11064 12366
rect 360 11942 10404 11984
rect 360 11706 402 11942
rect 638 11706 1202 11942
rect 1438 11706 4302 11942
rect 4538 11706 7402 11942
rect 7638 11706 10126 11942
rect 10362 11706 10404 11942
rect 360 11664 10404 11706
rect -300 10444 11064 10486
rect -300 10208 -258 10444
rect -22 10208 2752 10444
rect 2988 10208 5852 10444
rect 6088 10208 8952 10444
rect 9188 10208 10786 10444
rect 11022 10208 11064 10444
rect -300 10166 11064 10208
rect -1620 9794 12384 9836
rect -1620 9558 -918 9794
rect -682 9558 2102 9794
rect 2338 9558 5202 9794
rect 5438 9558 8302 9794
rect 8538 9558 11446 9794
rect 11682 9558 12384 9794
rect -1620 9516 12384 9558
rect -300 8894 11064 8936
rect -300 8658 402 8894
rect 638 8658 1202 8894
rect 1438 8658 4302 8894
rect 4538 8658 7402 8894
rect 7638 8658 10126 8894
rect 10362 8658 11064 8894
rect -300 8616 11064 8658
rect -1620 8244 12384 8286
rect -1620 8008 -1578 8244
rect -1342 8008 3652 8244
rect 3888 8008 6752 8244
rect 6988 8008 12106 8244
rect 12342 8008 12384 8244
rect -1620 7966 12384 8008
rect -300 7344 11064 7386
rect -300 7108 -258 7344
rect -22 7108 2752 7344
rect 2988 7108 5852 7344
rect 6088 7108 8952 7344
rect 9188 7108 10786 7344
rect 11022 7108 11064 7344
rect -300 7066 11064 7108
rect -1620 6694 12384 6736
rect -1620 6458 -918 6694
rect -682 6458 2102 6694
rect 2338 6458 5202 6694
rect 5438 6458 8302 6694
rect 8538 6458 11446 6694
rect 11682 6458 12384 6694
rect -1620 6416 12384 6458
rect -300 5794 11064 5836
rect -300 5558 402 5794
rect 638 5558 4302 5794
rect 4538 5558 7402 5794
rect 7638 5558 10126 5794
rect 10362 5558 11064 5794
rect -300 5516 11064 5558
rect -1620 5144 12384 5186
rect -1620 4908 -1578 5144
rect -1342 4908 1878 5144
rect 2114 4908 2678 5144
rect 2914 4908 6752 5144
rect 6988 4908 12106 5144
rect 12342 4908 12384 5144
rect -1620 4866 12384 4908
rect -300 4244 11064 4286
rect -300 4008 -258 4244
rect -22 4008 5852 4244
rect 6088 4008 8952 4244
rect 9188 4008 10786 4244
rect 11022 4008 11064 4244
rect -300 3966 11064 4008
rect -1620 3594 12384 3636
rect -1620 3358 -918 3594
rect -682 3358 1478 3594
rect 1714 3358 2278 3594
rect 2514 3358 3078 3594
rect 3314 3358 5202 3594
rect 5438 3358 8302 3594
rect 8538 3358 11446 3594
rect 11682 3358 12384 3594
rect -1620 3316 12384 3358
rect -300 2694 11064 2736
rect -300 2458 402 2694
rect 638 2458 4302 2694
rect 4538 2458 7402 2694
rect 7638 2458 10126 2694
rect 10362 2458 11064 2694
rect -300 2416 11064 2458
rect 360 1894 10404 1936
rect 360 1658 402 1894
rect 638 1658 1202 1894
rect 1438 1658 4302 1894
rect 4538 1658 7402 1894
rect 7638 1658 10126 1894
rect 10362 1658 10404 1894
rect 360 1616 10404 1658
rect -300 1234 11064 1276
rect -300 998 -258 1234
rect -22 998 2752 1234
rect 2988 998 5852 1234
rect 6088 998 8952 1234
rect 9188 998 10786 1234
rect 11022 998 11064 1234
rect -300 956 11064 998
rect -960 574 11724 616
rect -960 338 -918 574
rect -682 338 2102 574
rect 2338 338 5202 574
rect 5438 338 8302 574
rect 8538 338 11446 574
rect 11682 338 11724 574
rect -960 296 11724 338
rect -1620 -86 12384 -44
rect -1620 -322 -1578 -86
rect -1342 -322 3652 -86
rect 3888 -322 6752 -86
rect 6988 -322 12106 -86
rect 12342 -322 12384 -86
rect -1620 -364 12384 -322
use gpio_logic_high  gpio_logic_high
timestamp 1633363087
transform 1 0 1196 0 1 2480
box -208 -248 2622 2920
use sky130_fd_sc_hd__decap_4  FILLER_1_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 4324 0 1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_4  FILLER_0_37
timestamp 1631720020
transform 1 0 4324 0 -1 2720
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_32 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 4048 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_0
timestamp 1631720020
transform 1 0 4048 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_1_41 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 4692 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_0_41
timestamp 1631720020
transform 1 0 4692 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _108_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 4784 0 1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _096_
timestamp 1631720020
transform 1 0 4784 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_4  FILLER_2_37
timestamp 1631720020
transform 1 0 4324 0 -1 3808
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_2
timestamp 1631720020
transform 1 0 4048 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _103_
timestamp 1631720020
transform 1 0 4692 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_4
timestamp 1631720020
transform 1 0 4048 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _104_
timestamp 1631720020
transform 1 0 4784 0 1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_3_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 4324 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _044_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 4508 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_6
timestamp 1631720020
transform 1 0 4048 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_4_37
timestamp 1631720020
transform 1 0 4324 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _105_
timestamp 1631720020
transform 1 0 4416 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _045_
timestamp 1631720020
transform 1 0 6348 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_8
timestamp 1631720020
transform 1 0 4048 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _107_
timestamp 1631720020
transform 1 0 4600 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_5_61
timestamp 1631720020
transform 1 0 6532 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _043_
timestamp 1631720020
transform 1 0 4324 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_58 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 6716 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_34
timestamp 1631720020
transform 1 0 6716 0 1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_1_73 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 7636 0 1 2720
box -38 -48 774 592
use sky130_fd_sc_hd__conb_1  const_source $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 7360 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _057_
timestamp 1631720020
transform 1 0 7084 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__inv_2  _072_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 6808 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_59
timestamp 1631720020
transform 1 0 9384 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_0_85 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8740 0 -1 2720
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_91
timestamp 1631720020
transform 1 0 9292 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_1_81
timestamp 1631720020
transform 1 0 8372 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _081_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8740 0 1 2720
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8556 0 1 2720
box -38 -48 222 592
use sky130_fd_sc_hd__dfrtp_2  _094_
timestamp 1631720020
transform 1 0 6808 0 -1 2720
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_35
timestamp 1631720020
transform 1 0 9292 0 -1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _095_
timestamp 1631720020
transform 1 0 6624 0 -1 3808
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_2_89
timestamp 1631720020
transform 1 0 9108 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_2_92
timestamp 1631720020
transform 1 0 9384 0 -1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _056_
timestamp 1631720020
transform 1 0 8832 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _055_
timestamp 1631720020
transform 1 0 8556 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_36
timestamp 1631720020
transform 1 0 6716 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_3_76
timestamp 1631720020
transform 1 0 7912 0 1 3808
box -38 -48 590 592
use sky130_fd_sc_hd__decap_12  FILLER_3_64 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 6808 0 1 3808
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_3_82
timestamp 1631720020
transform 1 0 8464 0 1 3808
box -38 -48 130 592
use sky130_fd_sc_hd__mux2_1  _080_
timestamp 1631720020
transform 1 0 8740 0 1 3808
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_0
timestamp 1631720020
transform 1 0 8556 0 1 3808
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_37
timestamp 1631720020
transform 1 0 9292 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_4_83
timestamp 1631720020
transform 1 0 8556 0 -1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _091_
timestamp 1631720020
transform 1 0 6624 0 -1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_2  FILLER_4_92
timestamp 1631720020
transform 1 0 9384 0 -1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__nand2b_2  _073_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8648 0 -1 4896
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_38
timestamp 1631720020
transform 1 0 6716 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_5_67
timestamp 1631720020
transform 1 0 7084 0 1 4896
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_5_92
timestamp 1631720020
transform 1 0 9384 0 1 4896
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _042_
timestamp 1631720020
transform 1 0 6808 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _059_
timestamp 1631720020
transform 1 0 9108 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _092_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 7176 0 1 4896
box -38 -48 1970 592
use sky130_fd_sc_hd__decap_3  PHY_33
timestamp 1631720020
transform -1 0 9844 0 -1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_1
timestamp 1631720020
transform -1 0 9844 0 1 2720
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_3
timestamp 1631720020
transform -1 0 9844 0 -1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_5
timestamp 1631720020
transform -1 0 9844 0 1 3808
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_7
timestamp 1631720020
transform -1 0 9844 0 -1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_9
timestamp 1631720020
transform -1 0 9844 0 1 4896
box -38 -48 314 592
use sky130_fd_sc_hd__fill_1  FILLER_0_93
timestamp 1631720020
transform 1 0 9476 0 -1 2720
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_40
timestamp 1631720020
transform 1 0 3588 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_7_23
timestamp 1631720020
transform 1 0 3036 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_12
timestamp 1631720020
transform 1 0 920 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_7_15
timestamp 1631720020
transform 1 0 2300 0 1 5984
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_7_3
timestamp 1631720020
transform 1 0 1196 0 1 5984
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_7_30
timestamp 1631720020
transform 1 0 3680 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_0_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 3312 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_8_15
timestamp 1631720020
transform 1 0 2300 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_14
timestamp 1631720020
transform 1 0 920 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_8_3
timestamp 1631720020
transform 1 0 1196 0 -1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__einvp_8  gpio_in_buf $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 2576 0 -1 7072
box -38 -48 1694 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_44
timestamp 1631720020
transform 1 0 3588 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_16
timestamp 1631720020
transform 1 0 920 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_9_15
timestamp 1631720020
transform 1 0 2300 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_9_3
timestamp 1631720020
transform 1 0 1196 0 1 7072
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_9_30
timestamp 1631720020
transform 1 0 3680 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_9_27
timestamp 1631720020
transform 1 0 3404 0 1 7072
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_18
timestamp 1631720020
transform 1 0 920 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_8  FILLER_10_27
timestamp 1631720020
transform 1 0 3404 0 -1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_10_15
timestamp 1631720020
transform 1 0 2300 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_10_3
timestamp 1631720020
transform 1 0 1196 0 -1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_11_30
timestamp 1631720020
transform 1 0 3680 0 1 8160
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_47
timestamp 1631720020
transform 1 0 3588 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  PHY_20
timestamp 1631720020
transform 1 0 920 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_11_3
timestamp 1631720020
transform 1 0 1196 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_11_15
timestamp 1631720020
transform 1 0 2300 0 1 8160
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_11_27
timestamp 1631720020
transform 1 0 3404 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_10
timestamp 1631720020
transform 1 0 4048 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _076_
timestamp 1631720020
transform 1 0 3772 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _048_
timestamp 1631720020
transform 1 0 4048 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_41
timestamp 1631720020
transform 1 0 6256 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_7_59
timestamp 1631720020
transform 1 0 6348 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _047_
timestamp 1631720020
transform 1 0 6532 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _041_
timestamp 1631720020
transform 1 0 6256 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _106_
timestamp 1631720020
transform 1 0 4324 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _102_
timestamp 1631720020
transform 1 0 4324 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _089_
timestamp 1631720020
transform 1 0 6440 0 1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_43
timestamp 1631720020
transform 1 0 6164 0 -1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _109_
timestamp 1631720020
transform 1 0 4232 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _049_
timestamp 1631720020
transform 1 0 6532 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _046_
timestamp 1631720020
transform 1 0 6256 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfrtp_2  _101_
timestamp 1631720020
transform 1 0 4140 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _088_
timestamp 1631720020
transform 1 0 6072 0 1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _050_
timestamp 1631720020
transform 1 0 3864 0 1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_46
timestamp 1631720020
transform 1 0 6164 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_10_35
timestamp 1631720020
transform 1 0 4140 0 -1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _099_
timestamp 1631720020
transform 1 0 4232 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _085_
timestamp 1631720020
transform 1 0 6256 0 -1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__fill_1  FILLER_11_34
timestamp 1631720020
transform 1 0 4048 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _100_
timestamp 1631720020
transform 1 0 4140 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__dfrtp_2  _086_
timestamp 1631720020
transform 1 0 6072 0 1 8160
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _061_
timestamp 1631720020
transform 1 0 6808 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _060_
timestamp 1631720020
transform 1 0 7084 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_39
timestamp 1631720020
transform 1 0 9292 0 -1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_42
timestamp 1631720020
transform 1 0 8924 0 1 5984
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_6_92
timestamp 1631720020
transform 1 0 9384 0 -1 5984
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _062_
timestamp 1631720020
transform 1 0 9016 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _058_
timestamp 1631720020
transform 1 0 8648 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _052_
timestamp 1631720020
transform 1 0 8372 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _063_
timestamp 1631720020
transform 1 0 9292 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _093_
timestamp 1631720020
transform 1 0 7360 0 -1 5984
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _051_
timestamp 1631720020
transform 1 0 6808 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _090_
timestamp 1631720020
transform 1 0 7084 0 -1 7072
box -38 -48 1970 592
use sky130_fd_sc_hd__and2_2  _071_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 9016 0 -1 7072
box -38 -48 590 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_45
timestamp 1631720020
transform 1 0 8832 0 1 7072
box -38 -48 130 592
use sky130_fd_sc_hd__nand2b_2  _070_
timestamp 1631720020
transform 1 0 8924 0 1 7072
box -38 -48 682 592
use sky130_fd_sc_hd__ebufn_2  _083_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8004 0 1 7072
box -38 -48 866 592
use sky130_fd_sc_hd__fill_2  FILLER_10_79
timestamp 1631720020
transform 1 0 8188 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_10_92
timestamp 1631720020
transform 1 0 9384 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__mux2_1  _082_
timestamp 1631720020
transform -1 0 9384 0 -1 8160
box -38 -48 866 592
use sky130_fd_sc_hd__diode_2  ANTENNA_3
timestamp 1631720020
transform -1 0 8556 0 -1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_48
timestamp 1631720020
transform 1 0 8832 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_11_77
timestamp 1631720020
transform 1 0 8004 0 1 8160
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_11_92
timestamp 1631720020
transform 1 0 9384 0 1 8160
box -38 -48 222 592
use sky130_fd_sc_hd__or2_2  _039_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8924 0 1 8160
box -38 -48 498 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8096 0 1 8160
box -38 -48 774 592
use sky130_fd_sc_hd__buf_1  _XX1_
timestamp 1631720020
transform 1 0 9568 0 -1 7072
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_11
timestamp 1631720020
transform -1 0 9844 0 -1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_13
timestamp 1631720020
transform -1 0 9844 0 1 5984
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_19
timestamp 1631720020
transform -1 0 9844 0 -1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_21
timestamp 1631720020
transform -1 0 9844 0 1 8160
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_22
timestamp 1631720020
transform 1 0 920 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_12_3
timestamp 1631720020
transform 1 0 1196 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_15
timestamp 1631720020
transform 1 0 2300 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_12_27
timestamp 1631720020
transform 1 0 3404 0 -1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  PHY_24
timestamp 1631720020
transform 1 0 920 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_26
timestamp 1631720020
transform 1 0 920 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_13_3
timestamp 1631720020
transform 1 0 1196 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_3
timestamp 1631720020
transform 1 0 1196 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_13_15
timestamp 1631720020
transform 1 0 2300 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_15
timestamp 1631720020
transform 1 0 2300 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_50
timestamp 1631720020
transform 1 0 3588 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_13_30
timestamp 1631720020
transform 1 0 3680 0 1 9248
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_14_27
timestamp 1631720020
transform 1 0 3404 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_13_27
timestamp 1631720020
transform 1 0 3404 0 1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_28
timestamp 1631720020
transform 1 0 920 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_15_3
timestamp 1631720020
transform 1 0 1196 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_15_15
timestamp 1631720020
transform 1 0 2300 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_53
timestamp 1631720020
transform 1 0 3588 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_15_30
timestamp 1631720020
transform 1 0 3680 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_27
timestamp 1631720020
transform 1 0 3404 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__decap_3  PHY_30
timestamp 1631720020
transform 1 0 920 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_16_3
timestamp 1631720020
transform 1 0 1196 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_12  FILLER_16_15
timestamp 1631720020
transform 1 0 2300 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_55
timestamp 1631720020
transform 1 0 3588 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_12  FILLER_16_30
timestamp 1631720020
transform 1 0 3680 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_16_27
timestamp 1631720020
transform 1 0 3404 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_49
timestamp 1631720020
transform 1 0 6164 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__decap_6  FILLER_12_39
timestamp 1631720020
transform 1 0 4508 0 -1 9248
box -38 -48 590 592
use sky130_fd_sc_hd__dfrtp_2  _087_
timestamp 1631720020
transform 1 0 6256 0 -1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _068_
timestamp 1631720020
transform 1 0 5336 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _067_
timestamp 1631720020
transform 1 0 5612 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _064_
timestamp 1631720020
transform 1 0 5888 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  clkbuf_1_1_0_serial_clock
timestamp 1631720020
transform 1 0 5060 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_52
timestamp 1631720020
transform 1 0 6164 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_13_42
timestamp 1631720020
transform 1 0 4784 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  FILLER_14_51
timestamp 1631720020
transform 1 0 5612 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_12  FILLER_14_39
timestamp 1631720020
transform 1 0 4508 0 -1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_14_58
timestamp 1631720020
transform 1 0 6256 0 -1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__buf_1  _053_
timestamp 1631720020
transform 1 0 6348 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  _069_
timestamp 1631720020
transform 1 0 5888 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_16  clkbuf_0_serial_clock $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 5060 0 1 9248
box -38 -48 1878 592
use sky130_fd_sc_hd__decap_4  FILLER_15_54
timestamp 1631720020
transform 1 0 5888 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__decap_12  FILLER_15_42
timestamp 1631720020
transform 1 0 4784 0 1 10336
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_15_61
timestamp 1631720020
transform 1 0 6532 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _066_
timestamp 1631720020
transform 1 0 6256 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_4  FILLER_16_54
timestamp 1631720020
transform 1 0 5888 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_56
timestamp 1631720020
transform 1 0 6256 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_16_59
timestamp 1631720020
transform 1 0 6348 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__decap_12  FILLER_16_42
timestamp 1631720020
transform 1 0 4784 0 -1 11424
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_12_82
timestamp 1631720020
transform 1 0 8464 0 -1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_12_92
timestamp 1631720020
transform 1 0 9384 0 -1 9248
box -38 -48 222 592
use sky130_fd_sc_hd__buf_1  _040_
timestamp 1631720020
transform 1 0 8188 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__mux2_1  _079_
timestamp 1631720020
transform 1 0 8556 0 -1 9248
box -38 -48 866 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_51
timestamp 1631720020
transform 1 0 8832 0 1 9248
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _098_
timestamp 1631720020
transform 1 0 6900 0 1 9248
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _054_
timestamp 1631720020
transform 1 0 9292 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__dfstp_2  _084_
timestamp 1631720020
transform 1 0 7360 0 -1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold3
timestamp 1631720020
transform 1 0 6624 0 -1 10336
box -38 -48 774 592
use sky130_fd_sc_hd__nor2b_2  _075_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8924 0 1 9248
box -38 -48 682 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_54
timestamp 1631720020
transform 1 0 8832 0 1 10336
box -38 -48 130 592
use sky130_fd_sc_hd__dfrtp_2  _097_
timestamp 1631720020
transform -1 0 8832 0 1 10336
box -38 -48 1970 592
use sky130_fd_sc_hd__buf_1  _065_
timestamp 1631720020
transform 1 0 9292 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__diode_2  ANTENNA_2
timestamp 1631720020
transform -1 0 6900 0 1 10336
box -38 -48 222 592
use sky130_fd_sc_hd__buf_2  _077_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1631720020
transform 1 0 8924 0 1 10336
box -38 -48 406 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  PHY_57
timestamp 1631720020
transform 1 0 8924 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_1  FILLER_16_67
timestamp 1631720020
transform 1 0 7084 0 -1 11424
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_16_92
timestamp 1631720020
transform 1 0 9384 0 -1 11424
box -38 -48 222 592
use sky130_fd_sc_hd__inv_2  _074_
timestamp 1631720020
transform 1 0 7176 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold2
timestamp 1631720020
transform 1 0 8188 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__dlygate4sd3_1  hold4
timestamp 1631720020
transform 1 0 7452 0 -1 11424
box -38 -48 774 592
use sky130_fd_sc_hd__buf_2  _078_
timestamp 1631720020
transform 1 0 9016 0 -1 11424
box -38 -48 406 592
use sky130_fd_sc_hd__decap_3  PHY_23
timestamp 1631720020
transform -1 0 9844 0 -1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_25
timestamp 1631720020
transform -1 0 9844 0 1 9248
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_29
timestamp 1631720020
transform -1 0 9844 0 1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_27
timestamp 1631720020
transform -1 0 9844 0 -1 10336
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_31
timestamp 1631720020
transform -1 0 9844 0 -1 11424
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  _XX2_
timestamp 1631720020
transform 1 0 9568 0 1 7072
box -38 -48 406 592
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 0 nsew signal tristate
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 1 nsew signal input
rlabel metal3 s 14000 2048 34000 2168 6 mgmt_gpio_out
port 2 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 3 nsew signal tristate
rlabel metal3 s 14000 2592 34000 2712 6 pad_gpio_ana_en
port 4 nsew signal tristate
rlabel metal3 s 14000 3136 34000 3256 6 pad_gpio_ana_pol
port 5 nsew signal tristate
rlabel metal3 s 14000 3544 34000 3664 6 pad_gpio_ana_sel
port 6 nsew signal tristate
rlabel metal3 s 14000 4088 34000 4208 6 pad_gpio_dm[0]
port 7 nsew signal tristate
rlabel metal3 s 14000 4632 34000 4752 6 pad_gpio_dm[1]
port 8 nsew signal tristate
rlabel metal3 s 14000 5040 34000 5160 6 pad_gpio_dm[2]
port 9 nsew signal tristate
rlabel metal3 s 14000 5584 34000 5704 6 pad_gpio_holdover
port 10 nsew signal tristate
rlabel metal3 s 14000 6128 34000 6248 6 pad_gpio_ib_mode_sel
port 11 nsew signal tristate
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_in
port 12 nsew signal input
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_inenb
port 13 nsew signal tristate
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_out
port 14 nsew signal tristate
rlabel metal3 s 14000 8032 34000 8152 6 pad_gpio_outenb
port 15 nsew signal tristate
rlabel metal3 s 14000 8576 34000 8696 6 pad_gpio_slow_sel
port 16 nsew signal tristate
rlabel metal3 s 14000 9120 34000 9240 6 pad_gpio_vtrip_sel
port 17 nsew signal tristate
rlabel metal3 s 14000 9528 34000 9648 6 resetn
port 18 nsew signal input
rlabel metal3 s 14000 10072 34000 10192 6 resetn_out
port 19 nsew signal tristate
rlabel metal3 s 14000 10616 34000 10736 6 serial_clock
port 20 nsew signal input
rlabel metal3 s 14000 11024 34000 11144 6 serial_clock_out
port 21 nsew signal tristate
rlabel metal3 s 14000 11568 34000 11688 6 serial_data_in
port 22 nsew signal input
rlabel metal3 s 14000 12112 34000 12232 6 serial_data_out
port 23 nsew signal tristate
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 24 nsew signal tristate
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 25 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 26 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 27 nsew signal tristate
rlabel metal4 s 7360 956 7680 12644 6 vccd
port 28 nsew power bidirectional
rlabel metal4 s 4260 956 4580 12644 6 vccd
port 29 nsew power bidirectional
rlabel metal4 s 1160 5632 1480 12644 6 vccd
port 30 nsew power bidirectional
rlabel metal4 s 10084 1616 10404 11984 6 vccd
port 31 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 32 nsew power bidirectional
rlabel metal4 s 1160 956 1480 2128 6 vccd
port 33 nsew power bidirectional
rlabel metal5 s 360 11664 10404 11984 6 vccd
port 34 nsew power bidirectional
rlabel metal5 s -300 8616 11064 8936 6 vccd
port 35 nsew power bidirectional
rlabel metal5 s -300 5516 11064 5836 6 vccd
port 36 nsew power bidirectional
rlabel metal5 s -300 2416 11064 2736 6 vccd
port 37 nsew power bidirectional
rlabel metal5 s 360 1616 10404 1936 6 vccd
port 38 nsew power bidirectional
rlabel metal4 s 10744 956 11064 12644 6 vssd
port 39 nsew ground bidirectional
rlabel metal4 s 8910 956 9230 12644 6 vssd
port 40 nsew ground bidirectional
rlabel metal4 s 5810 956 6130 12644 6 vssd
port 41 nsew ground bidirectional
rlabel metal4 s 2710 5632 3030 12644 6 vssd
port 42 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 43 nsew ground bidirectional
rlabel metal4 s 2710 956 3030 2128 6 vssd
port 44 nsew ground bidirectional
rlabel metal5 s -300 12324 11064 12644 6 vssd
port 45 nsew ground bidirectional
rlabel metal5 s -300 10166 11064 10486 6 vssd
port 46 nsew ground bidirectional
rlabel metal5 s -300 7066 11064 7386 6 vssd
port 47 nsew ground bidirectional
rlabel metal5 s -300 3966 11064 4286 6 vssd
port 48 nsew ground bidirectional
rlabel metal5 s -300 956 11064 1276 6 vssd
port 49 nsew ground bidirectional
rlabel metal4 s 8260 -364 8580 13964 6 vccd1
port 50 nsew power bidirectional
rlabel metal4 s 5160 -364 5480 13964 6 vccd1
port 51 nsew power bidirectional
rlabel metal4 s 2060 5680 2380 13964 6 vccd1
port 52 nsew power bidirectional
rlabel metal4 s 11404 296 11724 13304 6 vccd1
port 53 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 54 nsew power bidirectional
rlabel metal4 s 2060 -364 2380 2080 6 vccd1
port 55 nsew power bidirectional
rlabel metal5 s -960 12984 11724 13304 6 vccd1
port 56 nsew power bidirectional
rlabel metal5 s -1620 9516 12384 9836 6 vccd1
port 57 nsew power bidirectional
rlabel metal5 s -1620 6416 12384 6736 6 vccd1
port 58 nsew power bidirectional
rlabel metal5 s -1620 3316 12384 3636 6 vccd1
port 59 nsew power bidirectional
rlabel metal5 s -960 296 11724 616 6 vccd1
port 60 nsew power bidirectional
rlabel metal4 s 12064 -364 12384 13964 6 vssd1
port 61 nsew ground bidirectional
rlabel metal4 s 6710 -364 7030 13964 6 vssd1
port 62 nsew ground bidirectional
rlabel metal4 s 3610 5680 3930 13964 6 vssd1
port 63 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 64 nsew ground bidirectional
rlabel metal4 s 3610 -364 3930 2080 6 vssd1
port 65 nsew ground bidirectional
rlabel metal5 s -1620 13644 12384 13964 6 vssd1
port 66 nsew ground bidirectional
rlabel metal5 s -1620 7966 12384 8286 6 vssd1
port 67 nsew ground bidirectional
rlabel metal5 s -1620 4866 12384 5186 6 vssd1
port 68 nsew ground bidirectional
rlabel metal5 s -1620 -364 12384 -44 8 vssd1
port 69 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 34000 14000
<< end >>
