I* SPICE NETLIST
***************************************


***************************************

***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808692 2 3
**
R0 3 2 sky130_fd_pr__res_generic_po L=900 W=0.33 m=1
.ENDS


***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808687 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=1.96 PD=7.28 PS=14.56 NRD=0 NRS=0 m=1 sa=90000.2 sb=90004.3 a=1.26 p=14.36
XM1 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90000.7 sb=90003.9 a=1.26 p=14.36
XM2 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90001.1 sb=90003.4 a=1.26 p=14.36
XM3 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90001.6 sb=90002.9 a=1.26 p=14.36
XM4 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90002 sb=90002.5 a=1.26 p=14.36
XM5 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90002.5 sb=90002 a=1.26 p=14.36
XM6 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90002.9 sb=90001.6 a=1.26 p=14.36
XM7 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90003.4 sb=90001.1 a=1.26 p=14.36
XM8 4 3 2 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=90003.9 sb=90000.7 a=1.26 p=14.36
XM9 2 3 4 2 sky130_fd_pr__pfet_01v8 L=0.18 W=7 AD=1.96 AS=0.98 PD=14.56 PS=7.28 NRD=0 NRS=0 m=1 sa=90004.3 sb=90000.2 a=1.26 p=14.36
.ENDS
***************************************


***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808691 2 3
**
R0 3 2 sky130_fd_pr__res_generic_po L=200 W=0.33 m=1
.ENDS
***************************************


***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808704 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS

***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808695 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
.ENDS



***************************************
.SUBCKT sky130_fd_io__gnd2gnd_sub_dnwl 1 2
**
X0 1 2 sky130_fd_pr__model__parasitic__diode_ps2nw a=283.052 p=67.56 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gnd2gnd_120x2_lv_isosub VSUB VSSI VSS_N
**
XD0 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD1 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD2 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD3 VSS_N VSSI sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD4 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD5 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD6 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
XD7 VSSI VSS_N sky130_fd_pr__diode_pd2nw_05v5 AREA=22.5 m=1
X8 VSUB VSSI sky130_fd_io__gnd2gnd_sub_dnwl
X9 VSUB VSS_N sky130_fd_io__gnd2gnd_sub_dnwl
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808701 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808703 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808705 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=2.1 p=14.6 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808693 2
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
X1 2 2 sky130_fd_pr__diode_pw2nd_05v5 a=1.5 p=10.6 m=1
.ENDS
***************************************
**************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808688 3 4
**
*.SEEDPROM
R0 3 4 sky130_fd_pr__res_generic_po L=720 W=0.33 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808690 2 3
**
R0 3 2 sky130_fd_pr__res_generic_po L=300 W=0.33 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_power_lvc_wpad VSSD SRC_BDY_LVC2 SRC_BDY_LVC1 DRN_LVC1 VDDIO DRN_LVC2 BDY2_B2B P_CORE P_PAD
**
*.CALIBRE ISOLATED NETS: OGC_LVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
XM0 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM1 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM2 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM3 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM4 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90001.1 sb=90019.9 a=0.9 p=10.36
XM5 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM6 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM7 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM8 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM9 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM10 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90002.3 sb=90019.9 a=0.9 p=10.36
XM11 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM12 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=4 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=20 p=18
XM13 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM14 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM15 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM16 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM17 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90003.9 sb=90019.9 a=0.9 p=10.36
XM18 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM19 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM20 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM21 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM22 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM23 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM24 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM25 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM26 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM27 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90005.1 sb=90019.9 a=0.9 p=10.36
XM28 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM29 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM30 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM31 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM32 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM33 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM34 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM35 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM36 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM37 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90006.6 sb=90019.9 a=0.9 p=10.36
XM38 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM39 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM40 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM41 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM42 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM43 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM44 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90007.8 sb=90019.9 a=0.9 p=10.36
XM45 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM46 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM47 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM48 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM49 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM50 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM51 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM52 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM53 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM54 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90009.4 sb=90019.9 a=0.9 p=10.36
XM55 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM56 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM57 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM58 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM59 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM60 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM61 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM62 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM63 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM64 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90010.6 sb=90019.9 a=0.9 p=10.36
XM65 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM66 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM67 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM68 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM69 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM70 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM71 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM72 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=40 p=26
XM73 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM74 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM75 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM76 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM77 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90012.2 sb=90019.9 a=0.9 p=10.36
XM78 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM79 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM80 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90001.7 sb=90019.9 a=0.9 p=10.36
XM81 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM82 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM83 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM84 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM85 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM86 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM87 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM88 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM89 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90013.4 sb=90019.9 a=0.9 p=10.36
XM90 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM91 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM92 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90003.1 sb=90019.9 a=0.9 p=10.36
XM93 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM94 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM95 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM96 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM97 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM98 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM99 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM100 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM101 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90015 sb=90019.9 a=0.9 p=10.36
XM102 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM103 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM104 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM105 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM106 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM107 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM108 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90016.1 sb=90019.9 a=0.9 p=10.36
XM109 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM110 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM111 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90005.9 sb=90019.9 a=0.9 p=10.36
XM112 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM113 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM114 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM115 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM116 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM117 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM118 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM119 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM120 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90017.7 sb=90019.9 a=0.9 p=10.36
XM121 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM122 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM123 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90007.3 sb=90019.9 a=0.9 p=10.36
XM124 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM125 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM126 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM127 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM128 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM129 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM130 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM131 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM132 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90018.9 sb=90019.9 a=0.9 p=10.36
XM133 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM134 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM135 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=40 p=26
XM136 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM137 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM138 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM139 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM140 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM141 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM142 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM143 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM144 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM145 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM146 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM147 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM148 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90010.1 sb=90019.9 a=0.9 p=10.36
XM149 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM150 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM151 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM152 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM153 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM154 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM155 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM156 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM157 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM158 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM159 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM160 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90011.4 sb=90019.9 a=0.9 p=10.36
XM161 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM162 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM163 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM164 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM165 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM166 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM167 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM168 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM169 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM170 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM171 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM172 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM173 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM174 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM175 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM176 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM177 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM178 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM179 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90014.3 sb=90019.9 a=0.9 p=10.36
XM180 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM181 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM182 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM183 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM184 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM185 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM186 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM187 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM188 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM189 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM190 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM191 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90015.6 sb=90019.9 a=0.9 p=10.36
XM192 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM193 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM194 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM195 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM196 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM197 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM198 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM199 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM200 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM201 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM202 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM203 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4.00002e+06 a=40 p=26
XM204 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM205 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM206 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM207 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM208 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM209 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM210 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM211 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM212 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM213 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM214 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM215 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM216 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90018.5 sb=90019.9 a=0.9 p=10.36
XM217 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM218 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM219 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM220 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM221 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM222 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM223 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM224 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM225 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM226 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM227 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM228 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.8 sb=90019.9 a=0.9 p=10.36
XM229 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM230 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM231 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM232 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM233 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM234 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM235 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM236 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM237 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM238 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM239 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM240 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM241 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM242 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM243 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM244 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM245 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM246 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM247 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90019.8 a=0.9 p=10.36
XM248 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM249 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM250 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM251 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM252 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM253 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM254 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM255 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM256 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90018.9 a=0.9 p=10.36
XM257 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM258 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM259 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90018.5 a=0.9 p=10.36
XM260 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM261 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM262 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM263 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM264 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM265 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM266 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM267 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM268 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90017.7 a=0.9 p=10.36
XM269 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM270 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM271 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4.00001e+06 a=40 p=26
XM272 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM273 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM274 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM275 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM276 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM277 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM278 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM279 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM280 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM281 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90016.1 a=0.9 p=10.36
XM282 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM283 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM284 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90015.6 a=0.9 p=10.36
XM285 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM286 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM287 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM288 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM289 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM290 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM291 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM292 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM293 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90015 a=0.9 p=10.36
XM294 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM295 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM296 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90014.3 a=0.9 p=10.36
XM297 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM298 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM299 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM300 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM301 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM302 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM303 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM304 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM305 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90013.4 a=0.9 p=10.36
XM306 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM307 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM308 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM309 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM310 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM311 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM312 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90012.2 a=0.9 p=10.36
XM313 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM314 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM315 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90011.4 a=0.9 p=10.36
XM316 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM317 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM318 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM319 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM320 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM321 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM322 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM323 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM324 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90010.6 a=0.9 p=10.36
XM325 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM326 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM327 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90010.1 a=0.9 p=10.36
XM328 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM329 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM330 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM331 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM332 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM333 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM334 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM335 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM336 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90009.4 a=0.9 p=10.36
XM337 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM338 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM339 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=40 p=26
XM340 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM341 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM342 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM343 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM344 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM345 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM346 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM347 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM348 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM349 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90007.8 a=0.9 p=10.36
XM350 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM351 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM352 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90007.3 a=0.9 p=10.36
XM353 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM354 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM355 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM356 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM357 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM358 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM359 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM360 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM361 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90006.6 a=0.9 p=10.36
XM362 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM363 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM364 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90005.9 a=0.9 p=10.36
XM365 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM366 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM367 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM368 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM369 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM370 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM371 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM372 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM373 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90005.1 a=0.9 p=10.36
XM374 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM375 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM376 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM377 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM378 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM379 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM380 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90003.9 a=0.9 p=10.36
XM381 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM382 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM383 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90003.1 a=0.9 p=10.36
XM384 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM385 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM386 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM387 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM388 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM389 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM390 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM391 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM392 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90002.3 a=0.9 p=10.36
XM393 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM394 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM395 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90001.7 a=0.9 p=10.36
XM396 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM397 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM398 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM399 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM400 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM401 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM402 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM403 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM404 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90001.1 a=0.9 p=10.36
XM405 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM406 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM407 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=40 p=26
XM408 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM409 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM410 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM411 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM412 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
X413 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1
X414 SRC_BDY_LVC2 VDDIO condiode a=1e-06 p=0.004 m=1
X415 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1
X416 VSSD DRN_LVC1 sky130_fd_pr__model__parasitic__diode_ps2nw a=108.41 p=46.58 m=1
X417 VSSD DRN_LVC2 sky130_fd_pr__model__parasitic__diode_ps2nw a=108.41 p=46.58 m=1
X418 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn a=10516.3 p=468.87 m=1
X419 SRC_BDY_LVC2 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=4115.42 p=264.63 m=1
X420 SRC_BDY_LVC1 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=5703.29 p=340.89 m=1
R421 DRN_LVC1 21 sky130_fd_pr__res_generic_po L=1950 W=0.33 m=1
R422 P_CORE P_PAD 0.01 short m=1
X423 27 DRN_LVC2 sky130_fd_pr__res_bent_po__example_55959141808692
X424 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X425 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X426 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X427 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X616 23 26 sky130_fd_pr__res_bent_po__example_55959141808691
X622 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808704
X623 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808695
X630 VSSD BDY2_B2B SRC_BDY_LVC1 sky130_fd_io__gnd2gnd_120x2_lv_isosub
X631 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808701
X632 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X633 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X634 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X635 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X636 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X637 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X638 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X639 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808705
X640 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808693
X642 22 26 sky130_fd_pr__res_bent_po__example_55959141808688
X643 27 22 sky130_fd_pr__res_bent_po__example_55959141808690
.ENDS
***************************************
.SUBCKT sky130_ef_io__vccd_lvc_clamped2_pad VSSD VSSA VSSIO VCCD VDDIO VCCD_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSIO VCCD VDDIO VCCD VSSA VCCD VCCD_PAD sky130_fd_io__top_power_lvc_wpad
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808669 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=470 W=0.33 m=1
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 2 3
**
*.SEEDPROM
XM0 2 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=2e+06 sb=2e+06 a=20 p=18
.ENDS
***************************************
.SUBCKT sky130_fd_io__sio_clamp_pcap_4x5 2 3
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664
.ENDS
***************************************
.SUBCKT sky130_fd_io__esd_rcclamp_nfetcap 2 3
**
*.SEEDPROM
XM0 2 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 sa=4e+06 sb=4e+06 a=40 p=26
.ENDS

***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808677 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 sa=250000 sb=250011 a=3.5 p=15
XM1 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250001 sb=250010 a=3.5 p=15
XM2 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250002 sb=250009 a=3.5 p=15
XM3 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250002 sb=250009 a=3.5 p=15
XM4 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250003 sb=250008 a=3.5 p=15
XM5 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250004 sb=250007 a=3.5 p=15
XM6 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250005 sb=250006 a=3.5 p=15
XM7 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250005 sb=250005 a=3.5 p=15
XM8 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250006 sb=250005 a=3.5 p=15
XM9 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250007 sb=250004 a=3.5 p=15
XM10 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250008 sb=250003 a=3.5 p=15
XM11 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250009 sb=250002 a=3.5 p=15
XM12 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250009 sb=250002 a=3.5 p=15
XM13 2 3 4 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250010 sb=250001 a=3.5 p=15
XM14 4 3 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=250011 sb=250000 a=3.5 p=15
.ENDS
***************************************
.SUBCKT ICV_8 2 3
**
*.SEEDPROM
X0 2 3 sky130_fd_io__esd_rcclamp_nfetcap
X1 2 3 sky130_fd_io__esd_rcclamp_nfetcap
.ENDS
***************************************



***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808668 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=700 W=0.33 m=1
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808665 2 3 4
**
*.SEEDPROM
XM0 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 sa=250000 sb=250020 a=3.5 p=15
XM1 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250001 sb=250020 a=3.5 p=15
XM2 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250002 sb=250020 a=3.5 p=15
XM3 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250002 sb=250020 a=3.5 p=15
XM4 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250003 sb=250020 a=3.5 p=15
XM5 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250004 sb=250020 a=3.5 p=15
XM6 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250005 sb=250020 a=3.5 p=15
XM7 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250005 sb=250020 a=3.5 p=15
XM8 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250006 sb=250020 a=3.5 p=15
XM9 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250007 sb=250020 a=3.5 p=15
XM10 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250008 sb=250020 a=3.5 p=15
XM11 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250009 sb=250020 a=3.5 p=15
XM12 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250009 sb=250020 a=3.5 p=15
XM13 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250010 sb=250020 a=3.5 p=15
XM14 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250011 sb=250020 a=3.5 p=15
XM15 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250012 sb=250020 a=3.5 p=15
XM16 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250012 sb=250020 a=3.5 p=15
XM17 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250013 sb=250020 a=3.5 p=15
XM18 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250014 sb=250020 a=3.5 p=15
XM19 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250015 sb=250020 a=3.5 p=15
XM20 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250016 sb=250020 a=3.5 p=15
XM21 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250016 sb=250020 a=3.5 p=15
XM22 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250017 sb=250020 a=3.5 p=15
XM23 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250018 sb=250020 a=3.5 p=15
XM24 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250019 sb=250020 a=3.5 p=15
XM25 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250019 a=3.5 p=15
XM26 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250018 a=3.5 p=15
XM27 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250017 a=3.5 p=15
XM28 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250016 a=3.5 p=15
XM29 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250016 a=3.5 p=15
XM30 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250015 a=3.5 p=15
XM31 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250014 a=3.5 p=15
XM32 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250013 a=3.5 p=15
XM33 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250012 a=3.5 p=15
XM34 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250012 a=3.5 p=15
XM35 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250011 a=3.5 p=15
XM36 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250010 a=3.5 p=15
XM37 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250009 a=3.5 p=15
XM38 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250009 a=3.5 p=15
XM39 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250008 a=3.5 p=15
XM40 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250007 a=3.5 p=15
XM41 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250006 a=3.5 p=15
XM42 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250005 a=3.5 p=15
XM43 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250005 a=3.5 p=15
XM44 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250004 a=3.5 p=15
XM45 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250003 a=3.5 p=15
XM46 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250002 a=3.5 p=15
XM47 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250002 a=3.5 p=15
XM48 4 3 2 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250001 a=3.5 p=15
XM49 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=250020 sb=250000 a=3.5 p=15
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_55959141808667 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=1550 W=0.33 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_ground_hvc_wpad VSSD SRC_BDY_HVC DRN_HVC VDDIO G_CORE G_PAD
**
*.CALIBRE ISOLATED NETS: OGC_HVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
XM0 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM1 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM2 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM3 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250001 sb=250020 a=5 p=21
XM4 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM5 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM6 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM7 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250003 sb=250020 a=5 p=21
XM8 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM9 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM10 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM11 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250006 sb=250020 a=5 p=21
XM12 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM13 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM14 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM15 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250008 sb=250020 a=5 p=21
XM16 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM17 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM18 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM19 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM20 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM21 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM22 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250010 sb=250020 a=5 p=21
XM23 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM24 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM25 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM26 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM27 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM28 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM29 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250012 sb=250020 a=5 p=21
XM30 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM31 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM32 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM33 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM34 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM35 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM36 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250015 sb=250020 a=5 p=21
XM37 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM38 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM39 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM40 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM41 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM42 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM43 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250017 sb=250020 a=5 p=21
XM44 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM45 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM46 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM47 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM48 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM49 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM50 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250020 a=5 p=21
XM51 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM52 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM53 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM54 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM55 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM56 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM57 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250020 a=5 p=21
XM58 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM59 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM60 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM61 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM62 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM63 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM64 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250020 a=5 p=21
XM65 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM66 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM67 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM68 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM69 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM70 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM71 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250020 a=5 p=21
XM72 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM73 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM74 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM75 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM76 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM77 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM78 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250020 a=5 p=21
XM79 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM80 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM81 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM82 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM83 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM84 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM85 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250020 a=5 p=21
XM86 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM87 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM88 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM89 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM90 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM91 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM92 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250017 a=5 p=21
XM93 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM94 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM95 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM96 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM97 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM98 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM99 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250015 a=5 p=21
XM100 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM101 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM102 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM103 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM104 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM105 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM106 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250012 a=5 p=21
XM107 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM108 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM109 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM110 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM111 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM112 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM113 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250010 a=5 p=21
XM114 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM115 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM116 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM117 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM118 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM119 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM120 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250008 a=5 p=21
XM121 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM122 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM123 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM124 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM125 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM126 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM127 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250006 a=5 p=21
XM128 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM129 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM130 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM131 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM132 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM133 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM134 DRN_HVC 19 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250003 a=5 p=21
XM135 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM136 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM137 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM138 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM139 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM140 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM141 SRC_BDY_HVC 19 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250001 a=5 p=21
X142 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X143 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X144 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X145 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X146 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=126.883 p=0 m=1
X147 VSSD DRN_HVC sky130_fd_pr__model__parasitic__diode_ps2nw a=376.949 p=101.73 m=1
X148 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn a=10358.7 p=619.08 m=1
X149 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=137.463 p=47.72 m=1
X150 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=8184.99 p=443.22 m=1
X151 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=1172.63 p=163 m=1
R152 G_CORE G_PAD 0.01 short m=1
X153 18 20 sky130_fd_pr__res_bent_po__example_55959141808669
X225 SRC_BDY_HVC 18 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664
X226 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X227 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X228 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X229 SRC_BDY_HVC 18 sky130_fd_io__sio_clamp_pcap_4x5
X230 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap
X231 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap
X232 SRC_BDY_HVC 18 sky130_fd_io__esd_rcclamp_nfetcap
X233 SRC_BDY_HVC 18 19 sky130_fd_pr__nfet_01v8__example_55959141808677
X234 SRC_BDY_HVC 18 ICV_8
X235 SRC_BDY_HVC 18 ICV_8
X236 SRC_BDY_HVC 18 ICV_8
X237 SRC_BDY_HVC 18 ICV_8
X238 SRC_BDY_HVC 18 ICV_8
X239 SRC_BDY_HVC 18 ICV_8
X247 DRN_HVC 21 sky130_fd_pr__res_bent_po__example_55959141808668
X248 DRN_HVC 18 19 sky130_fd_pr__pfet_01v8__example_55959141808665
X249 21 20 sky130_fd_pr__res_bent_po__example_55959141808667
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssio_hvc_clamped_pad VSSD VDDIO VSSIO VSSIO_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VDDIO_Q
X0 VSSD VSSIO VDDIO VDDIO VSSIO VSSIO_PAD sky130_fd_io__top_ground_hvc_wpad
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssa_hvc_clamped_pad VSSD VDDIO VSSA VDDA VSSA_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSA VDDA VDDIO VSSA VSSA_PAD sky130_fd_io__top_ground_hvc_wpad
.ENDS
***************************************
.SUBCKT ICV_13 1 16 115 193 195 199 206 207 212 213 214 215
**
X0 1 193 16 199 195 212 sky130_ef_io__vccd_lvc_clamped2_pad
X1 1 115 16 207 195 215 sky130_ef_io__vccd_lvc_clamped2_pad
X2 1 195 16 213 sky130_ef_io__vssio_hvc_clamped_pad
X3 1 195 115 206 214 sky130_ef_io__vssa_hvc_clamped_pad
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_power_hvc_wpadv2 VSSD SRC_BDY_HVC DRN_HVC VDDIO P_CORE P_PAD
**
*.CALIBRE ISOLATED NETS: OGC_HVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
XM0 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM1 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM2 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM3 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250001 sb=250020 a=5 p=21
XM4 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM5 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM6 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM7 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250003 sb=250020 a=5 p=21
XM8 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM9 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM10 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM11 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250006 sb=250020 a=5 p=21
XM12 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM13 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM14 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM15 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250008 sb=250020 a=5 p=21
XM16 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM17 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM18 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM19 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250001 sb=250020 a=10 p=41
XM20 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM21 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM22 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250010 sb=250020 a=5 p=21
XM23 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM24 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM25 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM26 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250003 sb=250020 a=10 p=41
XM27 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM28 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM29 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250012 sb=250020 a=5 p=21
XM30 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM31 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM32 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM33 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250006 sb=250020 a=10 p=41
XM34 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM35 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM36 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250015 sb=250020 a=5 p=21
XM37 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM38 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM39 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM40 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250008 sb=250020 a=10 p=41
XM41 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM42 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM43 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250017 sb=250020 a=5 p=21
XM44 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM45 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM46 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM47 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250010 sb=250020 a=10 p=41
XM48 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM49 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM50 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250020 a=5 p=21
XM51 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM52 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM53 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM54 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250012 sb=250020 a=10 p=41
XM55 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM56 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM57 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250020 a=5 p=21
XM58 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM59 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM60 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM61 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250015 sb=250020 a=10 p=41
XM62 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM63 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM64 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250020 a=5 p=21
XM65 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM66 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM67 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM68 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250017 sb=250020 a=10 p=41
XM69 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM70 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM71 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250020 a=5 p=21
XM72 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM73 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM74 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM75 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM76 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM77 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250020 a=10 p=41
XM78 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250020 a=5 p=21
XM79 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM80 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM81 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM82 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM83 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM84 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250020 a=10 p=41
XM85 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250020 a=5 p=21
XM86 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM87 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM88 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM89 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM90 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM91 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250017 a=10 p=41
XM92 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250017 a=5 p=21
XM93 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM94 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM95 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM96 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM97 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM98 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250015 a=10 p=41
XM99 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250015 a=5 p=21
XM100 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM101 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM102 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM103 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM104 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM105 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250012 a=10 p=41
XM106 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250012 a=5 p=21
XM107 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM108 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM109 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM110 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM111 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM112 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250010 a=10 p=41
XM113 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250010 a=5 p=21
XM114 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM115 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM116 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM117 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM118 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM119 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250008 a=10 p=41
XM120 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250008 a=5 p=21
XM121 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM122 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM123 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM124 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM125 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM126 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250006 a=10 p=41
XM127 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250006 a=5 p=21
XM128 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM129 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM130 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM131 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM132 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM133 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 sa=250020 sb=250003 a=10 p=41
XM134 DRN_HVC 21 SRC_BDY_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 sa=250020 sb=250003 a=5 p=21
XM135 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM136 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM137 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM138 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM139 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM140 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 sa=250020 sb=250001 a=10 p=41
XM141 SRC_BDY_HVC 21 DRN_HVC SRC_BDY_HVC sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 sa=250020 sb=250001 a=5 p=21
X142 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X143 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X144 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X145 SRC_BDY_HVC VDDIO condiode a=1e-06 p=0.004 m=1
X146 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=126.766 p=0 m=1
X147 VSSD DRN_HVC sky130_fd_pr__model__parasitic__diode_ps2nw a=369.745 p=100.13 m=1
X148 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn a=10358.7 p=619.08 m=1
X149 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=137.463 p=47.72 m=1
X150 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=8184.99 p=443.22 m=1
X151 SRC_BDY_HVC VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=1172.63 p=163 m=1
R152 P_CORE P_PAD 0.01 short m=1
X153 19 20 sky130_fd_pr__res_bent_po__example_55959141808669
X225 SRC_BDY_HVC 19 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664
X226 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X227 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X228 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X229 SRC_BDY_HVC 19 sky130_fd_io__sio_clamp_pcap_4x5
X230 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap
X231 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap
X232 SRC_BDY_HVC 19 sky130_fd_io__esd_rcclamp_nfetcap
X233 SRC_BDY_HVC 19 21 sky130_fd_pr__nfet_01v8__example_55959141808677
X234 SRC_BDY_HVC 19 ICV_8
X235 SRC_BDY_HVC 19 ICV_8
X236 SRC_BDY_HVC 19 ICV_8
X237 SRC_BDY_HVC 19 ICV_8
X238 SRC_BDY_HVC 19 ICV_8
X239 SRC_BDY_HVC 19 ICV_8
X247 DRN_HVC 18 sky130_fd_pr__res_bent_po__example_55959141808668
X248 DRN_HVC 19 21 sky130_fd_pr__pfet_01v8__example_55959141808665
X249 18 20 sky130_fd_pr__res_bent_po__example_55959141808667
.ENDS
***************************************
.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad VSSD VSSIO VDDIO VDDIO_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
X0 VSSD VSSIO VDDIO VDDIO VDDIO VDDIO_PAD sky130_fd_io__top_power_hvc_wpadv2
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
.SUBCKT ICV_14 1 3 16
**
X0 1 3 16 38 sky130_ef_io__vddio_hvc_clamped_pad
.ENDS
***************************************
.SUBCKT sky130_ef_io__vdda_hvc_clamped_pad VSSD VSSA VDDIO VDDA VDDA_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VCCD VSSIO VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSA VDDA VDDIO VDDA VDDA_PAD sky130_fd_io__top_power_hvc_wpadv2
.ENDS
***************************************
.SUBCKT ICV_15 1 142 191 192 229 239 248 249
**
X0 1 191 229 239 248 sky130_ef_io__vssa_hvc_clamped_pad
X1 1 192 191 142 249 sky130_ef_io__vdda_hvc_clamped_pad
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_ground_lvc_wpad VSSD SRC_BDY_LVC2 SRC_BDY_LVC1 DRN_LVC1 VDDIO DRN_LVC2 BDY2_B2B G_CORE G_PAD
**
*.CALIBRE ISOLATED NETS: OGC_LVC VCCHIB VCCD VDDA VSSIO VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
XM0 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM1 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM2 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM3 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM4 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90001.1 sb=90019.9 a=0.9 p=10.36
XM5 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM6 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM7 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM8 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM9 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM10 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90002.3 sb=90019.9 a=0.9 p=10.36
XM11 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM12 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=4 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=20 p=18
XM13 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM14 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM15 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM16 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM17 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90003.9 sb=90019.9 a=0.9 p=10.36
XM18 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90001.1 sb=90019.9 a=1.26 p=14.36
XM19 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM20 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM21 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM22 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM23 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM24 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM25 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM26 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM27 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90005.1 sb=90019.9 a=0.9 p=10.36
XM28 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90002.3 sb=90019.9 a=1.26 p=14.36
XM29 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM30 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM31 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM32 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM33 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM34 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM35 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM36 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM37 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90006.6 sb=90019.9 a=0.9 p=10.36
XM38 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90003.9 sb=90019.9 a=1.26 p=14.36
XM39 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM40 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM41 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM42 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM43 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM44 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90007.8 sb=90019.9 a=0.9 p=10.36
XM45 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90005.1 sb=90019.9 a=1.26 p=14.36
XM46 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM47 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM48 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM49 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM50 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM51 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM52 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM53 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM54 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90009.4 sb=90019.9 a=0.9 p=10.36
XM55 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90006.6 sb=90019.9 a=1.26 p=14.36
XM56 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM57 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM58 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM59 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM60 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM61 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM62 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM63 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM64 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90010.6 sb=90019.9 a=0.9 p=10.36
XM65 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90007.8 sb=90019.9 a=1.26 p=14.36
XM66 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM67 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM68 SRC_BDY_LVC2 23 25 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM69 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM70 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM71 SRC_BDY_LVC1 21 24 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=2.3975 AS=4.76 PD=7.685 PS=15.36 NRD=6.936 NRS=6.852 m=1 sa=90000.6 sb=90019.9 a=1.26 p=14.36
XM72 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=40 p=26
XM73 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM74 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM75 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM76 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM77 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90012.2 sb=90019.9 a=0.9 p=10.36
XM78 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90009.4 sb=90019.9 a=1.26 p=14.36
XM79 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM80 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90001.7 sb=90019.9 a=0.9 p=10.36
XM81 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90001.7 sb=90019.9 a=1.26 p=14.36
XM82 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM83 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM84 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM85 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM86 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM87 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM88 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM89 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90013.4 sb=90019.9 a=0.9 p=10.36
XM90 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90010.6 sb=90019.9 a=1.26 p=14.36
XM91 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM92 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90003.1 sb=90019.9 a=0.9 p=10.36
XM93 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90003.1 sb=90019.9 a=1.26 p=14.36
XM94 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM95 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM96 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM97 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM98 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM99 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM100 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM101 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90015 sb=90019.9 a=0.9 p=10.36
XM102 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90012.2 sb=90019.9 a=1.26 p=14.36
XM103 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM104 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM105 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM106 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM107 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM108 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90016.1 sb=90019.9 a=0.9 p=10.36
XM109 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90013.4 sb=90019.9 a=1.26 p=14.36
XM110 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM111 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90005.9 sb=90019.9 a=0.9 p=10.36
XM112 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90005.9 sb=90019.9 a=1.26 p=14.36
XM113 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM114 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM115 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM116 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM117 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM118 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM119 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM120 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90017.7 sb=90019.9 a=0.9 p=10.36
XM121 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90015 sb=90019.9 a=1.26 p=14.36
XM122 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM123 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90007.3 sb=90019.9 a=0.9 p=10.36
XM124 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90007.3 sb=90019.9 a=1.26 p=14.36
XM125 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM126 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM127 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM128 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM129 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM130 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM131 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM132 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90018.9 sb=90019.9 a=0.9 p=10.36
XM133 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90016.2 sb=90019.9 a=1.26 p=14.36
XM134 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM135 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=40 p=26
XM136 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM137 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM138 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM139 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM140 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=2.3975 PD=7.28 PS=7.685 NRD=0 NRS=0 m=1 sa=4e+06 sb=4.00002e+06 a=56 p=30
XM141 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM142 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM143 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM144 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM145 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM146 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90017.7 sb=90019.9 a=1.26 p=14.36
XM147 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM148 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90010.1 sb=90019.9 a=0.9 p=10.36
XM149 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90010.1 sb=90019.9 a=1.26 p=14.36
XM150 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM151 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM152 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM153 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM154 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM155 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM156 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM157 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM158 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90018.9 sb=90019.9 a=1.26 p=14.36
XM159 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM160 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90011.4 sb=90019.9 a=0.9 p=10.36
XM161 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90011.4 sb=90019.9 a=1.26 p=14.36
XM162 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM163 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM164 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM165 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM166 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM167 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM168 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM169 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM170 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM171 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM172 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM173 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM174 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM175 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM176 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM177 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM178 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM179 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90014.3 sb=90019.9 a=0.9 p=10.36
XM180 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90014.3 sb=90019.9 a=1.26 p=14.36
XM181 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM182 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM183 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM184 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM185 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM186 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM187 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM188 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM189 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM190 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM191 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90015.6 sb=90019.9 a=0.9 p=10.36
XM192 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90015.6 sb=90019.9 a=1.26 p=14.36
XM193 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM194 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM195 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM196 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM197 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM198 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM199 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM200 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM201 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM202 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM203 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4.00002e+06 a=40 p=26
XM204 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM205 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM206 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM207 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM208 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00002e+06 a=56 p=30
XM209 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM210 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM211 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM212 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM213 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM214 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM215 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM216 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90018.5 sb=90019.9 a=0.9 p=10.36
XM217 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90018.5 sb=90019.9 a=1.26 p=14.36
XM218 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM219 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM220 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM221 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM222 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM223 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM224 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM225 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM226 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM227 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM228 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.8 sb=90019.9 a=0.9 p=10.36
XM229 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.8 sb=90019.9 a=1.26 p=14.36
XM230 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM231 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM232 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM233 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM234 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM235 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM236 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM237 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM238 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM239 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM240 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM241 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM242 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM243 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM244 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90019.9 a=0.9 p=10.36
XM245 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM246 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90019.9 a=1.26 p=14.36
XM247 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90019.8 a=0.9 p=10.36
XM248 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM249 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM250 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM251 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90019.8 a=1.26 p=14.36
XM252 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM253 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM254 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM255 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM256 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90018.9 a=0.9 p=10.36
XM257 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM258 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90018.9 a=1.26 p=14.36
XM259 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90018.5 a=0.9 p=10.36
XM260 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM261 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM262 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM263 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90018.5 a=1.26 p=14.36
XM264 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM265 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM266 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM267 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM268 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90017.7 a=0.9 p=10.36
XM269 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM270 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90017.7 a=1.26 p=14.36
XM271 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4.00001e+06 a=40 p=26
XM272 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM273 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM274 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM275 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM276 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00001e+06 sb=4.00001e+06 a=56 p=30
XM277 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM278 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM279 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM280 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM281 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90016.1 a=0.9 p=10.36
XM282 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM283 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90016.2 a=1.26 p=14.36
XM284 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90015.6 a=0.9 p=10.36
XM285 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM286 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM287 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM288 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90015.6 a=1.26 p=14.36
XM289 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM290 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM291 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM292 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM293 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90015 a=0.9 p=10.36
XM294 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM295 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90015 a=1.26 p=14.36
XM296 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90014.3 a=0.9 p=10.36
XM297 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM298 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM299 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM300 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90014.3 a=1.26 p=14.36
XM301 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM302 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM303 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM304 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM305 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90013.4 a=0.9 p=10.36
XM306 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM307 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90013.4 a=1.26 p=14.36
XM308 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM309 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM310 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM311 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM312 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90012.2 a=0.9 p=10.36
XM313 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM314 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90012.2 a=1.26 p=14.36
XM315 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90011.4 a=0.9 p=10.36
XM316 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM317 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM318 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM319 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90011.4 a=1.26 p=14.36
XM320 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM321 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM322 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM323 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM324 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90010.6 a=0.9 p=10.36
XM325 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM326 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90010.6 a=1.26 p=14.36
XM327 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90010.1 a=0.9 p=10.36
XM328 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM329 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM330 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM331 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90010.1 a=1.26 p=14.36
XM332 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM333 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM334 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM335 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM336 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90009.4 a=0.9 p=10.36
XM337 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM338 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90009.4 a=1.26 p=14.36
XM339 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=40 p=26
XM340 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM341 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM342 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM343 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM344 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM345 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM346 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM347 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM348 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM349 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90007.8 a=0.9 p=10.36
XM350 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM351 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90007.8 a=1.26 p=14.36
XM352 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90007.3 a=0.9 p=10.36
XM353 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM354 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM355 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM356 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90007.3 a=1.26 p=14.36
XM357 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM358 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM359 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM360 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM361 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90006.6 a=0.9 p=10.36
XM362 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM363 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90006.6 a=1.26 p=14.36
XM364 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90005.9 a=0.9 p=10.36
XM365 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM366 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM367 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM368 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90005.9 a=1.26 p=14.36
XM369 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM370 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM371 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM372 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM373 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90005.1 a=0.9 p=10.36
XM374 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM375 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90005.1 a=1.26 p=14.36
XM376 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM377 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM378 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM379 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM380 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90003.9 a=0.9 p=10.36
XM381 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM382 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90003.9 a=1.26 p=14.36
XM383 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.925 AS=5.625 PD=6.17 PS=12.25 NRD=6.6 NRS=19.788 m=1 sa=90019.9 sb=90003.1 a=0.9 p=10.36
XM384 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM385 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM386 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM387 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=4.095 AS=7.875 PD=8.17 PS=16.25 NRD=4.704 NRS=14.136 m=1 sa=90019.9 sb=90003.1 a=1.26 p=14.36
XM388 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM389 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM390 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM391 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM392 DRN_LVC2 25 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.525 AS=2.5 PD=6.01 PS=11 NRD=4.68 NRS=4.8 m=1 sa=90019.9 sb=90002.3 a=0.9 p=10.36
XM393 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM394 DRN_LVC1 24 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.535 AS=3.5 PD=8.01 PS=15 NRD=3.336 NRS=3.42 m=1 sa=90019.9 sb=90002.3 a=1.26 p=14.36
XM395 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=5.625 AS=2.925 PD=12.25 PS=6.17 NRD=19.788 NRS=6.6 m=1 sa=90019.9 sb=90001.7 a=0.9 p=10.36
XM396 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM397 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM398 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM399 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=7.875 AS=4.095 PD=16.25 PS=8.17 NRD=14.136 NRS=4.704 m=1 sa=90019.9 sb=90001.7 a=1.26 p=14.36
XM400 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM401 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM402 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM403 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM404 SRC_BDY_LVC2 25 DRN_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=0.18 W=5 AD=2.5 AS=2.525 PD=11 PS=6.01 NRD=4.8 NRS=4.68 m=1 sa=90019.9 sb=90001.1 a=0.9 p=10.36
XM405 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM406 SRC_BDY_LVC1 24 DRN_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=0.18 W=7 AD=3.5 AS=3.535 PD=15 PS=8.01 NRD=3.42 NRS=3.336 m=1 sa=90019.9 sb=90001.1 a=1.26 p=14.36
XM407 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=40 p=26
XM408 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM409 SRC_BDY_LVC2 23 SRC_BDY_LVC2 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM410 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM411 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
XM412 SRC_BDY_LVC1 21 SRC_BDY_LVC1 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8 L=8 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=4.00002e+06 sb=4e+06 a=56 p=30
X413 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1
X414 SRC_BDY_LVC2 VDDIO condiode a=1e-06 p=0.004 m=1
X415 SRC_BDY_LVC1 VDDIO condiode a=1e-06 p=0.004 m=1
X416 VSSD DRN_LVC1 sky130_fd_pr__model__parasitic__diode_ps2nw a=108.41 p=46.58 m=1
X417 VSSD DRN_LVC2 sky130_fd_pr__model__parasitic__diode_ps2nw a=108.41 p=46.58 m=1
X418 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2dn a=10516.3 p=468.87 m=1
X419 SRC_BDY_LVC2 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=4115.42 p=264.63 m=1
X420 SRC_BDY_LVC1 VDDIO sky130_fd_pr__model__parasitic__diode_pw2dn a=5703.29 p=340.89 m=1
R421 DRN_LVC1 21 sky130_fd_pr__res_generic_po L=1950 W=0.33 m=1
R422 G_CORE G_PAD 0.01 short m=1
X423 27 DRN_LVC2 sky130_fd_pr__res_bent_po__example_55959141808692
X424 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X425 DRN_LVC1 21 24 sky130_fd_pr__pfet_01v8__example_55959141808687
X426 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X427 DRN_LVC2 23 25 sky130_fd_pr__pfet_01v8__example_55959141808687
X616 23 26 sky130_fd_pr__res_bent_po__example_55959141808691
X622 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808704
X623 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808695
X630 VSSD BDY2_B2B SRC_BDY_LVC1 sky130_fd_io__gnd2gnd_120x2_lv_isosub
X631 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808701
X632 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X633 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X634 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808703
X635 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X636 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X637 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X638 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808705
X639 SRC_BDY_LVC1 sky130_fd_pr__nfet_01v8__example_55959141808705
X640 SRC_BDY_LVC2 sky130_fd_pr__nfet_01v8__example_55959141808693
X642 22 26 sky130_fd_pr__res_bent_po__example_55959141808688
X643 27 22 sky130_fd_pr__res_bent_po__example_55959141808690
.ENDS
***************************************
.SUBCKT sky130_ef_io__vssd_lvc_clamped2_pad VSSD VSSA VSSIO VCCD VDDIO VSSD_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSIO VCCD VDDIO VCCD VSSA VSSD VSSD_PAD sky130_fd_io__top_ground_lvc_wpad
.ENDS
***************************************
.SUBCKT ICV_16 1 2 3 6 7 8 9 12 13 14 15 16
**
X0 1 9 6 8 15 sky130_ef_io__vdda_hvc_clamped_pad
X1 1 7 6 2 17 sky130_ef_io__vdda_hvc_clamped_pad
X2 1 9 3 12 6 14 sky130_ef_io__vssd_lvc_clamped2_pad
X3 1 7 3 13 6 16 sky130_ef_io__vssd_lvc_clamped2_pad
.ENDS
***************************************
.SUBCKT ICV_17 1 68 132 176 233 241
**
X0 1 176 132 233 329 sky130_ef_io__vssa_hvc_clamped_pad
X1 1 68 176 241 sky130_ef_io__vddio_hvc_clamped_pad
.ENDS
***************************************
.SUBCKT ICV_18 1 3 8 26 30 42 43
**
X0 1 8 3 88 sky130_ef_io__vssio_hvc_clamped_pad
X1 1 8 26 30 42 sky130_ef_io__vssa_hvc_clamped_pad
X2 1 26 8 30 43 sky130_ef_io__vdda_hvc_clamped_pad
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2o_cdns_55959141808653 2 3
**
R0 2 6 0.01 short m=1
R1 7 3 0.01 short m=1
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808652 2 3
**
R0 2 6 0.01 short m=1
R1 6 3 0.01 short m=1
.ENDS
***************************************


***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180838 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=10.2 W=0.5 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180864 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=1.5 W=0.8 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180859 2 3
**
R0 2 6 0.01 short m=1
R1 6 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__res250only_small PAD ROUT
**
R0 PAD 6 sky130_fd_pr__res_generic_po L=0.17 W=2 m=1
R1 6 7 sky130_fd_pr__res_generic_po L=10.07 W=2 m=1
R2 7 ROUT sky130_fd_pr__res_generic_po L=0.17 W=2 m=1
R3 PAD 6 0.01 short m=1
R4 7 ROUT 0.01 short m=1
R5 PAD 6 0.01 short m=1
R6 7 ROUT 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180862 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=6 W=0.8 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180863 2 3
**
R0 2 3 sky130_fd_pr__res_generic_po L=12 W=0.8 m=1
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 2 3
**
R0 2 6 0.01 short m=1
R1 7 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_p_em1c_cdns_55959141808753 2
**
R0 2 5 0.01 short m=1
R1 2 6 0.01 short m=1
.ENDS
***************************************
.SUBCKT ICV_20 2 3
**
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X1 2 sky130_fd_io__xres_p_em1c_cdns_55959141808753
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808754 2 3
**
*.SEEDPROM
R0 2 3 sky130_fd_pr__res_generic_nd L=14 W=0.5 m=1
.ENDS
***************************************
.SUBCKT ICV_21 2 3 4 5
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754
X1 4 5 sky130_fd_pr__res_generic_nd__example_55959141808754
.ENDS
***************************************
.SUBCKT ICV_22 2 3 4 5 6 7 8 9
**
*.SEEDPROM
X0 4 2 3 5 ICV_21
X1 8 6 7 9 ICV_21
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 2 3
**
R0 2 6 0.01 short m=1
R1 7 3 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 2
**
R0 2 5 0.01 short m=1
R1 2 6 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 2
**
R0 2 5 0.01 short m=1
R1 2 6 0.01 short m=1
.ENDS
***************************************


***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 1
**
R0 1 4 0.01 short m=1
R1 1 5 0.01 short m=1
.ENDS
***************************************
.SUBCKT ICV_25 2 3 4
**
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X1 4 sky130_fd_io__xres_p_em1c_cdns_55959141808753
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 1 2
**
R0 2 5 0.01 short m=1
R1 6 1 0.01 short m=1
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808755 2 3
**
*.SEEDPROM
R0 2 3 sky130_fd_pr__res_generic_nd L=47 W=0.5 m=1
.ENDS
***************************************
.SUBCKT ICV_26 2 3 4
**
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754
X1 4 2 sky130_fd_pr__res_generic_nd__example_55959141808755
.ENDS
***************************************
.SUBCKT ICV_27 2 3
**
*.SEEDPROM
X0 2 2 sky130_fd_pr__res_generic_nd__example_55959141808754
X1 2 3 sky130_fd_pr__res_generic_nd__example_55959141808755
.ENDS
***************************************
.SUBCKT ICV_28 2 3 4 5 6
**
*.SEEDPROM
X0 3 4 2 ICV_26
X1 5 6 ICV_27
.ENDS
***************************************
.SUBCKT ICV_29 2 3 4 5 6 7 8 9 10 11
**
*.SEEDPROM
X0 2 4 6 5 3 ICV_28
X1 7 9 11 10 8 ICV_28
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres2v2_rcfilter_lpfv2 1 VCC_IO 3 4 5 6 7 8 9 10 11 12 13 IN
**
XM0 1 3 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=28 p=22
XM1 1 4 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=28 p=22
XM2 1 5 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22
XM3 1 6 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22
XM4 1 7 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM5 1 8 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM6 1 9 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM7 1 10 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM8 1 11 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22
XM9 1 11 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22
XM10 1 12 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2e+06 a=28 p=22
XM11 1 13 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=4 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2e+06 a=28 p=22
XM12 VCC_IO 3 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=28 p=22
XM13 VCC_IO 4 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2e+06 sb=2.00002e+06 a=28 p=22
XM14 VCC_IO 5 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22
XM15 VCC_IO 6 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22
XM16 VCC_IO 7 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM17 VCC_IO 8 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM18 VCC_IO 9 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM19 VCC_IO 10 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22
XM20 VCC_IO 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22
XM21 VCC_IO 11 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22
XM22 VCC_IO 12 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2e+06 a=28 p=22
XM23 VCC_IO 13 VCC_IO VCC_IO sky130_fd_pr__pfet_g5v0d10v5 L=4 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 sa=2.00002e+06 sb=2e+06 a=28 p=22
X24 1 8 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X25 1 7 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X26 1 6 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X27 1 5 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X28 1 4 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X29 1 3 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X30 1 15 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X31 1 16 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X32 1 17 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X33 1 18 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X34 1 19 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X35 1 20 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X36 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X37 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X38 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X39 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X40 1 3 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X41 1 9 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X42 1 15 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X43 1 16 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X44 1 17 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X45 1 18 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X46 1 19 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X47 1 20 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X48 1 21 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X49 1 22 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X50 1 23 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X51 1 24 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X52 1 25 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X53 1 26 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X54 1 27 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X55 1 28 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X56 1 29 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X57 1 30 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X58 1 31 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X59 1 32 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X60 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X61 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X62 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X63 1 1 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X64 1 3 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X65 1 9 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X66 1 15 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X67 1 16 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X68 1 17 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X69 1 18 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X70 1 19 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X71 1 20 sky130_fd_pr__diode_pw2nd_05v5 a=15.5025 p=62.01 m=1
X72 1 38 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X73 1 39 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X74 1 37 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X75 1 40 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X76 1 36 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X77 1 41 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X78 1 35 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X79 1 42 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X80 1 34 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X81 1 43 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X82 1 33 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X83 1 44 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X84 1 45 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X85 1 10 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X86 1 46 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X87 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X88 1 47 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X89 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X90 1 48 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X91 1 12 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X92 1 49 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X93 1 13 sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X94 1 50 sky130_fd_pr__diode_pw2nd_05v5 a=12.0235 p=48.594 m=1
X95 1 IN sky130_fd_pr__diode_pw2nd_05v5 a=12.024 p=48.596 m=1
X96 1 33 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X97 1 34 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X98 1 35 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X99 1 36 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X100 1 37 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X101 1 38 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X102 1 13 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X103 1 12 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X104 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X105 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X106 1 10 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X107 1 9 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X108 1 33 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X109 1 34 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X110 1 35 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X111 1 36 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X112 1 37 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X113 1 38 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X114 1 IN sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X115 1 13 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X116 1 12 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X117 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X118 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X119 1 10 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X120 1 44 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X121 1 33 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X122 1 43 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X123 1 34 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X124 1 42 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X125 1 35 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X126 1 41 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X127 1 36 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X128 1 40 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X129 1 37 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X130 1 39 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X131 1 38 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X132 1 IN sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X133 1 50 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X134 1 13 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X135 1 49 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X136 1 12 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X137 1 48 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X138 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X139 1 47 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X140 1 11 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X141 1 46 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X142 1 10 sky130_fd_pr__diode_pw2nd_05v5 a=3.7735 p=15.594 m=1
X143 1 45 sky130_fd_pr__diode_pw2nd_05v5 a=3.774 p=15.596 m=1
X144 1 VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=501.44 p=125.96 m=1
X164 20 32 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X165 8 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X166 7 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X167 6 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X168 5 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X169 3 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X170 9 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X171 12 49 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X172 11 47 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X173 9 45 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757
X174 15 sky130_fd_io__xres_p_em1c_cdns_55959141808753
X175 IN sky130_fd_io__xres_p_em1c_cdns_55959141808753
X176 12 sky130_fd_io__xres_p_em1c_cdns_55959141808753
X177 11 sky130_fd_io__xres_p_em1c_cdns_55959141808753
X178 33 44 ICV_20
X179 34 43 ICV_20
X180 35 42 ICV_20
X181 36 41 ICV_20
X182 37 40 ICV_20
X183 38 39 ICV_20
X184 13 50 ICV_20
X185 11 48 ICV_20
X186 10 46 ICV_20
X187 34 43 34 34 33 44 33 33 ICV_22
X188 36 41 36 36 35 42 35 35 ICV_22
X189 38 39 38 38 37 40 37 37 ICV_22
X190 12 13 49 13 13 IN 50 IN ICV_22
X191 11 11 47 11 11 12 48 12 ICV_22
X192 9 10 45 10 10 11 46 11 ICV_22
X193 1 7 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X194 1 6 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X195 1 5 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X196 1 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X197 13 12 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X198 12 11 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X199 11 10 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X200 10 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758
X201 3 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760
X202 11 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760
X203 9 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761
X204 4 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761
X218 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X219 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X220 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X221 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759
X222 8 21 1 ICV_25
X223 7 22 1 ICV_25
X224 6 23 1 ICV_25
X225 5 24 1 ICV_25
X226 4 25 3 ICV_25
X227 3 26 9 ICV_25
X228 15 27 16 ICV_25
X229 16 28 17 ICV_25
X230 17 29 18 ICV_25
X231 18 30 19 ICV_25
X232 19 31 20 ICV_25
X233 1 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756
X234 1 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756
X235 32 20 IN ICV_26
X236 15 45 ICV_27
X237 13 31 19 20 50 ICV_28
X238 38 39 21 1 8 37 40 22 1 7 ICV_29
X239 36 41 23 1 6 35 42 24 1 5 ICV_29
X240 34 43 25 3 4 33 44 26 9 3 ICV_29
X241 10 46 27 16 15 11 47 28 17 16 ICV_29
X242 11 48 29 18 17 12 49 30 19 18 ICV_29
.ENDS


***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808767 2 3 4 5
**
*.SEEDPROM
XM0 5 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
.ENDS


***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808764 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808779 1 2 3 4
**
XM0 4 2 3 1 sky130_fd_pr__nfet_05v0_nvt L=0.9 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 sa=450000 sb=450000 a=0.9 p=3.8
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808777 1 2 3
**
XM0 3 2 1 1 sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=3 AD=0.84 AS=0.795 PD=6.56 PS=6.53 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
.ENDS

***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808784 2 3 4
**
*.SEEDPROM
XM0 2 3 4 2 sky130_fd_pr__pfet_g5v0d10v5 L=0.8 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=0.8 p=3.6
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term NBODY NWELLRING GATE VGND IN 7
**
*.SEEDPROM
XM0 IN GATE VGND NBODY sky130_fd_pr__esd_nfet_g5v0d10v5 L=0.6 W=5.4 AD=3.65486 AS=3.65486 PD=11.6192 PS=11.6192 NRD=8.436 NRS=9.2796 m=1 sa=300000 sb=300000 a=3.24 p=12
R1 NWELLRING 7 0.01 short m=1
R2 NBODY 51 0.01 short m=1
.ENDS
***************************************

***************************************
.SUBCKT sky130_fd_io__gpio_buf_localesdv2 VGND VCC_IO VTRIP_SEL_H OUT_H 5
**
*.SEEDPROM
XM0 OUT_VT VTRIP_SEL_H OUT_H VGND sky130_fd_pr__nfet_g5v0d10v5 L=1 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 sa=500000 sb=500000 a=3 p=8
X1 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=8.5092 p=29.27 m=1
X2 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=8.5092 p=29.27 m=1
X3 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=8.5092 p=29.27 m=1
X4 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=8.5092 p=29.27 m=1
X5 VGND VCC_IO sky130_fd_pr__model__parasitic__diode_ps2nw a=5.1688 p=17.34 m=1
X6 5 OUT_H sky130_fd_io__res250only_small
X7 VGND VCC_IO VGND VGND OUT_VT 8 sky130_fd_io__signal_5_sym_hv_local_5term
X8 VGND VCC_IO VGND VGND OUT_H 10 sky130_fd_io__signal_5_sym_hv_local_5term
X9 VGND VCC_IO VGND OUT_VT VCC_IO 7 sky130_fd_io__signal_5_sym_hv_local_5term
X10 VGND VCC_IO VGND OUT_H VCC_IO 9 sky130_fd_io__signal_5_sym_hv_local_5term
.ENDS


***************************************
.SUBCKT sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 1 2 VCC_IO 4 5 6 7 8 9 10 11 12 13 14
**
*.SEEDPROM
XM0 14 4 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 sa=300002 sb=300020 a=3 p=11.2
XM1 14 4 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 sa=300002 sb=300020 a=3 p=11.2
XM2 2 4 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300004 sb=300020 a=3 p=11.2
XM3 2 4 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300004 sb=300020 a=3 p=11.2
XM4 14 4 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300007 sb=300020 a=3 p=11.2
XM5 14 4 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300007 sb=300020 a=3 p=11.2
XM6 2 4 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300009 sb=300020 a=3 p=11.2
XM7 2 4 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300009 sb=300020 a=3 p=11.2
XM8 14 5 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300011 sb=300020 a=3 p=11.2
XM9 14 5 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300011 sb=300020 a=3 p=11.2
XM10 2 5 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300014 sb=300020 a=3 p=11.2
XM11 2 5 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300014 sb=300020 a=3 p=11.2
XM12 14 5 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300016 sb=300020 a=3 p=11.2
XM13 14 5 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300016 sb=300020 a=3 p=11.2
XM14 2 6 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300019 sb=300020 a=3 p=11.2
XM15 2 6 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300019 sb=300020 a=3 p=11.2
XM16 14 6 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM17 14 6 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM18 2 6 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM19 2 6 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM20 14 7 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM21 14 7 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM22 2 7 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM23 2 7 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM24 14 7 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM25 14 7 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM26 2 8 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM27 2 8 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM28 14 9 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM29 14 9 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM30 2 9 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM31 2 9 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM32 14 9 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM33 14 9 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM34 2 10 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM35 2 10 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM36 14 10 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM37 14 10 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM38 2 10 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM39 2 10 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300020 a=3 p=11.2
XM40 14 10 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300018 a=3 p=11.2
XM41 14 10 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300018 a=3 p=11.2
XM42 2 10 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300016 a=3 p=11.2
XM43 2 10 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300016 a=3 p=11.2
XM44 14 10 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300013 a=3 p=11.2
XM45 14 10 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300013 a=3 p=11.2
XM46 2 11 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300011 a=3 p=11.2
XM47 2 11 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300011 a=3 p=11.2
XM48 14 12 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300008 a=3 p=11.2
XM49 14 12 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300008 a=3 p=11.2
XM50 2 13 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300006 a=3 p=11.2
XM51 2 13 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300006 a=3 p=11.2
XM52 14 13 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300003 a=3 p=11.2
XM53 14 13 2 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 sa=300020 sb=300003 a=3 p=11.2
XM54 2 13 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 sa=300020 sb=300002 a=3 p=11.2
XM55 2 13 14 2 sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 sa=300020 sb=300002 a=3 p=11.2
X56 1 VCC_IO sky130_fd_pr__model__parasitic__diode_ps2dn a=1791.37 p=197.77 m=1
X57 2 VCC_IO sky130_fd_pr__model__parasitic__diode_pw2dn a=1558.74 p=186.49 m=1
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_xres4v2 1 TIE_LO_ESD VGND_IO VCC_IO PD_H[2] PD_H[3] 7 8
**
*.SEEDPROM
X0 VGND_IO VCC_IO condiode a=1e-06 p=0.004 m=1
X1 PD_H[3] 7 sky130_fd_io__tk_em2o_cdns_55959141808653
X2 PD_H[2] 7 sky130_fd_io__tk_em2o_cdns_55959141808653
X3 PD_H[3] 15 sky130_fd_io__tk_em2o_cdns_55959141808653
X4 TIE_LO_ESD 15 sky130_fd_io__tk_em2o_cdns_55959141808653
X5 PD_H[3] 14 sky130_fd_io__tk_em2o_cdns_55959141808653
X6 TIE_LO_ESD 14 sky130_fd_io__tk_em2o_cdns_55959141808653
X7 PD_H[2] 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X8 TIE_LO_ESD 13 sky130_fd_io__tk_em2o_cdns_55959141808653
X9 PD_H[2] 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X10 TIE_LO_ESD 12 sky130_fd_io__tk_em2o_cdns_55959141808653
X11 PD_H[2] 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X12 TIE_LO_ESD 11 sky130_fd_io__tk_em2o_cdns_55959141808653
X13 PD_H[2] 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X14 TIE_LO_ESD 10 sky130_fd_io__tk_em2o_cdns_55959141808653
X15 PD_H[2] 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X16 PD_H[3] 9 sky130_fd_io__tk_em2o_cdns_55959141808653
X17 TIE_LO_ESD 7 sky130_fd_io__tk_em2s_cdns_55959141808652
X18 PD_H[2] 15 sky130_fd_io__tk_em2s_cdns_55959141808652
X19 PD_H[2] 14 sky130_fd_io__tk_em2s_cdns_55959141808652
X20 PD_H[3] 13 sky130_fd_io__tk_em2s_cdns_55959141808652
X21 PD_H[3] 12 sky130_fd_io__tk_em2s_cdns_55959141808652
X22 PD_H[3] 11 sky130_fd_io__tk_em2s_cdns_55959141808652
X23 PD_H[3] 10 sky130_fd_io__tk_em2s_cdns_55959141808652
X24 TIE_LO_ESD 9 sky130_fd_io__tk_em2s_cdns_55959141808652
X25 TIE_LO_ESD VGND_IO sky130_fd_pr__res_generic_po__example_5595914180838
X26 1 VGND_IO VCC_IO 9 10 11 12 13 PD_H[2] PD_H[3] 14 15 7 8 sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2
.ENDS
***************************************
.SUBCKT ICV_1 VSSD VDDIO VCCHIB VDDIO_Q ENABLE_H EN_VDDIO_SIG_H INP_SEL_H ENABLE_VDDIO PAD PULLUP_H DISABLE_PULLUP_H PAD_A_ESD_H VSSIO FILT_IN_H XRES_H_N TIE_WEAK_HI_H
**
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VCCD VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
XM0 VSSD ENABLE_VDDIO 36 VSSD sky130_fd_pr__nfet_01v8 L=0.15 W=0.74 AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 m=1 sa=75000.2 sb=75000.3 a=0.111 p=1.78
XM1 61 34 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 sa=300000 sb=300001 a=0.42 p=2.6
XM2 54 ENABLE_H 61 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 sa=300001 sb=300000 a=0.42 p=2.6
XM3 35 54 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.42 p=2.6
XM4 33 39 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM5 VSSD 39 33 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM6 32 37 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM7 VSSD 37 32 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM8 64 37 62 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 sa=400000 sb=400007 a=4 p=11.6
XM9 62 37 64 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400001 sb=400006 a=4 p=11.6
XM10 64 37 62 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400002 sb=400005 a=4 p=11.6
XM11 62 37 64 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400003 sb=400004 a=4 p=11.6
XM12 VSSD 30 62 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400004 sb=400003 a=4 p=11.6
XM13 62 30 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400005 sb=400002 a=4 p=11.6
XM14 37 30 62 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=400006 sb=400001 a=4 p=11.6
XM15 62 30 37 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 sa=400007 sb=400000 a=4 p=11.6
XM16 62 37 57 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.8 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 sa=400000 sb=400000 a=4 p=11.6
XM17 VSSD 31 52 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=0.5 p=3
XM18 52 31 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=250001 sb=250001 a=0.5 p=3
XM19 VSSD 31 52 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=0.5 p=3
XM20 43 71 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM21 VSSD 71 43 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM22 71 DISABLE_PULLUP_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM23 VSSD DISABLE_PULLUP_H 71 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM24 VSSD 41 63 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 sa=500000 sb=500000 a=0.42 p=2.84
XM25 63 42 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=1 p=4
XM26 44 42 63 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=1 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=1 p=4
XM27 41 44 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.5 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=0.5 p=3
XM28 40 INP_SEL_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300007 a=0.42 p=2.6
XM29 VSSD INP_SEL_H 40 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300006 a=0.42 p=2.6
XM30 34 EN_VDDIO_SIG_H VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300005 a=0.42 p=2.6
XM31 VSSD EN_VDDIO_SIG_H 34 VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300004 a=0.42 p=2.6
XM32 XRES_H_N 72 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.42 p=2.6
XM33 VSSD 72 XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300004 sb=300003 a=0.42 p=2.6
XM34 XRES_H_N 72 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300005 sb=300002 a=0.42 p=2.6
XM35 VSSD 72 XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300006 sb=300001 a=0.42 p=2.6
XM36 72 41 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300007 sb=300000 a=0.42 p=2.6
XM37 XRES_H_N 72 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.42 p=2.6
XM38 VSSD 72 XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.42 p=2.6
XM39 XRES_H_N 72 VSSD VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.42 p=2.6
XM40 VSSD 72 XRES_H_N VSSD sky130_fd_pr__nfet_g5v0d10v5 L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.42 p=2.6
XM41 24 35 60 VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=10 AD=2.8 AS=2.8 PD=20.56 PS=20.56 NRD=0 NRS=0 m=1 sa=450000 sb=450000 a=9 p=21.8
XM42 VSSD VSSD VSSD VSSD sky130_fd_pr__nfet_05v0_nvt L=0.9 W=10 AD=2.8 AS=2.65 PD=20.56 PS=20.53 NRD=0 NRS=0 m=1 sa=450000 sb=450000 a=9 p=21.8
XM43 VCCHIB ENABLE_VDDIO 36 VCCHIB sky130_fd_pr__pfet_01v8_hvt L=0.15 W=1.12 AD=0.3864 AS=0.3304 PD=2.93 PS=2.83 NRD=10.5395 NRS=1.7533 m=1 sa=75000.2 sb=75000.3 a=0.168 p=2.54
XM44 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 sa=300002 sb=300020 a=3 p=11.2
XM45 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 sa=300002 sb=300020 a=3 p=11.2
XM46 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300004 sb=300020 a=3 p=11.2
XM47 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300004 sb=300020 a=3 p=11.2
XM48 VDDIO_Q 32 33 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=0.21 p=1.84
XM49 32 33 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=0.42 AD=0.1176 AS=0.0588 PD=1.4 PS=0.7 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=0.21 p=1.84
XM50 54 34 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM51 54 34 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300001 a=0.6 p=3.2
XM52 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300007 sb=300020 a=3 p=11.2
XM53 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300007 sb=300020 a=3 p=11.2
XM54 VDDIO_Q ENABLE_H 54 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM55 VDDIO_Q ENABLE_H 54 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300000 a=0.6 p=3.2
XM56 VDDIO_Q 31 52 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.84 PD=3.28 PS=6.56 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=1.5 p=7
XM57 52 31 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 sa=250001 sb=250001 a=1.5 p=7
XM58 VDDIO_Q 31 52 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=1.5 p=7
XM59 VDDIO_Q 32 31 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.795 AS=0.84 PD=6.53 PS=6.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
XM60 35 54 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM61 35 54 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300000 a=0.6 p=3.2
XM62 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300009 sb=300020 a=3 p=11.2
XM63 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300009 sb=300020 a=3 p=11.2
XM64 VDDIO_Q ENABLE_H 55 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=1.4 PD=10.53 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=2.5 p=11
XM65 51 30 37 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=2.5 p=11
XM66 56 35 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM67 51 34 56 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM68 VDDIO_Q 34 57 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM69 58 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM70 VCCHIB 36 59 VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250001 a=2.5 p=11
XM71 60 36 VCCHIB VCCHIB sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250000 a=2.5 p=11
XM72 25 37 39 25 sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=2.5 p=11
XM73 45 37 39 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM74 26 34 45 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250001 a=2.5 p=11
XM75 VDDIO_Q 35 26 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM76 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300012 sb=300020 a=3 p=11.2
XM77 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300012 sb=300020 a=3 p=11.2
XM78 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300014 sb=300020 a=3 p=11.2
XM79 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300014 sb=300020 a=3 p=11.2
XM80 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300017 sb=300020 a=3 p=11.2
XM81 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300017 sb=300020 a=3 p=11.2
XM82 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300019 sb=300020 a=3 p=11.2
XM83 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300019 sb=300020 a=3 p=11.2
XM84 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM85 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM86 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM87 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM88 53 41 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=1 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 sa=500000 sb=500000 a=0.42 p=2.84
XM89 29 43 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 sa=250000 sb=250002 a=2.5 p=11
XM90 40 INP_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300007 a=0.6 p=3.2
XM91 VDDIO_Q INP_SEL_H 40 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300006 a=0.6 p=3.2
XM92 34 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300005 a=0.6 p=3.2
XM93 VDDIO_Q EN_VDDIO_SIG_H 34 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300004 a=0.6 p=3.2
XM94 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.6 p=3.2
XM95 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300003 a=0.6 p=3.2
XM96 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300002 a=0.6 p=3.2
XM97 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300001 a=0.6 p=3.2
XM98 72 41 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300007 sb=300000 a=0.6 p=3.2
XM99 VDDIO 43 29 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250001 sb=250002 a=2.5 p=11
XM100 53 42 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 AD=0.42 AS=0.84 PD=3.28 PS=6.56 NRD=0 NRS=0 m=1 sa=500000 sb=500001 a=3 p=8
XM101 44 42 53 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=1 W=3 AD=0.84 AS=0.42 PD=6.56 PS=3.28 NRD=0 NRS=0 m=1 sa=500001 sb=500000 a=3 p=8
XM102 41 44 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 sa=250000 sb=250000 a=1.5 p=7
XM103 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM104 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM105 29 43 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250001 a=2.5 p=11
XM106 40 INP_SEL_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300007 a=0.6 p=3.2
XM107 VDDIO_Q INP_SEL_H 40 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300006 a=0.6 p=3.2
XM108 34 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300005 a=0.6 p=3.2
XM109 VDDIO_Q EN_VDDIO_SIG_H 34 VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300004 a=0.6 p=3.2
XM110 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300003 a=0.6 p=3.2
XM111 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300004 sb=300003 a=0.6 p=3.2
XM112 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300005 sb=300002 a=0.6 p=3.2
XM113 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300006 sb=300001 a=0.6 p=3.2
XM114 72 41 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300007 sb=300000 a=0.6 p=3.2
XM115 43 71 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM116 VDDIO 71 43 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM117 71 DISABLE_PULLUP_H VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM118 VDDIO DISABLE_PULLUP_H 71 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM119 VDDIO 43 29 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 sa=250002 sb=250000 a=2.5 p=11
XM120 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM121 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM122 43 71 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM123 VDDIO 71 43 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM124 71 DISABLE_PULLUP_H VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM125 VDDIO DISABLE_PULLUP_H 71 VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM126 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM127 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM128 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM129 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 sa=300000 sb=300003 a=0.6 p=3.2
XM130 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM131 VDDIO 27 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM132 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM133 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300001 sb=300002 a=0.6 p=3.2
XM134 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM135 XRES_H_N 72 VDDIO_Q VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 sa=300002 sb=300001 a=0.6 p=3.2
XM136 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM137 VDDIO_Q 72 XRES_H_N VDDIO_Q sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 sa=300003 sb=300000 a=0.6 p=3.2
XM138 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM139 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM140 VDDIO 46 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM141 VDDIO 46 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM142 PAD 46 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM143 PAD 46 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM144 VDDIO 46 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM145 VDDIO 46 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM146 PAD 47 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM147 PAD 47 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM148 VDDIO 47 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM149 VDDIO 47 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300020 a=3 p=11.2
XM150 PAD 47 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300018 a=3 p=11.2
XM151 PAD 47 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300018 a=3 p=11.2
XM152 VDDIO 48 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300016 a=3 p=11.2
XM153 VDDIO 48 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300016 a=3 p=11.2
XM154 PAD 48 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300013 a=3 p=11.2
XM155 PAD 48 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300013 a=3 p=11.2
XM156 VDDIO 48 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300011 a=3 p=11.2
XM157 VDDIO 48 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300011 a=3 p=11.2
XM158 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300008 a=3 p=11.2
XM159 PAD 27 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300008 a=3 p=11.2
XM160 VDDIO 49 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300006 a=3 p=11.2
XM161 VDDIO 49 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300006 a=3 p=11.2
XM162 PAD 50 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300003 a=3 p=11.2
XM163 PAD 50 VDDIO VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 sa=300020 sb=300003 a=3 p=11.2
XM164 VDDIO 50 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 sa=300020 sb=300002 a=3 p=11.2
XM165 VDDIO 50 PAD VDDIO sky130_fd_pr__pfet_g5v0d10v5 L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 sa=300020 sb=300002 a=3 p=11.2
X166 VSSD 56 sky130_fd_pr__diode_pw2nd_11v0 a=156.97 p=1082.84 m=1
X167 VSSD 51 sky130_fd_pr__diode_pw2nd_11v0 a=156.981 p=1082.92 m=1
X168 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=16.2631 p=16.27 m=1
X169 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw a=15.5 p=17.4 m=1
X170 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=96.7627 p=49.03 m=1
X171 VSSD 24 sky130_fd_pr__model__parasitic__diode_ps2nw a=23.8226 p=21.54 m=1
X172 VSSD 25 sky130_fd_pr__model__parasitic__diode_ps2nw a=21.9076 p=21.04 m=1
X173 VSSD VCCHIB sky130_fd_pr__model__parasitic__diode_ps2nw a=4.2823 p=8.33 m=1
X174 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=108.48 p=83.5 m=1
X175 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=40.2643 p=30.01 m=1
X176 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=32.0172 p=25.17 m=1
X177 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=36.4812 p=24.46 m=1
X178 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=15.7043 p=15.95 m=1
X179 VSSD VDDIO_Q sky130_fd_pr__model__parasitic__diode_ps2nw a=16.8897 p=16.63 m=1
X180 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=1473.41 p=184.25 m=1
X181 VSSD VDDIO sky130_fd_pr__model__parasitic__diode_ps2nw a=735.037 p=170.75 m=1
R182 56 51 sky130_fd_pr__res_generic_nd__hv L=1077.19 W=0.29 m=1
R183 28 29 sky130_fd_pr__res_generic_po L=50 W=0.8 m=1
R184 VDDIO 38 sky130_fd_pr__res_generic_po L=50 W=0.8 m=1
R185 45 26 sky130_fd_pr__res_generic_po L=713.695 W=0.4 m=1
R186 65 91 0.01 short m=1
R187 91 67 0.01 short m=1
R188 67 93 0.01 short m=1
R189 94 70 0.01 short m=1
R190 73 97 0.01 short m=1
R191 98 74 0.01 short m=1
X192 27 46 sky130_fd_io__tk_em2o_cdns_55959141808653
X193 27 46 sky130_fd_io__tk_em2o_cdns_55959141808653
X194 27 47 sky130_fd_io__tk_em2o_cdns_55959141808653
X195 27 47 sky130_fd_io__tk_em2o_cdns_55959141808653
X196 27 48 sky130_fd_io__tk_em2o_cdns_55959141808653
X197 27 48 sky130_fd_io__tk_em2o_cdns_55959141808653
X198 27 49 sky130_fd_io__tk_em2o_cdns_55959141808653
X199 27 49 sky130_fd_io__tk_em2o_cdns_55959141808653
X200 27 50 sky130_fd_io__tk_em2o_cdns_55959141808653
X201 27 50 sky130_fd_io__tk_em2o_cdns_55959141808653
X210 27 46 sky130_fd_io__tk_em2s_cdns_55959141808652
X211 27 47 sky130_fd_io__tk_em2s_cdns_55959141808652
X212 27 48 sky130_fd_io__tk_em2s_cdns_55959141808652
X213 27 49 sky130_fd_io__tk_em2s_cdns_55959141808652
X214 27 50 sky130_fd_io__tk_em2s_cdns_55959141808652
X241 27 VDDIO sky130_fd_pr__res_generic_po__example_5595914180838
X242 66 PULLUP_H sky130_fd_pr__res_generic_po__example_5595914180864
X243 68 66 sky130_fd_pr__res_generic_po__example_5595914180864
X244 69 68 sky130_fd_pr__res_generic_po__example_5595914180864
X245 65 69 sky130_fd_pr__res_generic_po__example_5595914180864
X246 78 75 sky130_fd_pr__res_generic_po__example_5595914180864
X247 76 77 sky130_fd_pr__res_generic_po__example_5595914180864
X248 79 78 sky130_fd_pr__res_generic_po__example_5595914180864
X249 77 79 sky130_fd_pr__res_generic_po__example_5595914180864
X250 66 PULLUP_H sky130_fd_io__tk_em1s_cdns_5595914180859
X251 68 66 sky130_fd_io__tk_em1s_cdns_5595914180859
X252 69 68 sky130_fd_io__tk_em1s_cdns_5595914180859
X253 65 69 sky130_fd_io__tk_em1s_cdns_5595914180859
X254 74 76 sky130_fd_io__tk_em1s_cdns_5595914180859
X255 78 75 sky130_fd_io__tk_em1s_cdns_5595914180859
X256 76 77 sky130_fd_io__tk_em1s_cdns_5595914180859
X257 77 79 sky130_fd_io__tk_em1s_cdns_5595914180859
X258 79 78 sky130_fd_io__tk_em1s_cdns_5595914180859
X259 PAD PAD_A_ESD_H sky130_fd_io__res250only_small
X260 TIE_WEAK_HI_H 75 sky130_fd_io__res250only_small
X261 67 65 sky130_fd_pr__res_bent_po__example_5595914180862
X262 70 67 sky130_fd_pr__res_bent_po__example_5595914180862
X263 74 73 sky130_fd_pr__res_bent_po__example_5595914180862
X264 76 74 sky130_fd_pr__res_bent_po__example_5595914180862
X265 70 28 sky130_fd_pr__res_bent_po__example_5595914180863
X266 73 38 sky130_fd_pr__res_bent_po__example_5595914180863
X269 VSSD VDDIO_Q 80 42 81 82 83 84 85 86 87 88 89 92 sky130_fd_io__xres2v2_rcfilter_lpfv2
X301 VDDIO_Q INP_SEL_H 52 92 sky130_fd_pr__pfet_01v8__example_55959141808767
X302 VDDIO_Q 40 92 FILT_IN_H sky130_fd_pr__pfet_01v8__example_55959141808767
X303 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd
X304 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd
X305 VSSD 40 52 92 sky130_fd_pr__nfet_01v8__example_55959141808764
X306 VSSD INP_SEL_H 92 FILT_IN_H sky130_fd_pr__nfet_01v8__example_55959141808764
X307 VSSD 30 64 58 sky130_fd_pr__nfet_01v8__example_55959141808779
X308 VSSD 35 59 25 sky130_fd_pr__nfet_01v8__example_55959141808779
X309 VSSD 32 31 sky130_fd_pr__nfet_01v8__example_55959141808777
X310 VSSD 37 39 sky130_fd_pr__nfet_01v8__example_55959141808777
X311 VSSD ENABLE_H 55 sky130_fd_pr__nfet_01v8__example_55959141808777
X327 24 24 24 sky130_fd_pr__pfet_01v8__example_55959141808784
X328 24 30 37 sky130_fd_pr__pfet_01v8__example_55959141808784
X348 VSSD VDDIO VSSD 30 PAD sky130_fd_io__gpio_buf_localesdv2
X351 VSSD 99 VSSIO VDDIO 99 99 90 PAD sky130_fd_io__gpio_pddrvr_strong_xres4v2
.ENDS
***************************************
.SUBCKT ICV_2 VSSD VSSIO VCCD VDDIO VSSD_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSD VCCD VDDIO VCCD VSSIO VSSD VSSD_PAD sky130_fd_io__top_ground_lvc_wpad
.ENDS
***************************************
.SUBCKT ICV_3 VSSD VSSIO VCCD VDDIO VCCD_PAD
**
*.CALIBRE ISOLATED NETS: VCCHIB VDDA VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VDDIO_Q
X0 VSSD VSSD VSSD VCCD VDDIO VCCD VSSIO VCCD VCCD_PAD sky130_fd_io__top_power_lvc_wpad
.ENDS
***************************************
.SUBCKT chip_io   mprj_io_oeb[24] mprj_io_ib_mode_sel[24] mprj_io_vtrip_sel[24] mprj_io_out[24] mprj_io_holdover[24] mprj_io_dm[74] mprj_io_analog_sel[24] mprj_io_hldh_n[24] mprj_io_enh[24] mprj_io_inp_dis[24] mprj_io_analog_pol[24] mprj_io_dm[72] mprj_io_analog_en[24] mprj_io_dm[73] mprj_analog_io[17] mprj_io_slow_sel[24] mprj_io_in[24] porb_h mprj_io_oeb[23] mprj_io_ib_mode_sel[23]
+ mprj_io_vtrip_sel[23] mprj_io_out[23] mprj_io_holdover[23] mprj_io_dm[71] mprj_io_analog_sel[23] mprj_io_hldh_n[23] mprj_io_enh[23] mprj_io_inp_dis[23] mprj_io_analog_pol[23] mprj_io_dm[69] mprj_io_analog_en[23] mprj_io_dm[70] mprj_analog_io[16] mprj_io_slow_sel[23] mprj_io_in[23] mprj_io_oeb[22] mprj_io_ib_mode_sel[22] mprj_io_vtrip_sel[22] mprj_io_out[22] mprj_io_holdover[22]
+ mprj_io_dm[68] mprj_io_analog_sel[22] mprj_io_hldh_n[22] mprj_io_enh[22] mprj_io_inp_dis[22] mprj_io_analog_pol[22] mprj_io_dm[66] mprj_io_analog_en[22] mprj_io_dm[67] mprj_analog_io[15] mprj_io_slow_sel[22] mprj_io_in[22] mprj_io_oeb[21] mprj_io_ib_mode_sel[21] mprj_io_vtrip_sel[21] mprj_io_out[21] mprj_io_holdover[21] mprj_io_dm[65] mprj_io_analog_sel[21] mprj_io_hldh_n[21]
+ mprj_io_enh[21] mprj_io_inp_dis[21] mprj_io_analog_pol[21] mprj_io_dm[63] mprj_io_analog_en[21] mprj_io_dm[64] mprj_analog_io[14] mprj_io_slow_sel[21] mprj_io_in[21] mprj_io_oeb[20] mprj_io_ib_mode_sel[20] mprj_io_vtrip_sel[20] mprj_io_out[20] mprj_io_holdover[20] mprj_io_dm[62] mprj_io_analog_sel[20] mprj_io_hldh_n[20] mprj_io_enh[20] mprj_io_inp_dis[20] mprj_io_analog_pol[20]
+ mprj_io_dm[60] mprj_io_analog_en[20] mprj_io_dm[61] mprj_analog_io[13] mprj_io_slow_sel[20] mprj_io_in[20] mprj_io_oeb[19] mprj_io_ib_mode_sel[19] mprj_io_vtrip_sel[19] mprj_io_out[19] mprj_io_holdover[19] mprj_io_dm[59] mprj_io_analog_sel[19] mprj_io_hldh_n[19] mprj_io_enh[19] mprj_io_inp_dis[19] mprj_io_analog_pol[19] mprj_io_dm[57] mprj_io_analog_en[19] mprj_io_dm[58]
+ mprj_analog_io[12] mprj_io_slow_sel[19] mprj_io_in[19] mprj_io_oeb[18] mprj_io_ib_mode_sel[18] mprj_io_vtrip_sel[18] mprj_io_out[18] mprj_io_holdover[18] mprj_io_dm[56] mprj_io_analog_sel[18] mprj_io_hldh_n[18] mprj_io_enh[18] mprj_io_inp_dis[18] mprj_io_analog_pol[18] mprj_io_dm[54] mprj_io_analog_en[18] mprj_io_dm[55] mprj_analog_io[11] mprj_io_slow_sel[18] mprj_io_in[18]
+ mprj_io_oeb[17] mprj_io_ib_mode_sel[17] mprj_io_vtrip_sel[17] mprj_io_out[17] mprj_io_holdover[17] mprj_io_dm[53] mprj_io_analog_sel[17] mprj_io_hldh_n[17] mprj_io_enh[17] mprj_io_inp_dis[17] mprj_io_analog_pol[17] mprj_io_dm[51] mprj_io_analog_en[17] mprj_io_dm[52] mprj_analog_io[10] mprj_io_slow_sel[17] mprj_io_in[17] mprj_io_oeb[16] mprj_io_ib_mode_sel[16] mprj_io_vtrip_sel[16]
+ mprj_io_out[16] mprj_io_holdover[16] mprj_io_dm[50] mprj_io_analog_sel[16] mprj_io_hldh_n[16] mprj_io_enh[16] mprj_io_inp_dis[16] mprj_io_analog_pol[16] mprj_io_dm[48] mprj_io_analog_en[16] mprj_io_dm[49] mprj_analog_io[9] mprj_io_slow_sel[16] mprj_io_in[16] mprj_io_oeb[15] mprj_io_ib_mode_sel[15] mprj_io_vtrip_sel[15] mprj_io_out[15] mprj_io_holdover[15] mprj_io_dm[47]
+ mprj_io_analog_sel[15] mprj_io_hldh_n[15] mprj_io_enh[15] mprj_io_inp_dis[15] mprj_io_analog_pol[15] mprj_io_dm[45] mprj_io_analog_en[15] mprj_io_dm[46] mprj_analog_io[8] mprj_io_slow_sel[15] mprj_io_in[15] mprj_io_in[14] mprj_io_slow_sel[14] mprj_analog_io[7] mprj_io_dm[43] mprj_io_analog_en[14] mprj_io_dm[42] mprj_io_analog_pol[14] mprj_io_inp_dis[14] mprj_io_enh[14]
+ mprj_io_hldh_n[14] mprj_io_analog_sel[14] mprj_io_dm[44] mprj_io_holdover[14] mprj_io_out[14] mprj_io_vtrip_sel[14] mprj_io_ib_mode_sel[14] mprj_io_oeb[14] mprj_io_in[13] mprj_io_slow_sel[13] mprj_analog_io[6] mprj_io_dm[40] mprj_io_analog_en[13] mprj_io_dm[39] mprj_io_analog_pol[13] mprj_io_inp_dis[13] mprj_io_enh[13] mprj_io_hldh_n[13] mprj_io_analog_sel[13] mprj_io_dm[41]
+ mprj_io_holdover[13] mprj_io_out[13] mprj_io_vtrip_sel[13] mprj_io_ib_mode_sel[13] mprj_io_oeb[13] mprj_io_oeb[31] mprj_io_ib_mode_sel[31] mprj_io_vtrip_sel[31] mprj_io_out[31] mprj_io_holdover[31] mprj_io_dm[95] mprj_io_analog_sel[31] mprj_io_hldh_n[31] mprj_io_enh[31] mprj_io_inp_dis[31] mprj_io_analog_pol[31] mprj_io_dm[93] mprj_io_analog_en[31] mprj_io_dm[94] mprj_analog_io[24]
+ mprj_io_slow_sel[31] mprj_io_in[31] mprj_io_oeb[30] mprj_io_ib_mode_sel[30] mprj_io_vtrip_sel[30] mprj_io_out[30] mprj_io_holdover[30] mprj_io_dm[92] mprj_io_analog_sel[30] mprj_io_hldh_n[30] mprj_io_enh[30] mprj_io_inp_dis[30] mprj_io_analog_pol[30] mprj_io_dm[90] mprj_io_analog_en[30] mprj_io_dm[91] mprj_analog_io[23] mprj_io_slow_sel[30] mprj_io_in[30] mprj_io_oeb[29]
+ mprj_io_ib_mode_sel[29] mprj_io_vtrip_sel[29] mprj_io_out[29] mprj_io_holdover[29] mprj_io_dm[89] mprj_io_analog_sel[29] mprj_io_hldh_n[29] mprj_io_enh[29] mprj_io_inp_dis[29] mprj_io_analog_pol[29] mprj_io_dm[87] mprj_io_analog_en[29] mprj_io_dm[88] mprj_analog_io[22] mprj_io_slow_sel[29] mprj_io_in[29] mprj_io_oeb[28] mprj_io_ib_mode_sel[28] mprj_io_vtrip_sel[28] mprj_io_out[28]
+ mprj_io_holdover[28] mprj_io_dm[86] mprj_io_analog_sel[28] mprj_io_hldh_n[28] mprj_io_enh[28] mprj_io_inp_dis[28] mprj_io_analog_pol[28] mprj_io_dm[84] mprj_io_analog_en[28] mprj_io_dm[85] mprj_analog_io[21] mprj_io_slow_sel[28] mprj_io_in[28] mprj_io_oeb[27] mprj_io_ib_mode_sel[27] mprj_io_vtrip_sel[27] mprj_io_out[27] mprj_io_holdover[27] mprj_io_dm[83] mprj_io_analog_sel[27]
+ mprj_io_hldh_n[27] mprj_io_enh[27] mprj_io_inp_dis[27] mprj_io_analog_pol[27] mprj_io_dm[81] mprj_io_analog_en[27] mprj_io_dm[82] mprj_analog_io[20] mprj_io_slow_sel[27] mprj_io_in[27] mprj_io_oeb[26] mprj_io_ib_mode_sel[26] mprj_io_vtrip_sel[26] mprj_io_out[26] mprj_io_holdover[26] mprj_io_dm[80] mprj_io_analog_sel[26] mprj_io_hldh_n[26] mprj_io_enh[26] mprj_io_inp_dis[26]
+ mprj_io_analog_pol[26] mprj_io_dm[78] mprj_io_analog_en[26] mprj_io_dm[79] mprj_analog_io[19] mprj_io_slow_sel[26] mprj_io_in[26] mprj_io_oeb[25] mprj_io_ib_mode_sel[25] mprj_io_vtrip_sel[25] mprj_io_out[25] mprj_io_holdover[25] mprj_io_dm[77] mprj_io_analog_sel[25] mprj_io_hldh_n[25] mprj_io_enh[25] mprj_io_inp_dis[25] mprj_io_analog_pol[25] mprj_io_dm[75] mprj_io_analog_en[25]
+ mprj_io_dm[76] mprj_analog_io[18] mprj_io_slow_sel[25] mprj_io_in[25] mprj_io_in[7] mprj_io_slow_sel[7] mprj_analog_io[0] mprj_io_dm[22] mprj_io_analog_en[7] mprj_io_dm[21] mprj_io_analog_pol[7] mprj_io_inp_dis[7] mprj_io_enh[7] mprj_io_hldh_n[7] mprj_io_analog_sel[7] mprj_io_dm[23] mprj_io_holdover[7] mprj_io_out[7] mprj_io_vtrip_sel[7] mprj_io_ib_mode_sel[7]
+ mprj_io_oeb[7] mprj_io_in[8] mprj_io_slow_sel[8] mprj_analog_io[1] mprj_io_dm[25] mprj_io_analog_en[8] mprj_io_dm[24] mprj_io_analog_pol[8] mprj_io_inp_dis[8] mprj_io_enh[8] mprj_io_hldh_n[8] mprj_io_analog_sel[8] mprj_io_dm[26] mprj_io_holdover[8] mprj_io_out[8] mprj_io_vtrip_sel[8] mprj_io_ib_mode_sel[8] mprj_io_oeb[8] mprj_io_in[9] mprj_io_slow_sel[9]
+ mprj_analog_io[2] mprj_io_dm[28] mprj_io_analog_en[9] mprj_io_dm[27] mprj_io_analog_pol[9] mprj_io_inp_dis[9] mprj_io_enh[9] mprj_io_hldh_n[9] mprj_io_analog_sel[9] mprj_io_dm[29] mprj_io_holdover[9] mprj_io_out[9] mprj_io_vtrip_sel[9] mprj_io_ib_mode_sel[9] mprj_io_oeb[9] mprj_io_in[10] mprj_io_slow_sel[10] mprj_analog_io[3] mprj_io_dm[31] mprj_io_analog_en[10]
+ mprj_io_dm[30] mprj_io_analog_pol[10] mprj_io_inp_dis[10] mprj_io_enh[10] mprj_io_hldh_n[10] mprj_io_analog_sel[10] mprj_io_dm[32] mprj_io_holdover[10] mprj_io_out[10] mprj_io_vtrip_sel[10] mprj_io_ib_mode_sel[10] mprj_io_oeb[10] mprj_io_in[11] mprj_io_slow_sel[11] mprj_analog_io[4] mprj_io_dm[34] mprj_io_analog_en[11] mprj_io_dm[33] mprj_io_analog_pol[11] mprj_io_inp_dis[11]
+ mprj_io_enh[11] mprj_io_hldh_n[11] mprj_io_analog_sel[11] mprj_io_dm[35] mprj_io_holdover[11] mprj_io_out[11] mprj_io_vtrip_sel[11] mprj_io_ib_mode_sel[11] mprj_io_oeb[11] mprj_io_in[12] mprj_io_slow_sel[12] mprj_analog_io[5] mprj_io_dm[37] mprj_io_analog_en[12] mprj_io_dm[36] mprj_io_analog_pol[12] mprj_io_inp_dis[12] mprj_io_enh[12] mprj_io_hldh_n[12] mprj_io_analog_sel[12]
+ mprj_io_dm[38] mprj_io_holdover[12] mprj_io_out[12] mprj_io_vtrip_sel[12] mprj_io_ib_mode_sel[12] mprj_io_oeb[12] mprj_io_oeb[37] mprj_io_ib_mode_sel[37] mprj_io_vtrip_sel[37] mprj_io_out[37] mprj_io_holdover[37] mprj_io_dm[113] mprj_io_analog_sel[37] mprj_io_hldh_n[37] mprj_io_enh[37] mprj_io_inp_dis[37] mprj_io_analog_pol[37] mprj_io_dm[111] mprj_io_analog_en[37] mprj_io_dm[112]
+ mprj_io_slow_sel[37] mprj_io_in[37] mprj_io_oeb[36] mprj_io_ib_mode_sel[36] mprj_io_vtrip_sel[36] mprj_io_out[36] mprj_io_holdover[36] mprj_io_dm[110] mprj_io_analog_sel[36] mprj_io_hldh_n[36] mprj_io_enh[36] mprj_io_inp_dis[36] mprj_io_analog_pol[36] mprj_io_dm[108] mprj_io_analog_en[36] mprj_io_dm[109] mprj_io_slow_sel[36] mprj_io_in[36] mprj_io_oeb[35] mprj_io_ib_mode_sel[35]
+ mprj_io_vtrip_sel[35] mprj_io_out[35] mprj_io_holdover[35] mprj_io_dm[107] mprj_io_analog_sel[35] mprj_io_hldh_n[35] mprj_io_enh[35] mprj_io_inp_dis[35] mprj_io_analog_pol[35] mprj_io_dm[105] mprj_io_analog_en[35] mprj_io_dm[106] mprj_analog_io[28] mprj_io_slow_sel[35] mprj_io_in[35] mprj_io_oeb[34] mprj_io_ib_mode_sel[34] mprj_io_vtrip_sel[34] mprj_io_out[34] mprj_io_holdover[34]
+ mprj_io_dm[104] mprj_io_analog_sel[34] mprj_io_hldh_n[34] mprj_io_enh[34] mprj_io_inp_dis[34] mprj_io_analog_pol[34] mprj_io_dm[102] mprj_io_analog_en[34] mprj_io_dm[103] mprj_analog_io[27] mprj_io_slow_sel[34] mprj_io_in[34] mprj_io_oeb[33] mprj_io_ib_mode_sel[33] mprj_io_vtrip_sel[33] mprj_io_out[33] mprj_io_holdover[33] mprj_io_dm[101] mprj_io_analog_sel[33] mprj_io_hldh_n[33]
+ mprj_io_enh[33] mprj_io_inp_dis[33] mprj_io_analog_pol[33] mprj_io_dm[99] mprj_io_analog_en[33] mprj_io_dm[100] mprj_analog_io[26] mprj_io_slow_sel[33] mprj_io_in[33] mprj_io_oeb[32] mprj_io_ib_mode_sel[32] mprj_io_vtrip_sel[32] mprj_io_out[32] mprj_io_holdover[32] mprj_io_dm[98] mprj_io_analog_sel[32] mprj_io_hldh_n[32] mprj_io_enh[32] mprj_io_inp_dis[32] mprj_io_analog_pol[32]
+ mprj_io_dm[96] mprj_io_analog_en[32] mprj_io_dm[97] mprj_analog_io[25] mprj_io_slow_sel[32] mprj_io_in[32] mprj_io_in[0] mprj_io_slow_sel[0] mprj_io_dm[1] mprj_io_analog_en[0] mprj_io_dm[0] mprj_io_analog_pol[0] mprj_io_inp_dis[0] mprj_io_enh[0] mprj_io_hldh_n[0] mprj_io_analog_sel[0] mprj_io_dm[2] mprj_io_holdover[0] mprj_io_out[0] mprj_io_vtrip_sel[0]
+ mprj_io_ib_mode_sel[0] mprj_io_oeb[0] mprj_io_in[1] mprj_io_slow_sel[1] mprj_io_dm[4] mprj_io_analog_en[1] mprj_io_dm[3] mprj_io_analog_pol[1] mprj_io_inp_dis[1] mprj_io_enh[1] mprj_io_hldh_n[1] mprj_io_analog_sel[1] mprj_io_dm[5] mprj_io_holdover[1] mprj_io_out[1] mprj_io_vtrip_sel[1] mprj_io_ib_mode_sel[1] mprj_io_oeb[1] mprj_io_in[2] mprj_io_slow_sel[2]
+ mprj_io_dm[7] mprj_io_analog_en[2] mprj_io_dm[6] mprj_io_analog_pol[2] mprj_io_inp_dis[2] mprj_io_enh[2] mprj_io_hldh_n[2] mprj_io_analog_sel[2] mprj_io_dm[8] mprj_io_holdover[2] mprj_io_out[2] mprj_io_vtrip_sel[2] mprj_io_ib_mode_sel[2] mprj_io_oeb[2] mprj_io_in[3] mprj_io_slow_sel[3] mprj_io_dm[10] mprj_io_analog_en[3] mprj_io_dm[9] mprj_io_analog_pol[3]
+ mprj_io_inp_dis[3] mprj_io_enh[3] mprj_io_hldh_n[3] mprj_io_analog_sel[3] mprj_io_dm[11] mprj_io_holdover[3] mprj_io_out[3] mprj_io_vtrip_sel[3] mprj_io_ib_mode_sel[3] mprj_io_oeb[3] mprj_io_in[4] mprj_io_slow_sel[4] mprj_io_dm[13] mprj_io_analog_en[4] mprj_io_dm[12] mprj_io_analog_pol[4] mprj_io_inp_dis[4] mprj_io_enh[4] mprj_io_hldh_n[4] mprj_io_analog_sel[4]
+ mprj_io_dm[14] mprj_io_holdover[4] mprj_io_out[4] mprj_io_vtrip_sel[4] mprj_io_ib_mode_sel[4] mprj_io_oeb[4] mprj_io_in[5] mprj_io_slow_sel[5] mprj_io_dm[16] mprj_io_analog_en[5] mprj_io_dm[15] mprj_io_analog_pol[5] mprj_io_inp_dis[5] mprj_io_enh[5] mprj_io_hldh_n[5] mprj_io_analog_sel[5] mprj_io_dm[17] mprj_io_holdover[5] mprj_io_out[5] mprj_io_vtrip_sel[5]
+ mprj_io_ib_mode_sel[5] mprj_io_oeb[5] mprj_io_in[6] mprj_io_slow_sel[6] mprj_io_dm[19] mprj_io_analog_en[6] mprj_io_dm[18] mprj_io_analog_pol[6] mprj_io_inp_dis[6] mprj_io_enh[6] mprj_io_hldh_n[6] mprj_io_analog_sel[6] mprj_io_dm[20] mprj_io_holdover[6] mprj_io_out[6] mprj_io_vtrip_sel[6] mprj_io_ib_mode_sel[6] mprj_io_oeb[6] clock_core por
+ flash_csb_ieb_core flash_csb_core flash_csb_oeb_core flash_clk_ieb_core flash_clk_core flash_clk_oeb_core flash_io0_di_core flash_io0_ieb_core flash_io0_do_core flash_io0_oeb_core flash_io1_di_core flash_io1_ieb_core flash_io1_do_core flash_io1_oeb_core gpio_in_core gpio_mode0_core gpio_inenb_core gpio_mode1_core gpio_out_core gpio_outenb_core
+ resetb_core_h mprj_io[24] vccd2_pad mprj_io[23] mprj_io[22] mprj_io[21] mprj_io[20] mprj_io[19] vssio_pad mprj_io[18] mprj_io[17] mprj_io[16] vssa1_pad mprj_io[15] vccd1_pad mprj_io[14] mprj_io[13] mprj_io[31] mprj_io[30] mprj_io[29]
+ mprj_io[28] mprj_io[27] mprj_io[26] mprj_io[25] vssa2_pad vdda1_pad mprj_io[7] mprj_io[8] mprj_io[9] mprj_io[10] mprj_io[11] mprj_io[12] vssd2_pad vdda2_pad vssd1_pad mprj_io[37] mprj_io[36] mprj_io[35] mprj_io[34] mprj_io[33]
+ mprj_io[32] vddio_pad mprj_io[0] mprj_io[1] mprj_io[2] mprj_io[3] mprj_io[4] mprj_io[5] mprj_io[6] vssa_pad clock flash_csb flash_clk flash_io0 flash_io1 gpio vdda_pad resetb vssd_pad vccd_pad
**
X0 1 193 sky130_fd_pr__model__parasitic__diode_ps2nw a=57.3765 p=0 m=1
X1 1 2 175 669 193 673 330 674 vccd2_pad vssio_pad vssa1_pad vccd1_pad ICV_13
X2 1 2 193 ICV_14
X3 1 330 193 175 669 672 vssa2_pad vdda1_pad ICV_15
X4 1 330 2 193 175 672 669 673 674 vssd2_pad vdda2_pad vssd1_pad ICV_16
X5 1 2 175 193 330 vddio_pad ICV_17
X6 1 2 193 675 676 vssa_pad vdda_pad ICV_18
X7 1 193 174 193 porb_h 2 2 174 resetb 2 2 645 2 2 resetb_core_h 645 ICV_1
X8 1 2 174 193 vssd_pad ICV_2
X9 1 2 174 193 vccd_pad ICV_3
.ENDS
***************************************
