*---------------------------------------------------------------------------
* SPDX-FileCopyrightText: 2020 Efabless Corporation
* Licensed under the Apache License, Version 2.0 (the "License");
* you may not use this file except in compliance with the License.
* You may obtain a copy of the License at
*
*     https://www.apache.org/licenses/LICENSE-2.0
*
* Unless required by applicable law or agreed to in writing, software
* distributed under the License is distributed on an "AS IS" BASIS,
* WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
* See the License for the specific language governing permissions and
* limitations under the License.
*
* SPDX-License-Identifier: Apache-2.0
*---------------------------------------------------------------------------
* All-digital Frequency-locked loop
*---------------------------------------------------------------------------
* To make this simulatable, the circuit is broken into the ring oscillator
* and controller, separately, with the controller converted into an xspice
* model.
*
* For simplicity, the DCO mode has been removed, so no external trim with
* multiplexer.  Also no multiplexer on the internal reset.
*---------------------------------------------------------------------------

.include "digital_pll_controller.xspice"
.include "ring_osc2x13.spice"

.subckt digital_pll vdd vss reset osc clockp1 clockp0 div4 div3 div2 div1 div0

X0 vdd vss clockp0 div0 div1 div2 div3 div4 osc reset trim0 trim1 trim2 trim3
+ trim4 trim5 trim6 trim7 trim8 trim9 trim10 trim11 trim12 trim13 trim14
+ trim15 trim16 trim17 trim18 trim19 trim20 trim21 trim22 trim23 trim24
+ trim25 digital_pll_controller

X1 vdd vss clockp0 clockp1 reset trim0 trim1 trim2 trim3 trim4 trim5 trim6 trim7
+ trim8 trim9 trim10 trim11 trim12 trim13 trim14 trim15 trim16 trim17 trim18
+ trim19 trim20 trim21 trim22 trim23 trim24 trim25 ring_osc2x13

.ends


