* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2o_cdns_55959141808653 2 3
** N=7 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=260 $Y=0 $D=283
R1 7 3 0.01 m=1 $[short] $X=1770 $Y=0 $D=283
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808202
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808657
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em2s_cdns_55959141808652 2 3
** N=6 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=260 $Y=0 $D=283
R1 6 3 0.01 m=1 $[short] $X=1770 $Y=0 $D=283
.ENDS
***************************************
.SUBCKT ICV_1
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180838 2 3
** N=6 EP=2 IP=0 FDC=1
R0 2 3 L=10.2 W=0.5 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_po__example_5595914180864 2 3
** N=8 EP=2 IP=0 FDC=1
R0 2 3 L=1.5 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_em1s_cdns_5595914180859 2 3
** N=6 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=260 $Y=0 $D=282
R1 6 3 0.01 m=1 $[short] $X=1770 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__res250only_small PAD ROUT
** N=32 EP=2 IP=0 FDC=7
R0 PAD 6 L=0.17 W=2 m=1 mult=1 model="mrp1" $[mrp1] $X=300 $Y=10 $D=257
R1 6 7 L=10.07 W=2 m=1 mult=1 model="mrp1" $[mrp1] $X=640 $Y=10 $D=257
R2 7 ROUT L=0.17 W=2 m=1 mult=1 model="mrp1" $[mrp1] $X=10880 $Y=10 $D=257
R3 PAD 6 0.01 m=1 $[short] $X=380 $Y=0 $D=281
R4 7 ROUT 0.01 m=1 $[short] $X=10960 $Y=0 $D=281
R5 PAD 6 0.01 m=1 $[short] $X=380 $Y=5 $D=282
R6 7 ROUT 0.01 m=1 $[short] $X=10960 $Y=5 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180862 2 3
** N=8 EP=2 IP=0 FDC=1
R0 2 3 L=6 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_bent_po__example_5595914180863 2 3
** N=8 EP=2 IP=0 FDC=1
R0 2 3 L=12 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=0 $Y=0 $D=257
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808616
** N=39 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x4
** N=74 EP=0 IP=44 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: IN OUT
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 2 3
** N=7 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=130 $Y=0 $D=282
R1 7 3 0.01 m=1 $[short] $X=280 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_p_em1c_cdns_55959141808753 2
** N=6 EP=1 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 2 6 0.01 m=1 $[short] $X=160 $Y=250 $D=282
.ENDS
***************************************
.SUBCKT ICV_2 2 3
** N=7 EP=2 IP=9 FDC=4
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=0 0 0 0 $X=0 $Y=0
X1 2 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=-10 -770 0 0 $X=-10 $Y=-770
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808754 2 3
** N=5 EP=2 IP=0 FDC=1
*.SEEDPROM
R0 2 3 L=14 W=0.5 m=1 $[mrdn] $X=0 $Y=0 $D=253
.ENDS
***************************************
.SUBCKT ICV_3 2 3 4 5
** N=9 EP=4 IP=10 FDC=2
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=14000 -770 1 180 $X=-340 $Y=-900
X1 4 5 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=0 0 0 0 $X=-340 $Y=-130
.ENDS
***************************************
.SUBCKT ICV_4 2 3 4 5 6 7 8 9
** N=17 EP=8 IP=18 FDC=4
*.SEEDPROM
X0 4 2 3 5 ICV_3 $T=0 -1540 0 0 $X=-340 $Y=-2440
X1 8 6 7 9 ICV_3 $T=0 0 0 0 $X=-340 $Y=-900
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 2 3
** N=7 EP=2 IP=0 FDC=2
R0 2 6 0.01 m=1 $[short] $X=130 $Y=0 $D=282
R1 7 3 0.01 m=1 $[short] $X=280 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 2
** N=6 EP=1 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 2 6 0.01 m=1 $[short] $X=160 $Y=640 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 2
** N=6 EP=1 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 2 6 0.01 m=1 $[short] $X=160 $Y=250 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808700
** N=21 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_55959141808338
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808559
** N=21 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808666
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808337
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__via_pol1__example_55959141808273
** N=13 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_5
** N=3 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT ICV_6
** N=5 EP=0 IP=6 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 1
** N=5 EP=1 IP=0 FDC=2
R0 1 4 0.01 m=1 $[short] $X=160 $Y=0 $D=282
R1 1 5 0.01 m=1 $[short] $X=160 $Y=280 $D=282
.ENDS
***************************************
.SUBCKT ICV_7 2 3 4
** N=8 EP=3 IP=9 FDC=4
X0 2 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=0 0 0 0 $X=0 $Y=0
X1 4 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=-10 770 0 0 $X=-10 $Y=770
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 1 2
** N=6 EP=2 IP=0 FDC=2
R0 2 5 0.01 m=1 $[short] $X=130 $Y=0 $D=282
R1 6 1 0.01 m=1 $[short] $X=280 $Y=0 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__res_generic_nd__example_55959141808755 2 3
** N=5 EP=2 IP=0 FDC=1
*.SEEDPROM
R0 2 3 L=47 W=0.5 m=1 $[mrdn] $X=0 $Y=0 $D=253
.ENDS
***************************************
.SUBCKT ICV_8 2 3 4
** N=8 EP=3 IP=10 FDC=2
*.SEEDPROM
X0 2 3 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=0 0 0 0 $X=-340 $Y=-130
X1 4 2 sky130_fd_pr__res_generic_nd__example_55959141808755 $T=-47510 0 0 0 $X=-47850 $Y=-130
.ENDS
***************************************
.SUBCKT ICV_9 2 3
** N=7 EP=2 IP=10 FDC=2
*.SEEDPROM
X0 2 2 sky130_fd_pr__res_generic_nd__example_55959141808754 $T=0 0 0 0 $X=-340 $Y=-130
X1 2 3 sky130_fd_pr__res_generic_nd__example_55959141808755 $T=14510 0 0 0 $X=14170 $Y=-130
.ENDS
***************************************
.SUBCKT ICV_10 2 3 4 5 6
** N=14 EP=5 IP=15 FDC=4
*.SEEDPROM
X0 3 4 2 ICV_8 $T=0 0 0 0 $X=-47850 $Y=-130
X1 5 6 ICV_9 $T=14000 770 1 180 $X=-47850 $Y=640
.ENDS
***************************************
.SUBCKT ICV_11 2 3 4 5 6 7 8 9 10 11
** N=27 EP=10 IP=28 FDC=8
*.SEEDPROM
X0 2 4 6 5 3 ICV_10 $T=0 0 0 0 $X=-47850 $Y=-130
X1 7 9 11 10 8 ICV_10 $T=0 1540 0 0 $X=-47850 $Y=1410
.ENDS
***************************************
.SUBCKT sky130_fd_io__xres2v2_rcfilter_lpfv2 1 VCC_IO 3 4 5 6 7 8 9 10 11 12 13 IN
** N=5540 EP=14 IP=608 FDC=361
M0 1 3 1 1 nhv L=4 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=2725 $Y=11605 $D=49
M1 1 4 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=7005 $Y=11605 $D=49
M2 1 5 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=11285 $Y=11605 $D=49
M3 1 6 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=15565 $Y=11605 $D=49
M4 1 7 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=19845 $Y=11605 $D=49
M5 1 8 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=24125 $Y=11605 $D=49
M6 1 9 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=28405 $Y=11605 $D=49
M7 1 10 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=32685 $Y=11605 $D=49
M8 1 11 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=36965 $Y=11605 $D=49
M9 1 11 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=41245 $Y=11605 $D=49
M10 1 12 1 1 nhv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=45525 $Y=11605 $D=49
M11 1 13 1 1 nhv L=4 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=49805 $Y=11605 $D=49
M12 VCC_IO 3 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=2625 $Y=21435 $D=109
M13 VCC_IO 4 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=6905 $Y=21435 $D=109
M14 VCC_IO 5 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=11185 $Y=21435 $D=109
M15 VCC_IO 6 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00001e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=15465 $Y=21435 $D=109
M16 VCC_IO 7 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=19745 $Y=21435 $D=109
M17 VCC_IO 8 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=24025 $Y=21435 $D=109
M18 VCC_IO 9 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=28305 $Y=21435 $D=109
M19 VCC_IO 10 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00002e+06 a=28 p=22 mult=1 $X=32585 $Y=21435 $D=109
M20 VCC_IO 11 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=36865 $Y=21435 $D=109
M21 VCC_IO 11 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2.00001e+06 a=28 p=22 mult=1 $X=41145 $Y=21435 $D=109
M22 VCC_IO 12 VCC_IO VCC_IO phv L=4 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=45425 $Y=21435 $D=109
M23 VCC_IO 13 VCC_IO VCC_IO phv L=4 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=1.75 sa=2.00002e+06 sb=2e+06 a=28 p=22 mult=1 $X=49705 $Y=21435 $D=109
X24 1 8 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=815 $D=181
X25 1 7 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=2355 $D=181
X26 1 6 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=3895 $D=181
X27 1 5 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=5435 $D=181
X28 1 4 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=6975 $D=181
X29 1 3 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=8515 $D=181
X30 1 15 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=31330 $D=181
X31 1 16 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=32870 $D=181
X32 1 17 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=34410 $D=181
X33 1 18 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=35950 $D=181
X34 1 19 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=37490 $D=181
X35 1 20 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=2360 $Y=39030 $D=181
X36 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=1585 $D=181
X37 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=3125 $D=181
X38 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=4665 $D=181
X39 1 1 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=6205 $D=181
X40 1 3 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=7745 $D=181
X41 1 9 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=9285 $D=181
X42 1 15 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=30560 $D=181
X43 1 16 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=32100 $D=181
X44 1 17 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=33640 $D=181
X45 1 18 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=35180 $D=181
X46 1 19 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=36720 $D=181
X47 1 20 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=2360 $Y=38260 $D=181
X48 1 21 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=815 $D=181
X49 1 22 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=2355 $D=181
X50 1 23 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=3895 $D=181
X51 1 24 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=5435 $D=181
X52 1 25 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=6975 $D=181
X53 1 26 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=8515 $D=181
X54 1 27 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=31330 $D=181
X55 1 28 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=32870 $D=181
X56 1 29 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=34410 $D=181
X57 1 30 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=35950 $D=181
X58 1 31 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=37490 $D=181
X59 1 32 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9912 $Y=39030 $D=181
X60 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=1585 $D=181
X61 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=3125 $D=181
X62 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=4665 $D=181
X63 1 1 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=6205 $D=181
X64 1 3 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=7745 $D=181
X65 1 9 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=9285 $D=181
X66 1 15 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=30560 $D=181
X67 1 16 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=32100 $D=181
X68 1 17 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=33640 $D=181
X69 1 18 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=35180 $D=181
X70 1 19 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=36720 $D=181
X71 1 20 Dpar a=15.5025 p=62.01 m=1 $[ndiode] $X=9913 $Y=38260 $D=181
X72 1 38 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=815 $D=181
X73 1 39 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=1585 $D=181
X74 1 37 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=2355 $D=181
X75 1 40 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=3125 $D=181
X76 1 36 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=3895 $D=181
X77 1 41 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=4665 $D=181
X78 1 35 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=5435 $D=181
X79 1 42 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=6205 $D=181
X80 1 34 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=6975 $D=181
X81 1 43 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=7745 $D=181
X82 1 33 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=8515 $D=181
X83 1 44 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=9285 $D=181
X84 1 45 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=30560 $D=181
X85 1 10 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=31330 $D=181
X86 1 46 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=32100 $D=181
X87 1 11 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=32870 $D=181
X88 1 47 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=33640 $D=181
X89 1 11 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=34410 $D=181
X90 1 48 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=35180 $D=181
X91 1 12 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=35950 $D=181
X92 1 49 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=36720 $D=181
X93 1 13 Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=37490 $D=181
X94 1 50 Dpar a=12.0235 p=48.594 m=1 $[ndiode] $X=40923 $Y=38260 $D=181
X95 1 IN Dpar a=12.024 p=48.596 m=1 $[ndiode] $X=40922 $Y=39030 $D=181
X96 1 33 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=10735 $D=181
X97 1 34 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=12275 $D=181
X98 1 35 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=13815 $D=181
X99 1 36 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=15355 $D=181
X100 1 37 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=16895 $D=181
X101 1 38 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=18435 $D=181
X102 1 13 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=21405 $D=181
X103 1 12 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=22945 $D=181
X104 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=24485 $D=181
X105 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=26025 $D=181
X106 1 10 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=27565 $D=181
X107 1 9 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=58090 $Y=29105 $D=181
X108 1 33 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=11505 $D=181
X109 1 34 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=13045 $D=181
X110 1 35 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=14585 $D=181
X111 1 36 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=16125 $D=181
X112 1 37 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=17665 $D=181
X113 1 38 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=19205 $D=181
X114 1 IN Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=20635 $D=181
X115 1 13 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=22175 $D=181
X116 1 12 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=23715 $D=181
X117 1 11 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=25255 $D=181
X118 1 11 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=26795 $D=181
X119 1 10 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=58090 $Y=28335 $D=181
X120 1 44 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=10735 $D=181
X121 1 33 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=11505 $D=181
X122 1 43 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=12275 $D=181
X123 1 34 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=13045 $D=181
X124 1 42 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=13815 $D=181
X125 1 35 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=14585 $D=181
X126 1 41 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=15355 $D=181
X127 1 36 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=16125 $D=181
X128 1 40 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=16895 $D=181
X129 1 37 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=17665 $D=181
X130 1 39 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=18435 $D=181
X131 1 38 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=19205 $D=181
X132 1 IN Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=20635 $D=181
X133 1 50 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=21405 $D=181
X134 1 13 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=22175 $D=181
X135 1 49 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=22945 $D=181
X136 1 12 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=23715 $D=181
X137 1 48 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=24485 $D=181
X138 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=25255 $D=181
X139 1 47 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=26025 $D=181
X140 1 11 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=26795 $D=181
X141 1 46 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=27565 $D=181
X142 1 10 Dpar a=3.7735 p=15.594 m=1 $[ndiode] $X=65643 $Y=28335 $D=181
X143 1 45 Dpar a=3.774 p=15.596 m=1 $[ndiode] $X=65642 $Y=29105 $D=181
X144 1 VCC_IO Dpar a=501.44 p=125.96 m=1 $[nwdiode] $X=1350 $Y=20095 $D=191
X145 20 32 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=16535 39150 0 0 $X=16535 $Y=39150
X146 8 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 935 0 0 $X=54510 $Y=935
X147 7 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 2475 0 0 $X=54510 $Y=2475
X148 6 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 4015 0 0 $X=54510 $Y=4015
X149 5 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 5555 0 0 $X=54510 $Y=5555
X150 3 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=54510 8635 0 0 $X=54510 $Y=8635
X151 9 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=71780 29485 0 180 $X=71360 $Y=29225
X152 12 49 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=72265 23325 1 0 $X=72265 $Y=23065
X153 11 47 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=72265 26405 1 0 $X=72265 $Y=26145
X154 9 45 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808757 $T=72265 29485 1 0 $X=72265 $Y=29225
X155 15 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=16525 30680 0 0 $X=16525 $Y=30680
X156 IN sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=72255 21015 1 0 $X=72255 $Y=20755
X157 12 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=72255 24095 1 0 $X=72255 $Y=23835
X158 11 sky130_fd_io__xres_p_em1c_cdns_55959141808753 $T=72255 27175 1 0 $X=72255 $Y=26915
X159 33 44 ICV_2 $T=72265 11115 1 0 $X=72255 $Y=10855
X160 34 43 ICV_2 $T=72265 12655 1 0 $X=72255 $Y=12395
X161 35 42 ICV_2 $T=72265 14195 1 0 $X=72255 $Y=13935
X162 36 41 ICV_2 $T=72265 15735 1 0 $X=72255 $Y=15475
X163 37 40 ICV_2 $T=72265 17275 1 0 $X=72255 $Y=17015
X164 38 39 ICV_2 $T=72265 18815 1 0 $X=72255 $Y=18555
X165 13 50 ICV_2 $T=72265 21785 1 0 $X=72255 $Y=21525
X166 11 48 ICV_2 $T=72265 24865 1 0 $X=72255 $Y=24605
X167 10 46 ICV_2 $T=72265 27945 1 0 $X=72255 $Y=27685
X168 34 43 34 34 33 44 33 33 ICV_4 $T=72640 11235 0 180 $X=58300 $Y=10605
X169 36 41 36 36 35 42 35 35 ICV_4 $T=72640 14315 0 180 $X=58300 $Y=13685
X170 38 39 38 38 37 40 37 37 ICV_4 $T=72640 17395 0 180 $X=58300 $Y=16765
X171 12 13 49 13 13 IN 50 IN ICV_4 $T=58640 21135 1 0 $X=58300 $Y=20505
X172 11 11 47 11 11 12 48 12 ICV_4 $T=58640 24215 1 0 $X=58300 $Y=23585
X173 9 10 45 10 10 11 46 11 ICV_4 $T=58640 27295 1 0 $X=58300 $Y=26665
X174 1 7 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 2025 0 90 $X=2330 $Y=2025
X175 1 6 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 3565 0 90 $X=2330 $Y=3565
X176 1 5 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 5100 0 90 $X=2330 $Y=5100
X177 1 4 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=2980 6640 0 90 $X=2330 $Y=6640
X178 13 12 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 22600 1 90 $X=58060 $Y=22600
X179 12 11 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 24140 1 90 $X=58060 $Y=24140
X180 11 10 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 27220 1 90 $X=58060 $Y=27220
X181 10 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808758 $T=58060 28760 1 90 $X=58060 $Y=28760
X182 3 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 $T=2980 8155 0 90 $X=2330 $Y=8155
X183 11 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808760 $T=58060 25680 1 90 $X=58060 $Y=25680
X184 9 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 $T=29530 9405 0 0 $X=29530 $Y=9405
X185 4 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808761 $T=54470 7095 0 0 $X=54470 $Y=7095
X218 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=15570 6585 0 90 $X=15280 $Y=6585
X219 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=24130 5045 0 90 $X=23840 $Y=5045
X220 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=28410 3505 0 90 $X=28120 $Y=3505
X221 1 sky130_fd_io__xres_tk_p_em1c_cdns_55959141808759 $T=32690 1965 0 90 $X=32400 $Y=1965
X222 8 21 1 ICV_7 $T=16535 935 0 0 $X=16525 $Y=935
X223 7 22 1 ICV_7 $T=16535 2475 0 0 $X=16525 $Y=2475
X224 6 23 1 ICV_7 $T=16535 4015 0 0 $X=16525 $Y=4015
X225 5 24 1 ICV_7 $T=16535 5555 0 0 $X=16525 $Y=5555
X226 4 25 3 ICV_7 $T=16535 7095 0 0 $X=16525 $Y=7095
X227 3 26 9 ICV_7 $T=16535 8635 0 0 $X=16525 $Y=8635
X228 15 27 16 ICV_7 $T=16535 31450 0 0 $X=16525 $Y=31450
X229 16 28 17 ICV_7 $T=16535 32990 0 0 $X=16525 $Y=32990
X230 17 29 18 ICV_7 $T=16535 34530 0 0 $X=16525 $Y=34530
X231 18 30 19 ICV_7 $T=16535 36070 0 0 $X=16525 $Y=36070
X232 19 31 20 ICV_7 $T=16535 37610 0 0 $X=16525 $Y=37610
X233 1 9 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 $T=7010 9665 0 90 $X=6720 $Y=9665
X234 1 3 sky130_fd_io__xres_tk_p_em1o_cdns_55959141808756 $T=11290 8125 0 90 $X=11000 $Y=8125
X235 32 20 IN ICV_8 $T=16910 39030 1 180 $X=2570 $Y=38900
X236 15 45 ICV_9 $T=2910 30560 0 0 $X=2570 $Y=30430
X237 13 31 19 20 50 ICV_10 $T=16910 37490 1 180 $X=2570 $Y=37360
X238 38 39 21 1 8 37 40 22 1 7 ICV_11 $T=16910 815 1 180 $X=2570 $Y=685
X239 36 41 23 1 6 35 42 24 1 5 ICV_11 $T=16910 3895 1 180 $X=2570 $Y=3765
X240 34 43 25 3 4 33 44 26 9 3 ICV_11 $T=16910 6975 1 180 $X=2570 $Y=6845
X241 10 46 27 16 15 11 47 28 17 16 ICV_11 $T=16910 31330 1 180 $X=2570 $Y=31200
X242 11 48 29 18 17 12 49 30 19 18 ICV_11 $T=16910 34410 1 180 $X=2570 $Y=34280
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808243
** N=5 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808723
** N=13 EP=0 IP=10 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_5595914180848
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180849
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808371
** N=15 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x1
** N=31 EP=0 IP=24 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VGND VPWR OUT
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__pfet_highvoltage__example_55959141808421
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__hvsbt_inv_x2
** N=44 EP=0 IP=28 FDC=0
*.SEEDPROM
*.CALIBRE ISOLATED NETS: VGND VPWR IN OUT
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808719
** N=11 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808720
** N=24 EP=0 IP=22 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180829
** N=31 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808767 2 3 4 5
** N=26 EP=4 IP=22 FDC=1
*.SEEDPROM
M0 5 3 4 2 phv L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=0 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_fd_io__tk_tie_r_out_esd A B
** N=8 EP=2 IP=6 FDC=1
X0 A B sky130_fd_pr__res_generic_po__example_5595914180838 $T=1000 1095 0 0 $X=730 $Y=1095
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808765
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808764 1 2 3 4
** N=9 EP=4 IP=4 FDC=1
M0 4 2 3 1 nhv L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808779 1 2 3 4
** N=15 EP=4 IP=10 FDC=1
M0 4 2 3 1 nhvnative L=0.9 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 r=1.11111 sa=450000 sb=450000 a=0.9 p=3.8 mult=1 $X=0 $Y=0 $D=59
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808777 1 2 3
** N=16 EP=3 IP=2 FDC=1
M0 3 2 1 1 nhv L=0.5 W=3 AD=0.84 AS=0.795 PD=6.56 PS=6.53 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_5595914180827
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808233
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808778
** N=53 EP=0 IP=48 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd2__example_55959141808449
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808784 2 3 4
** N=9 EP=3 IP=6 FDC=1
*.SEEDPROM
M0 2 3 4 2 phv L=0.8 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 r=1.25 sa=400000 sb=400000 a=0.8 p=3.6 mult=1 $X=0 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_559591418085
** N=16 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808783
** N=11 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfm1sd__example_55959141808782
** N=10 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808786
** N=35 EP=0 IP=33 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808787
** N=36 EP=0 IP=34 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808151
** N=30 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808148
** N=17 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808150
** N=20 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__tpl1__example_55959141808149
** N=11 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808158
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__signal_5_sym_hv_local_5term NBODY NWELLRING GATE VGND IN 7
** N=101 EP=6 IP=102 FDC=3
*.SEEDPROM
M0 IN GATE VGND NBODY nhvesd L=0.6 W=5.4 AD=3.65486 AS=3.65486 PD=11.6192 PS=11.6192 NRD=8.436 NRS=9.2796 m=1 r=9 sa=300000 sb=300000 a=3.24 p=12 mult=1 $X=3675 $Y=3360 $D=129
R1 NWELLRING 7 0.01 m=1 $[short] $X=1015 $Y=330 $D=282
R2 NBODY 51 0.01 m=1 $[short] $X=2665 $Y=330 $D=282
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_5595914180819
** N=10 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_buf_localesdv2 VGND VCC_IO VTRIP_SEL_H OUT_H 5
** N=179 EP=5 IP=209 FDC=25
*.SEEDPROM
M0 OUT_VT VTRIP_SEL_H OUT_H VGND nhv L=1 W=3 AD=0.795 AS=0.795 PD=6.53 PS=6.53 NRD=0 NRS=0 m=1 r=3 sa=500000 sb=500000 a=3 p=8 mult=1 $X=16175 $Y=17310 $D=49
X1 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=1460 $Y=1770 $D=190
X2 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=1460 $Y=12530 $D=190
X3 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=8055 $Y=1770 $D=190
X4 VGND VCC_IO Dpar a=8.5092 p=29.27 m=1 $[nwdiode] $X=8055 $Y=12530 $D=190
X5 VGND VCC_IO Dpar a=5.1688 p=17.34 m=1 $[nwdiode] $X=14650 $Y=15810 $D=190
X6 5 OUT_H sky130_fd_io__res250only_small $T=17545 -185 0 90 $X=15525 $Y=-185
X7 VGND VCC_IO VGND VGND OUT_VT 8 sky130_fd_io__signal_5_sym_hv_local_5term $T=8335 690 1 180 $X=380 $Y=690
X8 VGND VCC_IO VGND VGND OUT_H 10 sky130_fd_io__signal_5_sym_hv_local_5term $T=8335 23570 0 180 $X=380 $Y=11450
X9 VGND VCC_IO VGND OUT_VT VCC_IO 7 sky130_fd_io__signal_5_sym_hv_local_5term $T=6975 690 0 0 $X=6975 $Y=690
X10 VGND VCC_IO VGND OUT_H VCC_IO 9 sky130_fd_io__signal_5_sym_hv_local_5term $T=6975 23570 1 0 $X=6975 $Y=11450
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpm1s2__example_55959141808659
** N=44 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__pfet_01v8__example_55959141808658
** N=36 EP=0 IP=26 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808646
** N=29 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808647
** N=4 EP=0 IP=1 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd2__example_55959141808378
** N=16 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpm1s2__example_55959141808649
** N=43 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_12
** N=2 EP=0 IP=4 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808650
** N=4 EP=0 IP=1 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 1 2 VCC_IO 4 5 6 7 8 9 10 11 12 13 14
** N=3678 EP=14 IP=101 FDC=58
*.SEEDPROM
M0 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4620 $Y=7285 $D=49
M1 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.425 PD=6.55 PS=11.37 NRD=10.374 NRS=8.7666 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4620 $Y=15290 $D=49
M2 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6770 $Y=7285 $D=49
M3 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6770 $Y=15290 $D=49
M4 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9580 $Y=7285 $D=49
M5 14 4 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9580 $Y=15290 $D=49
M6 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11730 $Y=7285 $D=49
M7 2 4 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11730 $Y=15290 $D=49
M8 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300011 sb=300020 a=3 p=11.2 mult=1 $X=14540 $Y=7285 $D=49
M9 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300011 sb=300020 a=3 p=11.2 mult=1 $X=14540 $Y=15290 $D=49
M10 2 5 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16690 $Y=7285 $D=49
M11 2 5 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16690 $Y=15290 $D=49
M12 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300016 sb=300020 a=3 p=11.2 mult=1 $X=19500 $Y=7285 $D=49
M13 14 5 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300016 sb=300020 a=3 p=11.2 mult=1 $X=19500 $Y=15290 $D=49
M14 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21650 $Y=7285 $D=49
M15 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21650 $Y=15290 $D=49
M16 14 6 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=24460 $Y=7285 $D=49
M17 14 6 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=24460 $Y=15290 $D=49
M18 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26610 $Y=7285 $D=49
M19 2 6 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26610 $Y=15290 $D=49
M20 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=29420 $Y=7285 $D=49
M21 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=29420 $Y=15290 $D=49
M22 2 7 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31570 $Y=7285 $D=49
M23 2 7 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31570 $Y=15290 $D=49
M24 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=34380 $Y=7285 $D=49
M25 14 7 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=34380 $Y=15290 $D=49
M26 2 8 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=36530 $Y=7285 $D=49
M27 2 8 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=36530 $Y=15290 $D=49
M28 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=39340 $Y=7285 $D=49
M29 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=39340 $Y=15290 $D=49
M30 2 9 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=41490 $Y=7285 $D=49
M31 2 9 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=41490 $Y=15290 $D=49
M32 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=44300 $Y=7285 $D=49
M33 14 9 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=44300 $Y=15290 $D=49
M34 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=46450 $Y=7285 $D=49
M35 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=46450 $Y=15290 $D=49
M36 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=49260 $Y=7285 $D=49
M37 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=49260 $Y=15290 $D=49
M38 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=51410 $Y=7285 $D=49
M39 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=51410 $Y=15290 $D=49
M40 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=54220 $Y=7285 $D=49
M41 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=54220 $Y=15290 $D=49
M42 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=56370 $Y=7285 $D=49
M43 2 10 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=56370 $Y=15290 $D=49
M44 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=59180 $Y=7285 $D=49
M45 14 10 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=59180 $Y=15290 $D=49
M46 2 11 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=61330 $Y=7285 $D=49
M47 2 11 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=61330 $Y=15290 $D=49
M48 14 12 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=64140 $Y=7285 $D=49
M49 14 12 2 2 nhv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=64140 $Y=15290 $D=49
M50 2 13 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=66290 $Y=7285 $D=49
M51 2 13 14 2 nhv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=66290 $Y=15290 $D=49
M52 14 13 2 2 nhv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=69100 $Y=7285 $D=49
M53 14 13 2 2 nhv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=10.374 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=69100 $Y=15290 $D=49
M54 2 13 14 2 nhv L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70890 $Y=7285 $D=49
M55 2 13 14 2 nhv L=0.6 W=5 AD=3.425 AS=2.975 PD=11.37 PS=6.19 NRD=8.7666 NRS=10.374 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70890 $Y=15290 $D=49
X56 1 VCC_IO Dpar a=1791.37 p=197.77 m=1 $[dnwdiode_psub] $X=440 $Y=2895 $D=193
X57 2 VCC_IO Dpar a=1558.74 p=186.49 m=1 $[dnwdiode_pw] $X=2345 $Y=3925 $D=194
.ENDS
***************************************
.SUBCKT sky130_fd_io__gpio_pddrvr_strong_xres4v2 1 TIE_LO_ESD 3 VCC_IO PD_H[2] PD_H[3] 7 8
** N=70 EP=8 IP=140 FDC=109
X0 3 VCC_IO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=6380 $Y=37555 $D=150
X1 1 VCC_IO Dpar a=57.3765 p=0 m=1 $[nwdiode] $X=-515 $Y=14600 $D=189
X2 PD_H[3] 7 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=3275 5230 1 90 $X=3275 $Y=5230
X3 PD_H[2] 7 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=4480 5230 1 90 $X=4480 $Y=5230
X4 PD_H[3] 15 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=8470 5230 0 90 $X=7820 $Y=5230
X5 TIE_LO_ESD 15 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=9885 5230 0 90 $X=9235 $Y=5230
X6 PD_H[3] 14 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=16120 5230 0 90 $X=15470 $Y=5230
X7 TIE_LO_ESD 14 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=17535 5230 0 90 $X=16885 $Y=5230
X8 PD_H[2] 13 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=34665 5230 0 90 $X=34015 $Y=5230
X9 TIE_LO_ESD 13 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=38965 5230 0 90 $X=38315 $Y=5230
X10 PD_H[2] 12 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=43175 5230 0 90 $X=42525 $Y=5230
X11 TIE_LO_ESD 12 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=47475 5230 0 90 $X=46825 $Y=5230
X12 PD_H[2] 11 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=50575 5230 0 90 $X=49925 $Y=5230
X13 TIE_LO_ESD 11 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=54875 5230 0 90 $X=54225 $Y=5230
X14 PD_H[2] 10 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=57290 5230 0 90 $X=56640 $Y=5230
X15 TIE_LO_ESD 10 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=61590 5230 0 90 $X=60940 $Y=5230
X16 PD_H[2] 9 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=64460 5230 0 90 $X=63810 $Y=5230
X17 PD_H[3] 9 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=66610 5230 0 90 $X=65960 $Y=5230
X18 TIE_LO_ESD 7 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=2065 5230 1 90 $X=2065 $Y=5230
X19 PD_H[2] 15 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=6950 5230 0 90 $X=6300 $Y=5230
X20 PD_H[2] 14 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=14600 5230 0 90 $X=13950 $Y=5230
X21 PD_H[3] 13 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=36815 5230 0 90 $X=36165 $Y=5230
X22 PD_H[3] 12 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=45325 5230 0 90 $X=44675 $Y=5230
X23 PD_H[3] 11 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=52725 5230 0 90 $X=52075 $Y=5230
X24 PD_H[3] 10 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=59440 5230 0 90 $X=58790 $Y=5230
X25 TIE_LO_ESD 9 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=68760 5230 0 90 $X=68110 $Y=5230
X26 TIE_LO_ESD 3 sky130_fd_pr__res_generic_po__example_5595914180838 $T=2320 46835 0 0 $X=2050 $Y=46835
X27 1 3 VCC_IO 9 10 11 12 13 PD_H[2] PD_H[3] 14 15 7 8 sky130_fd_io__nfet_con_diff_wo_abt_270_xres4v2 $T=75440 42045 0 180 $X=-515 $Y=14600
.ENDS
***************************************
.SUBCKT sky130_fd_io__top_xres4v2 VSSD VDDIO VCCHIB VDDIO_Q ENABLE_H EN_VDDIO_SIG_H INP_SEL_H ENABLE_VDDIO PAD PULLUP_H DISABLE_PULLUP_H PAD_A_ESD_H VSSIO FILT_IN_H TIE_LO_ESD XRES_H_N TIE_HI_ESD TIE_WEAK_HI_H VCCD VDDA
+ VSWITCH VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q
** N=38667 EP=25 IP=1572 FDC=777
M0 VSSD ENABLE_VDDIO 19 VSSD nshort L=0.15 W=0.74 AD=0.2627 AS=0.2109 PD=2.19 PS=2.05 NRD=11.34 NRS=0 m=1 r=4.93333 sa=75000.2 sb=75000.3 a=0.111 p=1.78 mult=1 $X=16840 $Y=40175 $D=9
M1 47 15 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=13.8396 NRS=0 m=1 r=1.16667 sa=300000 sb=300001 a=0.42 p=2.6 mult=1 $X=8460 $Y=7500 $D=49
M2 40 ENABLE_H 47 VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=13.8396 m=1 r=1.16667 sa=300001 sb=300000 a=0.42 p=2.6 mult=1 $X=9340 $Y=7500 $D=49
M3 17 40 VSSD VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.1855 PD=1.93 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300000 a=0.42 p=2.6 mult=1 $X=10845 $Y=7500 $D=49
M4 14 22 VSSD VSSD nhv L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250002 a=2.5 p=11 mult=1 $X=15285 $Y=20910 $D=49
M5 VSSD 22 14 VSSD nhv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250002 a=2.5 p=11 mult=1 $X=15285 $Y=21690 $D=49
M6 13 20 VSSD VSSD nhv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250001 a=2.5 p=11 mult=1 $X=15285 $Y=22470 $D=49
M7 VSSD 20 13 VSSD nhv L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250000 a=2.5 p=11 mult=1 $X=15285 $Y=23250 $D=49
M8 50 20 48 VSSD nhv L=0.8 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=6.25 sa=400000 sb=400007 a=4 p=11.6 mult=1 $X=15315 $Y=28245 $D=49
M9 48 20 50 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400001 sb=400006 a=4 p=11.6 mult=1 $X=15315 $Y=29325 $D=49
M10 50 20 48 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400002 sb=400005 a=4 p=11.6 mult=1 $X=15315 $Y=30405 $D=49
M11 48 20 50 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400003 sb=400004 a=4 p=11.6 mult=1 $X=15315 $Y=31485 $D=49
M12 VSSD 11 48 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400004 sb=400003 a=4 p=11.6 mult=1 $X=15315 $Y=32565 $D=49
M13 48 11 VSSD VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400005 sb=400002 a=4 p=11.6 mult=1 $X=15315 $Y=33645 $D=49
M14 20 11 48 VSSD nhv L=0.8 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400006 sb=400001 a=4 p=11.6 mult=1 $X=15315 $Y=34725 $D=49
M15 48 11 20 VSSD nhv L=0.8 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=6.25 sa=400007 sb=400000 a=4 p=11.6 mult=1 $X=15315 $Y=35805 $D=49
M16 48 20 43 VSSD nhv L=0.8 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 r=6.25 sa=400000 sb=400000 a=4 p=11.6 mult=1 $X=15315 $Y=37540 $D=49
M17 VSSD 12 37 VSSD nhv L=0.5 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 r=2 sa=250000 sb=250002 a=0.5 p=3 mult=1 $X=21425 $Y=21690 $D=49
M18 37 12 VSSD VSSD nhv L=0.5 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=2 sa=250001 sb=250001 a=0.5 p=3 mult=1 $X=21425 $Y=22470 $D=49
M19 VSSD 12 37 VSSD nhv L=0.5 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=2 sa=250002 sb=250000 a=0.5 p=3 mult=1 $X=21425 $Y=23250 $D=49
M20 28 59 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300003 a=0.42 p=2.6 mult=1 $X=27755 $Y=29045 $D=49
M21 VSSD 59 28 VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300001 sb=300002 a=0.42 p=2.6 mult=1 $X=27755 $Y=29925 $D=49
M22 59 DISABLE_PULLUP_H VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300002 sb=300001 a=0.42 p=2.6 mult=1 $X=27755 $Y=30805 $D=49
M23 VSSD DISABLE_PULLUP_H 59 VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300000 a=0.42 p=2.6 mult=1 $X=27755 $Y=31685 $D=49
M24 VSSD 26 49 VSSD nhv L=1 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 r=0.42 sa=500000 sb=500000 a=0.42 p=2.84 mult=1 $X=30440 $Y=14450 $D=49
M25 49 27 VSSD VSSD nhv L=1 W=1 AD=0.14 AS=0.28 PD=1.28 PS=2.56 NRD=0 NRS=0 m=1 r=1 sa=500000 sb=500001 a=1 p=4 mult=1 $X=30720 $Y=9780 $D=49
M26 29 27 49 VSSD nhv L=1 W=1 AD=0.28 AS=0.14 PD=2.56 PS=1.28 NRD=0 NRS=0 m=1 r=1 sa=500001 sb=500000 a=1 p=4 mult=1 $X=30720 $Y=11060 $D=49
M27 26 29 VSSD VSSD nhv L=0.5 W=1 AD=0.28 AS=0.28 PD=2.56 PS=2.56 NRD=0 NRS=0 m=1 r=2 sa=250000 sb=250000 a=0.5 p=3 mult=1 $X=30720 $Y=12990 $D=49
M28 23 INP_SEL_H VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300007 a=0.42 p=2.6 mult=1 $X=31240 $Y=17710 $D=49
M29 VSSD INP_SEL_H 23 VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300001 sb=300006 a=0.42 p=2.6 mult=1 $X=31240 $Y=18590 $D=49
M30 15 EN_VDDIO_SIG_H VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300002 sb=300005 a=0.42 p=2.6 mult=1 $X=31240 $Y=19470 $D=49
M31 VSSD EN_VDDIO_SIG_H 15 VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300004 a=0.42 p=2.6 mult=1 $X=31240 $Y=20350 $D=49
M32 XRES_H_N 60 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300003 a=0.42 p=2.6 mult=1 $X=31240 $Y=21230 $D=49
M33 VSSD 60 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300004 sb=300003 a=0.42 p=2.6 mult=1 $X=31240 $Y=22110 $D=49
M34 XRES_H_N 60 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300005 sb=300002 a=0.42 p=2.6 mult=1 $X=31240 $Y=22990 $D=49
M35 VSSD 60 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300006 sb=300001 a=0.42 p=2.6 mult=1 $X=31240 $Y=23870 $D=49
M36 60 26 VSSD VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300007 sb=300000 a=0.42 p=2.6 mult=1 $X=31240 $Y=24750 $D=49
M37 XRES_H_N 60 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.1855 PD=0.98 PS=1.93 NRD=0 NRS=0 m=1 r=1.16667 sa=300000 sb=300003 a=0.42 p=2.6 mult=1 $X=35355 $Y=4770 $D=49
M38 VSSD 60 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300001 sb=300002 a=0.42 p=2.6 mult=1 $X=36235 $Y=4770 $D=49
M39 XRES_H_N 60 VSSD VSSD nhv L=0.6 W=0.7 AD=0.098 AS=0.098 PD=0.98 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300002 sb=300001 a=0.42 p=2.6 mult=1 $X=37115 $Y=4770 $D=49
M40 VSSD 60 XRES_H_N VSSD nhv L=0.6 W=0.7 AD=0.1855 AS=0.098 PD=1.93 PS=0.98 NRD=0 NRS=0 m=1 r=1.16667 sa=300003 sb=300000 a=0.42 p=2.6 mult=1 $X=37995 $Y=4770 $D=49
M41 4 17 46 VSSD nhvnative L=0.9 W=10 AD=2.8 AS=2.8 PD=20.56 PS=20.56 NRD=0 NRS=0 m=1 r=11.1111 sa=450000 sb=450000 a=9 p=21.8 mult=1 $X=21675 $Y=26745 $D=59
M42 VSSD VSSD VSSD VSSD nhvnative L=0.9 W=10 AD=2.8 AS=2.65 PD=20.56 PS=20.53 NRD=0 NRS=0 m=1 r=11.1111 sa=450000 sb=450000 a=9 p=21.8 mult=1 $X=23490 $Y=26745 $D=59
M43 VCCHIB ENABLE_VDDIO 19 VCCHIB phighvt L=0.15 W=1.12 AD=0.3864 AS=0.3304 PD=2.93 PS=2.83 NRD=10.5395 NRS=1.7533 m=1 r=7.46667 sa=75000.2 sb=75000.3 a=0.168 p=2.54 mult=1 $X=14990 $Y=40185 $D=89
M44 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4065 $Y=107610 $D=109
M45 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=4.325 PD=6.55 PS=11.73 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300002 sb=300020 a=3 p=11.2 mult=1 $X=4065 $Y=115610 $D=109
M46 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6215 $Y=107610 $D=109
M47 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300004 sb=300020 a=3 p=11.2 mult=1 $X=6215 $Y=115610 $D=109
M48 VDDIO_Q 13 14 VDDIO_Q phv L=0.5 W=0.42 AD=0.0588 AS=0.1176 PD=0.7 PS=1.4 NRD=0 NRS=0 m=1 r=0.84 sa=250000 sb=250001 a=0.21 p=1.84 mult=1 $X=7410 $Y=24400 $D=109
M49 13 14 VDDIO_Q VDDIO_Q phv L=0.5 W=0.42 AD=0.1176 AS=0.0588 PD=1.4 PS=0.7 NRD=0 NRS=0 m=1 r=0.84 sa=250001 sb=250000 a=0.21 p=1.84 mult=1 $X=7410 $Y=25180 $D=109
M50 40 15 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300001 a=0.6 p=3.2 mult=1 $X=8460 $Y=4170 $D=109
M51 40 15 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300001 a=0.6 p=3.2 mult=1 $X=8460 $Y=5510 $D=109
M52 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9025 $Y=107610 $D=109
M53 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300007 sb=300020 a=3 p=11.2 mult=1 $X=9025 $Y=115610 $D=109
M54 VDDIO_Q ENABLE_H 40 VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300000 a=0.6 p=3.2 mult=1 $X=9340 $Y=4170 $D=109
M55 VDDIO_Q ENABLE_H 40 VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300000 a=0.6 p=3.2 mult=1 $X=9340 $Y=5510 $D=109
M56 VDDIO_Q 12 37 VDDIO_Q phv L=0.5 W=3 AD=0.42 AS=0.84 PD=3.28 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250002 a=1.5 p=7 mult=1 $X=7095 $Y=19975 $D=109
M57 37 12 VDDIO_Q VDDIO_Q phv L=0.5 W=3 AD=0.42 AS=0.42 PD=3.28 PS=3.28 NRD=0 NRS=0 m=1 r=6 sa=250001 sb=250001 a=1.5 p=7 mult=1 $X=7095 $Y=20755 $D=109
M58 VDDIO_Q 12 37 VDDIO_Q phv L=0.5 W=3 AD=0.795 AS=0.42 PD=6.53 PS=3.28 NRD=0 NRS=0 m=1 r=6 sa=250002 sb=250000 a=1.5 p=7 mult=1 $X=7095 $Y=21535 $D=109
M59 VDDIO_Q 13 12 VDDIO_Q phv L=0.5 W=3 AD=0.795 AS=0.84 PD=6.53 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=7095 $Y=22950 $D=109
M60 17 40 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300000 a=0.6 p=3.2 mult=1 $X=10845 $Y=4170 $D=109
M61 17 40 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.265 PD=2.53 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300000 a=0.6 p=3.2 mult=1 $X=10845 $Y=5510 $D=109
M62 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11175 $Y=107610 $D=109
M63 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300009 sb=300020 a=3 p=11.2 mult=1 $X=11175 $Y=115610 $D=109
M64 VDDIO_Q ENABLE_H 41 VDDIO_Q phv L=0.5 W=5 AD=1.325 AS=1.4 PD=10.53 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=29660 $D=109
M65 36 11 20 VDDIO_Q phv L=0.5 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=31460 $D=109
M66 42 17 VDDIO_Q VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250001 a=2.5 p=11 mult=1 $X=6920 $Y=32875 $D=109
M67 36 15 42 VDDIO_Q phv L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=33655 $D=109
M68 VDDIO_Q 15 43 VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250001 a=2.5 p=11 mult=1 $X=6920 $Y=35115 $D=109
M69 44 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q phv L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=35895 $D=109
M70 VCCHIB 19 45 VCCHIB phv L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250001 a=2.5 p=11 mult=1 $X=6920 $Y=39685 $D=109
M71 46 19 VCCHIB VCCHIB phv L=0.5 W=5 AD=1.4 AS=0.7 PD=10.56 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250000 a=2.5 p=11 mult=1 $X=6920 $Y=40465 $D=109
M72 5 20 22 5 phv L=0.5 W=5 AD=1.4 AS=1.4 PD=10.56 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250000 a=2.5 p=11 mult=1 $X=7095 $Y=15515 $D=109
M73 30 20 22 VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=1.4 PD=5.28 PS=10.56 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250002 a=2.5 p=11 mult=1 $X=7095 $Y=26635 $D=109
M74 7 15 30 VDDIO_Q phv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250001 a=2.5 p=11 mult=1 $X=7095 $Y=27415 $D=109
M75 VDDIO_Q 17 7 VDDIO_Q phv L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250000 a=2.5 p=11 mult=1 $X=7095 $Y=28195 $D=109
M76 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300012 sb=300020 a=3 p=11.2 mult=1 $X=13985 $Y=107610 $D=109
M77 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300012 sb=300020 a=3 p=11.2 mult=1 $X=13985 $Y=115610 $D=109
M78 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16135 $Y=107610 $D=109
M79 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300014 sb=300020 a=3 p=11.2 mult=1 $X=16135 $Y=115610 $D=109
M80 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300017 sb=300020 a=3 p=11.2 mult=1 $X=18945 $Y=107610 $D=109
M81 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300017 sb=300020 a=3 p=11.2 mult=1 $X=18945 $Y=115610 $D=109
M82 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21095 $Y=107610 $D=109
M83 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300019 sb=300020 a=3 p=11.2 mult=1 $X=21095 $Y=115610 $D=109
M84 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=23905 $Y=107610 $D=109
M85 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=23905 $Y=115610 $D=109
M86 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26055 $Y=107610 $D=109
M87 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=26055 $Y=115610 $D=109
M88 38 26 VDDIO_Q VDDIO_Q phv L=1 W=0.42 AD=0.1176 AS=0.1176 PD=1.4 PS=1.4 NRD=0 NRS=0 m=1 r=0.42 sa=500000 sb=500000 a=0.42 p=2.84 mult=1 $X=26705 $Y=14610 $D=109
M89 10 28 VDDIO VDDIO phv L=0.5 W=5 AD=0.7 AS=1.325 PD=5.28 PS=10.53 NRD=0 NRS=0 m=1 r=10 sa=250000 sb=250002 a=2.5 p=11 mult=1 $X=27850 $Y=35625 $D=109
M90 23 INP_SEL_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300007 a=0.6 p=3.2 mult=1 $X=27910 $Y=17710 $D=109
M91 VDDIO_Q INP_SEL_H 23 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300006 a=0.6 p=3.2 mult=1 $X=27910 $Y=18590 $D=109
M92 15 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300005 a=0.6 p=3.2 mult=1 $X=27910 $Y=19470 $D=109
M93 VDDIO_Q EN_VDDIO_SIG_H 15 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300004 a=0.6 p=3.2 mult=1 $X=27910 $Y=20350 $D=109
M94 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300003 a=0.6 p=3.2 mult=1 $X=27910 $Y=21230 $D=109
M95 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300004 sb=300003 a=0.6 p=3.2 mult=1 $X=27910 $Y=22110 $D=109
M96 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300005 sb=300002 a=0.6 p=3.2 mult=1 $X=27910 $Y=22990 $D=109
M97 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300006 sb=300001 a=0.6 p=3.2 mult=1 $X=27910 $Y=23870 $D=109
M98 60 26 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300007 sb=300000 a=0.6 p=3.2 mult=1 $X=27910 $Y=24750 $D=109
M99 VDDIO 28 10 VDDIO phv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250001 sb=250002 a=2.5 p=11 mult=1 $X=28630 $Y=35625 $D=109
M100 38 27 VDDIO_Q VDDIO_Q phv L=1 W=3 AD=0.42 AS=0.84 PD=3.28 PS=6.56 NRD=0 NRS=0 m=1 r=3 sa=500000 sb=500001 a=3 p=8 mult=1 $X=26420 $Y=9780 $D=109
M101 29 27 38 VDDIO_Q phv L=1 W=3 AD=0.84 AS=0.42 PD=6.56 PS=3.28 NRD=0 NRS=0 m=1 r=3 sa=500001 sb=500000 a=3 p=8 mult=1 $X=26420 $Y=11060 $D=109
M102 26 29 VDDIO_Q VDDIO_Q phv L=0.5 W=3 AD=0.84 AS=0.84 PD=6.56 PS=6.56 NRD=0 NRS=0 m=1 r=6 sa=250000 sb=250000 a=1.5 p=7 mult=1 $X=26420 $Y=12990 $D=109
M103 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=28865 $Y=107610 $D=109
M104 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=28865 $Y=115610 $D=109
M105 10 28 VDDIO VDDIO phv L=0.5 W=5 AD=0.7 AS=0.7 PD=5.28 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250001 a=2.5 p=11 mult=1 $X=29410 $Y=35625 $D=109
M106 23 INP_SEL_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300007 a=0.6 p=3.2 mult=1 $X=29250 $Y=17710 $D=109
M107 VDDIO_Q INP_SEL_H 23 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300006 a=0.6 p=3.2 mult=1 $X=29250 $Y=18590 $D=109
M108 15 EN_VDDIO_SIG_H VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300005 a=0.6 p=3.2 mult=1 $X=29250 $Y=19470 $D=109
M109 VDDIO_Q EN_VDDIO_SIG_H 15 VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300004 a=0.6 p=3.2 mult=1 $X=29250 $Y=20350 $D=109
M110 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300003 a=0.6 p=3.2 mult=1 $X=29250 $Y=21230 $D=109
M111 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300004 sb=300003 a=0.6 p=3.2 mult=1 $X=29250 $Y=22110 $D=109
M112 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300005 sb=300002 a=0.6 p=3.2 mult=1 $X=29250 $Y=22990 $D=109
M113 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300006 sb=300001 a=0.6 p=3.2 mult=1 $X=29250 $Y=23870 $D=109
M114 60 26 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300007 sb=300000 a=0.6 p=3.2 mult=1 $X=29250 $Y=24750 $D=109
M115 28 59 VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=29445 $Y=29045 $D=109
M116 VDDIO 59 28 VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=29445 $Y=29925 $D=109
M117 59 DISABLE_PULLUP_H VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=29445 $Y=30805 $D=109
M118 VDDIO DISABLE_PULLUP_H 59 VDDIO phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=29445 $Y=31685 $D=109
M119 VDDIO 28 10 VDDIO phv L=0.5 W=5 AD=1.325 AS=0.7 PD=10.53 PS=5.28 NRD=0 NRS=0 m=1 r=10 sa=250002 sb=250000 a=2.5 p=11 mult=1 $X=30190 $Y=35625 $D=109
M120 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31015 $Y=107610 $D=109
M121 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=31015 $Y=115610 $D=109
M122 28 59 VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=30785 $Y=29045 $D=109
M123 VDDIO 59 28 VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=30785 $Y=29925 $D=109
M124 59 DISABLE_PULLUP_H VDDIO VDDIO phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=30785 $Y=30805 $D=109
M125 VDDIO DISABLE_PULLUP_H 59 VDDIO phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=30785 $Y=31685 $D=109
M126 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=33825 $Y=107610 $D=109
M127 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=33825 $Y=115610 $D=109
M128 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=35355 $Y=1440 $D=109
M129 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.265 PD=1.28 PS=2.53 NRD=0 NRS=0 m=1 r=1.66667 sa=300000 sb=300003 a=0.6 p=3.2 mult=1 $X=35355 $Y=2780 $D=109
M130 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=35975 $Y=107610 $D=109
M131 VDDIO 8 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=35975 $Y=115610 $D=109
M132 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=36235 $Y=1440 $D=109
M133 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300001 sb=300002 a=0.6 p=3.2 mult=1 $X=36235 $Y=2780 $D=109
M134 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=37115 $Y=1440 $D=109
M135 XRES_H_N 60 VDDIO_Q VDDIO_Q phv L=0.6 W=1 AD=0.14 AS=0.14 PD=1.28 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300002 sb=300001 a=0.6 p=3.2 mult=1 $X=37115 $Y=2780 $D=109
M136 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=37995 $Y=1440 $D=109
M137 VDDIO_Q 60 XRES_H_N VDDIO_Q phv L=0.6 W=1 AD=0.265 AS=0.14 PD=2.53 PS=1.28 NRD=0 NRS=0 m=1 r=1.66667 sa=300003 sb=300000 a=0.6 p=3.2 mult=1 $X=37995 $Y=2780 $D=109
M138 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=38785 $Y=107610 $D=109
M139 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=38785 $Y=115610 $D=109
M140 VDDIO 31 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=40935 $Y=107610 $D=109
M141 VDDIO 31 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=40935 $Y=115610 $D=109
M142 PAD 31 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=43745 $Y=107610 $D=109
M143 PAD 31 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=43745 $Y=115610 $D=109
M144 VDDIO 31 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=45895 $Y=107610 $D=109
M145 VDDIO 31 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=45895 $Y=115610 $D=109
M146 PAD 32 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=48705 $Y=107610 $D=109
M147 PAD 32 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=48705 $Y=115610 $D=109
M148 VDDIO 32 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=50855 $Y=107610 $D=109
M149 VDDIO 32 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300020 a=3 p=11.2 mult=1 $X=50855 $Y=115610 $D=109
M150 PAD 32 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=53665 $Y=107610 $D=109
M151 PAD 32 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300018 a=3 p=11.2 mult=1 $X=53665 $Y=115610 $D=109
M152 VDDIO 33 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=55815 $Y=107610 $D=109
M153 VDDIO 33 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300016 a=3 p=11.2 mult=1 $X=55815 $Y=115610 $D=109
M154 PAD 33 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=58625 $Y=107610 $D=109
M155 PAD 33 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300013 a=3 p=11.2 mult=1 $X=58625 $Y=115610 $D=109
M156 VDDIO 33 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=60775 $Y=107610 $D=109
M157 VDDIO 33 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300011 a=3 p=11.2 mult=1 $X=60775 $Y=115610 $D=109
M158 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=63585 $Y=107610 $D=109
M159 PAD 8 VDDIO VDDIO phv L=0.6 W=5 AD=3.875 AS=3.775 PD=6.55 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300008 a=3 p=11.2 mult=1 $X=63585 $Y=115610 $D=109
M160 VDDIO 34 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=65735 $Y=107610 $D=109
M161 VDDIO 34 PAD VDDIO phv L=0.6 W=5 AD=3.775 AS=3.875 PD=11.51 PS=6.55 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300006 a=3 p=11.2 mult=1 $X=65735 $Y=115610 $D=109
M162 PAD 35 VDDIO VDDIO phv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=68545 $Y=107610 $D=109
M163 PAD 35 VDDIO VDDIO phv L=0.6 W=5 AD=2.975 AS=3.775 PD=6.19 PS=11.51 NRD=17.381 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300003 a=3 p=11.2 mult=1 $X=68545 $Y=115610 $D=109
M164 VDDIO 35 PAD VDDIO phv L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70335 $Y=107610 $D=109
M165 VDDIO 35 PAD VDDIO phv L=0.6 W=5 AD=4.3 AS=2.975 PD=11.72 PS=6.19 NRD=17.19 NRS=17.381 m=1 r=8.33333 sa=300020 sb=300002 a=3 p=11.2 mult=1 $X=70335 $Y=115610 $D=109
X166 VSSD 42 Dpar a=156.97 p=1082.84 m=1 $[ndiode_h] $X=8720 $Y=183570 $D=182
X167 VSSD 36 Dpar a=156.981 p=1082.92 m=1 $[ndiode_h] $X=8720 $Y=189310 $D=182
X168 VSSD VDDIO_Q Dpar a=16.2631 p=16.27 m=1 $[nwdiode] $X=7655 $Y=3340 $D=191
X169 VSSD VCCHIB Dpar a=15.5 p=17.4 m=1 $[nwdiode] $X=6050 $Y=39075 $D=191
X170 VSSD VDDIO_Q Dpar a=96.7627 p=49.03 m=1 $[nwdiode] $X=6050 $Y=19410 $D=191
X171 VSSD 4 Dpar a=23.8226 p=21.54 m=1 $[nwdiode] $X=6220 $Y=9200 $D=191
X172 VSSD 5 Dpar a=21.9076 p=21.04 m=1 $[nwdiode] $X=6220 $Y=14310 $D=191
X173 VSSD VCCHIB Dpar a=4.2823 p=8.33 m=1 $[nwdiode] $X=14430 $Y=39555 $D=191
X174 VSSD VDDIO Dpar a=108.48 p=83.5 m=1 $[nwdiode] $X=5010 $Y=47395 $D=191
X175 VSSD VDDIO_Q Dpar a=40.2643 p=30.01 m=1 $[nwdiode] $X=20935 $Y=9430 $D=191
X176 VSSD VDDIO_Q Dpar a=32.0172 p=25.17 m=1 $[nwdiode] $X=27040 $Y=17115 $D=191
X177 VSSD VDDIO Dpar a=36.4812 p=24.46 m=1 $[nwdiode] $X=26670 $Y=34430 $D=191
X178 VSSD VDDIO Dpar a=15.7043 p=15.95 m=1 $[nwdiode] $X=29110 $Y=28450 $D=191
X179 VSSD VDDIO_Q Dpar a=16.8897 p=16.63 m=1 $[nwdiode] $X=34550 $Y=610 $D=191
X180 VSSD VDDIO Dpar a=1473.41 p=184.25 m=1 $[nwdiode] $X=1735 $Y=102850 $D=191
X181 VSSD VDDIO Dpar a=735.037 p=170.75 m=1 $[nwdiode] $X=-330 $Y=130665 $D=191
R182 42 36 L=1077.19 W=0.29 m=1 $[mrdn_hv] $X=8720 $Y=183570 $D=254
R183 9 10 L=50 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=5800 $Y=45140 $D=257
R184 VDDIO 21 L=50 W=0.8 m=1 mult=1 model="mrp1" $[mrp1] $X=13810 $Y=131810 $D=257
R185 30 7 L=713.695 W=0.4 m=1 mult=1 model="mrp1" $[mrp1] $X=3520 $Y=87005 $D=257
R186 51 81 0.01 m=1 $[short] $X=11385 $Y=43760 $D=282
R187 81 54 0.01 m=1 $[short] $X=11575 $Y=43760 $D=282
R188 54 83 0.01 m=1 $[short] $X=18125 $Y=43760 $D=282
R189 84 57 0.01 m=1 $[short] $X=18315 $Y=43760 $D=282
R190 61 89 0.01 m=1 $[short] $X=45905 $Y=129760 $D=282
R191 90 62 0.01 m=1 $[short] $X=47415 $Y=129760 $D=282
X192 8 31 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=44185 96810 1 90 $X=44185 $Y=96810
X193 8 31 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=45395 96810 1 90 $X=45395 $Y=96810
X194 8 32 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=52095 96810 1 90 $X=52095 $Y=96810
X195 8 32 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=54480 96810 1 90 $X=54480 $Y=96810
X196 8 33 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=59920 96455 1 90 $X=59920 $Y=96455
X197 8 33 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=61125 96455 1 90 $X=61125 $Y=96455
X198 8 34 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=65335 101140 1 90 $X=65335 $Y=101140
X199 8 34 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=67745 101140 1 90 $X=67745 $Y=101140
X200 8 35 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=70030 101140 1 90 $X=70030 $Y=101140
X201 8 35 sky130_fd_io__tk_em2o_cdns_55959141808653 $T=71215 101140 1 90 $X=71215 $Y=101140
X210 8 31 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=46570 96810 1 90 $X=46570 $Y=96810
X211 8 32 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=53305 96810 1 90 $X=53305 $Y=96810
X212 8 33 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=58710 96455 1 90 $X=58710 $Y=96455
X213 8 34 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=66560 101140 1 90 $X=66560 $Y=101140
X214 8 35 sky130_fd_io__tk_em2s_cdns_55959141808652 $T=68805 101140 1 90 $X=68805 $Y=101140
X241 8 VDDIO sky130_fd_pr__res_generic_po__example_5595914180838 $T=60050 98360 0 0 $X=59780 $Y=98360
X242 53 PULLUP_H sky130_fd_pr__res_generic_po__example_5595914180864 $T=8510 43145 0 180 $X=6740 $Y=42345
X243 55 53 sky130_fd_pr__res_generic_po__example_5595914180864 $T=11435 43145 0 180 $X=9665 $Y=42345
X244 56 55 sky130_fd_pr__res_generic_po__example_5595914180864 $T=14215 42335 1 180 $X=12445 $Y=42335
X245 51 56 sky130_fd_pr__res_generic_po__example_5595914180864 $T=17140 42335 1 180 $X=15370 $Y=42335
X246 66 63 sky130_fd_pr__res_generic_po__example_5595914180864 $T=57830 133080 1 180 $X=56060 $Y=133080
X247 64 65 sky130_fd_pr__res_generic_po__example_5595914180864 $T=56430 130495 1 0 $X=56160 $Y=129695
X248 67 66 sky130_fd_pr__res_generic_po__example_5595914180864 $T=60755 133080 1 180 $X=58985 $Y=133080
X249 65 67 sky130_fd_pr__res_generic_po__example_5595914180864 $T=59355 130495 1 0 $X=59085 $Y=129695
X250 53 PULLUP_H sky130_fd_io__tk_em1s_cdns_5595914180859 $T=8820 43070 0 180 $X=6780 $Y=42410
X251 55 53 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=11620 43070 0 180 $X=9580 $Y=42410
X252 56 55 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=14565 42410 1 180 $X=12525 $Y=42410
X253 51 56 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=17470 42410 1 180 $X=15430 $Y=42410
X254 62 64 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=52355 130420 1 0 $X=52355 $Y=129760
X255 66 63 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=58180 133155 1 180 $X=56140 $Y=133155
X256 64 65 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=56245 130420 1 0 $X=56245 $Y=129760
X257 65 67 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=59045 130420 1 0 $X=59045 $Y=129760
X258 67 66 sky130_fd_io__tk_em1s_cdns_5595914180859 $T=61085 133155 1 180 $X=59045 $Y=133155
X259 PAD PAD_A_ESD_H sky130_fd_io__res250only_small $T=5710 1135 0 0 $X=5710 $Y=1135
X260 TIE_WEAK_HI_H 63 sky130_fd_io__res250only_small $T=66435 137450 0 180 $X=55085 $Y=135430
X261 54 51 sky130_fd_pr__res_bent_po__example_5595914180862 $T=11875 43685 1 180 $X=5605 $Y=43685
X262 57 54 sky130_fd_pr__res_bent_po__example_5595914180862 $T=18585 43685 1 180 $X=12315 $Y=43685
X263 62 61 sky130_fd_pr__res_bent_po__example_5595914180862 $T=49010 130505 0 180 $X=42740 $Y=129705
X264 64 62 sky130_fd_pr__res_bent_po__example_5595914180862 $T=55720 130505 0 180 $X=49450 $Y=129705
X265 57 9 sky130_fd_pr__res_bent_po__example_5595914180863 $T=19445 44485 1 0 $X=19175 $Y=43685
X266 61 21 sky130_fd_pr__res_bent_po__example_5595914180863 $T=52600 133880 0 180 $X=40330 $Y=133080
X269 VSSD VDDIO_Q 69 27 70 71 72 73 74 75 76 77 78 82 sky130_fd_io__xres2v2_rcfilter_lpfv2 $T=73595 4860 0 90 $X=33055 $Y=6020
X301 VDDIO_Q INP_SEL_H 37 82 sky130_fd_pr__pfet_01v8__example_55959141808767 $T=21265 10040 1 90 $X=20935 $Y=9430
X302 VDDIO_Q 23 82 FILT_IN_H sky130_fd_pr__pfet_01v8__example_55959141808767 $T=21265 11470 1 90 $X=20935 $Y=10860
X303 VSSIO TIE_LO_ESD sky130_fd_io__tk_tie_r_out_esd $T=17060 2635 0 0 $X=17450 $Y=3730
X304 VDDIO TIE_HI_ESD sky130_fd_io__tk_tie_r_out_esd $T=17060 3875 0 0 $X=17450 $Y=4970
X305 VSSD 23 37 82 sky130_fd_pr__nfet_01v8__example_55959141808764 $T=20005 10040 0 90 $X=16825 $Y=9580
X306 VSSD INP_SEL_H 82 FILT_IN_H sky130_fd_pr__nfet_01v8__example_55959141808764 $T=20005 11470 0 90 $X=16825 $Y=11010
X307 VSSD 11 50 44 sky130_fd_pr__nfet_01v8__example_55959141808779 $T=13635 35115 1 90 $X=13455 $Y=34655
X308 VSSD 17 45 5 sky130_fd_pr__nfet_01v8__example_55959141808779 $T=16525 17790 1 270 $X=15345 $Y=16430
X309 VSSD 13 12 sky130_fd_pr__nfet_01v8__example_55959141808777 $T=18315 20005 1 270 $X=15135 $Y=19045
X310 VSSD 20 22 sky130_fd_pr__nfet_01v8__example_55959141808777 $T=18390 25165 1 270 $X=15210 $Y=24205
X311 VSSD ENABLE_H 41 sky130_fd_pr__nfet_01v8__example_55959141808777 $T=18390 26580 1 270 $X=15210 $Y=25620
X327 4 4 4 sky130_fd_pr__pfet_01v8__example_55959141808784 $T=8380 11155 1 270 $X=7050 $Y=9745
X328 4 11 20 sky130_fd_pr__pfet_01v8__example_55959141808784 $T=10910 10355 0 90 $X=9580 $Y=9745
X348 VSSD VDDIO VSSD 11 PAD sky130_fd_io__gpio_buf_localesdv2 $T=4630 70965 1 0 $X=4923 $Y=47395
X351 VSSD 92 VSSIO VDDIO 92 92 80 PAD sky130_fd_io__gpio_pddrvr_strong_xres4v2 $T=0 184810 1 0 $X=-515 $Y=137270
.ENDS
***************************************
