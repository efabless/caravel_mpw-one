* SPICE NETLIST
***************************************

.SUBCKT drainOnly g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808671
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808672
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808673 2 3 4
** N=4 EP=3 IP=12 FDC=22
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
M18 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=41400 $Y=0 $D=49
M19 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=43410 $Y=0 $D=49
M20 4 3 2 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=46000 $Y=0 $D=49
M21 2 3 4 2 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=48010 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808663
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2 2 3 4
** N=5 EP=3 IP=26 FDC=22
*.SEEDPROM
X0 2 3 4 sky130_fd_pr__nfet_01v8__example_55959141808673 $T=0 0 0 0 $X=-1575 $Y=-180
.ENDS
***************************************
.SUBCKT ICV_3 2 3 4
** N=5 EP=3 IP=26 FDC=22
*.SEEDPROM
X0 2 3 4 sky130_fd_pr__nfet_01v8__example_55959141808673 $T=0 0 0 0 $X=-1575 $Y=-180
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808670 1 2 3
** N=3 EP=3 IP=10 FDC=18
M0 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 3 2 1 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 1 2 3 1 nhv L=0.5 W=20 m=1 r=40 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_4 2 3 4
** N=5 EP=3 IP=21 FDC=18
*.SEEDPROM
X9 2 3 4 sky130_fd_pr__nfet_01v8__example_55959141808670 $T=0 0 0 0 $X=-1575 $Y=-180
.ENDS
***************************************
.SUBCKT ICV_5 2 3 4
** N=5 EP=3 IP=21 FDC=18
*.SEEDPROM
X9 2 3 4 sky130_fd_pr__nfet_01v8__example_55959141808670 $T=0 0 0 0 $X=-1575 $Y=-180
.ENDS
***************************************
.SUBCKT ICV_6 2 3 4
** N=4 EP=3 IP=21 FDC=18
*.SEEDPROM
X9 2 3 4 sky130_fd_pr__nfet_01v8__example_55959141808670 $T=0 0 0 0 $X=-1575 $Y=-180
.ENDS
***************************************
.SUBCKT ICV_7 2 3 4
** N=10 EP=3 IP=26 FDC=22
*.SEEDPROM
X0 2 3 4 sky130_fd_pr__nfet_01v8__example_55959141808673 $T=0 0 0 0 $X=-1575 $Y=-180
.ENDS
***************************************
.SUBCKT ICV_8
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_9
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_10
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_11
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_12
** N=10 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_13
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_14
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808676
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808675
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808662
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15 2 3 4
** N=5 EP=3 IP=4 FDC=3
*.SEEDPROM
M0 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-64395 $D=49
M1 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-62385 $D=49
M2 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-59795 $D=49
.ENDS
***************************************
.SUBCKT ICV_16
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_17
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_5595914180851
** N=1 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 1 2
** N=2 EP=2 IP=2 FDC=1
M0 1 2 1 1 nhv L=4 W=5 m=1 r=1.25 a=20 p=18 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_io__sio_clamp_pcap_4x5 1 2
** N=2 EP=2 IP=2 FDC=1
X0 1 2 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=1145 720 0 0 $X=700 $Y=540
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808679
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808678
** N=2 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 2 4 5
** N=8 EP=3 IP=22 FDC=10
*.SEEDPROM
M0 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-66335 $D=49
M1 5 4 2 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-65555 $D=49
M2 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-64775 $D=49
M3 5 4 2 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-63995 $D=49
M4 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-63215 $D=49
M5 5 4 2 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-62435 $D=49
M6 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-61655 $D=49
M7 5 4 2 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-60875 $D=49
M8 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-60095 $D=49
X9 2 4 sky130_fd_io__sio_clamp_pcap_4x5 $T=25830 -68720 0 90 $X=19080 $Y=-68720
.ENDS
***************************************
.SUBCKT sky130_fd_io__esd_rcclamp_nfetcap 2 3
** N=4 EP=2 IP=2 FDC=1
*.SEEDPROM
M0 2 3 2 2 nhv L=8 W=5 m=1 r=0.625 a=40 p=26 mult=1 $X=895 $Y=630 $D=49
.ENDS
***************************************
.SUBCKT ICV_19 2 4
** N=7 EP=2 IP=12 FDC=3
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=7080 -68470 0 90 $X=420 $Y=-68720
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=13300 -68470 0 90 $X=6640 $Y=-68720
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=19520 -68470 0 90 $X=12860 $Y=-68720
.ENDS
***************************************
.SUBCKT ICV_20 2 3 4
** N=5 EP=3 IP=8 FDC=4
*.SEEDPROM
M0 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-57785 $D=49
M1 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-55195 $D=49
M2 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-53185 $D=49
M3 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-50595 $D=49
.ENDS
***************************************
.SUBCKT ICV_21 2 4 5
** N=8 EP=3 IP=12 FDC=5
*.SEEDPROM
M0 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-58535 $D=49
M1 5 4 2 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-57755 $D=49
M2 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-56975 $D=49
M3 5 4 2 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-56195 $D=49
M4 2 4 5 2 nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30545 $Y=-55415 $D=49
.ENDS
***************************************
.SUBCKT ICV_22 2 4
** N=7 EP=2 IP=12 FDC=3
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=7080 -58710 0 90 $X=420 $Y=-58960
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=13300 -58710 0 90 $X=6640 $Y=-58960
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=19520 -58710 0 90 $X=12860 $Y=-58960
.ENDS
***************************************
.SUBCKT ICV_23 2 3 4
** N=5 EP=3 IP=6 FDC=4
*.SEEDPROM
M0 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-48585 $D=49
M1 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-45995 $D=49
M2 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-43985 $D=49
M3 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-41395 $D=49
.ENDS
***************************************
.SUBCKT ICV_24
** N=8 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_25 2 4
** N=7 EP=2 IP=12 FDC=3
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=7080 -48950 0 90 $X=420 $Y=-49200
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=13300 -48950 0 90 $X=6640 $Y=-49200
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=19520 -48950 0 90 $X=12860 $Y=-49200
.ENDS
***************************************
.SUBCKT ICV_26 2 3 4
** N=5 EP=3 IP=15 FDC=10
*.SEEDPROM
M0 2 4 3 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=17895 $Y=183145 $D=49
M1 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=20485 $Y=183145 $D=49
M2 2 4 3 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=22495 $Y=183145 $D=49
M3 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=25085 $Y=183145 $D=49
M4 2 4 3 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=27095 $Y=183145 $D=49
M5 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=29685 $Y=183145 $D=49
M6 2 4 3 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=31695 $Y=183145 $D=49
M7 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=34285 $Y=183145 $D=49
M8 2 4 3 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=36295 $Y=183145 $D=49
M9 3 4 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=38885 $Y=183145 $D=49
.ENDS
***************************************
.SUBCKT ICV_27
** N=5 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_28
** N=4 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_29
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_30 2 4
** N=7 EP=2 IP=24 FDC=6
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=29430 7080 0 180 $X=19390 $Y=420
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=29430 13300 0 180 $X=19390 $Y=6640
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=29430 19520 0 180 $X=19390 $Y=12860
X3 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=39190 7080 0 180 $X=29150 $Y=420
X4 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=39190 13300 0 180 $X=29150 $Y=6640
X5 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=39190 19520 0 180 $X=29150 $Y=12860
.ENDS
***************************************
.SUBCKT ICV_31 2 3 6
** N=7 EP=3 IP=1 FDC=1
*.SEEDPROM
M0 3 6 2 2 nhv L=0.5 W=10 m=1 r=20 a=5 p=21 mult=1 $X=183145 $Y=-16385 $D=49
.ENDS
***************************************
.SUBCKT ICV_32
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_33
** N=7 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_34
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_35
** N=12 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_36
** N=9 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_37
** N=6 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808336
** N=2 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808666
** N=3 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_38
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_39
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_40
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_41
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1 2 3 4
** N=7 EP=3 IP=16 FDC=50
*.SEEDPROM
M0 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=0 $Y=0 $D=109
M1 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=780 $Y=0 $D=109
M2 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=1560 $Y=0 $D=109
M3 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=2340 $Y=0 $D=109
M4 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=3120 $Y=0 $D=109
M5 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=3900 $Y=0 $D=109
M6 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=4680 $Y=0 $D=109
M7 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=5460 $Y=0 $D=109
M8 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=6240 $Y=0 $D=109
M9 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=7020 $Y=0 $D=109
M10 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=7800 $Y=0 $D=109
M11 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=8580 $Y=0 $D=109
M12 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=9360 $Y=0 $D=109
M13 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=10140 $Y=0 $D=109
M14 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=10920 $Y=0 $D=109
M15 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=11700 $Y=0 $D=109
M16 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=12480 $Y=0 $D=109
M17 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=13260 $Y=0 $D=109
M18 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=14040 $Y=0 $D=109
M19 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=14820 $Y=0 $D=109
M20 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=15600 $Y=0 $D=109
M21 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=16380 $Y=0 $D=109
M22 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=17160 $Y=0 $D=109
M23 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=17940 $Y=0 $D=109
M24 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=18720 $Y=0 $D=109
M25 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=19500 $Y=0 $D=109
M26 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=20280 $Y=0 $D=109
M27 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=21060 $Y=0 $D=109
M28 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=21840 $Y=0 $D=109
M29 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=22620 $Y=0 $D=109
M30 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=23400 $Y=0 $D=109
M31 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=24180 $Y=0 $D=109
M32 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=24960 $Y=0 $D=109
M33 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=25740 $Y=0 $D=109
M34 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=26520 $Y=0 $D=109
M35 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=27300 $Y=0 $D=109
M36 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=28080 $Y=0 $D=109
M37 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=28860 $Y=0 $D=109
M38 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=29640 $Y=0 $D=109
M39 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=30420 $Y=0 $D=109
M40 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=31200 $Y=0 $D=109
M41 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=31980 $Y=0 $D=109
M42 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=32760 $Y=0 $D=109
M43 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=33540 $Y=0 $D=109
M44 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=34320 $Y=0 $D=109
M45 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=35100 $Y=0 $D=109
M46 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=35880 $Y=0 $D=109
M47 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=36660 $Y=0 $D=109
M48 4 3 2 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=37440 $Y=0 $D=109
M49 2 3 4 2 phv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=38220 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad VSSD VSSIO VDDIO 8 AMUXBUS_B 10 AMUXBUS_A 12 VSSIO_Q VSWITCH VSSA VCCHIB VCCD VDDA 19
** N=19 EP=15 IP=241 FDC=241
R0 VDDIO 19 0.01 m=1 $[short] $X=6670 $Y=103310 $D=269
M1 VSSIO 5 4 VSSIO nhv L=0.5 W=7 m=1 r=14 a=3.5 p=15 mult=1 $X=58815 $Y=30545 $D=49
X2 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=19700 $D=150
X3 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=43275 $D=150
X4 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=64770 $Y=38800 $D=150
X5 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=68375 $Y=195640 $D=150
R6 6 5 L=470 W=0.33 m=1 $[mrp1] $X=70725 $Y=39980 $D=250
R7 7 VDDIO L=700 W=0.33 m=1 $[mrp1] $X=9500 $Y=72320 $D=250
R8 7 6 L=1550 W=0.33 m=1 $[mrp1] $X=1070 $Y=41405 $D=250
X9 VSSD VDDIO Dpar a=126.766 p=0 m=1 $[nwdiode] $X=8835 $Y=41140 $D=183
X10 VSSIO VDDIO Dpar a=8184.99 p=443.22 m=1 $[dnwdiode_pw] $X=10695 $Y=43000 $D=188
X11 VSSIO VDDIO Dpar a=1172.63 p=163 m=1 $[dnwdiode_pw] $X=13380 $Y=170 $D=188
X12 VSSIO VDDIO Dpar a=137.463 p=47.72 m=1 $[dnwdiode_pw] $X=53530 $Y=29360 $D=188
X13 VSSD VDDIO Dpar a=10358.7 p=619.08 m=1 $[dnwdiode_psub] $X=9500 $Y=131800 $D=187
X14 VSSD VDDIO Dpar a=369.745 p=100.13 m=1 $[nwdiode] $X=5200 $Y=26890 $D=185
X15 VSSIO 4 VDDIO ICV_2 $T=15885 160145 0 0 $X=14310 $Y=159965
X16 VSSIO 4 VDDIO ICV_3 $T=15885 137145 0 0 $X=14310 $Y=136965
X17 VSSIO 4 VDDIO ICV_4 $T=25085 114145 0 0 $X=23510 $Y=113965
X18 VSSIO 4 VDDIO ICV_5 $T=25085 91145 0 0 $X=23510 $Y=90965
X19 VSSIO 4 VDDIO ICV_6 $T=25085 68145 0 0 $X=23510 $Y=67965
X20 VSSIO 4 VDDIO ICV_7 $T=15885 45145 0 0 $X=14310 $Y=44965
X28 VSSIO VDDIO 4 ICV_15 $T=0 0 0 90 $X=59000 $Y=157100
X31 VSSIO 5 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=61815 25110 0 180 $X=57370 $Y=19930
X32 VSSIO 5 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 7170 0 180 $X=13630 $Y=420
X33 VSSIO 5 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 13390 0 180 $X=13630 $Y=6640
X34 VSSIO 5 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 19610 0 180 $X=13630 $Y=12860
X35 VSSIO 5 4 ICV_18 $T=0 0 0 90 $X=59000 $Y=19080
X36 VSSIO 5 ICV_19 $T=0 0 0 90 $X=58430 $Y=-2035
X37 VSSIO VDDIO 4 ICV_20 $T=0 0 0 90 $X=48900 $Y=157325
X38 VSSIO 5 4 ICV_21 $T=0 0 0 90 $X=48900 $Y=19600
X39 VSSIO 5 ICV_22 $T=0 0 0 90 $X=48670 $Y=-2035
X40 VSSIO VDDIO 4 ICV_23 $T=0 0 0 90 $X=39700 $Y=157325
X42 VSSIO 5 ICV_25 $T=0 0 0 90 $X=38910 $Y=-2035
X43 VSSIO VDDIO 4 ICV_26 $T=0 0 0 0 $X=16700 $Y=157325
X47 VSSIO 5 ICV_30 $T=0 0 0 0 $X=16700 $Y=-2035
X48 VSSIO VDDIO 4 ICV_31 $T=0 0 0 90 $X=0 $Y=157100
X55 VDDIO 5 4 ICV_1 $T=6340 27765 0 0 $X=5745 $Y=27435
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
*.CALIBRE WARNING OPEN Open circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
