* NGSPICE file created from mgmt_protect.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_1 abstract view
.subckt sky130_fd_sc_hd__and2_1 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2b_1 abstract view
.subckt sky130_fd_sc_hd__and2b_1 A_N B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_8 abstract view
.subckt sky130_fd_sc_hd__inv_8 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_8 abstract view
.subckt sky130_fd_sc_hd__buf_8 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for mprj2_logic_high abstract view
.subckt mprj2_logic_high HI vccd2 vssd2
.ends

* Black-box entry subcircuit for mprj_logic_high abstract view
.subckt mprj_logic_high HI[0] HI[100] HI[101] HI[102] HI[103] HI[104] HI[105] HI[106]
+ HI[107] HI[108] HI[109] HI[10] HI[110] HI[111] HI[112] HI[113] HI[114] HI[115] HI[116]
+ HI[117] HI[118] HI[119] HI[11] HI[120] HI[121] HI[122] HI[123] HI[124] HI[125] HI[126]
+ HI[127] HI[128] HI[129] HI[12] HI[130] HI[131] HI[132] HI[133] HI[134] HI[135] HI[136]
+ HI[137] HI[138] HI[139] HI[13] HI[140] HI[141] HI[142] HI[143] HI[144] HI[145] HI[146]
+ HI[147] HI[148] HI[149] HI[14] HI[150] HI[151] HI[152] HI[153] HI[154] HI[155] HI[156]
+ HI[157] HI[158] HI[159] HI[15] HI[160] HI[161] HI[162] HI[163] HI[164] HI[165] HI[166]
+ HI[167] HI[168] HI[169] HI[16] HI[170] HI[171] HI[172] HI[173] HI[174] HI[175] HI[176]
+ HI[177] HI[178] HI[179] HI[17] HI[180] HI[181] HI[182] HI[183] HI[184] HI[185] HI[186]
+ HI[187] HI[188] HI[189] HI[18] HI[190] HI[191] HI[192] HI[193] HI[194] HI[195] HI[196]
+ HI[197] HI[198] HI[199] HI[19] HI[1] HI[200] HI[201] HI[202] HI[203] HI[204] HI[205]
+ HI[206] HI[207] HI[208] HI[209] HI[20] HI[210] HI[211] HI[212] HI[213] HI[214] HI[215]
+ HI[216] HI[217] HI[218] HI[219] HI[21] HI[220] HI[221] HI[222] HI[223] HI[224] HI[225]
+ HI[226] HI[227] HI[228] HI[229] HI[22] HI[230] HI[231] HI[232] HI[233] HI[234] HI[235]
+ HI[236] HI[237] HI[238] HI[239] HI[23] HI[240] HI[241] HI[242] HI[243] HI[244] HI[245]
+ HI[246] HI[247] HI[248] HI[249] HI[24] HI[250] HI[251] HI[252] HI[253] HI[254] HI[255]
+ HI[256] HI[257] HI[258] HI[259] HI[25] HI[260] HI[261] HI[262] HI[263] HI[264] HI[265]
+ HI[266] HI[267] HI[268] HI[269] HI[26] HI[270] HI[271] HI[272] HI[273] HI[274] HI[275]
+ HI[276] HI[277] HI[278] HI[279] HI[27] HI[280] HI[281] HI[282] HI[283] HI[284] HI[285]
+ HI[286] HI[287] HI[288] HI[289] HI[28] HI[290] HI[291] HI[292] HI[293] HI[294] HI[295]
+ HI[296] HI[297] HI[298] HI[299] HI[29] HI[2] HI[300] HI[301] HI[302] HI[303] HI[304]
+ HI[305] HI[306] HI[307] HI[308] HI[309] HI[30] HI[310] HI[311] HI[312] HI[313] HI[314]
+ HI[315] HI[316] HI[317] HI[318] HI[319] HI[31] HI[320] HI[321] HI[322] HI[323] HI[324]
+ HI[325] HI[326] HI[327] HI[328] HI[329] HI[32] HI[330] HI[331] HI[332] HI[333] HI[334]
+ HI[335] HI[336] HI[337] HI[338] HI[339] HI[33] HI[340] HI[341] HI[342] HI[343] HI[344]
+ HI[345] HI[346] HI[347] HI[348] HI[349] HI[34] HI[350] HI[351] HI[352] HI[353] HI[354]
+ HI[355] HI[356] HI[357] HI[358] HI[359] HI[35] HI[360] HI[361] HI[362] HI[363] HI[364]
+ HI[365] HI[366] HI[367] HI[368] HI[369] HI[36] HI[370] HI[371] HI[372] HI[373] HI[374]
+ HI[375] HI[376] HI[377] HI[378] HI[379] HI[37] HI[380] HI[381] HI[382] HI[383] HI[384]
+ HI[385] HI[386] HI[387] HI[388] HI[389] HI[38] HI[390] HI[391] HI[392] HI[393] HI[394]
+ HI[395] HI[396] HI[397] HI[398] HI[399] HI[39] HI[3] HI[400] HI[401] HI[402] HI[403]
+ HI[404] HI[405] HI[406] HI[407] HI[408] HI[409] HI[40] HI[410] HI[411] HI[412] HI[413]
+ HI[414] HI[415] HI[416] HI[417] HI[418] HI[419] HI[41] HI[420] HI[421] HI[422] HI[423]
+ HI[424] HI[425] HI[426] HI[427] HI[428] HI[429] HI[42] HI[430] HI[431] HI[432] HI[433]
+ HI[434] HI[435] HI[436] HI[437] HI[438] HI[439] HI[43] HI[440] HI[441] HI[442] HI[443]
+ HI[444] HI[445] HI[446] HI[447] HI[448] HI[449] HI[44] HI[450] HI[451] HI[452] HI[453]
+ HI[454] HI[455] HI[456] HI[457] HI[458] HI[459] HI[45] HI[460] HI[461] HI[46] HI[47]
+ HI[48] HI[49] HI[4] HI[50] HI[51] HI[52] HI[53] HI[54] HI[55] HI[56] HI[57] HI[58]
+ HI[59] HI[5] HI[60] HI[61] HI[62] HI[63] HI[64] HI[65] HI[66] HI[67] HI[68] HI[69]
+ HI[6] HI[70] HI[71] HI[72] HI[73] HI[74] HI[75] HI[76] HI[77] HI[78] HI[79] HI[7]
+ HI[80] HI[81] HI[82] HI[83] HI[84] HI[85] HI[86] HI[87] HI[88] HI[89] HI[8] HI[90]
+ HI[91] HI[92] HI[93] HI[94] HI[95] HI[96] HI[97] HI[98] HI[99] HI[9] vccd1 vssd1
.ends

* Black-box entry subcircuit for mgmt_protect_hv abstract view
.subckt mgmt_protect_hv mprj2_vdd_logic1 mprj_vdd_logic1 vccd vssd vdda1 vssa1 vdda2
+ vssa2
.ends

.subckt mgmt_protect caravel_clk caravel_clk2 caravel_rstn la_data_in_core[0] la_data_in_core[100]
+ la_data_in_core[101] la_data_in_core[102] la_data_in_core[103] la_data_in_core[104]
+ la_data_in_core[105] la_data_in_core[106] la_data_in_core[107] la_data_in_core[108]
+ la_data_in_core[109] la_data_in_core[10] la_data_in_core[110] la_data_in_core[111]
+ la_data_in_core[112] la_data_in_core[113] la_data_in_core[114] la_data_in_core[115]
+ la_data_in_core[116] la_data_in_core[117] la_data_in_core[118] la_data_in_core[119]
+ la_data_in_core[11] la_data_in_core[120] la_data_in_core[121] la_data_in_core[122]
+ la_data_in_core[123] la_data_in_core[124] la_data_in_core[125] la_data_in_core[126]
+ la_data_in_core[127] la_data_in_core[12] la_data_in_core[13] la_data_in_core[14]
+ la_data_in_core[15] la_data_in_core[16] la_data_in_core[17] la_data_in_core[18]
+ la_data_in_core[19] la_data_in_core[1] la_data_in_core[20] la_data_in_core[21] la_data_in_core[22]
+ la_data_in_core[23] la_data_in_core[24] la_data_in_core[25] la_data_in_core[26]
+ la_data_in_core[27] la_data_in_core[28] la_data_in_core[29] la_data_in_core[2] la_data_in_core[30]
+ la_data_in_core[31] la_data_in_core[32] la_data_in_core[33] la_data_in_core[34]
+ la_data_in_core[35] la_data_in_core[36] la_data_in_core[37] la_data_in_core[38]
+ la_data_in_core[39] la_data_in_core[3] la_data_in_core[40] la_data_in_core[41] la_data_in_core[42]
+ la_data_in_core[43] la_data_in_core[44] la_data_in_core[45] la_data_in_core[46]
+ la_data_in_core[47] la_data_in_core[48] la_data_in_core[49] la_data_in_core[4] la_data_in_core[50]
+ la_data_in_core[51] la_data_in_core[52] la_data_in_core[53] la_data_in_core[54]
+ la_data_in_core[55] la_data_in_core[56] la_data_in_core[57] la_data_in_core[58]
+ la_data_in_core[59] la_data_in_core[5] la_data_in_core[60] la_data_in_core[61] la_data_in_core[62]
+ la_data_in_core[63] la_data_in_core[64] la_data_in_core[65] la_data_in_core[66]
+ la_data_in_core[67] la_data_in_core[68] la_data_in_core[69] la_data_in_core[6] la_data_in_core[70]
+ la_data_in_core[71] la_data_in_core[72] la_data_in_core[73] la_data_in_core[74]
+ la_data_in_core[75] la_data_in_core[76] la_data_in_core[77] la_data_in_core[78]
+ la_data_in_core[79] la_data_in_core[7] la_data_in_core[80] la_data_in_core[81] la_data_in_core[82]
+ la_data_in_core[83] la_data_in_core[84] la_data_in_core[85] la_data_in_core[86]
+ la_data_in_core[87] la_data_in_core[88] la_data_in_core[89] la_data_in_core[8] la_data_in_core[90]
+ la_data_in_core[91] la_data_in_core[92] la_data_in_core[93] la_data_in_core[94]
+ la_data_in_core[95] la_data_in_core[96] la_data_in_core[97] la_data_in_core[98]
+ la_data_in_core[99] la_data_in_core[9] la_data_in_mprj[0] la_data_in_mprj[100] la_data_in_mprj[101]
+ la_data_in_mprj[102] la_data_in_mprj[103] la_data_in_mprj[104] la_data_in_mprj[105]
+ la_data_in_mprj[106] la_data_in_mprj[107] la_data_in_mprj[108] la_data_in_mprj[109]
+ la_data_in_mprj[10] la_data_in_mprj[110] la_data_in_mprj[111] la_data_in_mprj[112]
+ la_data_in_mprj[113] la_data_in_mprj[114] la_data_in_mprj[115] la_data_in_mprj[116]
+ la_data_in_mprj[117] la_data_in_mprj[118] la_data_in_mprj[119] la_data_in_mprj[11]
+ la_data_in_mprj[120] la_data_in_mprj[121] la_data_in_mprj[122] la_data_in_mprj[123]
+ la_data_in_mprj[124] la_data_in_mprj[125] la_data_in_mprj[126] la_data_in_mprj[127]
+ la_data_in_mprj[12] la_data_in_mprj[13] la_data_in_mprj[14] la_data_in_mprj[15]
+ la_data_in_mprj[16] la_data_in_mprj[17] la_data_in_mprj[18] la_data_in_mprj[19]
+ la_data_in_mprj[1] la_data_in_mprj[20] la_data_in_mprj[21] la_data_in_mprj[22] la_data_in_mprj[23]
+ la_data_in_mprj[24] la_data_in_mprj[25] la_data_in_mprj[26] la_data_in_mprj[27]
+ la_data_in_mprj[28] la_data_in_mprj[29] la_data_in_mprj[2] la_data_in_mprj[30] la_data_in_mprj[31]
+ la_data_in_mprj[32] la_data_in_mprj[33] la_data_in_mprj[34] la_data_in_mprj[35]
+ la_data_in_mprj[36] la_data_in_mprj[37] la_data_in_mprj[38] la_data_in_mprj[39]
+ la_data_in_mprj[3] la_data_in_mprj[40] la_data_in_mprj[41] la_data_in_mprj[42] la_data_in_mprj[43]
+ la_data_in_mprj[44] la_data_in_mprj[45] la_data_in_mprj[46] la_data_in_mprj[47]
+ la_data_in_mprj[48] la_data_in_mprj[49] la_data_in_mprj[4] la_data_in_mprj[50] la_data_in_mprj[51]
+ la_data_in_mprj[52] la_data_in_mprj[53] la_data_in_mprj[54] la_data_in_mprj[55]
+ la_data_in_mprj[56] la_data_in_mprj[57] la_data_in_mprj[58] la_data_in_mprj[59]
+ la_data_in_mprj[5] la_data_in_mprj[60] la_data_in_mprj[61] la_data_in_mprj[62] la_data_in_mprj[63]
+ la_data_in_mprj[64] la_data_in_mprj[65] la_data_in_mprj[66] la_data_in_mprj[67]
+ la_data_in_mprj[68] la_data_in_mprj[69] la_data_in_mprj[6] la_data_in_mprj[70] la_data_in_mprj[71]
+ la_data_in_mprj[72] la_data_in_mprj[73] la_data_in_mprj[74] la_data_in_mprj[75]
+ la_data_in_mprj[76] la_data_in_mprj[77] la_data_in_mprj[78] la_data_in_mprj[79]
+ la_data_in_mprj[7] la_data_in_mprj[80] la_data_in_mprj[81] la_data_in_mprj[82] la_data_in_mprj[83]
+ la_data_in_mprj[84] la_data_in_mprj[85] la_data_in_mprj[86] la_data_in_mprj[87]
+ la_data_in_mprj[88] la_data_in_mprj[89] la_data_in_mprj[8] la_data_in_mprj[90] la_data_in_mprj[91]
+ la_data_in_mprj[92] la_data_in_mprj[93] la_data_in_mprj[94] la_data_in_mprj[95]
+ la_data_in_mprj[96] la_data_in_mprj[97] la_data_in_mprj[98] la_data_in_mprj[99]
+ la_data_in_mprj[9] la_data_out_core[0] la_data_out_core[100] la_data_out_core[101]
+ la_data_out_core[102] la_data_out_core[103] la_data_out_core[104] la_data_out_core[105]
+ la_data_out_core[106] la_data_out_core[107] la_data_out_core[108] la_data_out_core[109]
+ la_data_out_core[10] la_data_out_core[110] la_data_out_core[111] la_data_out_core[112]
+ la_data_out_core[113] la_data_out_core[114] la_data_out_core[115] la_data_out_core[116]
+ la_data_out_core[117] la_data_out_core[118] la_data_out_core[119] la_data_out_core[11]
+ la_data_out_core[120] la_data_out_core[121] la_data_out_core[122] la_data_out_core[123]
+ la_data_out_core[124] la_data_out_core[125] la_data_out_core[126] la_data_out_core[127]
+ la_data_out_core[12] la_data_out_core[13] la_data_out_core[14] la_data_out_core[15]
+ la_data_out_core[16] la_data_out_core[17] la_data_out_core[18] la_data_out_core[19]
+ la_data_out_core[1] la_data_out_core[20] la_data_out_core[21] la_data_out_core[22]
+ la_data_out_core[23] la_data_out_core[24] la_data_out_core[25] la_data_out_core[26]
+ la_data_out_core[27] la_data_out_core[28] la_data_out_core[29] la_data_out_core[2]
+ la_data_out_core[30] la_data_out_core[31] la_data_out_core[32] la_data_out_core[33]
+ la_data_out_core[34] la_data_out_core[35] la_data_out_core[36] la_data_out_core[37]
+ la_data_out_core[38] la_data_out_core[39] la_data_out_core[3] la_data_out_core[40]
+ la_data_out_core[41] la_data_out_core[42] la_data_out_core[43] la_data_out_core[44]
+ la_data_out_core[45] la_data_out_core[46] la_data_out_core[47] la_data_out_core[48]
+ la_data_out_core[49] la_data_out_core[4] la_data_out_core[50] la_data_out_core[51]
+ la_data_out_core[52] la_data_out_core[53] la_data_out_core[54] la_data_out_core[55]
+ la_data_out_core[56] la_data_out_core[57] la_data_out_core[58] la_data_out_core[59]
+ la_data_out_core[5] la_data_out_core[60] la_data_out_core[61] la_data_out_core[62]
+ la_data_out_core[63] la_data_out_core[64] la_data_out_core[65] la_data_out_core[66]
+ la_data_out_core[67] la_data_out_core[68] la_data_out_core[69] la_data_out_core[6]
+ la_data_out_core[70] la_data_out_core[71] la_data_out_core[72] la_data_out_core[73]
+ la_data_out_core[74] la_data_out_core[75] la_data_out_core[76] la_data_out_core[77]
+ la_data_out_core[78] la_data_out_core[79] la_data_out_core[7] la_data_out_core[80]
+ la_data_out_core[81] la_data_out_core[82] la_data_out_core[83] la_data_out_core[84]
+ la_data_out_core[85] la_data_out_core[86] la_data_out_core[87] la_data_out_core[88]
+ la_data_out_core[89] la_data_out_core[8] la_data_out_core[90] la_data_out_core[91]
+ la_data_out_core[92] la_data_out_core[93] la_data_out_core[94] la_data_out_core[95]
+ la_data_out_core[96] la_data_out_core[97] la_data_out_core[98] la_data_out_core[99]
+ la_data_out_core[9] la_data_out_mprj[0] la_data_out_mprj[100] la_data_out_mprj[101]
+ la_data_out_mprj[102] la_data_out_mprj[103] la_data_out_mprj[104] la_data_out_mprj[105]
+ la_data_out_mprj[106] la_data_out_mprj[107] la_data_out_mprj[108] la_data_out_mprj[109]
+ la_data_out_mprj[10] la_data_out_mprj[110] la_data_out_mprj[111] la_data_out_mprj[112]
+ la_data_out_mprj[113] la_data_out_mprj[114] la_data_out_mprj[115] la_data_out_mprj[116]
+ la_data_out_mprj[117] la_data_out_mprj[118] la_data_out_mprj[119] la_data_out_mprj[11]
+ la_data_out_mprj[120] la_data_out_mprj[121] la_data_out_mprj[122] la_data_out_mprj[123]
+ la_data_out_mprj[124] la_data_out_mprj[125] la_data_out_mprj[126] la_data_out_mprj[127]
+ la_data_out_mprj[12] la_data_out_mprj[13] la_data_out_mprj[14] la_data_out_mprj[15]
+ la_data_out_mprj[16] la_data_out_mprj[17] la_data_out_mprj[18] la_data_out_mprj[19]
+ la_data_out_mprj[1] la_data_out_mprj[20] la_data_out_mprj[21] la_data_out_mprj[22]
+ la_data_out_mprj[23] la_data_out_mprj[24] la_data_out_mprj[25] la_data_out_mprj[26]
+ la_data_out_mprj[27] la_data_out_mprj[28] la_data_out_mprj[29] la_data_out_mprj[2]
+ la_data_out_mprj[30] la_data_out_mprj[31] la_data_out_mprj[32] la_data_out_mprj[33]
+ la_data_out_mprj[34] la_data_out_mprj[35] la_data_out_mprj[36] la_data_out_mprj[37]
+ la_data_out_mprj[38] la_data_out_mprj[39] la_data_out_mprj[3] la_data_out_mprj[40]
+ la_data_out_mprj[41] la_data_out_mprj[42] la_data_out_mprj[43] la_data_out_mprj[44]
+ la_data_out_mprj[45] la_data_out_mprj[46] la_data_out_mprj[47] la_data_out_mprj[48]
+ la_data_out_mprj[49] la_data_out_mprj[4] la_data_out_mprj[50] la_data_out_mprj[51]
+ la_data_out_mprj[52] la_data_out_mprj[53] la_data_out_mprj[54] la_data_out_mprj[55]
+ la_data_out_mprj[56] la_data_out_mprj[57] la_data_out_mprj[58] la_data_out_mprj[59]
+ la_data_out_mprj[5] la_data_out_mprj[60] la_data_out_mprj[61] la_data_out_mprj[62]
+ la_data_out_mprj[63] la_data_out_mprj[64] la_data_out_mprj[65] la_data_out_mprj[66]
+ la_data_out_mprj[67] la_data_out_mprj[68] la_data_out_mprj[69] la_data_out_mprj[6]
+ la_data_out_mprj[70] la_data_out_mprj[71] la_data_out_mprj[72] la_data_out_mprj[73]
+ la_data_out_mprj[74] la_data_out_mprj[75] la_data_out_mprj[76] la_data_out_mprj[77]
+ la_data_out_mprj[78] la_data_out_mprj[79] la_data_out_mprj[7] la_data_out_mprj[80]
+ la_data_out_mprj[81] la_data_out_mprj[82] la_data_out_mprj[83] la_data_out_mprj[84]
+ la_data_out_mprj[85] la_data_out_mprj[86] la_data_out_mprj[87] la_data_out_mprj[88]
+ la_data_out_mprj[89] la_data_out_mprj[8] la_data_out_mprj[90] la_data_out_mprj[91]
+ la_data_out_mprj[92] la_data_out_mprj[93] la_data_out_mprj[94] la_data_out_mprj[95]
+ la_data_out_mprj[96] la_data_out_mprj[97] la_data_out_mprj[98] la_data_out_mprj[99]
+ la_data_out_mprj[9] la_iena_mprj[0] la_iena_mprj[100] la_iena_mprj[101] la_iena_mprj[102]
+ la_iena_mprj[103] la_iena_mprj[104] la_iena_mprj[105] la_iena_mprj[106] la_iena_mprj[107]
+ la_iena_mprj[108] la_iena_mprj[109] la_iena_mprj[10] la_iena_mprj[110] la_iena_mprj[111]
+ la_iena_mprj[112] la_iena_mprj[113] la_iena_mprj[114] la_iena_mprj[115] la_iena_mprj[116]
+ la_iena_mprj[117] la_iena_mprj[118] la_iena_mprj[119] la_iena_mprj[11] la_iena_mprj[120]
+ la_iena_mprj[121] la_iena_mprj[122] la_iena_mprj[123] la_iena_mprj[124] la_iena_mprj[125]
+ la_iena_mprj[126] la_iena_mprj[127] la_iena_mprj[12] la_iena_mprj[13] la_iena_mprj[14]
+ la_iena_mprj[15] la_iena_mprj[16] la_iena_mprj[17] la_iena_mprj[18] la_iena_mprj[19]
+ la_iena_mprj[1] la_iena_mprj[20] la_iena_mprj[21] la_iena_mprj[22] la_iena_mprj[23]
+ la_iena_mprj[24] la_iena_mprj[25] la_iena_mprj[26] la_iena_mprj[27] la_iena_mprj[28]
+ la_iena_mprj[29] la_iena_mprj[2] la_iena_mprj[30] la_iena_mprj[31] la_iena_mprj[32]
+ la_iena_mprj[33] la_iena_mprj[34] la_iena_mprj[35] la_iena_mprj[36] la_iena_mprj[37]
+ la_iena_mprj[38] la_iena_mprj[39] la_iena_mprj[3] la_iena_mprj[40] la_iena_mprj[41]
+ la_iena_mprj[42] la_iena_mprj[43] la_iena_mprj[44] la_iena_mprj[45] la_iena_mprj[46]
+ la_iena_mprj[47] la_iena_mprj[48] la_iena_mprj[49] la_iena_mprj[4] la_iena_mprj[50]
+ la_iena_mprj[51] la_iena_mprj[52] la_iena_mprj[53] la_iena_mprj[54] la_iena_mprj[55]
+ la_iena_mprj[56] la_iena_mprj[57] la_iena_mprj[58] la_iena_mprj[59] la_iena_mprj[5]
+ la_iena_mprj[60] la_iena_mprj[61] la_iena_mprj[62] la_iena_mprj[63] la_iena_mprj[64]
+ la_iena_mprj[65] la_iena_mprj[66] la_iena_mprj[67] la_iena_mprj[68] la_iena_mprj[69]
+ la_iena_mprj[6] la_iena_mprj[70] la_iena_mprj[71] la_iena_mprj[72] la_iena_mprj[73]
+ la_iena_mprj[74] la_iena_mprj[75] la_iena_mprj[76] la_iena_mprj[77] la_iena_mprj[78]
+ la_iena_mprj[79] la_iena_mprj[7] la_iena_mprj[80] la_iena_mprj[81] la_iena_mprj[82]
+ la_iena_mprj[83] la_iena_mprj[84] la_iena_mprj[85] la_iena_mprj[86] la_iena_mprj[87]
+ la_iena_mprj[88] la_iena_mprj[89] la_iena_mprj[8] la_iena_mprj[90] la_iena_mprj[91]
+ la_iena_mprj[92] la_iena_mprj[93] la_iena_mprj[94] la_iena_mprj[95] la_iena_mprj[96]
+ la_iena_mprj[97] la_iena_mprj[98] la_iena_mprj[99] la_iena_mprj[9] la_oenb_core[0]
+ la_oenb_core[100] la_oenb_core[101] la_oenb_core[102] la_oenb_core[103] la_oenb_core[104]
+ la_oenb_core[105] la_oenb_core[106] la_oenb_core[107] la_oenb_core[108] la_oenb_core[109]
+ la_oenb_core[10] la_oenb_core[110] la_oenb_core[111] la_oenb_core[112] la_oenb_core[113]
+ la_oenb_core[114] la_oenb_core[115] la_oenb_core[116] la_oenb_core[117] la_oenb_core[118]
+ la_oenb_core[119] la_oenb_core[11] la_oenb_core[120] la_oenb_core[121] la_oenb_core[122]
+ la_oenb_core[123] la_oenb_core[124] la_oenb_core[125] la_oenb_core[126] la_oenb_core[127]
+ la_oenb_core[12] la_oenb_core[13] la_oenb_core[14] la_oenb_core[15] la_oenb_core[16]
+ la_oenb_core[17] la_oenb_core[18] la_oenb_core[19] la_oenb_core[1] la_oenb_core[20]
+ la_oenb_core[21] la_oenb_core[22] la_oenb_core[23] la_oenb_core[24] la_oenb_core[25]
+ la_oenb_core[26] la_oenb_core[27] la_oenb_core[28] la_oenb_core[29] la_oenb_core[2]
+ la_oenb_core[30] la_oenb_core[31] la_oenb_core[32] la_oenb_core[33] la_oenb_core[34]
+ la_oenb_core[35] la_oenb_core[36] la_oenb_core[37] la_oenb_core[38] la_oenb_core[39]
+ la_oenb_core[3] la_oenb_core[40] la_oenb_core[41] la_oenb_core[42] la_oenb_core[43]
+ la_oenb_core[44] la_oenb_core[45] la_oenb_core[46] la_oenb_core[47] la_oenb_core[48]
+ la_oenb_core[49] la_oenb_core[4] la_oenb_core[50] la_oenb_core[51] la_oenb_core[52]
+ la_oenb_core[53] la_oenb_core[54] la_oenb_core[55] la_oenb_core[56] la_oenb_core[57]
+ la_oenb_core[58] la_oenb_core[59] la_oenb_core[5] la_oenb_core[60] la_oenb_core[61]
+ la_oenb_core[62] la_oenb_core[63] la_oenb_core[64] la_oenb_core[65] la_oenb_core[66]
+ la_oenb_core[67] la_oenb_core[68] la_oenb_core[69] la_oenb_core[6] la_oenb_core[70]
+ la_oenb_core[71] la_oenb_core[72] la_oenb_core[73] la_oenb_core[74] la_oenb_core[75]
+ la_oenb_core[76] la_oenb_core[77] la_oenb_core[78] la_oenb_core[79] la_oenb_core[7]
+ la_oenb_core[80] la_oenb_core[81] la_oenb_core[82] la_oenb_core[83] la_oenb_core[84]
+ la_oenb_core[85] la_oenb_core[86] la_oenb_core[87] la_oenb_core[88] la_oenb_core[89]
+ la_oenb_core[8] la_oenb_core[90] la_oenb_core[91] la_oenb_core[92] la_oenb_core[93]
+ la_oenb_core[94] la_oenb_core[95] la_oenb_core[96] la_oenb_core[97] la_oenb_core[98]
+ la_oenb_core[99] la_oenb_core[9] la_oenb_mprj[0] la_oenb_mprj[100] la_oenb_mprj[101]
+ la_oenb_mprj[102] la_oenb_mprj[103] la_oenb_mprj[104] la_oenb_mprj[105] la_oenb_mprj[106]
+ la_oenb_mprj[107] la_oenb_mprj[108] la_oenb_mprj[109] la_oenb_mprj[10] la_oenb_mprj[110]
+ la_oenb_mprj[111] la_oenb_mprj[112] la_oenb_mprj[113] la_oenb_mprj[114] la_oenb_mprj[115]
+ la_oenb_mprj[116] la_oenb_mprj[117] la_oenb_mprj[118] la_oenb_mprj[119] la_oenb_mprj[11]
+ la_oenb_mprj[120] la_oenb_mprj[121] la_oenb_mprj[122] la_oenb_mprj[123] la_oenb_mprj[124]
+ la_oenb_mprj[125] la_oenb_mprj[126] la_oenb_mprj[127] la_oenb_mprj[12] la_oenb_mprj[13]
+ la_oenb_mprj[14] la_oenb_mprj[15] la_oenb_mprj[16] la_oenb_mprj[17] la_oenb_mprj[18]
+ la_oenb_mprj[19] la_oenb_mprj[1] la_oenb_mprj[20] la_oenb_mprj[21] la_oenb_mprj[22]
+ la_oenb_mprj[23] la_oenb_mprj[24] la_oenb_mprj[25] la_oenb_mprj[26] la_oenb_mprj[27]
+ la_oenb_mprj[28] la_oenb_mprj[29] la_oenb_mprj[2] la_oenb_mprj[30] la_oenb_mprj[31]
+ la_oenb_mprj[32] la_oenb_mprj[33] la_oenb_mprj[34] la_oenb_mprj[35] la_oenb_mprj[36]
+ la_oenb_mprj[37] la_oenb_mprj[38] la_oenb_mprj[39] la_oenb_mprj[3] la_oenb_mprj[40]
+ la_oenb_mprj[41] la_oenb_mprj[42] la_oenb_mprj[43] la_oenb_mprj[44] la_oenb_mprj[45]
+ la_oenb_mprj[46] la_oenb_mprj[47] la_oenb_mprj[48] la_oenb_mprj[49] la_oenb_mprj[4]
+ la_oenb_mprj[50] la_oenb_mprj[51] la_oenb_mprj[52] la_oenb_mprj[53] la_oenb_mprj[54]
+ la_oenb_mprj[55] la_oenb_mprj[56] la_oenb_mprj[57] la_oenb_mprj[58] la_oenb_mprj[59]
+ la_oenb_mprj[5] la_oenb_mprj[60] la_oenb_mprj[61] la_oenb_mprj[62] la_oenb_mprj[63]
+ la_oenb_mprj[64] la_oenb_mprj[65] la_oenb_mprj[66] la_oenb_mprj[67] la_oenb_mprj[68]
+ la_oenb_mprj[69] la_oenb_mprj[6] la_oenb_mprj[70] la_oenb_mprj[71] la_oenb_mprj[72]
+ la_oenb_mprj[73] la_oenb_mprj[74] la_oenb_mprj[75] la_oenb_mprj[76] la_oenb_mprj[77]
+ la_oenb_mprj[78] la_oenb_mprj[79] la_oenb_mprj[7] la_oenb_mprj[80] la_oenb_mprj[81]
+ la_oenb_mprj[82] la_oenb_mprj[83] la_oenb_mprj[84] la_oenb_mprj[85] la_oenb_mprj[86]
+ la_oenb_mprj[87] la_oenb_mprj[88] la_oenb_mprj[89] la_oenb_mprj[8] la_oenb_mprj[90]
+ la_oenb_mprj[91] la_oenb_mprj[92] la_oenb_mprj[93] la_oenb_mprj[94] la_oenb_mprj[95]
+ la_oenb_mprj[96] la_oenb_mprj[97] la_oenb_mprj[98] la_oenb_mprj[99] la_oenb_mprj[9]
+ mprj_adr_o_core[0] mprj_adr_o_core[10] mprj_adr_o_core[11] mprj_adr_o_core[12] mprj_adr_o_core[13]
+ mprj_adr_o_core[14] mprj_adr_o_core[15] mprj_adr_o_core[16] mprj_adr_o_core[17]
+ mprj_adr_o_core[18] mprj_adr_o_core[19] mprj_adr_o_core[1] mprj_adr_o_core[20] mprj_adr_o_core[21]
+ mprj_adr_o_core[22] mprj_adr_o_core[23] mprj_adr_o_core[24] mprj_adr_o_core[25]
+ mprj_adr_o_core[26] mprj_adr_o_core[27] mprj_adr_o_core[28] mprj_adr_o_core[29]
+ mprj_adr_o_core[2] mprj_adr_o_core[30] mprj_adr_o_core[31] mprj_adr_o_core[3] mprj_adr_o_core[4]
+ mprj_adr_o_core[5] mprj_adr_o_core[6] mprj_adr_o_core[7] mprj_adr_o_core[8] mprj_adr_o_core[9]
+ mprj_adr_o_user[0] mprj_adr_o_user[10] mprj_adr_o_user[11] mprj_adr_o_user[12] mprj_adr_o_user[13]
+ mprj_adr_o_user[14] mprj_adr_o_user[15] mprj_adr_o_user[16] mprj_adr_o_user[17]
+ mprj_adr_o_user[18] mprj_adr_o_user[19] mprj_adr_o_user[1] mprj_adr_o_user[20] mprj_adr_o_user[21]
+ mprj_adr_o_user[22] mprj_adr_o_user[23] mprj_adr_o_user[24] mprj_adr_o_user[25]
+ mprj_adr_o_user[26] mprj_adr_o_user[27] mprj_adr_o_user[28] mprj_adr_o_user[29]
+ mprj_adr_o_user[2] mprj_adr_o_user[30] mprj_adr_o_user[31] mprj_adr_o_user[3] mprj_adr_o_user[4]
+ mprj_adr_o_user[5] mprj_adr_o_user[6] mprj_adr_o_user[7] mprj_adr_o_user[8] mprj_adr_o_user[9]
+ mprj_cyc_o_core mprj_cyc_o_user mprj_dat_o_core[0] mprj_dat_o_core[10] mprj_dat_o_core[11]
+ mprj_dat_o_core[12] mprj_dat_o_core[13] mprj_dat_o_core[14] mprj_dat_o_core[15]
+ mprj_dat_o_core[16] mprj_dat_o_core[17] mprj_dat_o_core[18] mprj_dat_o_core[19]
+ mprj_dat_o_core[1] mprj_dat_o_core[20] mprj_dat_o_core[21] mprj_dat_o_core[22] mprj_dat_o_core[23]
+ mprj_dat_o_core[24] mprj_dat_o_core[25] mprj_dat_o_core[26] mprj_dat_o_core[27]
+ mprj_dat_o_core[28] mprj_dat_o_core[29] mprj_dat_o_core[2] mprj_dat_o_core[30] mprj_dat_o_core[31]
+ mprj_dat_o_core[3] mprj_dat_o_core[4] mprj_dat_o_core[5] mprj_dat_o_core[6] mprj_dat_o_core[7]
+ mprj_dat_o_core[8] mprj_dat_o_core[9] mprj_dat_o_user[0] mprj_dat_o_user[10] mprj_dat_o_user[11]
+ mprj_dat_o_user[12] mprj_dat_o_user[13] mprj_dat_o_user[14] mprj_dat_o_user[15]
+ mprj_dat_o_user[16] mprj_dat_o_user[17] mprj_dat_o_user[18] mprj_dat_o_user[19]
+ mprj_dat_o_user[1] mprj_dat_o_user[20] mprj_dat_o_user[21] mprj_dat_o_user[22] mprj_dat_o_user[23]
+ mprj_dat_o_user[24] mprj_dat_o_user[25] mprj_dat_o_user[26] mprj_dat_o_user[27]
+ mprj_dat_o_user[28] mprj_dat_o_user[29] mprj_dat_o_user[2] mprj_dat_o_user[30] mprj_dat_o_user[31]
+ mprj_dat_o_user[3] mprj_dat_o_user[4] mprj_dat_o_user[5] mprj_dat_o_user[6] mprj_dat_o_user[7]
+ mprj_dat_o_user[8] mprj_dat_o_user[9] mprj_sel_o_core[0] mprj_sel_o_core[1] mprj_sel_o_core[2]
+ mprj_sel_o_core[3] mprj_sel_o_user[0] mprj_sel_o_user[1] mprj_sel_o_user[2] mprj_sel_o_user[3]
+ mprj_stb_o_core mprj_stb_o_user mprj_we_o_core mprj_we_o_user user1_vcc_powergood
+ user1_vdd_powergood user2_vcc_powergood user2_vdd_powergood user_clock user_clock2
+ user_irq[0] user_irq[1] user_irq[2] user_irq_core[0] user_irq_core[1] user_irq_core[2]
+ user_irq_ena[0] user_irq_ena[1] user_irq_ena[2] user_reset user_resetn vccd vssd
+ vccd1 vssd1 vccd2 vssd2 vdda1 vssa1 vdda2 vssa2
XFILLER_3_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1788 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[34\]_A la_data_out_core[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[72\] la_iena_mprj[72] mprj_logic_high_inst/HI[402] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_2137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_501_ la_data_out_mprj[30] vssd vssd vccd vccd _501_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[50\] la_oenb_mprj[50] la_buf_enable\[50\]/B vssd vssd vccd vccd la_buf\[50\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_432_ mprj_adr_o_core[25] vssd vssd vccd vccd _432_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_363_ la_oenb_mprj[95] vssd vssd vccd vccd _363_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[36\] _507_/Y la_buf\[36\]/TE vssd vssd vccd vccd la_data_in_core[36] sky130_fd_sc_hd__einvp_8
XFILLER_35_1587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[108\] la_iena_mprj[108] mprj_logic_high_inst/HI[438] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[108\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_822 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[25\]_A la_data_out_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[25\] la_data_out_core[25] user_to_mprj_in_gates\[25\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[16\]_A la_data_out_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[100\]_A la_data_out_core[100] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_12_1373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_905 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_916 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_927 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_949 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_938 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[76\] _344_/Y mprj_logic_high_inst/HI[278] vssd vssd vccd
+ vccd la_oenb_core[76] sky130_fd_sc_hd__einvp_8
XFILLER_8_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[98\] la_oenb_mprj[98] la_buf_enable\[98\]/B vssd vssd vccd vccd la_buf\[98\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[24\] _463_/Y mprj_dat_buf\[24\]/TE vssd vssd vccd vccd mprj_dat_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_46_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[104\]_TE mprj_logic_high_inst/HI[306] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_415_ mprj_adr_o_core[8] vssd vssd vccd vccd _415_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_346_ la_oenb_mprj[78] vssd vssd vccd vccd _346_/Y sky130_fd_sc_hd__inv_2
XFILLER_48_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[122\]_A la_iena_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1758 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[4\] la_oenb_mprj[4] la_buf_enable\[4\]/B vssd vssd vccd vccd la_buf\[4\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[127\]_TE mprj_logic_high_inst/HI[329] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1658 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_A la_iena_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[35\] la_iena_mprj[35] mprj_logic_high_inst/HI[365] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[13\] la_oenb_mprj[13] la_buf_enable\[13\]/B vssd vssd vccd vccd la_buf\[13\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[41\]_TE la_buf\[41\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[26\]_TE mprj_logic_high_inst/HI[228] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[92\]_A_N la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[104\]_A la_iena_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[30\]_A_N la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[45\]_A_N la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[92\] la_data_out_core[92] user_to_mprj_in_gates\[92\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_44_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1862 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1822 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[49\]_TE mprj_logic_high_inst/HI[251] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[109\] _377_/Y mprj_logic_high_inst/HI[311] vssd vssd vccd
+ vccd la_oenb_core[109] sky130_fd_sc_hd__einvp_8
XFILLER_47_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[93\]_A la_iena_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_42 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_53 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[39\] _638_/Y mprj_logic_high_inst/HI[241] vssd vssd vccd
+ vccd la_oenb_core[39] sky130_fd_sc_hd__einvp_8
XFILLER_43_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_548 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_2033 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_2011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1120 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[13\]_TE mprj_dat_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__402__A mprj_we_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_A la_iena_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[62\] user_to_mprj_in_gates\[62\]/Y vssd vssd vccd vccd la_data_in_mprj[62]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[87\]_TE la_buf\[87\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[75\]_A la_iena_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_2075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[80\] la_oenb_mprj[80] la_buf_enable\[80\]/B vssd vssd vccd vccd la_buf\[80\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[66\]_A la_iena_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_594_ la_data_out_mprj[123] vssd vssd vccd vccd _594_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[66\] _537_/Y la_buf\[66\]/TE vssd vssd vccd vccd la_data_in_core[66] sky130_fd_sc_hd__einvp_8
XFILLER_45_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[122\] _593_/Y la_buf\[122\]/TE vssd vssd vccd vccd la_data_in_core[122] sky130_fd_sc_hd__einvp_8
XFILLER_6_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[57\]_A la_iena_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[55\] la_data_out_core[55] user_to_mprj_in_gates\[55\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_47_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[48\]_A la_iena_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[39\]_A la_iena_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_646_ la_oenb_mprj[47] vssd vssd vccd vccd _646_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_577_ la_data_out_mprj[106] vssd vssd vccd vccd _577_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[6\]_A _445_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_178 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[25\] user_to_mprj_in_gates\[25\]/Y vssd vssd vccd vccd la_data_in_mprj[25]
+ sky130_fd_sc_hd__inv_8
XFILLER_9_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[27\]_TE mprj_adr_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[95\]_A user_to_mprj_in_gates\[95\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[65\] la_iena_mprj[65] mprj_logic_high_inst/HI[395] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__500__A la_data_out_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1689 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_500_ la_data_out_mprj[29] vssd vssd vccd vccd _500_/Y sky130_fd_sc_hd__inv_2
X_431_ mprj_adr_o_core[24] vssd vssd vccd vccd _431_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[3\] _602_/Y mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd la_oenb_core[3] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[21\] _620_/Y mprj_logic_high_inst/HI[223] vssd vssd vccd
+ vccd la_oenb_core[21] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[43\] la_oenb_mprj[43] la_buf_enable\[43\]/B vssd vssd vccd vccd la_buf\[43\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_42_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_362_ la_oenb_mprj[94] vssd vssd vccd vccd _362_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[122\]_A _593_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[29\] _500_/Y la_buf\[29\]/TE vssd vssd vccd vccd la_data_in_core[29] sky130_fd_sc_hd__einvp_8
XFILLER_5_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__410__A mprj_adr_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1993 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_629_ la_oenb_mprj[30] vssd vssd vccd vccd _629_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[10\]_A user_to_mprj_in_gates\[10\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[18\] la_data_out_core[18] user_to_mprj_in_gates\[18\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[113\]_A _584_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_171 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[16\]_B user_to_mprj_in_gates\[16\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[82\]_TE mprj_logic_high_inst/HI[284] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_906 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_917 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_939 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_928 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_487 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[104\]_A _575_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[68\]_A user_to_mprj_in_gates\[68\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[69\] _337_/Y mprj_logic_high_inst/HI[271] vssd vssd vccd
+ vccd la_oenb_core[69] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[17\] _456_/Y mprj_dat_buf\[17\]/TE vssd vssd vccd vccd mprj_dat_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_414_ mprj_adr_o_core[7] vssd vssd vccd vccd _414_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[106\]_A user_to_mprj_in_gates\[106\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[120\] la_iena_mprj[120] mprj_logic_high_inst/HI[450] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[120\]/B sky130_fd_sc_hd__and2_1
X_345_ la_oenb_mprj[77] vssd vssd vccd vccd _345_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__405__A mprj_sel_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[59\]_A user_to_mprj_in_gates\[59\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[12\] _419_/Y mprj_adr_buf\[12\]/TE vssd vssd vccd vccd mprj_adr_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[126\] user_to_mprj_in_gates\[126\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[126] sky130_fd_sc_hd__inv_8
XANTENNA_la_buf_enable\[50\]_B la_buf_enable\[50\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[92\] user_to_mprj_in_gates\[92\]/Y vssd vssd vccd vccd la_data_in_mprj[92]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[122\]_B mprj_logic_high_inst/HI[452] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[41\]_B la_buf_enable\[41\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[113\]_B mprj_logic_high_inst/HI[443] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[28\] la_iena_mprj[28] mprj_logic_high_inst/HI[358] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[32\]_B la_buf_enable\[32\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[1\]_A la_iena_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[96\] _567_/Y la_buf\[96\]/TE vssd vssd vccd vccd la_data_in_core[96] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[1\] la_iena_mprj[1] mprj_logic_high_inst/HI[331] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[1\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[111\] la_oenb_mprj[111] la_buf_enable\[111\]/B vssd vssd vccd vccd
+ la_buf\[111\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_19_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[104\]_B mprj_logic_high_inst/HI[434] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[99\]_B la_buf_enable\[99\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[85\] la_data_out_core[85] user_to_mprj_in_gates\[85\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[23\]_B la_buf_enable\[23\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_298 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[14\]_B la_buf_enable\[14\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_1412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1110 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2023 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1121 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[7\] _478_/Y la_buf\[7\]/TE vssd vssd vccd vccd la_data_in_core[7] sky130_fd_sc_hd__einvp_8
XFILLER_4_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[11\] _482_/Y la_buf\[11\]/TE vssd vssd vccd vccd la_data_in_core[11] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[4\] _411_/Y mprj_adr_buf\[4\]/TE vssd vssd vccd vccd mprj_adr_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_43_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[84\]_B mprj_logic_high_inst/HI[414] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[55\] user_to_mprj_in_gates\[55\]/Y vssd vssd vccd vccd la_data_in_mprj[55]
+ sky130_fd_sc_hd__inv_8
XFILLER_43_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[117\]_TE mprj_logic_high_inst/HI[319] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[111\] la_data_out_core[111] user_to_mprj_in_gates\[111\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[111\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[75\]_B mprj_logic_high_inst/HI[405] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1019 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[1\]_A la_data_out_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[91\]_A_N la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[16\]_TE mprj_logic_high_inst/HI[218] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[95\] la_iena_mprj[95] mprj_logic_high_inst/HI[425] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/B sky130_fd_sc_hd__and2_1
XFILLER_14_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__503__A la_data_out_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[121\] _389_/Y mprj_logic_high_inst/HI[323] vssd vssd vccd
+ vccd la_oenb_core[121] sky130_fd_sc_hd__einvp_8
XFILLER_1_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_sel_buf\[2\] _405_/Y mprj_sel_buf\[2\]/TE vssd vssd vccd vccd mprj_sel_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1242 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[51\] _650_/Y mprj_logic_high_inst/HI[253] vssd vssd vccd
+ vccd la_oenb_core[51] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[73\] la_oenb_mprj[73] la_buf_enable\[73\]/B vssd vssd vccd vccd la_buf\[73\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[44\]_A_N la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_74 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_593_ la_data_out_mprj[122] vssd vssd vccd vccd _593_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[59\] _530_/Y la_buf\[59\]/TE vssd vssd vccd vccd la_data_in_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_34_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[59\]_A_N la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[115\] _586_/Y la_buf\[115\]/TE vssd vssd vccd vccd la_data_in_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_4_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__413__A mprj_adr_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[54\]_TE la_buf\[54\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[48\] la_data_out_core[48] user_to_mprj_in_gates\[48\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_15_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1700 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[10\] la_iena_mprj[10] mprj_logic_high_inst/HI[340] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[99\] _367_/Y mprj_logic_high_inst/HI[301] vssd vssd vccd
+ vccd la_oenb_core[99] sky130_fd_sc_hd__einvp_8
XFILLER_46_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_vdd_pwrgood mprj2_vdd_pwrgood/A vssd vssd vccd vccd user2_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_46_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[77\]_TE la_buf\[77\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_645_ la_oenb_mprj[46] vssd vssd vccd vccd _645_/Y sky130_fd_sc_hd__inv_2
X_576_ la_data_out_mprj[105] vssd vssd vccd vccd _576_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__408__A mprj_adr_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[18\] user_to_mprj_in_gates\[18\]/Y vssd vssd vccd vccd la_data_in_mprj[18]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[26\]_TE mprj_dat_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[58\] la_iena_mprj[58] mprj_logic_high_inst/HI[388] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_430_ mprj_adr_o_core[23] vssd vssd vccd vccd _430_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[14\] _613_/Y mprj_logic_high_inst/HI[216] vssd vssd vccd
+ vccd la_oenb_core[14] sky130_fd_sc_hd__einvp_8
X_361_ la_oenb_mprj[93] vssd vssd vccd vccd _361_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[36\] la_oenb_mprj[36] la_buf_enable\[36\]/B vssd vssd vccd vccd la_buf\[36\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_sel_buf\[0\]_TE mprj_sel_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_628_ la_oenb_mprj[29] vssd vssd vccd vccd _628_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_559_ la_data_out_mprj[88] vssd vssd vccd vccd _559_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__601__A la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_249 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_907 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_918 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_929 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__511__A la_data_out_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_205 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_413_ mprj_adr_o_core[6] vssd vssd vccd vccd _413_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[102\]_TE la_buf\[102\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_344_ la_oenb_mprj[76] vssd vssd vccd vccd _344_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[41\] _512_/Y la_buf\[41\]/TE vssd vssd vccd vccd la_data_in_core[41] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[113\] la_iena_mprj[113] mprj_logic_high_inst/HI[443] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[113\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[17\]_TE mprj_adr_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__421__A mprj_adr_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[1\]_TE mprj_adr_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[119\] user_to_mprj_in_gates\[119\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[119] sky130_fd_sc_hd__inv_8
XFILLER_2_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[85\] user_to_mprj_in_gates\[85\]/Y vssd vssd vccd vccd la_data_in_mprj[85]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[30\] la_data_out_core[30] user_to_mprj_in_gates\[30\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__331__A la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[5\]_TE mprj_dat_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_937 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__506__A la_data_out_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[81\] _349_/Y mprj_logic_high_inst/HI[283] vssd vssd vccd
+ vccd la_oenb_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_10_1868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[89\] _560_/Y la_buf\[89\]/TE vssd vssd vccd vccd la_data_in_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_0_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[104\] la_oenb_mprj[104] la_buf_enable\[104\]/B vssd vssd vccd vccd
+ la_buf\[104\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_19_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_775 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__416__A mprj_adr_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[78\] la_data_out_core[78] user_to_mprj_in_gates\[78\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_583 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[91\]_A la_data_out_core[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj2_pwrgood_A mprj2_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_366 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[40\] la_iena_mprj[40] mprj_logic_high_inst/HI[370] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[95\]_TE mprj_logic_high_inst/HI[297] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1111 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1100 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1122 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[82\]_A la_data_out_core[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[104\]_B la_buf_enable\[104\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[48\] user_to_mprj_in_gates\[48\]/Y vssd vssd vccd vccd la_data_in_mprj[48]
+ sky130_fd_sc_hd__inv_8
XFILLER_43_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[73\]_A la_data_out_core[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1576 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[104\] la_data_out_core[104] user_to_mprj_in_gates\[104\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[104\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2099 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[1\]_B user_to_mprj_in_gates\[1\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1621 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[64\]_A la_data_out_core[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[88\] la_iena_mprj[88] mprj_logic_high_inst/HI[418] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[114\] _382_/Y mprj_logic_high_inst/HI[316] vssd vssd vccd
+ vccd la_oenb_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_5_1210 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1232 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[44\] _643_/Y mprj_logic_high_inst/HI[246] vssd vssd vccd
+ vccd la_oenb_core[44] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[66\] la_oenb_mprj[66] la_buf_enable\[66\]/B vssd vssd vccd vccd la_buf\[66\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_irq_buffers\[2\] user_irq_gates\[2\]/Y vssd vssd vccd vccd user_irq[2] sky130_fd_sc_hd__inv_8
XFILLER_44_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_592_ la_data_out_mprj[121] vssd vssd vccd vccd _592_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1418 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[55\]_A la_data_out_core[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[108\] _579_/Y la_buf\[108\]/TE vssd vssd vccd vccd la_data_in_core[108] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[101\] user_to_mprj_in_gates\[101\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[101] sky130_fd_sc_hd__inv_8
XFILLER_3_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[5\]_A user_to_mprj_in_gates\[5\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[46\]_A la_data_out_core[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__604__A la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xmprj_dat_buf\[0\] _439_/Y mprj_dat_buf\[0\]/TE vssd vssd vccd vccd mprj_dat_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_2141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[37\]_A la_data_out_core[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[121\]_A la_data_out_core[121] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_21_394 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__514__A la_data_out_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1349 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1466 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_644_ la_oenb_mprj[45] vssd vssd vccd vccd _644_/Y sky130_fd_sc_hd__inv_2
XFILLER_5_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[71\] _542_/Y la_buf\[71\]/TE vssd vssd vccd vccd la_data_in_core[71] sky130_fd_sc_hd__einvp_8
XFILLER_17_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_575_ la_data_out_mprj[104] vssd vssd vccd vccd _575_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__424__A mprj_adr_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[28\]_A la_data_out_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1671 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[112\]_A la_data_out_core[112] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_47_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[21\]_TE la_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[60\] la_data_out_core[60] user_to_mprj_in_gates\[60\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_1642 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[90\]_A_N la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[19\]_A la_data_out_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[103\]_A la_data_out_core[103] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__334__A la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[43\]_A_N la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[58\]_A_N la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__509__A la_data_out_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_360_ la_oenb_mprj[92] vssd vssd vccd vccd _360_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[29\] la_oenb_mprj[29] la_buf_enable\[29\]/B vssd vssd vccd vccd la_buf\[29\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_42_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[29\]_TE mprj_logic_high_inst/HI[231] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__419__A mprj_adr_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_627_ la_oenb_mprj[28] vssd vssd vccd vccd _627_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_558_ la_data_out_mprj[87] vssd vssd vccd vccd _558_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_489_ la_data_out_mprj[18] vssd vssd vccd vccd _489_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[30\] user_to_mprj_in_gates\[30\]/Y vssd vssd vccd vccd la_data_in_mprj[30]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[1\]_B la_buf_enable\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[125\]_A la_iena_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_908 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_919 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[70\] la_iena_mprj[70] mprj_logic_high_inst/HI[400] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[116\]_A la_iena_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_412_ mprj_adr_o_core[5] vssd vssd vccd vccd _412_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_343_ la_oenb_mprj[75] vssd vssd vccd vccd _343_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[34\] _505_/Y la_buf\[34\]/TE vssd vssd vccd vccd la_data_in_core[34] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[106\] la_iena_mprj[106] mprj_logic_high_inst/HI[436] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[106\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[16\]_TE mprj_dat_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[107\]_A la_iena_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[78\] user_to_mprj_in_gates\[78\]/Y vssd vssd vccd vccd la_data_in_mprj[78]
+ sky130_fd_sc_hd__inv_8
XFILLER_20_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1739 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[23\] la_data_out_core[23] user_to_mprj_in_gates\[23\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__612__A la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__522__A la_data_out_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[74\] _342_/Y mprj_logic_high_inst/HI[276] vssd vssd vccd
+ vccd la_oenb_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_2_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[96\] la_oenb_mprj[96] la_buf_enable\[96\]/B vssd vssd vccd vccd la_buf\[96\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[22\] _461_/Y mprj_dat_buf\[22\]/TE vssd vssd vccd vccd mprj_dat_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[96\]_A la_iena_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[20\]_A la_iena_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__432__A mprj_adr_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[87\]_A la_iena_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__607__A la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[11\]_A la_iena_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[2\] la_oenb_mprj[2] la_buf_enable\[2\]/B vssd vssd vccd vccd la_buf\[2\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__342__A la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1607 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[78\]_A la_iena_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[33\] la_iena_mprj[33] mprj_logic_high_inst/HI[363] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/B sky130_fd_sc_hd__and2_1
XPHY_502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__517__A la_data_out_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1112 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1101 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1123 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_216 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[11\] la_oenb_mprj[11] la_buf_enable\[11\]/B vssd vssd vccd vccd la_buf\[11\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[69\]_A la_iena_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__427__A mprj_adr_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_562 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[90\] la_data_out_core[90] user_to_mprj_in_gates\[90\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_44_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1377 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__337__A la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1953 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[107\] _375_/Y mprj_logic_high_inst/HI[309] vssd vssd vccd
+ vccd la_oenb_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_40_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_660_ la_oenb_mprj[61] vssd vssd vccd vccd _660_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_591_ la_data_out_mprj[120] vssd vssd vccd vccd _591_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[37\] _636_/Y mprj_logic_high_inst/HI[239] vssd vssd vccd
+ vccd la_oenb_core[37] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[59\] la_oenb_mprj[59] la_buf_enable\[59\]/B vssd vssd vccd vccd la_buf\[59\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[40\]_A user_to_mprj_in_gates\[40\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[60\] user_to_mprj_in_gates\[60\]/Y vssd vssd vccd vccd la_data_in_mprj[60]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1828 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1374 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[85\]_TE mprj_logic_high_inst/HI[287] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__620__A la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[31\]_A user_to_mprj_in_gates\[31\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1130 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[98\]_A user_to_mprj_in_gates\[98\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[71\]_A _542_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__530__A la_data_out_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[22\]_A user_to_mprj_in_gates\[22\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_643_ la_oenb_mprj[44] vssd vssd vccd vccd _643_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_484 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[64\] _535_/Y la_buf\[64\]/TE vssd vssd vccd vccd la_data_in_core[64] sky130_fd_sc_hd__einvp_8
X_574_ la_data_out_mprj[103] vssd vssd vccd vccd _574_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_159 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[125\]_A _596_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_845 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[89\]_A user_to_mprj_in_gates\[89\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_1525 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[120\] _591_/Y la_buf\[120\]/TE vssd vssd vccd vccd la_data_in_core[120] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[28\] _435_/Y mprj_adr_buf\[28\]/TE vssd vssd vccd vccd mprj_adr_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[80\]_B la_buf_enable\[80\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__440__A mprj_dat_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[53\] la_data_out_core[53] user_to_mprj_in_gates\[53\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_buffers\[13\]_A user_to_mprj_in_gates\[13\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[116\]_A _587_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__615__A la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[19\]_B user_to_mprj_in_gates\[19\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__350__A la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1598 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[107\]_A _578_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__525__A la_data_out_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_826 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[44\]_A _515_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_899 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[127\] la_oenb_mprj[127] la_buf_enable\[127\]/B vssd vssd vccd vccd
+ la_buf\[127\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_24_1963 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_626_ la_oenb_mprj[27] vssd vssd vccd vccd _626_/Y sky130_fd_sc_hd__inv_2
X_557_ la_data_out_mprj[86] vssd vssd vccd vccd _557_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_44_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_488_ la_data_out_mprj[17] vssd vssd vccd vccd _488_/Y sky130_fd_sc_hd__inv_2
XANTENNA__435__A mprj_adr_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[23\] user_to_mprj_in_gates\[23\]/Y vssd vssd vccd vccd la_data_in_mprj[23]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[53\]_B la_buf_enable\[53\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[125\]_B mprj_logic_high_inst/HI[455] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_909 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_1_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__345__A la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[26\]_A _497_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[44\]_B la_buf_enable\[44\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[63\] la_iena_mprj[63] mprj_logic_high_inst/HI[393] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[116\]_B mprj_logic_high_inst/HI[446] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[1\] _600_/Y mprj_logic_high_inst/HI[203] vssd vssd vccd
+ vccd la_oenb_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_2_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[41\] la_oenb_mprj[41] la_buf_enable\[41\]/B vssd vssd vccd vccd la_buf\[41\]/TE
+ sky130_fd_sc_hd__and2b_1
X_411_ mprj_adr_o_core[4] vssd vssd vccd vccd _411_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_342_ la_oenb_mprj[74] vssd vssd vccd vccd _342_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[27\] _498_/Y la_buf\[27\]/TE vssd vssd vccd vccd la_data_in_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_46_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[35\]_B la_buf_enable\[35\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[4\]_A la_iena_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[107\]_B mprj_logic_high_inst/HI[437] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_609_ la_oenb_mprj[10] vssd vssd vccd vccd _609_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[42\]_A_N la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[16\] la_data_out_core[16] user_to_mprj_in_gates\[16\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1553 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[57\]_A_N la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[26\]_B la_buf_enable\[26\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[127\] la_data_out_core[127] user_to_mprj_in_gates\[127\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[127\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[19\]_TE mprj_logic_high_inst/HI[221] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_23_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[17\]_B la_buf_enable\[17\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[67\] _335_/Y mprj_logic_high_inst/HI[269] vssd vssd vccd
+ vccd la_oenb_core[67] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[89\] la_oenb_mprj[89] la_buf_enable\[89\]/B vssd vssd vccd vccd la_buf\[89\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[15\] _454_/Y mprj_dat_buf\[15\]/TE vssd vssd vccd vccd mprj_dat_o_user[15]
+ sky130_fd_sc_hd__einvp_8
XFILLER_47_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[2\]_TE la_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1748 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[10\] _417_/Y mprj_adr_buf\[10\]/TE vssd vssd vccd vccd mprj_adr_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[124\] user_to_mprj_in_gates\[124\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[124] sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[57\]_TE la_buf\[57\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[90\] user_to_mprj_in_gates\[90\]/Y vssd vssd vccd vccd la_data_in_mprj[90]
+ sky130_fd_sc_hd__inv_8
XFILLER_38_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__623__A la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[78\]_B mprj_logic_high_inst/HI[408] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[4\]_A la_data_out_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[26\] la_iena_mprj[26] mprj_logic_high_inst/HI[356] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/B sky130_fd_sc_hd__and2_1
XPHY_503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1113 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1102 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1124 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_279 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__533__A la_data_out_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[94\] _565_/Y la_buf\[94\]/TE vssd vssd vccd vccd la_data_in_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_19_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__443__A mprj_dat_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[83\] la_data_out_core[83] user_to_mprj_in_gates\[83\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[29\]_TE mprj_dat_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__618__A la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2068 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[8\]_TE mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1000 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__353__A la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2093 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_590_ la_data_out_mprj[119] vssd vssd vccd vccd _590_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__528__A la_data_out_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[5\] _476_/Y la_buf\[5\]/TE vssd vssd vccd vccd la_data_in_core[5] sky130_fd_sc_hd__einvp_8
XFILLER_6_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_pwrgood_A mprj_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_TE mprj_sel_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[2\] _409_/Y mprj_adr_buf\[2\]/TE vssd vssd vccd vccd mprj_adr_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__438__A mprj_adr_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[53\] user_to_mprj_in_gates\[53\]/Y vssd vssd vccd vccd la_data_in_mprj[53]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1593 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_319 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[10\]_A _449_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1943 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1217 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1587 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__348__A la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[93\] la_iena_mprj[93] mprj_logic_high_inst/HI[423] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[0\] _403_/Y mprj_sel_buf\[0\]/TE vssd vssd vccd vccd mprj_sel_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1329 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[71\] la_oenb_mprj[71] la_buf_enable\[71\]/B vssd vssd vccd vccd la_buf\[71\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_642_ la_oenb_mprj[43] vssd vssd vccd vccd _642_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_573_ la_data_out_mprj[102] vssd vssd vccd vccd _573_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[57\] _528_/Y la_buf\[57\]/TE vssd vssd vccd vccd la_data_in_core[57] sky130_fd_sc_hd__einvp_8
XFILLER_38_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[113\] _584_/Y la_buf\[113\]/TE vssd vssd vccd vccd la_data_in_core[113] sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_adr_buf\[4\]_TE mprj_adr_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[46\] la_data_out_core[46] user_to_mprj_in_gates\[46\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1462 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[52\]_TE mprj_logic_high_inst/HI[254] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__631__A la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[8\]_TE mprj_dat_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[8\] la_data_out_core[8] user_to_mprj_in_gates\[8\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[8\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_400 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_948 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1651 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[97\] _365_/Y mprj_logic_high_inst/HI[299] vssd vssd vccd
+ vccd la_oenb_core[97] sky130_fd_sc_hd__einvp_8
XANTENNA__541__A la_data_out_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[90\]_TE la_buf\[90\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_625_ la_oenb_mprj[26] vssd vssd vccd vccd _625_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[75\]_TE mprj_logic_high_inst/HI[277] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_556_ la_data_out_mprj[85] vssd vssd vccd vccd _556_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_948 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_487_ la_data_out_mprj[16] vssd vssd vccd vccd _487_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[16\] user_to_mprj_in_gates\[16\]/Y vssd vssd vccd vccd la_data_in_mprj[16]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_175 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__451__A mprj_dat_o_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__626__A la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__361__A la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[56\] la_iena_mprj[56] mprj_logic_high_inst/HI[386] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[98\]_TE mprj_logic_high_inst/HI[300] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_410_ mprj_adr_o_core[3] vssd vssd vccd vccd _410_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__536__A la_data_out_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_341_ la_oenb_mprj[73] vssd vssd vccd vccd _341_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[12\] _611_/Y mprj_logic_high_inst/HI[214] vssd vssd vccd
+ vccd la_oenb_core[12] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[34\] la_oenb_mprj[34] la_buf_enable\[34\]/B vssd vssd vccd vccd la_buf\[34\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[8\] user_to_mprj_in_gates\[8\]/Y vssd vssd vccd vccd la_data_in_mprj[8]
+ sky130_fd_sc_hd__inv_8
XFILLER_14_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_stb_buf _401_/Y mprj_stb_buf/TE vssd vssd vccd vccd mprj_stb_o_user sky130_fd_sc_hd__einvp_8
XFILLER_2_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_608_ la_oenb_mprj[9] vssd vssd vccd vccd _608_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__446__A mprj_dat_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_539_ la_data_out_mprj[68] vssd vssd vccd vccd _539_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_707 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_718 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__356__A la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_729 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[94\]_A la_data_out_core[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[85\]_A la_data_out_core[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[111\] la_iena_mprj[111] mprj_logic_high_inst/HI[441] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[111\]/B sky130_fd_sc_hd__and2_1
XPHY_1840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_adr_buf\[30\]_TE mprj_adr_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[117\] user_to_mprj_in_gates\[117\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[117] sky130_fd_sc_hd__inv_8
XFILLER_42_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[83\] user_to_mprj_in_gates\[83\]/Y vssd vssd vccd vccd la_data_in_mprj[83]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[76\]_A la_data_out_core[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1215 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_608 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[4\]_B user_to_mprj_in_gates\[4\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_504 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_515 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_526 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1114 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1103 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_537 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_548 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[19\] la_iena_mprj[19] mprj_logic_high_inst/HI[349] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/B sky130_fd_sc_hd__and2_1
XPHY_559 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1125 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[67\]_A la_data_out_core[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[41\]_A_N la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[56\]_A_N la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[87\] _558_/Y la_buf\[87\]/TE vssd vssd vccd vccd la_data_in_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_46_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[102\] la_oenb_mprj[102] la_buf_enable\[102\]/B vssd vssd vccd vccd
+ la_buf\[102\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_34_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[58\]_A la_data_out_core[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_578 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[24\]_TE la_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_991 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[76\] la_data_out_core[76] user_to_mprj_in_gates\[76\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[8\]_A user_to_mprj_in_gates\[8\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[49\]_A la_data_out_core[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__634__A la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_589 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_301 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_323 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_312 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_334 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_356 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_367 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_345 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[124\]_A la_data_out_core[124] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XPHY_389 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_378 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__544__A la_data_out_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[47\]_TE la_buf\[47\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_irq_ena_buf\[2\] user_irq_ena[2] user_irq_ena_buf\[2\]/B vssd vssd vccd vccd
+ user_irq_gates\[2\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[46\] user_to_mprj_in_gates\[46\]/Y vssd vssd vccd vccd la_data_in_mprj[46]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[115\]_A la_data_out_core[115] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__454__A mprj_dat_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_890 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1955 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__629__A la_oenb_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[102\] la_data_out_core[102] user_to_mprj_in_gates\[102\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[102\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1187 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[106\]_A la_data_out_core[106] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__364__A la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[86\] la_iena_mprj[86] mprj_logic_high_inst/HI[416] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_202 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[112\] _380_/Y mprj_logic_high_inst/HI[314] vssd vssd vccd
+ vccd la_oenb_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_48_228 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_641_ la_oenb_mprj[42] vssd vssd vccd vccd _641_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[42\] _641_/Y mprj_logic_high_inst/HI[244] vssd vssd vccd
+ vccd la_oenb_core[42] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[64\] la_oenb_mprj[64] la_buf_enable\[64\]/B vssd vssd vccd vccd la_buf\[64\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__539__A la_data_out_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_buffers\[0\] user_irq_gates\[0\]/Y vssd vssd vccd vccd user_irq[0] sky130_fd_sc_hd__inv_8
X_572_ la_data_out_mprj[101] vssd vssd vccd vccd _572_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_131 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_142 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_175 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_164 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_153 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_186 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_197 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[19\]_TE mprj_dat_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[106\] _577_/Y la_buf\[106\]/TE vssd vssd vccd vccd la_data_in_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_45_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__449__A mprj_dat_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[39\] la_data_out_core[39] user_to_mprj_in_gates\[39\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/Y sky130_fd_sc_hd__nand2_4
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[4\]_B la_buf_enable\[4\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_1523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__359__A la_oenb_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_879 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[119\]_A la_iena_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[120\]_TE mprj_logic_high_inst/HI[322] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
X_624_ la_oenb_mprj[25] vssd vssd vccd vccd _624_/Y sky130_fd_sc_hd__inv_2
X_555_ la_data_out_mprj[84] vssd vssd vccd vccd _555_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_486_ la_data_out_mprj[15] vssd vssd vccd vccd _486_/Y sky130_fd_sc_hd__inv_2
Xmprj_we_buf _402_/Y mprj_we_buf/TE vssd vssd vccd vccd mprj_we_o_user sky130_fd_sc_hd__einvp_8
XFILLER_9_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[50\]_A la_iena_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_pwrgood mprj_pwrgood/A vssd vssd vccd vccd user1_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_25_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[41\]_A la_iena_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__642__A la_oenb_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[49\] la_iena_mprj[49] mprj_logic_high_inst/HI[379] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_340_ la_oenb_mprj[72] vssd vssd vccd vccd _340_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[32\]_A la_iena_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[27\] la_oenb_mprj[27] la_buf_enable\[27\]/B vssd vssd vccd vccd la_buf\[27\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__552__A la_data_out_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1081 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[99\]_A la_iena_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[42\]_TE mprj_logic_high_inst/HI[244] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_607_ la_oenb_mprj[8] vssd vssd vccd vccd _607_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_538_ la_data_out_mprj[67] vssd vssd vccd vccd _538_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[23\]_A la_iena_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_469_ mprj_dat_o_core[30] vssd vssd vccd vccd _469_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_470 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__462__A mprj_dat_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[118\]_TE la_buf\[118\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1559 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__637__A la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_708 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_212 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[14\]_A la_iena_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_719 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__372__A la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__547__A la_data_out_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[1\]_A user_irq_ena[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_we_buf_A _402_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[85\]_B user_to_mprj_in_gates\[85\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_1852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[104\] la_iena_mprj[104] mprj_logic_high_inst/HI[434] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[104\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[32\] _503_/Y la_buf\[32\]/TE vssd vssd vccd vccd la_data_in_core[32] sky130_fd_sc_hd__einvp_8
XFILLER_10_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[70\]_A user_to_mprj_in_gates\[70\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[76\] user_to_mprj_in_gates\[76\]/Y vssd vssd vccd vccd la_data_in_mprj[76]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__457__A mprj_dat_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[21\] la_data_out_core[21] user_to_mprj_in_gates\[21\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_37_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[88\]_TE mprj_logic_high_inst/HI[290] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[9\] _448_/Y mprj_dat_buf\[9\]/TE vssd vssd vccd vccd mprj_dat_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_44_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1163 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__367__A la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_505 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_516 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1104 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_527 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_538 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_549 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1115 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[72\] _340_/Y mprj_logic_high_inst/HI[274] vssd vssd vccd
+ vccd la_oenb_core[72] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[94\] la_oenb_mprj[94] la_buf_enable\[94\]/B vssd vssd vccd vccd la_buf\[94\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[20\] _459_/Y mprj_dat_buf\[20\]/TE vssd vssd vccd vccd mprj_dat_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[52\]_A user_to_mprj_in_gates\[52\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1558 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[43\]_A user_to_mprj_in_gates\[43\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[69\] la_data_out_core[69] user_to_mprj_in_gates\[69\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_1_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[0\] la_oenb_mprj[0] la_buf_enable\[0\]/B vssd vssd vccd vccd la_buf\[0\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__650__A la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_38 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[34\]_A user_to_mprj_in_gates\[34\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[31\] la_iena_mprj[31] mprj_logic_high_inst/HI[361] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[20\]_TE mprj_adr_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_324 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_313 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_302 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_357 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_335 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_368 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_346 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[74\]_A _545_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_379 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[92\]_B la_buf_enable\[92\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__560__A la_data_out_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[25\]_A user_to_mprj_in_gates\[25\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[39\] user_to_mprj_in_gates\[39\]/Y vssd vssd vccd vccd la_data_in_mprj[39]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[65\]_A _536_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_880 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_891 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[83\]_B la_buf_enable\[83\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1691 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__470__A mprj_dat_o_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[16\]_A user_to_mprj_in_gates\[16\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1556 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[119\]_A _590_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__645__A la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[40\]_A_N la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[55\]_A_N la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__380__A la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[79\] la_iena_mprj[79] mprj_logic_high_inst/HI[409] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/B sky130_fd_sc_hd__and2_1
Xuser_to_mprj_oen_buffers\[105\] _373_/Y mprj_logic_high_inst/HI[307] vssd vssd vccd
+ vccd la_oenb_core[105] sky130_fd_sc_hd__einvp_8
X_640_ la_oenb_mprj[41] vssd vssd vccd vccd _640_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_571_ la_data_out_mprj[100] vssd vssd vccd vccd _571_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[35\] _634_/Y mprj_logic_high_inst/HI[237] vssd vssd vccd
+ vccd la_oenb_core[35] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[57\] la_oenb_mprj[57] la_buf_enable\[57\]/B vssd vssd vccd vccd la_buf\[57\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf\[14\]_TE la_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__555__A la_data_out_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_132 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_143 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_176 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_165 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_154 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_187 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_198 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[65\]_B la_buf_enable\[65\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_16_1697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_21_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__465__A mprj_dat_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[37\]_TE la_buf\[37\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1239 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_59 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__375__A la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_B la_buf_enable\[47\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[119\]_B mprj_logic_high_inst/HI[449] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_623_ la_oenb_mprj[24] vssd vssd vccd vccd _623_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_554_ la_data_out_mprj[83] vssd vssd vccd vccd _554_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[62\] _533_/Y la_buf\[62\]/TE vssd vssd vccd vccd la_data_in_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_45_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_485_ la_data_out_mprj[14] vssd vssd vccd vccd _485_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf\[5\]_TE la_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_12_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[38\]_B la_buf_enable\[38\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[26\] _433_/Y mprj_adr_buf\[26\]/TE vssd vssd vccd vccd mprj_adr_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[7\]_A la_iena_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[51\] la_data_out_core[51] user_to_mprj_in_gates\[51\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[29\]_B la_buf_enable\[29\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2044 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_622 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[125\] la_oenb_mprj[125] la_buf_enable\[125\]/B vssd vssd vccd vccd
+ la_buf\[125\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_20_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_606_ la_oenb_mprj[7] vssd vssd vccd vccd _606_/Y sky130_fd_sc_hd__inv_2
X_537_ la_data_out_mprj[66] vssd vssd vccd vccd _537_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[23\]_B mprj_logic_high_inst/HI[353] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_468_ mprj_dat_o_core[29] vssd vssd vccd vccd _468_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_399_ caravel_clk2 vssd vssd vccd vccd _399_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[21\] user_to_mprj_in_gates\[21\]/Y vssd vssd vccd vccd la_data_in_mprj[21]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[99\] la_data_out_core[99] user_to_mprj_in_gates\[99\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_709 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__653__A la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[61\] la_iena_mprj[61] mprj_logic_high_inst/HI[391] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[7\]_A la_data_out_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_ena_buf\[1\]_B user_irq_ena_buf\[1\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_736 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__563__A la_data_out_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[25\] _496_/Y la_buf\[25\]/TE vssd vssd vccd vccd la_data_in_core[25] sky130_fd_sc_hd__einvp_8
XFILLER_10_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[69\] user_to_mprj_in_gates\[69\]/Y vssd vssd vccd vccd la_data_in_mprj[69]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__473__A la_data_out_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[14\] la_data_out_core[14] user_to_mprj_in_gates\[14\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[125\] la_data_out_core[125] user_to_mprj_in_gates\[125\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[125\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__648__A la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_506 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_517 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1105 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_528 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_539 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1116 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__383__A la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[32\]_TE mprj_logic_high_inst/HI[234] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[65\] _333_/Y mprj_logic_high_inst/HI[267] vssd vssd vccd
+ vccd la_oenb_core[65] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[87\] la_oenb_mprj[87] la_buf_enable\[87\]/B vssd vssd vccd vccd la_buf\[87\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[13\] _452_/Y mprj_dat_buf\[13\]/TE vssd vssd vccd vccd mprj_dat_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__558__A la_data_out_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_547 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[7\]_TE mprj_adr_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[122\] user_to_mprj_in_gates\[122\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[122] sky130_fd_sc_hd__inv_8
XFILLER_26_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1666 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__468__A mprj_dat_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[70\]_TE la_buf\[70\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_dat_buf\[13\]_A _452_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__378__A la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_314 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_325 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_303 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[24\] la_iena_mprj[24] mprj_logic_high_inst/HI[354] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/B sky130_fd_sc_hd__and2_1
XPHY_358 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_336 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_347 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_369 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[92\] _563_/Y la_buf\[92\]/TE vssd vssd vccd vccd la_data_in_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_19_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[78\]_TE mprj_logic_high_inst/HI[280] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_vdd_pwrgood mprj_vdd_pwrgood/A vssd vssd vccd vccd user1_vdd_powergood sky130_fd_sc_hd__buf_8
XFILLER_21_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_870 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_881 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_892 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[81\] la_data_out_core[81] user_to_mprj_in_gates\[81\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_41_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1191 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[9\]_A_N la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_570_ la_data_out_mprj[99] vssd vssd vccd vccd _570_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[28\] _627_/Y mprj_logic_high_inst/HI[230] vssd vssd vccd
+ vccd la_oenb_core[28] sky130_fd_sc_hd__einvp_8
XPHY_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_133 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_166 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_155 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_144 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_177 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_199 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_188 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__571__A la_data_out_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[3\] _474_/Y la_buf\[3\]/TE vssd vssd vccd vccd la_data_in_core[3] sky130_fd_sc_hd__einvp_8
XFILLER_4_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[0\]_A user_irq_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1084 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[0\] _407_/Y mprj_adr_buf\[0\]/TE vssd vssd vccd vccd mprj_adr_o_user[0]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1708 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[51\] user_to_mprj_in_gates\[51\]/Y vssd vssd vccd vccd la_data_in_mprj[51]
+ sky130_fd_sc_hd__inv_8
XFILLER_23_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__481__A la_data_out_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[10\]_TE mprj_adr_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__656__A la_oenb_mprj[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[7\]_A _414_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__391__A la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_848 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[91\] la_iena_mprj[91] mprj_logic_high_inst/HI[421] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/B sky130_fd_sc_hd__and2_1
XFILLER_44_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_622_ la_oenb_mprj[23] vssd vssd vccd vccd _622_/Y sky130_fd_sc_hd__inv_2
XANTENNA__566__A la_data_out_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_553_ la_data_out_mprj[82] vssd vssd vccd vccd _553_/Y sky130_fd_sc_hd__inv_2
X_484_ la_data_out_mprj[13] vssd vssd vccd vccd _484_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[55\] _526_/Y la_buf\[55\]/TE vssd vssd vccd vccd la_data_in_core[55] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[127\] la_iena_mprj[127] mprj_logic_high_inst/HI[457] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[127\]/B sky130_fd_sc_hd__and2_1
XFILLER_18_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[19\] _426_/Y mprj_adr_buf\[19\]/TE vssd vssd vccd vccd mprj_adr_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[111\] _582_/Y la_buf\[111\]/TE vssd vssd vccd vccd la_data_in_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_10_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[99\] user_to_mprj_in_gates\[99\]/Y vssd vssd vccd vccd la_data_in_mprj[99]
+ sky130_fd_sc_hd__inv_8
XANTENNA__476__A la_data_out_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[54\]_A_N la_oenb_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[44\] la_data_out_core[44] user_to_mprj_in_gates\[44\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_35_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[69\]_A_N la_oenb_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[6\] la_data_out_core[6] user_to_mprj_in_gates\[6\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[6\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[30\]_A la_data_out_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1438 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1184 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_918 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__386__A la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[97\]_A la_data_out_core[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[95\] _363_/Y mprj_logic_high_inst/HI[297] vssd vssd vccd
+ vccd la_oenb_core[95] sky130_fd_sc_hd__einvp_8
XFILLER_46_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[21\]_A la_data_out_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[8\] la_iena_mprj[8] mprj_logic_high_inst/HI[338] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[8\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[118\] la_oenb_mprj[118] la_buf_enable\[118\]/B vssd vssd vccd vccd
+ la_buf\[118\]/TE sky130_fd_sc_hd__and2b_1
X_605_ la_oenb_mprj[6] vssd vssd vccd vccd _605_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_536_ la_data_out_mprj[65] vssd vssd vccd vccd _536_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[88\]_A la_data_out_core[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_467_ mprj_dat_o_core[28] vssd vssd vccd vccd _467_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_398_ caravel_clk vssd vssd vccd vccd _398_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[14\] user_to_mprj_in_gates\[14\]/Y vssd vssd vccd vccd la_data_in_mprj[14]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_A la_data_out_core[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1686 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_A la_data_out_core[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1267 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1245 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[54\] la_iena_mprj[54] mprj_logic_high_inst/HI[384] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_gates\[7\]_B user_to_mprj_in_gates\[7\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_oen_buffers\[10\] _609_/Y mprj_logic_high_inst/HI[212] vssd vssd vccd
+ vccd la_oenb_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_42_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[6\] user_to_mprj_in_gates\[6\]/Y vssd vssd vccd vccd la_data_in_mprj[6]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[32\] la_oenb_mprj[32] la_buf_enable\[32\]/B vssd vssd vccd vccd la_buf\[32\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_442 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[18\] _489_/Y la_buf\[18\]/TE vssd vssd vccd vccd la_data_in_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_10_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_519_ la_data_out_mprj[48] vssd vssd vccd vccd _519_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2004 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_2015 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[118\] la_data_out_core[118] user_to_mprj_in_gates\[118\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[118\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_507 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_518 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_529 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1106 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1117 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1042 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1020 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_939 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[58\] _657_/Y mprj_logic_high_inst/HI[260] vssd vssd vccd
+ vccd la_oenb_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_25_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_501 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[127\]_A la_data_out_core[127] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__574__A la_data_out_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[100\]_A la_iena_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[115\] user_to_mprj_in_gates\[115\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[115] sky130_fd_sc_hd__inv_8
XFILLER_26_1623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_buffers\[81\] user_to_mprj_in_gates\[81\]/Y vssd vssd vccd vccd la_data_in_mprj[81]
+ sky130_fd_sc_hd__inv_8
XFILLER_38_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[100\]_TE mprj_logic_high_inst/HI[302] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[118\]_A la_data_out_core[118] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__484__A la_data_out_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_2096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__659__A la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[109\]_A la_data_out_core[109] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XPHY_315 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_304 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__394__A la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_359 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_326 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_337 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[17\] la_iena_mprj[17] mprj_logic_high_inst/HI[347] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/B sky130_fd_sc_hd__and2_1
XPHY_348 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__569__A la_data_out_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[85\] _556_/Y la_buf\[85\]/TE vssd vssd vccd vccd la_data_in_core[85] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_oen_buffers\[123\]_TE mprj_logic_high_inst/HI[325] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_125 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[100\] la_oenb_mprj[100] la_buf_enable\[100\]/B vssd vssd vccd vccd
+ la_buf\[100\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_21_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[80\]_A la_iena_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_860 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_871 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_893 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_882 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_791 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[74\] la_data_out_core[74] user_to_mprj_in_gates\[74\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__479__A la_data_out_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[22\]_TE mprj_logic_high_inst/HI[224] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[71\]_A la_iena_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[7\]_B la_buf_enable\[7\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__389__A la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[62\]_A la_iena_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_134 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_813 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_167 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_156 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_145 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_178 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_189 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[60\]_TE la_buf\[60\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_ena_buf\[0\] user_irq_ena[0] user_irq_ena_buf\[0\]/B vssd vssd vccd vccd
+ user_irq_gates\[0\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_oen_buffers\[45\]_TE mprj_logic_high_inst/HI[247] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[53\]_A la_iena_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[44\] user_to_mprj_in_gates\[44\]/Y vssd vssd vccd vccd la_data_in_mprj[44]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_690 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_721 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_sel_buf\[1\]_A _404_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[100\] la_data_out_core[100] user_to_mprj_in_gates\[100\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[100\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[44\]_A la_iena_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[84\] la_iena_mprj[84] mprj_logic_high_inst/HI[414] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[110\] _378_/Y mprj_logic_high_inst/HI[312] vssd vssd vccd
+ vccd la_oenb_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_29_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[40\] _639_/Y mprj_logic_high_inst/HI[242] vssd vssd vccd
+ vccd la_oenb_core[40] sky130_fd_sc_hd__einvp_8
X_621_ la_oenb_mprj[22] vssd vssd vccd vccd _621_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[62\] la_oenb_mprj[62] la_buf_enable\[62\]/B vssd vssd vccd vccd la_buf\[62\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_552_ la_data_out_mprj[81] vssd vssd vccd vccd _552_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[35\]_A la_iena_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1764 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_483_ la_data_out_mprj[12] vssd vssd vccd vccd _483_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_974 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__582__A la_data_out_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[48\] _519_/Y la_buf\[48\]/TE vssd vssd vccd vccd la_data_in_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_31_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[104\] _575_/Y la_buf\[104\]/TE vssd vssd vccd vccd la_data_in_core[104] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[26\]_A la_iena_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[37\] la_data_out_core[37] user_to_mprj_in_gates\[37\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_16_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__492__A la_data_out_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1541 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_A_N la_oenb_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[17\]_A la_iena_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2072 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[88\] _356_/Y mprj_logic_high_inst/HI[290] vssd vssd vccd
+ vccd la_oenb_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_46_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[21\]_B user_to_mprj_in_gates\[21\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__577__A la_data_out_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_604_ la_oenb_mprj[5] vssd vssd vccd vccd _604_/Y sky130_fd_sc_hd__inv_2
X_535_ la_data_out_mprj[64] vssd vssd vccd vccd _535_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_466_ mprj_dat_o_core[27] vssd vssd vccd vccd _466_/Y sky130_fd_sc_hd__inv_2
X_397_ user_resetn vssd vssd vccd vccd user_reset sky130_fd_sc_hd__inv_2
XFILLER_43_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1102 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[31\] _438_/Y mprj_adr_buf\[31\]/TE vssd vssd vccd vccd mprj_adr_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_42 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[12\]_B user_to_mprj_in_gates\[12\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__487__A la_data_out_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[79\]_B user_to_mprj_in_gates\[79\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[100\]_A _571_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[47\] la_iena_mprj[47] mprj_logic_high_inst/HI[377] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_adr_buf\[23\]_TE mprj_adr_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[25\] la_oenb_mprj[25] la_buf_enable\[25\]/B vssd vssd vccd vccd la_buf\[25\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[102\]_A user_to_mprj_in_gates\[102\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[53\]_A_N la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_631 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[55\]_A user_to_mprj_in_gates\[55\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[68\]_A_N la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[95\]_A _566_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_518_ la_data_out_mprj[47] vssd vssd vccd vccd _518_/Y sky130_fd_sc_hd__inv_2
X_449_ mprj_dat_o_core[10] vssd vssd vccd vccd _449_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_351 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_508 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_519 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1107 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1118 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1076 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[37\]_A user_to_mprj_in_gates\[37\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[17\]_TE la_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_1757 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[100\]_B mprj_logic_high_inst/HI[430] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_1630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[95\]_B la_buf_enable\[95\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[102\] la_iena_mprj[102] mprj_logic_high_inst/HI[432] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[102\]/B sky130_fd_sc_hd__and2_1
XANTENNA__590__A la_data_out_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_251 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[30\] _501_/Y la_buf\[30\]/TE vssd vssd vccd vccd la_data_in_core[30] sky130_fd_sc_hd__einvp_8
XPHY_1696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[28\]_A user_to_mprj_in_gates\[28\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[108\] user_to_mprj_in_gates\[108\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[108] sky130_fd_sc_hd__inv_8
XFILLER_26_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[74\] user_to_mprj_in_gates\[74\]/Y vssd vssd vccd vccd la_data_in_mprj[74]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1453 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_B la_buf_enable\[86\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[7\] _446_/Y mprj_dat_buf\[7\]/TE vssd vssd vccd vccd mprj_dat_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[10\]_B la_buf_enable\[10\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_682 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_316 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_305 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_349 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_327 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_338 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_B la_buf_enable\[77\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[92\] la_oenb_mprj[92] la_buf_enable\[92\]/B vssd vssd vccd vccd la_buf\[92\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[70\] _338_/Y mprj_logic_high_inst/HI[272] vssd vssd vccd
+ vccd la_oenb_core[70] sky130_fd_sc_hd__einvp_8
XFILLER_47_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_115 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[78\] _549_/Y la_buf\[78\]/TE vssd vssd vccd vccd la_data_in_core[78] sky130_fd_sc_hd__einvp_8
XFILLER_21_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__585__A la_data_out_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[8\]_TE la_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[80\]_B mprj_logic_high_inst/HI[410] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_15_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_850 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_861 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_872 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_894 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_883 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_2100 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[67\] la_data_out_core[67] user_to_mprj_in_gates\[67\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__495__A la_data_out_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[71\]_B mprj_logic_high_inst/HI[401] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_33_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[59\]_B la_buf_enable\[59\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1025 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[62\]_B mprj_logic_high_inst/HI[392] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_40_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_157 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_135 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_146 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_179 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_168 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1774 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[53\]_B mprj_logic_high_inst/HI[383] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[37\] user_to_mprj_in_gates\[37\]/Y vssd vssd vccd vccd la_data_in_mprj[37]
+ sky130_fd_sc_hd__inv_8
XPHY_680 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_691 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_121 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[113\]_TE mprj_logic_high_inst/HI[315] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[77\] la_iena_mprj[77] mprj_logic_high_inst/HI[407] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_clk_buf_TE mprj_clk_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[103\] _371_/Y mprj_logic_high_inst/HI[305] vssd vssd vccd
+ vccd la_oenb_core[103] sky130_fd_sc_hd__einvp_8
X_620_ la_oenb_mprj[21] vssd vssd vccd vccd _620_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_551_ la_data_out_mprj[80] vssd vssd vccd vccd _551_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[30\]_A _437_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[33\] _632_/Y mprj_logic_high_inst/HI[235] vssd vssd vccd
+ vccd la_oenb_core[33] sky130_fd_sc_hd__einvp_8
XFILLER_6_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[55\] la_oenb_mprj[55] la_buf_enable\[55\]/B vssd vssd vccd vccd la_buf\[55\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_482_ la_data_out_mprj[11] vssd vssd vccd vccd _482_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[12\]_TE mprj_logic_high_inst/HI[214] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_592 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_A _428_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj2_vdd_pwrgood_A mprj2_vdd_pwrgood/A vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_290 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[35\]_TE mprj_logic_high_inst/HI[237] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[109\]_A_N la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[29\] _468_/Y mprj_dat_buf\[29\]/TE vssd vssd vccd vccd mprj_dat_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1777 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_603_ la_oenb_mprj[4] vssd vssd vccd vccd _603_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_534_ la_data_out_mprj[63] vssd vssd vccd vccd _534_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[60\] _531_/Y la_buf\[60\]/TE vssd vssd vccd vccd la_data_in_core[60] sky130_fd_sc_hd__einvp_8
XANTENNA__593__A la_data_out_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_465_ mprj_dat_o_core[26] vssd vssd vccd vccd _465_/Y sky130_fd_sc_hd__inv_2
X_396_ caravel_rstn vssd vssd vccd vccd _396_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[24\] _431_/Y mprj_adr_buf\[24\]/TE vssd vssd vccd vccd mprj_adr_o_user[24]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[9\] la_oenb_mprj[9] la_buf_enable\[9\]/B vssd vssd vccd vccd la_buf\[9\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_30_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[22\]_TE mprj_dat_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[18\] la_oenb_mprj[18] la_buf_enable\[18\]/B vssd vssd vccd vccd la_buf\[18\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_7_949 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_irq_gates\[1\] user_irq_core[1] user_irq_gates\[1\]/B vssd vssd vccd vccd user_irq_gates\[1\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_643 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_665 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__588__A la_data_out_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[123\] la_oenb_mprj[123] la_buf_enable\[123\]/B vssd vssd vccd vccd
+ la_buf\[123\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_24_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_500 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_24_1574 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[7\]_A_N la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_517_ la_data_out_mprj[46] vssd vssd vccd vccd _517_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_448_ mprj_dat_o_core[9] vssd vssd vccd vccd _448_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_379_ la_oenb_mprj[111] vssd vssd vccd vccd _379_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[97\] la_data_out_core[97] user_to_mprj_in_gates\[97\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__498__A la_data_out_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_509 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1108 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1119 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1769 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_333 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[23\] _494_/Y la_buf\[23\]/TE vssd vssd vccd vccd la_data_in_core[23] sky130_fd_sc_hd__einvp_8
XFILLER_32_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_484 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[67\] user_to_mprj_in_gates\[67\]/Y vssd vssd vccd vccd la_data_in_mprj[67]
+ sky130_fd_sc_hd__inv_8
XFILLER_33_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[12\] la_data_out_core[12] user_to_mprj_in_gates\[12\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_mprj_adr_buf\[13\]_TE mprj_adr_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[123\] la_data_out_core[123] user_to_mprj_in_gates\[123\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[123\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[52\]_A_N la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_306 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_317 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_328 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_339 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[67\]_A_N la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1945 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[63\] _331_/Y mprj_logic_high_inst/HI[265] vssd vssd vccd
+ vccd la_oenb_core[63] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[85\] la_oenb_mprj[85] la_buf_enable\[85\]/B vssd vssd vccd vccd la_buf\[85\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[11\] _450_/Y mprj_dat_buf\[11\]/TE vssd vssd vccd vccd mprj_dat_o_user[11]
+ sky130_fd_sc_hd__einvp_8
XFILLER_27_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[1\]_TE mprj_dat_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_840 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_851 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_862 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_895 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_884 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_873 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_32_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[127\] _598_/Y la_buf\[127\]/TE vssd vssd vccd vccd la_data_in_core[127] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[120\] user_to_mprj_in_gates\[120\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[120] sky130_fd_sc_hd__inv_8
XFILLER_2_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_653 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[60\]_A la_data_out_core[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[22\] la_iena_mprj[22] mprj_logic_high_inst/HI[352] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/B sky130_fd_sc_hd__and2_1
XFILLER_13_815 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_114 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_158 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_136 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_147 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_169 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[51\]_A la_data_out_core[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[90\] _561_/Y la_buf\[90\]/TE vssd vssd vccd vccd la_data_in_core[90] sky130_fd_sc_hd__einvp_8
XANTENNA__596__A la_data_out_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[91\]_TE mprj_logic_high_inst/HI[293] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1713 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_670 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_692 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_681 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[42\]_A la_data_out_core[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[33\]_A la_data_out_core[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_550_ la_data_out_mprj[79] vssd vssd vccd vccd _550_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_481_ la_data_out_mprj[10] vssd vssd vccd vccd _481_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[48\] la_oenb_mprj[48] la_buf_enable\[48\]/B vssd vssd vccd vccd la_buf\[48\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[26\] _625_/Y mprj_logic_high_inst/HI[228] vssd vssd vccd
+ vccd la_oenb_core[26] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[8\] _607_/Y mprj_logic_high_inst/HI[210] vssd vssd vccd
+ vccd la_oenb_core[8] sky130_fd_sc_hd__einvp_8
XFILLER_40_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_656 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[1\] _472_/Y la_buf\[1\]/TE vssd vssd vccd vccd la_data_in_core[1] sky130_fd_sc_hd__einvp_8
XFILLER_32_84 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[24\]_A la_data_out_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_442 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1565 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[15\]_A la_data_out_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1176 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_602_ la_oenb_mprj[3] vssd vssd vccd vccd _602_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_533_ la_data_out_mprj[62] vssd vssd vccd vccd _533_/Y sky130_fd_sc_hd__inv_2
X_464_ mprj_dat_o_core[25] vssd vssd vccd vccd _464_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[53\] _524_/Y la_buf\[53\]/TE vssd vssd vccd vccd la_data_in_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_14_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[125\] la_iena_mprj[125] mprj_logic_high_inst/HI[455] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[125\]/B sky130_fd_sc_hd__and2_1
XFILLER_9_424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_395_ la_oenb_mprj[127] vssd vssd vccd vccd _395_/Y sky130_fd_sc_hd__inv_2
XFILLER_43_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[17\] _424_/Y mprj_adr_buf\[17\]/TE vssd vssd vccd vccd mprj_adr_o_user[17]
+ sky130_fd_sc_hd__einvp_8
XFILLER_5_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2070 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[97\] user_to_mprj_in_gates\[97\]/Y vssd vssd vccd vccd la_data_in_mprj[97]
+ sky130_fd_sc_hd__inv_8
XFILLER_46_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[103\]_TE mprj_logic_high_inst/HI[305] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[42\] la_data_out_core[42] user_to_mprj_in_gates\[42\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[121\]_A la_iena_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[4\] la_data_out_core[4] user_to_mprj_in_gates\[4\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[4\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_43_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[112\]_A la_iena_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[93\] _361_/Y mprj_logic_high_inst/HI[295] vssd vssd vccd
+ vccd la_oenb_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_2_600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_655 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[126\]_TE mprj_logic_high_inst/HI[328] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[6\] la_iena_mprj[6] mprj_logic_high_inst/HI[336] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[6\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[116\] la_oenb_mprj[116] la_buf_enable\[116\]/B vssd vssd vccd vccd
+ la_buf\[116\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_2_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[103\]_A la_iena_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_516_ la_data_out_mprj[45] vssd vssd vccd vccd _516_/Y sky130_fd_sc_hd__inv_2
X_447_ mprj_dat_o_core[8] vssd vssd vccd vccd _447_/Y sky130_fd_sc_hd__inv_2
X_378_ la_oenb_mprj[110] vssd vssd vccd vccd _378_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[12\] user_to_mprj_in_gates\[12\]/Y vssd vssd vccd vccd la_data_in_mprj[12]
+ sky130_fd_sc_hd__inv_8
XFILLER_29_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[40\]_TE la_buf\[40\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_1157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[108\]_A_N la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1109 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1034 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[52\] la_iena_mprj[52] mprj_logic_high_inst/HI[382] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[92\]_A la_iena_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[4\] user_to_mprj_in_gates\[4\]/Y vssd vssd vccd vccd la_data_in_mprj[4]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[30\] la_oenb_mprj[30] la_buf_enable\[30\]/B vssd vssd vccd vccd la_buf\[30\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_24_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[16\] _487_/Y la_buf\[16\]/TE vssd vssd vccd vccd la_data_in_core[16] sky130_fd_sc_hd__einvp_8
XFILLER_13_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__599__A la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[9\] _416_/Y mprj_adr_buf\[9\]/TE vssd vssd vccd vccd mprj_adr_o_user[9]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[83\]_A la_iena_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2012 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[12\]_TE mprj_dat_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[116\] la_data_out_core[116] user_to_mprj_in_gates\[116\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[116\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_37_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[74\]_A la_iena_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_307 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_318 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_329 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[86\]_TE la_buf\[86\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[6\]_A_N la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_912 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[126\] _394_/Y mprj_logic_high_inst/HI[328] vssd vssd vccd
+ vccd la_oenb_core[126] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[56\] _655_/Y mprj_logic_high_inst/HI[258] vssd vssd vccd
+ vccd la_oenb_core[56] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[78\] la_oenb_mprj[78] la_buf_enable\[78\]/B vssd vssd vccd vccd la_buf\[78\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[65\]_A la_iena_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_830 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_841 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_852 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_863 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_896 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_885 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_874 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_772 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_750 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[113\] user_to_mprj_in_gates\[113\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[113] sky130_fd_sc_hd__inv_8
XFILLER_2_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[56\]_A la_iena_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_871 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[47\]_A la_iena_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_805 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_142 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_126 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_137 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_148 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[15\] la_iena_mprj[15] mprj_logic_high_inst/HI[345] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_159 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[83\] _554_/Y la_buf\[83\]/TE vssd vssd vccd vccd la_data_in_core[83] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[38\]_A la_iena_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_660 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_671 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_693 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_682 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[51\]_A_N la_oenb_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[72\] la_data_out_core[72] user_to_mprj_in_gates\[72\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[72\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[66\]_A_N la_oenb_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[29\]_A la_iena_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_819 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[19\]_A_N la_oenb_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[94\]_A user_to_mprj_in_gates\[94\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[111\]_TE la_buf\[111\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[26\]_TE mprj_adr_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_480_ la_data_out_mprj[9] vssd vssd vccd vccd _480_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[19\] _618_/Y mprj_logic_high_inst/HI[221] vssd vssd vccd
+ vccd la_oenb_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_0_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_624 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[121\]_A _592_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__400__A mprj_cyc_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[42\] user_to_mprj_in_gates\[42\]/Y vssd vssd vccd vccd la_data_in_mprj[42]
+ sky130_fd_sc_hd__inv_8
XFILLER_32_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_454 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_490 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1419 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[112\]_A _583_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[76\]_A user_to_mprj_in_gates\[76\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[15\]_B user_to_mprj_in_gates\[15\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[103\]_A _574_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[82\] la_iena_mprj[82] mprj_logic_high_inst/HI[412] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/B sky130_fd_sc_hd__and2_1
XFILLER_2_859 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[81\]_TE mprj_logic_high_inst/HI[283] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[60\] la_oenb_mprj[60] la_buf_enable\[60\]/B vssd vssd vccd vccd la_buf\[60\]/TE
+ sky130_fd_sc_hd__and2b_1
X_601_ la_oenb_mprj[2] vssd vssd vccd vccd _601_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_204 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_532_ la_data_out_mprj[61] vssd vssd vccd vccd _532_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_463_ mprj_dat_o_core[24] vssd vssd vccd vccd _463_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_394_ la_oenb_mprj[126] vssd vssd vccd vccd _394_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_988 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[46\] _517_/Y la_buf\[46\]/TE vssd vssd vccd vccd la_data_in_core[46] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[118\] la_iena_mprj[118] mprj_logic_high_inst/HI[448] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[118\]/B sky130_fd_sc_hd__and2_1
XFILLER_9_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[105\]_A user_to_mprj_in_gates\[105\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[58\]_A user_to_mprj_in_gates\[58\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[102\] _573_/Y la_buf\[102\]/TE vssd vssd vccd vccd la_data_in_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_7_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[35\] la_data_out_core[35] user_to_mprj_in_gates\[35\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[35\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[121\]_B mprj_logic_high_inst/HI[451] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[49\]_A user_to_mprj_in_gates\[49\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1217 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[89\]_A _560_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[112\]_B mprj_logic_high_inst/HI[442] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_1825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_936 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[86\] _354_/Y mprj_logic_high_inst/HI[288] vssd vssd vccd
+ vccd la_oenb_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[31\]_B la_buf_enable\[31\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_188 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[0\]_A la_iena_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[109\] la_oenb_mprj[109] la_buf_enable\[109\]/B vssd vssd vccd vccd
+ la_buf\[109\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_45_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_579 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_515_ la_data_out_mprj[44] vssd vssd vccd vccd _515_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_446_ mprj_dat_o_core[7] vssd vssd vccd vccd _446_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_377_ la_oenb_mprj[109] vssd vssd vccd vccd _377_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_B la_buf_enable\[22\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[89\]_B la_buf_enable\[89\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[13\]_B la_buf_enable\[13\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[45\] la_iena_mprj[45] mprj_logic_high_inst/HI[375] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_42 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[23\] la_oenb_mprj[23] la_buf_enable\[23\]/B vssd vssd vccd vccd la_buf\[23\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_19_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2052 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_429_ mprj_adr_o_core[22] vssd vssd vccd vccd _429_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[109\] la_data_out_core[109] user_to_mprj_in_gates\[109\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[109\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[74\]_B mprj_logic_high_inst/HI[404] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1211 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_319 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[0\]_A la_data_out_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_308 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[116\]_TE mprj_logic_high_inst/HI[318] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[119\] _387_/Y mprj_logic_high_inst/HI[321] vssd vssd vccd
+ vccd la_oenb_core[119] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[49\] _648_/Y mprj_logic_high_inst/HI[251] vssd vssd vccd
+ vccd la_oenb_core[49] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf\[30\]_TE la_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_820 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_831 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_842 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_853 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_897 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_886 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[15\]_TE mprj_logic_high_inst/HI[217] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_864 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_875 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[100\] la_iena_mprj[100] mprj_logic_high_inst/HI[430] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[100\]/B sky130_fd_sc_hd__and2_1
XFILLER_7_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1030 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__403__A mprj_sel_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[107\]_A_N la_oenb_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[106\] user_to_mprj_in_gates\[106\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[106] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[72\] user_to_mprj_in_gates\[72\]/Y vssd vssd vccd vccd la_data_in_mprj[72]
+ sky130_fd_sc_hd__inv_8
XFILLER_47_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[5\] _444_/Y mprj_dat_buf\[5\]/TE vssd vssd vccd vccd mprj_dat_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_44_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[53\]_TE la_buf\[53\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[38\]_TE mprj_logic_high_inst/HI[240] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_127 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_138 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_149 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[90\] la_oenb_mprj[90] la_buf_enable\[90\]/B vssd vssd vccd vccd la_buf\[90\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[76\] _547_/Y la_buf\[76\]/TE vssd vssd vccd vccd la_data_in_core[76] sky130_fd_sc_hd__einvp_8
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_146 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_661 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_650 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_694 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_672 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_683 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[76\]_TE la_buf\[76\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[65\] la_data_out_core[65] user_to_mprj_in_gates\[65\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[65\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_A_N la_oenb_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_791 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_dat_buf\[25\]_TE mprj_dat_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_117 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[4\]_TE mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_32_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_496 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_480 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[35\] user_to_mprj_in_gates\[35\]/Y vssd vssd vccd vccd la_data_in_mprj[35]
+ sky130_fd_sc_hd__inv_8
XPHY_491 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1090 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_544 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1910 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1342 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__501__A la_data_out_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[75\] la_iena_mprj[75] mprj_logic_high_inst/HI[405] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[101\] _369_/Y mprj_logic_high_inst/HI[303] vssd vssd vccd
+ vccd la_oenb_core[101] sky130_fd_sc_hd__einvp_8
X_600_ la_oenb_mprj[1] vssd vssd vccd vccd _600_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[31\] _630_/Y mprj_logic_high_inst/HI[233] vssd vssd vccd
+ vccd la_oenb_core[31] sky130_fd_sc_hd__einvp_8
X_531_ la_data_out_mprj[60] vssd vssd vccd vccd _531_/Y sky130_fd_sc_hd__inv_2
XFILLER_27_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[53\] la_oenb_mprj[53] la_buf_enable\[53\]/B vssd vssd vccd vccd la_buf\[53\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_462_ mprj_dat_o_core[23] vssd vssd vccd vccd _462_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[50\]_A_N la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_393_ la_oenb_mprj[125] vssd vssd vccd vccd _393_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[39\] _510_/Y la_buf\[39\]/TE vssd vssd vccd vccd la_data_in_core[39] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[65\]_A_N la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__411__A mprj_adr_o_core[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[18\]_A_N la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[28\] la_data_out_core[28] user_to_mprj_in_gates\[28\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[28\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1353 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[16\]_TE mprj_adr_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[0\]_A _407_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[0\]_TE mprj_adr_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2069 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[79\] _347_/Y mprj_logic_high_inst/HI[281] vssd vssd vccd
+ vccd la_oenb_core[79] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[27\] _466_/Y mprj_dat_buf\[27\]/TE vssd vssd vccd vccd mprj_dat_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_26_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[4\]_TE mprj_dat_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_514_ la_data_out_mprj[43] vssd vssd vccd vccd _514_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_445_ mprj_dat_o_core[6] vssd vssd vccd vccd _445_/Y sky130_fd_sc_hd__inv_2
X_376_ la_oenb_mprj[108] vssd vssd vccd vccd _376_/Y sky130_fd_sc_hd__inv_2
XANTENNA__406__A mprj_sel_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[22\] _429_/Y mprj_adr_buf\[22\]/TE vssd vssd vccd vccd mprj_adr_o_user[22]
+ sky130_fd_sc_hd__einvp_8
XFILLER_9_1538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[71\]_TE mprj_logic_high_inst/HI[273] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1014 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[7\] la_oenb_mprj[7] la_buf_enable\[7\]/B vssd vssd vccd vccd la_buf\[7\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[90\]_A la_data_out_core[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[38\] la_iena_mprj[38] mprj_logic_high_inst/HI[368] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/B sky130_fd_sc_hd__and2_1
XFILLER_15_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1802 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[16\] la_oenb_mprj[16] la_buf_enable\[16\]/B vssd vssd vccd vccd la_buf\[16\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[81\]_A la_data_out_core[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[121\] la_oenb_mprj[121] la_buf_enable\[121\]/B vssd vssd vccd vccd
+ la_buf\[121\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_43_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1468 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[94\]_TE mprj_logic_high_inst/HI[296] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[103\]_B la_buf_enable\[103\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_428_ mprj_adr_o_core[21] vssd vssd vccd vccd _428_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_359_ la_oenb_mprj[91] vssd vssd vccd vccd _359_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1356 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[72\]_A la_data_out_core[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[95\] la_data_out_core[95] user_to_mprj_in_gates\[95\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[95\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_2003 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_2036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_2069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[0\]_B user_to_mprj_in_gates\[0\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_309 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[63\]_A la_data_out_core[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1238 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_810 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_821 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_832 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_843 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_854 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_887 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_865 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_876 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_898 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[21\] _492_/Y la_buf\[21\]/TE vssd vssd vccd vccd la_data_in_core[21] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[54\]_A la_data_out_core[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_546 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1097 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[65\] user_to_mprj_in_gates\[65\]/Y vssd vssd vccd vccd la_data_in_mprj[65]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[10\] la_data_out_core[10] user_to_mprj_in_gates\[10\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[10\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[45\]_A la_data_out_core[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[121\] la_data_out_core[121] user_to_mprj_in_gates\[121\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[121\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_128 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_139 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[120\]_A la_data_out_core[120] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__504__A la_data_out_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[36\]_A la_data_out_core[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1248 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[61\] _660_/Y mprj_logic_high_inst/HI[263] vssd vssd vccd
+ vccd la_oenb_core[61] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[83\] la_oenb_mprj[83] la_buf_enable\[83\]/B vssd vssd vccd vccd la_buf\[83\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_48_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[69\] _540_/Y la_buf\[69\]/TE vssd vssd vccd vccd la_data_in_core[69] sky130_fd_sc_hd__einvp_8
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_640 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_662 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_651 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_695 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_673 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_684 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[111\]_A la_data_out_core[111] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_7_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[27\]_A la_data_out_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__414__A mprj_adr_o_core[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[125\] _596_/Y la_buf\[125\]/TE vssd vssd vccd vccd la_data_in_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_3_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[106\]_TE mprj_logic_high_inst/HI[308] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[58\] la_data_out_core[58] user_to_mprj_in_gates\[58\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[58\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_1627 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[102\]_A la_data_out_core[102] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_A la_data_out_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[20\]_TE la_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1907 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[20\] la_iena_mprj[20] mprj_logic_high_inst/HI[350] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[106\]_A_N la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_1067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__409__A mprj_adr_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_470 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_481 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[28\] user_to_mprj_in_gates\[28\]/Y vssd vssd vccd vccd la_data_in_mprj[28]
+ sky130_fd_sc_hd__inv_8
XPHY_492 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1091 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1080 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1281 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2007 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[43\]_TE la_buf\[43\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[0\]_B la_buf_enable\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[28\]_TE mprj_logic_high_inst/HI[230] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_A la_iena_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1873 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1704 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[68\] la_iena_mprj[68] mprj_logic_high_inst/HI[398] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[115\]_A la_iena_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_530_ la_data_out_mprj[59] vssd vssd vccd vccd _530_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1577 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[6\] _605_/Y mprj_logic_high_inst/HI[208] vssd vssd vccd
+ vccd la_oenb_core[6] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[24\] _623_/Y mprj_logic_high_inst/HI[226] vssd vssd vccd
+ vccd la_oenb_core[24] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[46\] la_oenb_mprj[46] la_buf_enable\[46\]/B vssd vssd vccd vccd la_buf\[46\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_14_913 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_461_ mprj_dat_o_core[22] vssd vssd vccd vccd _461_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_392_ la_oenb_mprj[124] vssd vssd vccd vccd _392_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_946 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[66\]_TE la_buf\[66\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[4\]_A_N la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[106\]_A la_iena_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_659_ la_oenb_mprj[60] vssd vssd vccd vccd _659_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[15\]_TE mprj_dat_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__602__A la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__512__A la_data_out_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[95\]_A la_iena_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_64 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_513_ la_data_out_mprj[42] vssd vssd vccd vccd _513_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_444_ mprj_dat_o_core[5] vssd vssd vccd vccd _444_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[51\] _522_/Y la_buf\[51\]/TE vssd vssd vccd vccd la_data_in_core[51] sky130_fd_sc_hd__einvp_8
XFILLER_14_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[123\] la_iena_mprj[123] mprj_logic_high_inst/HI[453] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[123\]/B sky130_fd_sc_hd__and2_1
X_375_ la_oenb_mprj[107] vssd vssd vccd vccd _375_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__422__A mprj_adr_o_core[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xmprj_adr_buf\[15\] _422_/Y mprj_adr_buf\[15\]/TE vssd vssd vccd vccd mprj_adr_o_user[15]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[95\] user_to_mprj_in_gates\[95\]/Y vssd vssd vccd vccd la_data_in_mprj[95]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[86\]_A la_iena_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1263 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[40\] la_data_out_core[40] user_to_mprj_in_gates\[40\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[40\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[10\]_A la_iena_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1471 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__332__A la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[2\] la_data_out_core[2] user_to_mprj_in_gates\[2\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[2\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_8_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1843 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[77\]_A la_iena_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[64\]_A_N la_oenb_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[79\]_A_N la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__507__A la_data_out_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1235 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1268 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[91\] _359_/Y mprj_logic_high_inst/HI[293] vssd vssd vccd
+ vccd la_oenb_core[91] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[17\]_A_N la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2021 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[99\] _570_/Y la_buf\[99\]/TE vssd vssd vccd vccd la_data_in_core[99] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[4\] la_iena_mprj[4] mprj_logic_high_inst/HI[334] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[4\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[68\]_A la_iena_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[114\] la_oenb_mprj[114] la_buf_enable\[114\]/B vssd vssd vccd vccd
+ la_buf\[114\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_33_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__417__A mprj_adr_o_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_427_ mprj_adr_o_core[20] vssd vssd vccd vccd _427_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_358_ la_oenb_mprj[90] vssd vssd vccd vccd _358_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[10\] user_to_mprj_in_gates\[10\]/Y vssd vssd vccd vccd la_data_in_mprj[10]
+ sky130_fd_sc_hd__inv_8
XFILLER_6_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[88\] la_data_out_core[88] user_to_mprj_in_gates\[88\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[88\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[59\]_A la_iena_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[29\]_TE mprj_adr_buf\[29\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[50\] la_iena_mprj[50] mprj_logic_high_inst/HI[380] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_800 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_811 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[2\] user_to_mprj_in_gates\[2\]/Y vssd vssd vccd vccd la_data_in_mprj[2]
+ sky130_fd_sc_hd__inv_8
XPHY_822 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_833 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_844 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_888 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_855 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_866 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_877 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_899 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_598 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[14\] _485_/Y la_buf\[14\]/TE vssd vssd vccd vccd la_data_in_core[14] sky130_fd_sc_hd__einvp_8
XFILLER_3_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[7\] _414_/Y mprj_adr_buf\[7\]/TE vssd vssd vccd vccd mprj_adr_o_user[7]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[58\] user_to_mprj_in_gates\[58\]/Y vssd vssd vccd vccd la_data_in_mprj[58]
+ sky130_fd_sc_hd__inv_8
XFILLER_18_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_mprj_dat_buf\[8\]_A _447_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_167 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__610__A la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[114\] la_data_out_core[114] user_to_mprj_in_gates\[114\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[114\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_129 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1205 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[98\] la_iena_mprj[98] mprj_logic_high_inst/HI[428] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf\[70\]_A _541_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[84\]_TE mprj_logic_high_inst/HI[286] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[124\] _392_/Y mprj_logic_high_inst/HI[326] vssd vssd vccd
+ vccd la_oenb_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_0_712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__520__A la_data_out_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[54\] _653_/Y mprj_logic_high_inst/HI[256] vssd vssd vccd
+ vccd la_oenb_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_48_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_226 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[76\] la_oenb_mprj[76] la_buf_enable\[76\]/B vssd vssd vccd vccd la_buf\[76\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_40_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_641 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_652 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_630 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_663 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_685 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_696 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_674 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[88\]_A user_to_mprj_in_gates\[88\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[118\] _589_/Y la_buf\[118\]/TE vssd vssd vccd vccd la_data_in_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_3_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[111\] user_to_mprj_in_gates\[111\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[111] sky130_fd_sc_hd__inv_8
XFILLER_3_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__430__A mprj_adr_o_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[12\]_A user_to_mprj_in_gates\[12\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[115\]_A _586_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__605__A la_oenb_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[18\]_B user_to_mprj_in_gates\[18\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__340__A la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_ena_buf\[13\] la_iena_mprj[13] mprj_logic_high_inst/HI[343] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf\[106\]_A _577_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__515__A la_data_out_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[61\]_B la_buf_enable\[61\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[81\] _552_/Y la_buf\[81\]/TE vssd vssd vccd vccd la_data_in_core[81] sky130_fd_sc_hd__einvp_8
XFILLER_40_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_914 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[108\]_A user_to_mprj_in_gates\[108\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_471 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_460 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__425__A mprj_adr_o_core[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_482 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_493 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1070 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1092 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1081 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2019 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[52\]_B la_buf_enable\[52\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[70\] la_data_out_core[70] user_to_mprj_in_gates\[70\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[70\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_41_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[124\]_B mprj_logic_high_inst/HI[454] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_clk_buf _398_/Y mprj_clk_buf/TE vssd vssd vccd vccd user_clock sky130_fd_sc_hd__einvp_8
XANTENNA__335__A la_oenb_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_2078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[43\]_B la_buf_enable\[43\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1131 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[115\]_B mprj_logic_high_inst/HI[445] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1681 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_460_ mprj_dat_o_core[21] vssd vssd vccd vccd _460_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[17\] _616_/Y mprj_logic_high_inst/HI[219] vssd vssd vccd
+ vccd la_oenb_core[17] sky130_fd_sc_hd__einvp_8
X_391_ la_oenb_mprj[123] vssd vssd vccd vccd _391_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_413 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[39\] la_oenb_mprj[39] la_buf_enable\[39\]/B vssd vssd vccd vccd la_buf\[39\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_41_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[34\]_B la_buf_enable\[34\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_2074 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[3\]_A la_iena_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[101\]_A _369_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[106\]_B mprj_logic_high_inst/HI[436] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_658_ la_oenb_mprj[59] vssd vssd vccd vccd _658_/Y sky130_fd_sc_hd__inv_2
X_589_ la_data_out_mprj[118] vssd vssd vccd vccd _589_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[40\] user_to_mprj_in_gates\[40\]/Y vssd vssd vccd vccd la_data_in_mprj[40]
+ sky130_fd_sc_hd__inv_8
XFILLER_38_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_290 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1219 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_12_1631 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[25\]_B la_buf_enable\[25\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[105\]_A_N la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[119\]_TE mprj_logic_high_inst/HI[321] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_17_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[16\]_B la_buf_enable\[16\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[80\] la_iena_mprj[80] mprj_logic_high_inst/HI[410] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/B sky130_fd_sc_hd__and2_1
XFILLER_11_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_512_ la_data_out_mprj[41] vssd vssd vccd vccd _512_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[33\]_TE la_buf\[33\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_443_ mprj_dat_o_core[4] vssd vssd vccd vccd _443_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[18\]_TE mprj_logic_high_inst/HI[220] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_374_ la_oenb_mprj[106] vssd vssd vccd vccd _374_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[44\] _515_/Y la_buf\[44\]/TE vssd vssd vccd vccd la_data_in_core[44] sky130_fd_sc_hd__einvp_8
XFILLER_9_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[116\] la_iena_mprj[116] mprj_logic_high_inst/HI[446] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[116\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_954 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[100\] _571_/Y la_buf\[100\]/TE vssd vssd vccd vccd la_data_in_core[100] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[86\]_B mprj_logic_high_inst/HI[416] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[88\] user_to_mprj_in_gates\[88\]/Y vssd vssd vccd vccd la_data_in_mprj[88]
+ sky130_fd_sc_hd__inv_8
XFILLER_40_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[33\] la_data_out_core[33] user_to_mprj_in_gates\[33\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[33\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[1\]_TE la_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__613__A la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[56\]_TE la_buf\[56\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_27_324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[3\]_A la_data_out_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1684 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[3\]_A_N la_oenb_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_19_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__523__A la_data_out_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[84\] _352_/Y mprj_logic_high_inst/HI[286] vssd vssd vccd
+ vccd la_oenb_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_46_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_968 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[68\]_B mprj_logic_high_inst/HI[398] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[107\] la_oenb_mprj[107] la_buf_enable\[107\]/B vssd vssd vccd vccd
+ la_buf\[107\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_18_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_426_ mprj_adr_o_core[19] vssd vssd vccd vccd _426_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_357_ la_oenb_mprj[89] vssd vssd vccd vccd _357_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__433__A mprj_adr_o_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[59\]_B mprj_logic_high_inst/HI[389] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__608__A la_oenb_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__343__A la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_927 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[28\]_TE mprj_dat_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[43\] la_iena_mprj[43] mprj_logic_high_inst/HI[373] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__518__A la_data_out_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_801 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_812 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_823 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_834 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_845 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_533 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_856 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[21\] la_oenb_mprj[21] la_buf_enable\[21\]/B vssd vssd vccd vccd la_buf\[21\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_867 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_878 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_889 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__428__A mprj_adr_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1578 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_409_ mprj_adr_o_core[2] vssd vssd vccd vccd _409_/Y sky130_fd_sc_hd__inv_2
XFILLER_15_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[63\]_A_N la_oenb_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[78\]_A_N la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[107\] la_data_out_core[107] user_to_mprj_in_gates\[107\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[107\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__338__A la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[16\]_A_N la_oenb_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_724 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[117\] _385_/Y mprj_logic_high_inst/HI[319] vssd vssd vccd
+ vccd la_oenb_core[117] sky130_fd_sc_hd__einvp_8
XFILLER_0_779 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[47\] _646_/Y mprj_logic_high_inst/HI[249] vssd vssd vccd
+ vccd la_oenb_core[47] sky130_fd_sc_hd__einvp_8
XFILLER_5_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[69\] la_oenb_mprj[69] la_buf_enable\[69\]/B vssd vssd vccd vccd la_buf\[69\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_16_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_620 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_831 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_642 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_653 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_631 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_664 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_686 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_842 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_675 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_697 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[104\] user_to_mprj_in_gates\[104\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[104] sky130_fd_sc_hd__inv_8
XFILLER_38_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[70\] user_to_mprj_in_gates\[70\]/Y vssd vssd vccd vccd la_data_in_mprj[70]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[19\]_TE mprj_adr_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__621__A la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[3\]_TE mprj_adr_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[3\] _442_/Y mprj_dat_buf\[3\]/TE vssd vssd vccd vccd mprj_dat_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_45_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__531__A la_data_out_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[74\] _545_/Y la_buf\[74\]/TE vssd vssd vccd vccd la_data_in_core[74] sky130_fd_sc_hd__einvp_8
XFILLER_43_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_926 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_461 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_450 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_483 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_472 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_494 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1071 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1060 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1082 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1093 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__441__A mprj_dat_o_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[63\] la_data_out_core[63] user_to_mprj_in_gates\[63\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[63\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_35_731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[74\]_TE mprj_logic_high_inst/HI[276] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__616__A la_oenb_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1047 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1301 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__351__A la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_241 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_425 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_390_ la_oenb_mprj[122] vssd vssd vccd vccd _390_/Y sky130_fd_sc_hd__inv_2
XFILLER_9_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__526__A la_data_out_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_668 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1424 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[97\]_TE mprj_logic_high_inst/HI[299] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1181 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_657_ la_oenb_mprj[58] vssd vssd vccd vccd _657_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_712 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_588_ la_data_out_mprj[117] vssd vssd vccd vccd _588_/Y sky130_fd_sc_hd__inv_2
XANTENNA__436__A mprj_adr_o_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[33\] user_to_mprj_in_gates\[33\]/Y vssd vssd vccd vccd la_data_in_mprj[33]
+ sky130_fd_sc_hd__inv_8
XPHY_291 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_280 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_12_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_907 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__346__A la_oenb_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[93\]_A la_data_out_core[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[73\] la_iena_mprj[73] mprj_logic_high_inst/HI[403] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_18_506 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[115\]_B la_buf_enable\[115\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_511_ la_data_out_mprj[40] vssd vssd vccd vccd _511_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[51\] la_oenb_mprj[51] la_buf_enable\[51\]/B vssd vssd vccd vccd la_buf\[51\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_2_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_442_ mprj_dat_o_core[3] vssd vssd vccd vccd _442_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_373_ la_oenb_mprj[105] vssd vssd vccd vccd _373_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[84\]_A la_data_out_core[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[37\] _508_/Y la_buf\[37\]/TE vssd vssd vccd vccd la_data_in_core[37] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[109\] la_iena_mprj[109] mprj_logic_high_inst/HI[439] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[109\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_2104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_443 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[26\] la_data_out_core[26] user_to_mprj_in_gates\[26\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[26\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_gates\[75\]_A la_data_out_core[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_196 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[3\]_B user_to_mprj_in_gates\[3\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[66\]_A la_data_out_core[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_269 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[77\] _345_/Y mprj_logic_high_inst/HI[279] vssd vssd vccd
+ vccd la_oenb_core[77] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[99\] la_oenb_mprj[99] la_buf_enable\[99\]/B vssd vssd vccd vccd la_buf\[99\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_46_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[25\] _464_/Y mprj_dat_buf\[25\]/TE vssd vssd vccd vccd mprj_dat_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_46_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_425_ mprj_adr_o_core[18] vssd vssd vccd vccd _425_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_356_ la_oenb_mprj[88] vssd vssd vccd vccd _356_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[104\]_A_N la_oenb_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2049 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1304 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[57\]_A la_data_out_core[57] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[20\] _427_/Y mprj_adr_buf\[20\]/TE vssd vssd vccd vccd mprj_adr_o_user[20]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[119\]_A_N la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[109\]_TE mprj_logic_high_inst/HI[311] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[7\]_A user_to_mprj_in_gates\[7\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_0_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_361 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_523 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_394 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[48\]_A la_data_out_core[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__624__A la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_534 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1546 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[5\] la_oenb_mprj[5] la_buf_enable\[5\]/B vssd vssd vccd vccd la_buf\[5\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_31_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[23\]_TE la_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1675 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[36\] la_iena_mprj[36] mprj_logic_high_inst/HI[366] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_802 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_42_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_78 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_813 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_824 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_835 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_846 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_857 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_868 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_879 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[39\]_A la_data_out_core[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[14\] la_oenb_mprj[14] la_buf_enable\[14\]/B vssd vssd vccd vccd la_buf\[14\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[123\]_A la_data_out_core[123] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_7_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__534__A la_data_out_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1922 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_623 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_408_ mprj_adr_o_core[1] vssd vssd vccd vccd _408_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[114\]_A la_data_out_core[114] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__444__A mprj_dat_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_898 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_339_ la_oenb_mprj[71] vssd vssd vccd vccd _339_/Y sky130_fd_sc_hd__inv_2
XFILLER_11_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[46\]_TE la_buf\[46\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[93\] la_data_out_core[93] user_to_mprj_in_gates\[93\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[93\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[2\]_A_N la_oenb_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__619__A la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[105\]_A la_data_out_core[105] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_36_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__354__A la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__529__A la_data_out_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_604 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_610 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_632 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_643 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_621 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_665 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_687 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_654 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_676 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_698 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_45_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__439__A mprj_dat_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[63\] user_to_mprj_in_gates\[63\]/Y vssd vssd vccd vccd la_data_in_mprj[63]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[18\]_TE mprj_dat_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1516 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[3\]_B la_buf_enable\[3\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[127\]_A la_iena_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__349__A la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_20_172 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[81\] la_oenb_mprj[81] la_buf_enable\[81\]/B vssd vssd vccd vccd la_buf\[81\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_27_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[118\]_A la_iena_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[62\]_A_N la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[67\] _538_/Y la_buf\[67\]/TE vssd vssd vccd vccd la_data_in_core[67] sky130_fd_sc_hd__einvp_8
XFILLER_16_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_462 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_440 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_451 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[77\]_A_N la_oenb_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1050 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_484 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_473 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_495 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1072 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1061 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1083 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1094 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[123\] _594_/Y la_buf\[123\]/TE vssd vssd vccd vccd la_data_in_core[123] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[15\]_A_N la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[109\]_A la_iena_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[56\] la_data_out_core[56] user_to_mprj_in_gates\[56\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[56\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[40\]_A la_iena_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1059 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__632__A la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1155 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1569 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_35_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[31\]_A la_iena_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__542__A la_data_out_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[98\]_A la_iena_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_656_ la_oenb_mprj[57] vssd vssd vccd vccd _656_/Y sky130_fd_sc_hd__inv_2
X_587_ la_data_out_mprj[116] vssd vssd vccd vccd _587_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[22\]_A la_iena_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_920 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_270 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_292 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_281 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[26\] user_to_mprj_in_gates\[26\]/Y vssd vssd vccd vccd la_data_in_mprj[26]
+ sky130_fd_sc_hd__inv_8
XANTENNA__452__A mprj_dat_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[89\]_A la_iena_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__627__A la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_234 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[13\]_A la_iena_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__362__A la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[66\] la_iena_mprj[66] mprj_logic_high_inst/HI[396] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_510_ la_data_out_mprj[39] vssd vssd vccd vccd _510_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_irq_ena_buf\[0\]_A user_irq_ena[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_441_ mprj_dat_o_core[2] vssd vssd vccd vccd _441_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[22\] _621_/Y mprj_logic_high_inst/HI[224] vssd vssd vccd
+ vccd la_oenb_core[22] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[4\] _603_/Y mprj_logic_high_inst/HI[206] vssd vssd vccd
+ vccd la_oenb_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_14_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__537__A la_data_out_mprj[66] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[44\] la_oenb_mprj[44] la_buf_enable\[44\]/B vssd vssd vccd vccd la_buf\[44\]/TE
+ sky130_fd_sc_hd__and2b_1
X_372_ la_oenb_mprj[104] vssd vssd vccd vccd _372_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_941 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2116 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1288 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__447__A mprj_dat_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_639_ la_oenb_mprj[40] vssd vssd vccd vccd _639_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[19\] la_data_out_core[19] user_to_mprj_in_gates\[19\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[19\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_1960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[60\]_A user_to_mprj_in_gates\[60\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__357__A la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[87\]_TE mprj_logic_high_inst/HI[289] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_79 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_1596 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[18\] _457_/Y mprj_dat_buf\[18\]/TE vssd vssd vccd vccd mprj_dat_o_user[18]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[51\]_A user_to_mprj_in_gates\[51\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1564 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_424_ mprj_adr_o_core[17] vssd vssd vccd vccd _424_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2006 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_355_ la_oenb_mprj[87] vssd vssd vccd vccd _355_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_ena_buf\[121\] la_iena_mprj[121] mprj_logic_high_inst/HI[451] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[121\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[13\] _420_/Y mprj_adr_buf\[13\]/TE vssd vssd vccd vccd mprj_adr_o_user[13]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[127\] user_to_mprj_in_gates\[127\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[127] sky130_fd_sc_hd__inv_8
XFILLER_9_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[93\] user_to_mprj_in_gates\[93\]/Y vssd vssd vccd vccd la_data_in_mprj[93]
+ sky130_fd_sc_hd__inv_8
XFILLER_46_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_874 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[82\]_A _553_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1558 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__640__A la_oenb_mprj[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[0\] la_data_out_core[0] user_to_mprj_in_gates\[0\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[0\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[33\]_A user_to_mprj_in_gates\[33\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[29\] la_iena_mprj[29] mprj_logic_high_inst/HI[359] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/B sky130_fd_sc_hd__and2_1
XPHY_803 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_814 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_825 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_836 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_847 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_858 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_869 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__550__A la_data_out_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[24\]_A user_to_mprj_in_gates\[24\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf\[97\] _568_/Y la_buf\[97\]/TE vssd vssd vccd vccd la_data_in_core[97] sky130_fd_sc_hd__einvp_8
XFILLER_4_1225 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[2\] la_iena_mprj[2] mprj_logic_high_inst/HI[332] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[2\]/B sky130_fd_sc_hd__and2_1
Xla_buf_enable\[112\] la_oenb_mprj[112] la_buf_enable\[112\]/B vssd vssd vccd vccd
+ la_buf\[112\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_46_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf\[127\]_A _598_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_811 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_800 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_407_ mprj_adr_o_core[0] vssd vssd vccd vccd _407_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_338_ la_oenb_mprj[70] vssd vssd vccd vccd _338_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[64\]_A _535_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1179 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_B la_buf_enable\[82\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__460__A mprj_dat_o_core[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[86\] la_data_out_core[86] user_to_mprj_in_gates\[86\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[86\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[15\]_A user_to_mprj_in_gates\[15\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf\[118\]_A _589_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__635__A la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1079 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_B la_buf_enable\[73\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__370__A la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[103\]_A_N la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[118\]_A_N la_oenb_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_600 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_611 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__545__A la_data_out_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[109\]_A _580_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[0\] user_to_mprj_in_gates\[0\]/Y vssd vssd vccd vccd la_data_in_mprj[0]
+ sky130_fd_sc_hd__inv_8
XPHY_633 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_644 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_622 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_666 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_677 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_655 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_688 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_699 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[12\] _483_/Y la_buf\[12\]/TE vssd vssd vccd vccd la_data_in_core[12] sky130_fd_sc_hd__einvp_8
Xla_buf\[8\] _479_/Y la_buf\[8\]/TE vssd vssd vccd vccd la_data_in_core[8] sky130_fd_sc_hd__einvp_8
XANTENNA_la_buf_enable\[64\]_B la_buf_enable\[64\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[5\] _412_/Y mprj_adr_buf\[5\]/TE vssd vssd vccd vccd mprj_adr_o_user[5]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[13\]_TE la_buf\[13\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[56\] user_to_mprj_in_gates\[56\]/Y vssd vssd vccd vccd la_data_in_mprj[56]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__455__A mprj_dat_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_490 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[55\]_B la_buf_enable\[55\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[127\]_B mprj_logic_high_inst/HI[457] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_gates\[112\] la_data_out_core[112] user_to_mprj_in_gates\[112\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[112\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_619 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__365__A la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_B la_buf_enable\[46\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_195 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[96\] la_iena_mprj[96] mprj_logic_high_inst/HI[426] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[122\] _390_/Y mprj_logic_high_inst/HI[324] vssd vssd vccd
+ vccd la_oenb_core[122] sky130_fd_sc_hd__einvp_8
Xmprj_sel_buf\[3\] _406_/Y mprj_sel_buf\[3\]/TE vssd vssd vccd vccd mprj_sel_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[118\]_B mprj_logic_high_inst/HI[448] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[52\] _651_/Y mprj_logic_high_inst/HI[254] vssd vssd vccd
+ vccd la_oenb_core[52] sky130_fd_sc_hd__einvp_8
XFILLER_5_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[74\] la_oenb_mprj[74] la_buf_enable\[74\]/B vssd vssd vccd vccd la_buf\[74\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_1228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_1386 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[1\]_A_N la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_430 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_441 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_452 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1040 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_485 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_474 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_463 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1073 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1062 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1051 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_496 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1095 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1084 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[37\]_B la_buf_enable\[37\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[116\] _587_/Y la_buf\[116\]/TE vssd vssd vccd vccd la_data_in_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_4_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[6\]_A la_iena_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[49\] la_data_out_core[49] user_to_mprj_in_gates\[49\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[49\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_35_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[4\]_TE la_buf\[4\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_B la_buf_enable\[28\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[59\]_TE la_buf\[59\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_6_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[11\] la_iena_mprj[11] mprj_logic_high_inst/HI[341] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[19\]_B la_buf_enable\[19\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1404 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1510 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_655_ la_oenb_mprj[56] vssd vssd vccd vccd _655_/Y sky130_fd_sc_hd__inv_2
X_586_ la_data_out_mprj[115] vssd vssd vccd vccd _586_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_260 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_293 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_282 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_271 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[19\] user_to_mprj_in_gates\[19\]/Y vssd vssd vccd vccd la_data_in_mprj[19]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[13\]_B mprj_logic_high_inst/HI[343] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA__643__A la_oenb_mprj[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1712 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[61\]_A_N la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[76\]_A_N la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[6\]_A la_data_out_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[59\] la_iena_mprj[59] mprj_logic_high_inst/HI[389] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/B sky130_fd_sc_hd__and2_1
XFILLER_46_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_541 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_irq_ena_buf\[0\]_B user_irq_ena_buf\[0\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_440_ mprj_dat_o_core[1] vssd vssd vccd vccd _440_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_371_ la_oenb_mprj[103] vssd vssd vccd vccd _371_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[37\] la_oenb_mprj[37] la_buf_enable\[37\]/B vssd vssd vccd vccd la_buf\[37\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[15\] _614_/Y mprj_logic_high_inst/HI[217] vssd vssd vccd
+ vccd la_oenb_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_39_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[14\]_A_N la_oenb_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__553__A la_data_out_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[29\]_A_N la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_638_ la_oenb_mprj[39] vssd vssd vccd vccd _638_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_569_ la_data_out_mprj[98] vssd vssd vccd vccd _569_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__463__A mprj_dat_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__638__A la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2090 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_1607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__373__A la_oenb_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__548__A la_data_out_mprj[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_423_ mprj_adr_o_core[16] vssd vssd vccd vccd _423_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_354_ la_oenb_mprj[86] vssd vssd vccd vccd _354_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[42\] _513_/Y la_buf\[42\]/TE vssd vssd vccd vccd la_data_in_core[42] sky130_fd_sc_hd__einvp_8
XFILLER_31_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[114\] la_iena_mprj[114] mprj_logic_high_inst/HI[444] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[114\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[31\]_TE mprj_logic_high_inst/HI[233] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1751 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_971 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[86\] user_to_mprj_in_gates\[86\]/Y vssd vssd vccd vccd la_data_in_mprj[86]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_625 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__458__A mprj_dat_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[31\] la_data_out_core[31] user_to_mprj_in_gates\[31\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[31\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_36_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_adr_buf\[6\]_TE mprj_adr_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_919 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1600 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__368__A la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_135 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_804 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_815 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_826 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[54\]_TE mprj_logic_high_inst/HI[256] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_837 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_848 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_859 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[82\] _350_/Y mprj_logic_high_inst/HI[284] vssd vssd vccd
+ vccd la_oenb_core[82] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[30\] _469_/Y mprj_dat_buf\[30\]/TE vssd vssd vccd vccd mprj_dat_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_606 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[105\] la_oenb_mprj[105] la_buf_enable\[105\]/B vssd vssd vccd vccd
+ la_buf\[105\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_33_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_864 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_91 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_406_ mprj_sel_o_core[3] vssd vssd vccd vccd _406_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_337_ la_oenb_mprj[69] vssd vssd vccd vccd _337_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1148 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[79\] la_data_out_core[79] user_to_mprj_in_gates\[79\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[79\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_37_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[92\]_TE la_buf\[92\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[77\]_TE mprj_logic_high_inst/HI[279] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1345 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__651__A la_oenb_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[41\] la_iena_mprj[41] mprj_logic_high_inst/HI[371] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/B sky130_fd_sc_hd__and2_1
XFILLER_28_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_cyc_buf_TE mprj_cyc_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_601 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_634 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_612 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_623 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_667 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_645 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_678 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_656 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_689 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__561__A la_data_out_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[49\] user_to_mprj_in_gates\[49\]/Y vssd vssd vccd vccd la_data_in_mprj[49]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_661 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__471__A la_data_out_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[105\] la_data_out_core[105] user_to_mprj_in_gates\[105\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[105\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1443 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__646__A la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj2_logic_high_inst mprj2_pwrgood/A vccd2 vssd2 mprj2_logic_high
XFILLER_25_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_141 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__381__A la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[89\] la_iena_mprj[89] mprj_logic_high_inst/HI[419] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[115\] _383_/Y mprj_logic_high_inst/HI[317] vssd vssd vccd
+ vccd la_oenb_core[115] sky130_fd_sc_hd__einvp_8
XFILLER_48_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[45\] _644_/Y mprj_logic_high_inst/HI[247] vssd vssd vccd
+ vccd la_oenb_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_5_1376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[67\] la_oenb_mprj[67] la_buf_enable\[67\]/B vssd vssd vccd vccd la_buf\[67\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__556__A la_data_out_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_431 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_442 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_453 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_420 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1030 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1041 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_486 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_475 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_464 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1074 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1063 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1052 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_497 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1096 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1085 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_rstn_buf_TE mprj_rstn_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[6\]_B mprj_logic_high_inst/HI[336] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[109\] _580_/Y la_buf\[109\]/TE vssd vssd vccd vccd la_data_in_core[109] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[102\] user_to_mprj_in_gates\[102\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[102] sky130_fd_sc_hd__inv_8
XFILLER_47_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__466__A mprj_dat_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[102\]_A_N la_oenb_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_494 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_2038 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[117\]_A_N la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[1\] _440_/Y mprj_dat_buf\[1\]/TE vssd vssd vccd vccd mprj_dat_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_logic_high_inst mprj_rstn_buf/TE la_buf_enable\[26\]/B la_buf_enable\[27\]/B
+ la_buf_enable\[28\]/B la_buf_enable\[29\]/B la_buf_enable\[30\]/B la_buf_enable\[31\]/B
+ la_buf_enable\[32\]/B la_buf_enable\[33\]/B la_buf_enable\[34\]/B la_buf_enable\[35\]/B
+ mprj_adr_buf\[0\]/TE la_buf_enable\[36\]/B la_buf_enable\[37\]/B la_buf_enable\[38\]/B
+ la_buf_enable\[39\]/B la_buf_enable\[40\]/B la_buf_enable\[41\]/B la_buf_enable\[42\]/B
+ la_buf_enable\[43\]/B la_buf_enable\[44\]/B la_buf_enable\[45\]/B mprj_adr_buf\[1\]/TE
+ la_buf_enable\[46\]/B la_buf_enable\[47\]/B la_buf_enable\[48\]/B la_buf_enable\[49\]/B
+ la_buf_enable\[50\]/B la_buf_enable\[51\]/B la_buf_enable\[52\]/B la_buf_enable\[53\]/B
+ la_buf_enable\[54\]/B la_buf_enable\[55\]/B mprj_adr_buf\[2\]/TE la_buf_enable\[56\]/B
+ la_buf_enable\[57\]/B la_buf_enable\[58\]/B la_buf_enable\[59\]/B la_buf_enable\[60\]/B
+ la_buf_enable\[61\]/B la_buf_enable\[62\]/B la_buf_enable\[63\]/B la_buf_enable\[64\]/B
+ la_buf_enable\[65\]/B mprj_adr_buf\[3\]/TE la_buf_enable\[66\]/B la_buf_enable\[67\]/B
+ la_buf_enable\[68\]/B la_buf_enable\[69\]/B la_buf_enable\[70\]/B la_buf_enable\[71\]/B
+ la_buf_enable\[72\]/B la_buf_enable\[73\]/B la_buf_enable\[74\]/B la_buf_enable\[75\]/B
+ mprj_adr_buf\[4\]/TE la_buf_enable\[76\]/B la_buf_enable\[77\]/B la_buf_enable\[78\]/B
+ la_buf_enable\[79\]/B la_buf_enable\[80\]/B la_buf_enable\[81\]/B la_buf_enable\[82\]/B
+ la_buf_enable\[83\]/B la_buf_enable\[84\]/B la_buf_enable\[85\]/B mprj_adr_buf\[5\]/TE
+ la_buf_enable\[86\]/B la_buf_enable\[87\]/B la_buf_enable\[88\]/B la_buf_enable\[89\]/B
+ la_buf_enable\[90\]/B la_buf_enable\[91\]/B la_buf_enable\[92\]/B la_buf_enable\[93\]/B
+ la_buf_enable\[94\]/B la_buf_enable\[95\]/B mprj_adr_buf\[6\]/TE la_buf_enable\[96\]/B
+ la_buf_enable\[97\]/B la_buf_enable\[98\]/B la_buf_enable\[99\]/B la_buf_enable\[100\]/B
+ la_buf_enable\[101\]/B la_buf_enable\[102\]/B la_buf_enable\[103\]/B la_buf_enable\[104\]/B
+ la_buf_enable\[105\]/B mprj_adr_buf\[7\]/TE la_buf_enable\[106\]/B la_buf_enable\[107\]/B
+ la_buf_enable\[108\]/B la_buf_enable\[109\]/B la_buf_enable\[110\]/B la_buf_enable\[111\]/B
+ la_buf_enable\[112\]/B la_buf_enable\[113\]/B la_buf_enable\[114\]/B la_buf_enable\[115\]/B
+ mprj_adr_buf\[8\]/TE la_buf_enable\[116\]/B la_buf_enable\[117\]/B la_buf_enable\[118\]/B
+ la_buf_enable\[119\]/B la_buf_enable\[120\]/B la_buf_enable\[121\]/B la_buf_enable\[122\]/B
+ la_buf_enable\[123\]/B la_buf_enable\[124\]/B la_buf_enable\[125\]/B mprj_adr_buf\[9\]/TE
+ mprj_clk_buf/TE la_buf_enable\[126\]/B la_buf_enable\[127\]/B mprj_logic_high_inst/HI[202]
+ mprj_logic_high_inst/HI[203] mprj_logic_high_inst/HI[204] mprj_logic_high_inst/HI[205]
+ mprj_logic_high_inst/HI[206] mprj_logic_high_inst/HI[207] mprj_logic_high_inst/HI[208]
+ mprj_logic_high_inst/HI[209] mprj_adr_buf\[10\]/TE mprj_logic_high_inst/HI[210]
+ mprj_logic_high_inst/HI[211] mprj_logic_high_inst/HI[212] mprj_logic_high_inst/HI[213]
+ mprj_logic_high_inst/HI[214] mprj_logic_high_inst/HI[215] mprj_logic_high_inst/HI[216]
+ mprj_logic_high_inst/HI[217] mprj_logic_high_inst/HI[218] mprj_logic_high_inst/HI[219]
+ mprj_adr_buf\[11\]/TE mprj_logic_high_inst/HI[220] mprj_logic_high_inst/HI[221]
+ mprj_logic_high_inst/HI[222] mprj_logic_high_inst/HI[223] mprj_logic_high_inst/HI[224]
+ mprj_logic_high_inst/HI[225] mprj_logic_high_inst/HI[226] mprj_logic_high_inst/HI[227]
+ mprj_logic_high_inst/HI[228] mprj_logic_high_inst/HI[229] mprj_adr_buf\[12\]/TE
+ mprj_logic_high_inst/HI[230] mprj_logic_high_inst/HI[231] mprj_logic_high_inst/HI[232]
+ mprj_logic_high_inst/HI[233] mprj_logic_high_inst/HI[234] mprj_logic_high_inst/HI[235]
+ mprj_logic_high_inst/HI[236] mprj_logic_high_inst/HI[237] mprj_logic_high_inst/HI[238]
+ mprj_logic_high_inst/HI[239] mprj_adr_buf\[13\]/TE mprj_logic_high_inst/HI[240]
+ mprj_logic_high_inst/HI[241] mprj_logic_high_inst/HI[242] mprj_logic_high_inst/HI[243]
+ mprj_logic_high_inst/HI[244] mprj_logic_high_inst/HI[245] mprj_logic_high_inst/HI[246]
+ mprj_logic_high_inst/HI[247] mprj_logic_high_inst/HI[248] mprj_logic_high_inst/HI[249]
+ mprj_adr_buf\[14\]/TE mprj_logic_high_inst/HI[250] mprj_logic_high_inst/HI[251]
+ mprj_logic_high_inst/HI[252] mprj_logic_high_inst/HI[253] mprj_logic_high_inst/HI[254]
+ mprj_logic_high_inst/HI[255] mprj_logic_high_inst/HI[256] mprj_logic_high_inst/HI[257]
+ mprj_logic_high_inst/HI[258] mprj_logic_high_inst/HI[259] mprj_adr_buf\[15\]/TE
+ mprj_logic_high_inst/HI[260] mprj_logic_high_inst/HI[261] mprj_logic_high_inst/HI[262]
+ mprj_logic_high_inst/HI[263] mprj_logic_high_inst/HI[264] mprj_logic_high_inst/HI[265]
+ mprj_logic_high_inst/HI[266] mprj_logic_high_inst/HI[267] mprj_logic_high_inst/HI[268]
+ mprj_logic_high_inst/HI[269] mprj_adr_buf\[16\]/TE mprj_logic_high_inst/HI[270]
+ mprj_logic_high_inst/HI[271] mprj_logic_high_inst/HI[272] mprj_logic_high_inst/HI[273]
+ mprj_logic_high_inst/HI[274] mprj_logic_high_inst/HI[275] mprj_logic_high_inst/HI[276]
+ mprj_logic_high_inst/HI[277] mprj_logic_high_inst/HI[278] mprj_logic_high_inst/HI[279]
+ mprj_adr_buf\[17\]/TE mprj_logic_high_inst/HI[280] mprj_logic_high_inst/HI[281]
+ mprj_logic_high_inst/HI[282] mprj_logic_high_inst/HI[283] mprj_logic_high_inst/HI[284]
+ mprj_logic_high_inst/HI[285] mprj_logic_high_inst/HI[286] mprj_logic_high_inst/HI[287]
+ mprj_logic_high_inst/HI[288] mprj_logic_high_inst/HI[289] mprj_adr_buf\[18\]/TE
+ mprj_logic_high_inst/HI[290] mprj_logic_high_inst/HI[291] mprj_logic_high_inst/HI[292]
+ mprj_logic_high_inst/HI[293] mprj_logic_high_inst/HI[294] mprj_logic_high_inst/HI[295]
+ mprj_logic_high_inst/HI[296] mprj_logic_high_inst/HI[297] mprj_logic_high_inst/HI[298]
+ mprj_logic_high_inst/HI[299] mprj_adr_buf\[19\]/TE mprj_clk2_buf/TE mprj_logic_high_inst/HI[300]
+ mprj_logic_high_inst/HI[301] mprj_logic_high_inst/HI[302] mprj_logic_high_inst/HI[303]
+ mprj_logic_high_inst/HI[304] mprj_logic_high_inst/HI[305] mprj_logic_high_inst/HI[306]
+ mprj_logic_high_inst/HI[307] mprj_logic_high_inst/HI[308] mprj_logic_high_inst/HI[309]
+ mprj_adr_buf\[20\]/TE mprj_logic_high_inst/HI[310] mprj_logic_high_inst/HI[311]
+ mprj_logic_high_inst/HI[312] mprj_logic_high_inst/HI[313] mprj_logic_high_inst/HI[314]
+ mprj_logic_high_inst/HI[315] mprj_logic_high_inst/HI[316] mprj_logic_high_inst/HI[317]
+ mprj_logic_high_inst/HI[318] mprj_logic_high_inst/HI[319] mprj_adr_buf\[21\]/TE
+ mprj_logic_high_inst/HI[320] mprj_logic_high_inst/HI[321] mprj_logic_high_inst/HI[322]
+ mprj_logic_high_inst/HI[323] mprj_logic_high_inst/HI[324] mprj_logic_high_inst/HI[325]
+ mprj_logic_high_inst/HI[326] mprj_logic_high_inst/HI[327] mprj_logic_high_inst/HI[328]
+ mprj_logic_high_inst/HI[329] mprj_adr_buf\[22\]/TE mprj_logic_high_inst/HI[330]
+ mprj_logic_high_inst/HI[331] mprj_logic_high_inst/HI[332] mprj_logic_high_inst/HI[333]
+ mprj_logic_high_inst/HI[334] mprj_logic_high_inst/HI[335] mprj_logic_high_inst/HI[336]
+ mprj_logic_high_inst/HI[337] mprj_logic_high_inst/HI[338] mprj_logic_high_inst/HI[339]
+ mprj_adr_buf\[23\]/TE mprj_logic_high_inst/HI[340] mprj_logic_high_inst/HI[341]
+ mprj_logic_high_inst/HI[342] mprj_logic_high_inst/HI[343] mprj_logic_high_inst/HI[344]
+ mprj_logic_high_inst/HI[345] mprj_logic_high_inst/HI[346] mprj_logic_high_inst/HI[347]
+ mprj_logic_high_inst/HI[348] mprj_logic_high_inst/HI[349] mprj_adr_buf\[24\]/TE
+ mprj_logic_high_inst/HI[350] mprj_logic_high_inst/HI[351] mprj_logic_high_inst/HI[352]
+ mprj_logic_high_inst/HI[353] mprj_logic_high_inst/HI[354] mprj_logic_high_inst/HI[355]
+ mprj_logic_high_inst/HI[356] mprj_logic_high_inst/HI[357] mprj_logic_high_inst/HI[358]
+ mprj_logic_high_inst/HI[359] mprj_adr_buf\[25\]/TE mprj_logic_high_inst/HI[360]
+ mprj_logic_high_inst/HI[361] mprj_logic_high_inst/HI[362] mprj_logic_high_inst/HI[363]
+ mprj_logic_high_inst/HI[364] mprj_logic_high_inst/HI[365] mprj_logic_high_inst/HI[366]
+ mprj_logic_high_inst/HI[367] mprj_logic_high_inst/HI[368] mprj_logic_high_inst/HI[369]
+ mprj_adr_buf\[26\]/TE mprj_logic_high_inst/HI[370] mprj_logic_high_inst/HI[371]
+ mprj_logic_high_inst/HI[372] mprj_logic_high_inst/HI[373] mprj_logic_high_inst/HI[374]
+ mprj_logic_high_inst/HI[375] mprj_logic_high_inst/HI[376] mprj_logic_high_inst/HI[377]
+ mprj_logic_high_inst/HI[378] mprj_logic_high_inst/HI[379] mprj_adr_buf\[27\]/TE
+ mprj_logic_high_inst/HI[380] mprj_logic_high_inst/HI[381] mprj_logic_high_inst/HI[382]
+ mprj_logic_high_inst/HI[383] mprj_logic_high_inst/HI[384] mprj_logic_high_inst/HI[385]
+ mprj_logic_high_inst/HI[386] mprj_logic_high_inst/HI[387] mprj_logic_high_inst/HI[388]
+ mprj_logic_high_inst/HI[389] mprj_adr_buf\[28\]/TE mprj_logic_high_inst/HI[390]
+ mprj_logic_high_inst/HI[391] mprj_logic_high_inst/HI[392] mprj_logic_high_inst/HI[393]
+ mprj_logic_high_inst/HI[394] mprj_logic_high_inst/HI[395] mprj_logic_high_inst/HI[396]
+ mprj_logic_high_inst/HI[397] mprj_logic_high_inst/HI[398] mprj_logic_high_inst/HI[399]
+ mprj_adr_buf\[29\]/TE mprj_cyc_buf/TE mprj_logic_high_inst/HI[400] mprj_logic_high_inst/HI[401]
+ mprj_logic_high_inst/HI[402] mprj_logic_high_inst/HI[403] mprj_logic_high_inst/HI[404]
+ mprj_logic_high_inst/HI[405] mprj_logic_high_inst/HI[406] mprj_logic_high_inst/HI[407]
+ mprj_logic_high_inst/HI[408] mprj_logic_high_inst/HI[409] mprj_adr_buf\[30\]/TE
+ mprj_logic_high_inst/HI[410] mprj_logic_high_inst/HI[411] mprj_logic_high_inst/HI[412]
+ mprj_logic_high_inst/HI[413] mprj_logic_high_inst/HI[414] mprj_logic_high_inst/HI[415]
+ mprj_logic_high_inst/HI[416] mprj_logic_high_inst/HI[417] mprj_logic_high_inst/HI[418]
+ mprj_logic_high_inst/HI[419] mprj_adr_buf\[31\]/TE mprj_logic_high_inst/HI[420]
+ mprj_logic_high_inst/HI[421] mprj_logic_high_inst/HI[422] mprj_logic_high_inst/HI[423]
+ mprj_logic_high_inst/HI[424] mprj_logic_high_inst/HI[425] mprj_logic_high_inst/HI[426]
+ mprj_logic_high_inst/HI[427] mprj_logic_high_inst/HI[428] mprj_logic_high_inst/HI[429]
+ mprj_dat_buf\[0\]/TE mprj_logic_high_inst/HI[430] mprj_logic_high_inst/HI[431] mprj_logic_high_inst/HI[432]
+ mprj_logic_high_inst/HI[433] mprj_logic_high_inst/HI[434] mprj_logic_high_inst/HI[435]
+ mprj_logic_high_inst/HI[436] mprj_logic_high_inst/HI[437] mprj_logic_high_inst/HI[438]
+ mprj_logic_high_inst/HI[439] mprj_dat_buf\[1\]/TE mprj_logic_high_inst/HI[440] mprj_logic_high_inst/HI[441]
+ mprj_logic_high_inst/HI[442] mprj_logic_high_inst/HI[443] mprj_logic_high_inst/HI[444]
+ mprj_logic_high_inst/HI[445] mprj_logic_high_inst/HI[446] mprj_logic_high_inst/HI[447]
+ mprj_logic_high_inst/HI[448] mprj_logic_high_inst/HI[449] mprj_dat_buf\[2\]/TE mprj_logic_high_inst/HI[450]
+ mprj_logic_high_inst/HI[451] mprj_logic_high_inst/HI[452] mprj_logic_high_inst/HI[453]
+ mprj_logic_high_inst/HI[454] mprj_logic_high_inst/HI[455] mprj_logic_high_inst/HI[456]
+ mprj_logic_high_inst/HI[457] user_irq_ena_buf\[0\]/B user_irq_ena_buf\[1\]/B mprj_dat_buf\[3\]/TE
+ user_irq_ena_buf\[2\]/B mprj_pwrgood/A mprj_dat_buf\[4\]/TE mprj_dat_buf\[5\]/TE
+ mprj_dat_buf\[6\]/TE mprj_dat_buf\[7\]/TE mprj_stb_buf/TE mprj_dat_buf\[8\]/TE mprj_dat_buf\[9\]/TE
+ mprj_dat_buf\[10\]/TE mprj_dat_buf\[11\]/TE mprj_dat_buf\[12\]/TE mprj_dat_buf\[13\]/TE
+ mprj_dat_buf\[14\]/TE mprj_dat_buf\[15\]/TE mprj_dat_buf\[16\]/TE mprj_dat_buf\[17\]/TE
+ mprj_we_buf/TE mprj_dat_buf\[18\]/TE mprj_dat_buf\[19\]/TE mprj_dat_buf\[20\]/TE
+ mprj_dat_buf\[21\]/TE mprj_dat_buf\[22\]/TE mprj_dat_buf\[23\]/TE mprj_dat_buf\[24\]/TE
+ mprj_dat_buf\[25\]/TE mprj_dat_buf\[26\]/TE mprj_dat_buf\[27\]/TE mprj_sel_buf\[0\]/TE
+ mprj_dat_buf\[28\]/TE mprj_dat_buf\[29\]/TE mprj_dat_buf\[30\]/TE mprj_dat_buf\[31\]/TE
+ la_buf_enable\[0\]/B la_buf_enable\[1\]/B la_buf_enable\[2\]/B la_buf_enable\[3\]/B
+ la_buf_enable\[4\]/B la_buf_enable\[5\]/B mprj_sel_buf\[1\]/TE la_buf_enable\[6\]/B
+ la_buf_enable\[7\]/B la_buf_enable\[8\]/B la_buf_enable\[9\]/B la_buf_enable\[10\]/B
+ la_buf_enable\[11\]/B la_buf_enable\[12\]/B la_buf_enable\[13\]/B la_buf_enable\[14\]/B
+ la_buf_enable\[15\]/B mprj_sel_buf\[2\]/TE la_buf_enable\[16\]/B la_buf_enable\[17\]/B
+ la_buf_enable\[18\]/B la_buf_enable\[19\]/B la_buf_enable\[20\]/B la_buf_enable\[21\]/B
+ la_buf_enable\[22\]/B la_buf_enable\[23\]/B la_buf_enable\[24\]/B la_buf_enable\[25\]/B
+ mprj_sel_buf\[3\]/TE vccd1 vssd1 mprj_logic_high
XFILLER_27_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__376__A la_oenb_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[96\]_A la_data_out_core[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1860 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1893 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2034 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[20\]_A la_data_out_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1416 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_654_ la_oenb_mprj[55] vssd vssd vccd vccd _654_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[72\] _543_/Y la_buf\[72\]/TE vssd vssd vccd vccd la_data_in_core[72] sky130_fd_sc_hd__einvp_8
XFILLER_29_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_38_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_585_ la_data_out_mprj[114] vssd vssd vccd vccd _585_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[87\]_A la_data_out_core[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_261 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_250 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1495 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_294 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_283 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_272 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[11\]_A la_data_out_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_325 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[61\] la_data_out_core[61] user_to_mprj_in_gates\[61\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[61\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1582 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[78\]_A la_data_out_core[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[26\]_TE la_buf\[26\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1664 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[0\]_A_N la_oenb_mprj[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[6\]_B user_to_mprj_in_gates\[6\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_39_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_370_ la_oenb_mprj[102] vssd vssd vccd vccd _370_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[69\]_A la_data_out_core[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_589 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_637_ la_oenb_mprj[38] vssd vssd vccd vccd _637_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_568_ la_data_out_mprj[97] vssd vssd vccd vccd _568_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_499_ la_data_out_mprj[28] vssd vssd vccd vccd _499_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[31\] user_to_mprj_in_gates\[31\]/Y vssd vssd vccd vccd la_data_in_mprj[31]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[49\]_TE la_buf\[49\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_781 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_774 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__654__A la_oenb_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1565 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[71\] la_iena_mprj[71] mprj_logic_high_inst/HI[401] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_422_ mprj_adr_o_core[15] vssd vssd vccd vccd _422_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[126\]_A la_data_out_core[126] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__564__A la_data_out_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_353_ la_oenb_mprj[85] vssd vssd vccd vccd _353_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf\[35\] _506_/Y la_buf\[35\]/TE vssd vssd vccd vccd la_data_in_core[35] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[107\] la_iena_mprj[107] mprj_logic_high_inst/HI[437] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[107\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_784 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_983 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1414 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1881 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[79\] user_to_mprj_in_gates\[79\]/Y vssd vssd vccd vccd la_data_in_mprj[79]
+ sky130_fd_sc_hd__inv_8
XFILLER_40_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1817 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[60\]_A_N la_oenb_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[117\]_A la_data_out_core[117] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_44_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__474__A la_data_out_mprj[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[24\] la_data_out_core[24] user_to_mprj_in_gates\[24\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[24\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf_enable\[75\]_A_N la_oenb_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1831 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[13\]_A_N la_oenb_mprj[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1853 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__649__A la_oenb_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[28\]_A_N la_oenb_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[108\]_A la_data_out_core[108] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__384__A la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_805 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_816 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_827 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_838 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_849 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1925 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[75\] _343_/Y mprj_logic_high_inst/HI[277] vssd vssd vccd
+ vccd la_oenb_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_8_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[97\] la_oenb_mprj[97] la_buf_enable\[97\]/B vssd vssd vccd vccd la_buf\[97\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_43_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[23\] _462_/Y mprj_dat_buf\[23\]/TE vssd vssd vccd vccd mprj_dat_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XFILLER_47_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__559__A la_data_out_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_405_ mprj_sel_o_core[2] vssd vssd vccd vccd _405_/Y sky130_fd_sc_hd__inv_2
XPHY_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_336_ la_oenb_mprj[68] vssd vssd vccd vccd _336_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__469__A mprj_dat_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1987 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[122\]_TE mprj_logic_high_inst/HI[324] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[70\]_A la_iena_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[3\] la_oenb_mprj[3] la_buf_enable\[3\]/B vssd vssd vccd vccd la_buf\[3\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[6\]_B la_buf_enable\[6\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__379__A la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[21\]_TE mprj_logic_high_inst/HI[223] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[34\] la_iena_mprj[34] mprj_logic_high_inst/HI[364] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_ena_buf\[61\]_A la_iena_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_602 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_635 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_613 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_624 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_646 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_668 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_657 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_679 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[12\] la_oenb_mprj[12] la_buf_enable\[12\]/B vssd vssd vccd vccd la_buf\[12\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_32_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xpowergood_check mprj2_vdd_pwrgood/A mprj_vdd_pwrgood/A vccd vssd vdda1 vssa1 vdda2
+ vssa2 mgmt_protect_hv
XFILLER_19_467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[52\]_A la_iena_mprj[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[91\] la_data_out_core[91] user_to_mprj_in_gates\[91\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[91\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[44\]_TE mprj_logic_high_inst/HI[246] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[0\]_A _403_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[43\]_A la_iena_mprj[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[108\] _376_/Y mprj_logic_high_inst/HI[310] vssd vssd vccd
+ vccd la_oenb_core[108] sky130_fd_sc_hd__einvp_8
XFILLER_5_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[38\] _637_/Y mprj_logic_high_inst/HI[240] vssd vssd vccd
+ vccd la_oenb_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_28_297 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[34\]_A la_iena_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_410 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_432 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_443 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_421 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1031 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1020 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_476 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_465 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_454 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1064 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1053 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1042 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__572__A la_data_out_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_487 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_498 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1075 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1097 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1086 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[1\]_A _440_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[67\]_TE mprj_logic_high_inst/HI[269] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1563 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_47_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[61\] user_to_mprj_in_gates\[61\]/Y vssd vssd vccd vccd la_data_in_mprj[61]
+ sky130_fd_sc_hd__inv_8
XFILLER_19_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[25\]_A la_iena_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__482__A la_data_out_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_dat_buf\[31\]_TE mprj_dat_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[90\]_A user_to_mprj_in_gates\[90\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__657__A la_oenb_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[16\]_A la_iena_mprj[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__392__A la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2046 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__567__A la_data_out_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_653_ la_oenb_mprj[54] vssd vssd vccd vccd _653_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[65\] _536_/Y la_buf\[65\]/TE vssd vssd vccd vccd la_data_in_core[65] sky130_fd_sc_hd__einvp_8
XFILLER_32_716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_584_ la_data_out_mprj[113] vssd vssd vccd vccd _584_/Y sky130_fd_sc_hd__inv_2
XPHY_251 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_240 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_295 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_262 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_284 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_273 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_81 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[121\] _592_/Y la_buf\[121\]/TE vssd vssd vccd vccd la_data_in_core[121] sky130_fd_sc_hd__einvp_8
Xmprj_adr_buf\[29\] _436_/Y mprj_adr_buf\[29\]/TE vssd vssd vccd vccd mprj_adr_o_user[29]
+ sky130_fd_sc_hd__einvp_8
XFILLER_10_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_672 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__477__A la_data_out_mprj[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[54\] la_data_out_core[54] user_to_mprj_in_gates\[54\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[54\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_760 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_15_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__387__A la_oenb_mprj[119] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[101\]_A user_to_mprj_in_gates\[101\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1691 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[54\]_A user_to_mprj_in_gates\[54\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[101\]_A_N la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_521 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_636_ la_oenb_mprj[37] vssd vssd vccd vccd _636_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_567_ la_data_out_mprj[96] vssd vssd vccd vccd _567_/Y sky130_fd_sc_hd__inv_2
XANTENNA_mprj_adr_buf\[22\]_TE mprj_adr_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[116\]_A_N la_oenb_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[94\]_A _565_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_498_ la_data_out_mprj[27] vssd vssd vccd vccd _498_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[24\] user_to_mprj_in_gates\[24\]/Y vssd vssd vccd vccd la_data_in_mprj[24]
+ sky130_fd_sc_hd__inv_8
XFILLER_8_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_buffers\[45\]_A user_to_mprj_in_gates\[45\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_373 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[85\]_A _556_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[36\]_A user_to_mprj_in_gates\[36\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[64\] la_iena_mprj[64] mprj_logic_high_inst/HI[394] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/B sky130_fd_sc_hd__and2_1
XFILLER_45_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_421_ mprj_adr_o_core[14] vssd vssd vccd vccd _421_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[42\] la_oenb_mprj[42] la_buf_enable\[42\]/B vssd vssd vccd vccd la_buf\[42\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[20\] _619_/Y mprj_logic_high_inst/HI[222] vssd vssd vccd
+ vccd la_oenb_core[20] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[2\] _601_/Y mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd la_oenb_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_41_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_352_ la_oenb_mprj[84] vssd vssd vccd vccd _352_/Y sky130_fd_sc_hd__inv_2
XFILLER_26_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[76\]_A _547_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[28\] _499_/Y la_buf\[28\]/TE vssd vssd vccd vccd la_data_in_core[28] sky130_fd_sc_hd__einvp_8
XANTENNA__580__A la_data_out_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_940 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_995 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[27\]_A user_to_mprj_in_gates\[27\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1022 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1724 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[16\]_TE la_buf\[16\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_619_ la_oenb_mprj[20] vssd vssd vccd vccd _619_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[67\]_A _538_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[17\] la_data_out_core[17] user_to_mprj_in_gates\[17\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[17\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_18_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__490__A la_data_out_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[18\]_A user_to_mprj_in_gates\[18\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1865 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_806 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_817 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_310 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[58\]_A _529_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_828 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_839 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2031 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[76\]_B la_buf_enable\[76\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1038 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[68\] _336_/Y mprj_logic_high_inst/HI[270] vssd vssd vccd
+ vccd la_oenb_core[68] sky130_fd_sc_hd__einvp_8
XFILLER_43_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[16\] _455_/Y mprj_dat_buf\[16\]/TE vssd vssd vccd vccd mprj_dat_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[39\]_TE la_buf\[39\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__575__A la_data_out_mprj[104] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_404_ mprj_sel_o_core[1] vssd vssd vccd vccd _404_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_335_ la_oenb_mprj[67] vssd vssd vccd vccd _335_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[67\]_B la_buf_enable\[67\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_adr_buf\[11\] _418_/Y mprj_adr_buf\[11\]/TE vssd vssd vccd vccd mprj_adr_o_user[11]
+ sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_buffers\[125\] user_to_mprj_in_gates\[125\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[125] sky130_fd_sc_hd__inv_8
XFILLER_46_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1944 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_buffers\[91\] user_to_mprj_in_gates\[91\]/Y vssd vssd vccd vccd la_data_in_mprj[91]
+ sky130_fd_sc_hd__inv_8
XFILLER_2_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__485__A la_data_out_mprj[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[70\]_B mprj_logic_high_inst/HI[400] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[7\]_TE la_buf\[7\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_la_buf_enable\[58\]_B la_buf_enable\[58\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1590 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__395__A la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[27\] la_iena_mprj[27] mprj_logic_high_inst/HI[357] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/B sky130_fd_sc_hd__and2_1
XPHY_603 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_614 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_625 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_636 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_658 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_647 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_669 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[95\] _566_/Y la_buf\[95\]/TE vssd vssd vccd vccd la_data_in_core[95] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[0\] la_iena_mprj[0] mprj_logic_high_inst/HI[330] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[0\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[110\] la_oenb_mprj[110] la_buf_enable\[110\]/B vssd vssd vccd vccd
+ la_buf\[110\]/TE sky130_fd_sc_hd__and2b_1
XANTENNA_la_buf_enable\[74\]_A_N la_oenb_mprj[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[89\]_A_N la_oenb_mprj[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_92 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[12\]_A_N la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1645 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[9\]_A la_iena_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1992 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_oen_buffers\[107\]_A _375_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[27\]_A_N la_oenb_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[84\] la_data_out_core[84] user_to_mprj_in_gates\[84\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[84\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_1785 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1478 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_154 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_400 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_433 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_444 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_411 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_422 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1032 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1021 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1010 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_477 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_466 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_455 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1065 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1054 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1043 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_488 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_499 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1076 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1098 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1087 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[6\] _477_/Y la_buf\[6\]/TE vssd vssd vccd vccd la_data_in_core[6] sky130_fd_sc_hd__einvp_8
XFILLER_7_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[10\] _481_/Y la_buf\[10\]/TE vssd vssd vccd vccd la_data_in_core[10] sky130_fd_sc_hd__einvp_8
XFILLER_4_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xmprj_adr_buf\[3\] _410_/Y mprj_adr_buf\[3\]/TE vssd vssd vccd vccd mprj_adr_o_user[3]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_we_buf_TE mprj_we_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_221 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_adr_buf\[20\]_A _427_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[54\] user_to_mprj_in_gates\[54\]/Y vssd vssd vccd vccd la_data_in_mprj[54]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[11\]_TE mprj_logic_high_inst/HI[213] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[110\] la_data_out_core[110] user_to_mprj_in_gates\[110\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[110\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[94\] la_iena_mprj[94] mprj_logic_high_inst/HI[424] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/B sky130_fd_sc_hd__and2_1
XFILLER_27_2058 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[120\] _388_/Y mprj_logic_high_inst/HI[322] vssd vssd vccd
+ vccd la_oenb_core[120] sky130_fd_sc_hd__einvp_8
XFILLER_46_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_sel_buf\[1\] _404_/Y mprj_sel_buf\[1\]/TE vssd vssd vccd vccd mprj_sel_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_1_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[9\]_A la_data_out_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[50\] _649_/Y mprj_logic_high_inst/HI[252] vssd vssd vccd
+ vccd la_oenb_core[50] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[72\] la_oenb_mprj[72] la_buf_enable\[72\]/B vssd vssd vccd vccd la_buf\[72\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_1_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_652_ la_oenb_mprj[53] vssd vssd vccd vccd _652_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_583_ la_data_out_mprj[112] vssd vssd vccd vccd _583_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[58\] _529_/Y la_buf\[58\]/TE vssd vssd vccd vccd la_data_in_core[58] sky130_fd_sc_hd__einvp_8
XFILLER_32_728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__583__A la_data_out_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_252 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_241 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_230 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_263 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[34\]_TE mprj_logic_high_inst/HI[236] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_285 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_274 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_93 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_296 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[114\] _585_/Y la_buf\[114\]/TE vssd vssd vccd vccd la_data_in_core[114] sky130_fd_sc_hd__einvp_8
XFILLER_4_684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[47\] la_data_out_core[47] user_to_mprj_in_gates\[47\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[47\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_35_599 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__493__A la_data_out_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_772 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[9\]_TE mprj_adr_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1272 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[9\] la_data_out_core[9] user_to_mprj_in_gates\[9\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[9\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_28_1644 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_38_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[72\]_TE la_buf\[72\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[98\] _366_/Y mprj_logic_high_inst/HI[300] vssd vssd vccd
+ vccd la_oenb_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_1_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__578__A la_data_out_mprj[107] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_635_ la_oenb_mprj[36] vssd vssd vccd vccd _635_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_566_ la_data_out_mprj[95] vssd vssd vccd vccd _566_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[21\]_TE mprj_dat_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_497_ la_data_out_mprj[26] vssd vssd vccd vccd _497_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1412 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[17\] user_to_mprj_in_gates\[17\]/Y vssd vssd vccd vccd la_data_in_mprj[17]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__488__A la_data_out_mprj[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_341 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__398__A caravel_clk vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[57\] la_iena_mprj[57] mprj_logic_high_inst/HI[387] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_18_319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_420_ mprj_adr_o_core[13] vssd vssd vccd vccd _420_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[13\] _612_/Y mprj_logic_high_inst/HI[215] vssd vssd vccd
+ vccd la_oenb_core[13] sky130_fd_sc_hd__einvp_8
X_351_ la_oenb_mprj[83] vssd vssd vccd vccd _351_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[35\] la_oenb_mprj[35] la_buf_enable\[35\]/B vssd vssd vccd vccd la_buf\[35\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[9\] user_to_mprj_in_gates\[9\]/Y vssd vssd vccd vccd la_data_in_mprj[9]
+ sky130_fd_sc_hd__inv_8
XFILLER_22_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_1736 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_618_ la_oenb_mprj[19] vssd vssd vccd vccd _618_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_549_ la_data_out_mprj[78] vssd vssd vccd vccd _549_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1877 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_807 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_818 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_829 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[100\]_A_N la_oenb_mprj[100] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[12\]_TE mprj_adr_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[115\]_A_N la_oenb_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_403_ mprj_sel_o_core[0] vssd vssd vccd vccd _403_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_61 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_14_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[40\] _511_/Y la_buf\[40\]/TE vssd vssd vccd vccd la_data_in_core[40] sky130_fd_sc_hd__einvp_8
X_334_ la_oenb_mprj[66] vssd vssd vccd vccd _334_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__591__A la_data_out_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[112\] la_iena_mprj[112] mprj_logic_high_inst/HI[442] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[112\]/B sky130_fd_sc_hd__and2_1
XFILLER_31_1139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[118\] user_to_mprj_in_gates\[118\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[118] sky130_fd_sc_hd__inv_8
XFILLER_26_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_irq_gates\[2\]_A user_irq_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1967 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[84\] user_to_mprj_in_gates\[84\]/Y vssd vssd vccd vccd la_data_in_mprj[84]
+ sky130_fd_sc_hd__inv_8
XFILLER_26_1989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_TE mprj_dat_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_119 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_46_38 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[9\]_A _416_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_604 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_615 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_626 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_637 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_659 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_648 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_30_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[80\] _348_/Y mprj_logic_high_inst/HI[282] vssd vssd vccd
+ vccd la_oenb_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_10_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[50\]_A la_data_out_core[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__586__A la_data_out_mprj[115] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[88\] _559_/Y la_buf\[88\]/TE vssd vssd vccd vccd la_data_in_core[88] sky130_fd_sc_hd__einvp_8
XFILLER_19_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[103\] la_oenb_mprj[103] la_buf_enable\[103\]/B vssd vssd vccd vccd
+ la_buf\[103\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_37_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[41\]_A la_data_out_core[41] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xuser_to_mprj_in_gates\[77\] la_data_out_core[77] user_to_mprj_in_gates\[77\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[77\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__496__A la_data_out_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[90\]_TE mprj_logic_high_inst/HI[292] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_199 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[32\]_A la_data_out_core[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[99\]_A la_data_out_core[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_401 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1635 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_434 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_412 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_423 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_40_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1000 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1022 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1011 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_467 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_445 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_456 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1033 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1055 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1044 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_478 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_489 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1077 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1099 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1066 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1088 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_800 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_84 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[23\]_A la_data_out_core[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1708 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[47\] user_to_mprj_in_gates\[47\]/Y vssd vssd vccd vccd la_data_in_mprj[47]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_990 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1307 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[14\]_A la_data_out_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_26_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1688 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[103\] la_data_out_core[103] user_to_mprj_in_gates\[103\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[103\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_43_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[73\]_A_N la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[87\] la_iena_mprj[87] mprj_logic_high_inst/HI[417] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf_enable\[88\]_A_N la_oenb_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_clk2_buf _399_/Y mprj_clk2_buf/TE vssd vssd vccd vccd user_clock2 sky130_fd_sc_hd__einvp_8
XFILLER_1_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[113\] _381_/Y mprj_logic_high_inst/HI[315] vssd vssd vccd
+ vccd la_oenb_core[113] sky130_fd_sc_hd__einvp_8
XFILLER_44_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[9\]_B user_to_mprj_in_gates\[9\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_A_N la_oenb_mprj[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_651_ la_oenb_mprj[52] vssd vssd vccd vccd _651_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[43\] _642_/Y mprj_logic_high_inst/HI[245] vssd vssd vccd
+ vccd la_oenb_core[43] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[65\] la_oenb_mprj[65] la_buf_enable\[65\]/B vssd vssd vccd vccd la_buf\[65\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_irq_buffers\[1\] user_irq_gates\[1\]/Y vssd vssd vccd vccd user_irq[1] sky130_fd_sc_hd__inv_8
XFILLER_40_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_582_ la_data_out_mprj[111] vssd vssd vccd vccd _582_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_247 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[26\]_A_N la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_220 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_242 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_231 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_253 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_286 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_275 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_264 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_965 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_297 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_497 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[107\] _578_/Y la_buf\[107\]/TE vssd vssd vccd vccd la_data_in_core[107] sky130_fd_sc_hd__einvp_8
XFILLER_4_696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[100\] user_to_mprj_in_gates\[100\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[100] sky130_fd_sc_hd__inv_8
XFILLER_27_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_A la_iena_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1852 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[102\]_TE mprj_logic_high_inst/HI[304] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[111\]_A la_iena_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_707 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2041 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_634_ la_oenb_mprj[35] vssd vssd vccd vccd _634_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__594__A la_data_out_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[70\] _541_/Y la_buf\[70\]/TE vssd vssd vccd vccd la_data_in_core[70] sky130_fd_sc_hd__einvp_8
X_565_ la_data_out_mprj[94] vssd vssd vccd vccd _565_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_496_ la_data_out_mprj[25] vssd vssd vccd vccd _496_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_ena_buf\[102\]_A la_iena_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_733 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1468 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[125\]_TE mprj_logic_high_inst/HI[327] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_397 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[24\]_TE mprj_logic_high_inst/HI[226] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[91\]_A la_iena_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_350_ la_oenb_mprj[82] vssd vssd vccd vccd _350_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[28\] la_oenb_mprj[28] la_buf_enable\[28\]/B vssd vssd vccd vccd la_buf\[28\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__589__A la_data_out_mprj[118] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[82\]_A la_iena_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_617_ la_oenb_mprj[18] vssd vssd vccd vccd _617_/Y sky130_fd_sc_hd__inv_2
X_548_ la_data_out_mprj[77] vssd vssd vccd vccd _548_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_479_ la_data_out_mprj[8] vssd vssd vccd vccd _479_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1688 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[62\]_TE la_buf\[62\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[47\]_TE mprj_logic_high_inst/HI[249] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__499__A la_data_out_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1889 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[73\]_A la_iena_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_808 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_819 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[9\]_B la_buf_enable\[9\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_2055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[11\]_TE mprj_dat_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[64\]_A la_iena_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_402_ mprj_we_o_core vssd vssd vccd vccd _402_/Y sky130_fd_sc_hd__inv_2
XPHY_40 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_73 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_333_ la_oenb_mprj[65] vssd vssd vccd vccd _333_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[85\]_TE la_buf\[85\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[33\] _504_/Y la_buf\[33\]/TE vssd vssd vccd vccd la_data_in_core[33] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[105\] la_iena_mprj[105] mprj_logic_high_inst/HI[435] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[105\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_1979 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[77\] user_to_mprj_in_gates\[77\]/Y vssd vssd vccd vccd la_data_in_mprj[77]
+ sky130_fd_sc_hd__inv_8
XFILLER_2_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[55\]_A la_iena_mprj[55] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[22\] la_data_out_core[22] user_to_mprj_in_gates\[22\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[22\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_20_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1641 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_9_371 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[3\]_A _406_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[46\]_A la_iena_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_605 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_616 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_638 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_838 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_649 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_627 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1140 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[73\] _341_/Y mprj_logic_high_inst/HI[275] vssd vssd vccd
+ vccd la_oenb_core[73] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[95\] la_oenb_mprj[95] la_buf_enable\[95\]/B vssd vssd vccd vccd la_buf\[95\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[21\] _460_/Y mprj_dat_buf\[21\]/TE vssd vssd vccd vccd mprj_dat_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[37\]_A la_iena_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_6_352 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[28\]_A la_iena_mprj[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[114\]_A_N la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[1\] la_oenb_mprj[1] la_buf_enable\[1\]/B vssd vssd vccd vccd la_buf\[1\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_buffers\[93\]_A user_to_mprj_in_gates\[93\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[19\]_A la_iena_mprj[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_278 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[32\] la_iena_mprj[32] mprj_logic_high_inst/HI[362] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/B sky130_fd_sc_hd__and2_1
XFILLER_37_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_435 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_424 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_402 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_413 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1001 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1023 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1012 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_468 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_446 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_457 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1034 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1056 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1045 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_479 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1078 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1067 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1089 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[10\] la_oenb_mprj[10] la_buf_enable\[10\]/B vssd vssd vccd vccd la_buf\[10\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_8_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[120\]_A _591_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_812 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__597__A la_data_out_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[25\]_TE mprj_adr_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_980 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_432 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_991 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[111\]_A _582_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1816 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[102\]_A _573_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[66\]_A user_to_mprj_in_gates\[66\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_347 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_358 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[106\] _374_/Y mprj_logic_high_inst/HI[308] vssd vssd vccd
+ vccd la_oenb_core[106] sky130_fd_sc_hd__einvp_8
XFILLER_44_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_650_ la_oenb_mprj[51] vssd vssd vccd vccd _650_/Y sky130_fd_sc_hd__inv_2
X_581_ la_data_out_mprj[110] vssd vssd vccd vccd _581_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[36\] _635_/Y mprj_logic_high_inst/HI[238] vssd vssd vccd
+ vccd la_oenb_core[36] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[58\] la_oenb_mprj[58] la_buf_enable\[58\]/B vssd vssd vccd vccd la_buf\[58\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_210 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_259 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_900 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_221 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_243 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_232 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_254 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_276 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_265 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_977 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_287 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_298 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_1054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[104\]_A user_to_mprj_in_gates\[104\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1639 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[57\]_A user_to_mprj_in_gates\[57\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[80\]_TE mprj_logic_high_inst/HI[282] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[19\]_TE la_buf\[19\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[97\]_A _568_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[120\]_B mprj_logic_high_inst/HI[450] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_796 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[48\]_A user_to_mprj_in_gates\[48\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[21\]_A _492_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[111\]_B mprj_logic_high_inst/HI[441] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[30\]_B la_buf_enable\[30\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_633_ la_oenb_mprj[34] vssd vssd vccd vccd _633_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_564_ la_data_out_mprj[93] vssd vssd vccd vccd _564_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[63\] _534_/Y la_buf\[63\]/TE vssd vssd vccd vccd la_data_in_core[63] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_ena_buf\[102\]_B mprj_logic_high_inst/HI[432] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_495_ la_data_out_mprj[24] vssd vssd vccd vccd _495_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_778 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_756 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[27\] _434_/Y mprj_adr_buf\[27\]/TE vssd vssd vccd vccd mprj_adr_o_user[27]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_461 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[21\]_B la_buf_enable\[21\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[52\] la_data_out_core[52] user_to_mprj_in_gates\[52\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[52\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1637 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[72\]_A_N la_oenb_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_321 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[87\]_A_N la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_23_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[88\]_B la_buf_enable\[88\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[10\]_A_N la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[25\]_A_N la_oenb_mprj[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[12\]_B la_buf_enable\[12\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[79\]_B la_buf_enable\[79\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1193 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[126\] la_oenb_mprj[126] la_buf_enable\[126\]/B vssd vssd vccd vccd
+ la_buf\[126\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_39_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_616_ la_oenb_mprj[17] vssd vssd vccd vccd _616_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_547_ la_data_out_mprj[76] vssd vssd vccd vccd _547_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_313 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_376 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_346 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_357 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_478_ la_data_out_mprj[7] vssd vssd vccd vccd _478_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[22\] user_to_mprj_in_gates\[22\]/Y vssd vssd vccd vccd la_data_in_mprj[22]
+ sky130_fd_sc_hd__inv_8
XFILLER_12_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1570 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[73\]_B mprj_logic_high_inst/HI[403] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_35_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_809 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2089 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1344 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[62\] la_iena_mprj[62] mprj_logic_high_inst/HI[392] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_401_ mprj_stb_o_core vssd vssd vccd vccd _401_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[0\] _599_/Y mprj_logic_high_inst/HI[202] vssd vssd vccd
+ vccd la_oenb_core[0] sky130_fd_sc_hd__einvp_8
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[40\] la_oenb_mprj[40] la_buf_enable\[40\]/B vssd vssd vccd vccd la_buf\[40\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_26_173 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_63 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_52 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_85 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_332_ la_oenb_mprj[64] vssd vssd vccd vccd _332_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[115\]_TE mprj_logic_high_inst/HI[317] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf\[26\] _497_/Y la_buf\[26\]/TE vssd vssd vccd vccd la_data_in_core[26] sky130_fd_sc_hd__einvp_8
XFILLER_6_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_1_250 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[55\]_B mprj_logic_high_inst/HI[385] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[15\] la_data_out_core[15] user_to_mprj_in_gates\[15\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[15\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_14_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[14\]_TE mprj_logic_high_inst/HI[216] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_383 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[126\] la_data_out_core[126] user_to_mprj_in_gates\[126\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[126\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_44_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1253 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_606 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_617 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_639 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_628 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1428 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1152 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_504 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[66\] _334_/Y mprj_logic_high_inst/HI[268] vssd vssd vccd
+ vccd la_oenb_core[66] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[88\] la_oenb_mprj[88] la_buf_enable\[88\]/B vssd vssd vccd vccd la_buf\[88\]/TE
+ sky130_fd_sc_hd__and2b_1
Xmprj_dat_buf\[14\] _453_/Y mprj_dat_buf\[14\]/TE vssd vssd vccd vccd mprj_dat_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_46_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_27_493 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_42_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_636 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1940 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_331 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_887 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1383 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1700 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_buffers\[123\] user_to_mprj_in_gates\[123\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[123] sky130_fd_sc_hd__inv_8
XFILLER_46_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[23\]_A _430_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2116 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_997 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[75\]_TE la_buf\[75\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[14\]_A _421_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[25\] la_iena_mprj[25] mprj_logic_high_inst/HI[355] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[25\]/B sky130_fd_sc_hd__and2_1
XFILLER_38_1659 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_425 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_403 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_414 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1002 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1013 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_436 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_447 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_458 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1035 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1024 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1046 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_469 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1068 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1057 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1079 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_139 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_824 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[93\] _564_/Y la_buf\[93\]/TE vssd vssd vccd vccd la_data_in_core[93] sky130_fd_sc_hd__einvp_8
XFILLER_21_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[24\]_TE mprj_dat_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_238 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_981 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_970 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[3\]_TE mprj_logic_high_inst/HI[205] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_992 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_11_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1243 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[82\] la_data_out_core[82] user_to_mprj_in_gates\[82\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[82\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_580_ la_data_out_mprj[109] vssd vssd vccd vccd _580_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[29\] _628_/Y mprj_logic_high_inst/HI[231] vssd vssd vccd
+ vccd la_oenb_core[29] sky130_fd_sc_hd__einvp_8
XPHY_200 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_222 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_211 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_233 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_912 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_255 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_244 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_277 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_266 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_288 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_299 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[4\] _475_/Y la_buf\[4\]/TE vssd vssd vccd vccd la_data_in_core[4] sky130_fd_sc_hd__einvp_8
XFILLER_4_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1364 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__401__A mprj_stb_o_core vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[113\]_A_N la_oenb_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xmprj_adr_buf\[1\] _408_/Y mprj_adr_buf\[1\]/TE vssd vssd vccd vccd mprj_adr_o_user[1]
+ sky130_fd_sc_hd__einvp_8
XFILLER_23_1725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_871 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[52\] user_to_mprj_in_gates\[52\]/Y vssd vssd vccd vccd la_data_in_mprj[52]
+ sky130_fd_sc_hd__inv_8
XFILLER_1_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_720 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_1231 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_11_1139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_28_1647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_6_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1342 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_mprj_adr_buf\[15\]_TE mprj_adr_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[92\] la_iena_mprj[92] mprj_logic_high_inst/HI[422] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[92\]/B sky130_fd_sc_hd__and2_1
XFILLER_0_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1207 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[70\] la_oenb_mprj[70] la_buf_enable\[70\]/B vssd vssd vccd vccd la_buf\[70\]/TE
+ sky130_fd_sc_hd__and2b_1
X_632_ la_oenb_mprj[33] vssd vssd vccd vccd _632_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_563_ la_data_out_mprj[92] vssd vssd vccd vccd _563_/Y sky130_fd_sc_hd__inv_2
X_494_ la_data_out_mprj[23] vssd vssd vccd vccd _494_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[56\] _527_/Y la_buf\[56\]/TE vssd vssd vccd vccd la_data_in_core[56] sky130_fd_sc_hd__einvp_8
XFILLER_38_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_591 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_713 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_245 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[112\] _583_/Y la_buf\[112\]/TE vssd vssd vccd vccd la_data_in_core[112] sky130_fd_sc_hd__einvp_8
XFILLER_5_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_473 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_1183 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_25_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_TE mprj_dat_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1627 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[45\] la_data_out_core[45] user_to_mprj_in_gates\[45\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[45\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_39_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[7\] la_data_out_core[7] user_to_mprj_in_gates\[7\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[7\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_24_2009 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_333 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[70\]_TE mprj_logic_high_inst/HI[272] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[96\] _364_/Y mprj_logic_high_inst/HI[298] vssd vssd vccd
+ vccd la_oenb_core[96] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_gates\[80\]_A la_data_out_core[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[9\] la_iena_mprj[9] mprj_logic_high_inst/HI[339] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[9\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xla_buf_enable\[119\] la_oenb_mprj[119] la_buf_enable\[119\]/B vssd vssd vccd vccd
+ la_buf\[119\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_344 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_615_ la_oenb_mprj[16] vssd vssd vccd vccd _615_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_546_ la_data_out_mprj[75] vssd vssd vccd vccd _546_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_477_ la_data_out_mprj[6] vssd vssd vccd vccd _477_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[15\] user_to_mprj_in_gates\[15\]/Y vssd vssd vccd vccd la_data_in_mprj[15]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_gates\[71\]_A la_data_out_core[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[93\]_TE mprj_logic_high_inst/HI[295] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_2002 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1009 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[62\]_A la_data_out_core[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj2_pwrgood mprj2_pwrgood/A vssd vssd vccd vccd user2_vcc_powergood sky130_fd_sc_hd__buf_8
XFILLER_8_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[55\] la_iena_mprj[55] mprj_logic_high_inst/HI[385] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[55\]/B sky130_fd_sc_hd__and2_1
XFILLER_42_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_400_ mprj_cyc_o_core vssd vssd vccd vccd _400_/Y sky130_fd_sc_hd__inv_2
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_152 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_64 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_331_ la_oenb_mprj[63] vssd vssd vccd vccd _331_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[11\] _610_/Y mprj_logic_high_inst/HI[213] vssd vssd vccd
+ vccd la_oenb_core[11] sky130_fd_sc_hd__einvp_8
XPHY_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_185 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_97 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[33\] la_oenb_mprj[33] la_buf_enable\[33\]/B vssd vssd vccd vccd la_buf\[33\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_in_buffers\[7\] user_to_mprj_in_gates\[7\]/Y vssd vssd vccd vccd la_data_in_mprj[7]
+ sky130_fd_sc_hd__inv_8
XFILLER_35_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[71\]_A_N la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1554 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[53\]_A la_data_out_core[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[19\] _490_/Y la_buf\[19\]/TE vssd vssd vccd vccd la_data_in_core[19] sky130_fd_sc_hd__einvp_8
XFILLER_6_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[86\]_A_N la_oenb_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_929 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_24_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_620 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[24\]_A_N la_oenb_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_529_ la_data_out_mprj[58] vssd vssd vccd vccd _529_/Y sky130_fd_sc_hd__inv_2
XFILLER_32_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1318 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_395 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[39\]_A_N la_oenb_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[44\]_A la_data_out_core[44] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1149 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_29_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1508 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_gates\[119\] la_data_out_core[119] user_to_mprj_in_gates\[119\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[119\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_607 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_618 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_629 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_133 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_gates\[35\]_A la_data_out_core[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1186 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1121 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[59\] _658_/Y mprj_logic_high_inst/HI[261] vssd vssd vccd
+ vccd la_oenb_core[59] sky130_fd_sc_hd__einvp_8
XFILLER_46_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_409 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[110\] la_iena_mprj[110] mprj_logic_high_inst/HI[440] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[110\]/B sky130_fd_sc_hd__and2_1
XPHY_1740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_851 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_1751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[26\]_A la_data_out_core[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[110\]_A la_data_out_core[110] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_7_899 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__404__A mprj_sel_o_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[116\] user_to_mprj_in_gates\[116\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[116] sky130_fd_sc_hd__inv_8
XFILLER_46_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[82\] user_to_mprj_in_gates\[82\]/Y vssd vssd vccd vccd la_data_in_mprj[82]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[17\]_A la_data_out_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_gates\[101\]_A la_data_out_core[101] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_31_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2070 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_2092 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1485 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_28_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_426 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_404 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_415 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1003 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1014 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[18\] la_iena_mprj[18] mprj_logic_high_inst/HI[348] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[18\]/B sky130_fd_sc_hd__and2_1
XPHY_437 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_448 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_459 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1036 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1025 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1047 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1069 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1058 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_14_1682 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[86\] _557_/Y la_buf\[86\]/TE vssd vssd vccd vccd la_data_in_core[86] sky130_fd_sc_hd__einvp_8
XFILLER_5_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[101\] la_oenb_mprj[101] la_buf_enable\[101\]/B vssd vssd vccd vccd
+ la_buf\[101\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_21_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_971 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_960 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_993 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_982 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_478 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1818 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[75\] la_data_out_core[75] user_to_mprj_in_gates\[75\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[75\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_ena_buf\[123\]_A la_iena_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1224 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1292 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[27\]_TE mprj_logic_high_inst/HI[229] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_512 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_515 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_A la_iena_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_201 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_223 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_212 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_234 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_924 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_256 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_245 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_267 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_445 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1012 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_53 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_289 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_405 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_278 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_ena_buf\[1\] user_irq_ena[1] user_irq_ena_buf\[1\]/B vssd vssd vccd vccd
+ user_irq_gates\[1\]/B sky130_fd_sc_hd__and2_1
XFILLER_10_1376 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_883 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_A la_iena_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[45\] user_to_mprj_in_gates\[45\]/Y vssd vssd vccd vccd la_data_in_mprj[45]
+ sky130_fd_sc_hd__inv_8
XFILLER_15_272 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_790 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[65\]_TE la_buf\[65\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1709 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[101\] la_data_out_core[101] user_to_mprj_in_gates\[101\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[101\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_26_526 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_26_537 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1354 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[14\]_TE mprj_dat_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[85\] la_iena_mprj[85] mprj_logic_high_inst/HI[415] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[85\]/B sky130_fd_sc_hd__and2_1
XANTENNA__502__A la_data_out_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[111\] _379_/Y mprj_logic_high_inst/HI[313] vssd vssd vccd
+ vccd la_oenb_core[111] sky130_fd_sc_hd__einvp_8
XFILLER_40_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[94\]_A la_iena_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_631_ la_oenb_mprj[32] vssd vssd vccd vccd _631_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[41\] _640_/Y mprj_logic_high_inst/HI[243] vssd vssd vccd
+ vccd la_oenb_core[41] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[63\] la_oenb_mprj[63] la_buf_enable\[63\]/B vssd vssd vccd vccd la_buf\[63\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_45_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_22_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_562_ la_data_out_mprj[91] vssd vssd vccd vccd _562_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_493_ la_data_out_mprj[22] vssd vssd vccd vccd _493_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[88\]_TE la_buf\[88\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_725 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf\[49\] _520_/Y la_buf\[49\]/TE vssd vssd vccd vccd la_data_in_core[49] sky130_fd_sc_hd__einvp_8
XFILLER_12_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_257 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__412__A mprj_adr_o_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[105\] _576_/Y la_buf\[105\]/TE vssd vssd vccd vccd la_data_in_core[105] sky130_fd_sc_hd__einvp_8
XFILLER_39_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[85\]_A la_iena_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[38\] la_data_out_core[38] user_to_mprj_in_gates\[38\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[38\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1549 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_A la_iena_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1263 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[112\]_A_N la_oenb_mprj[112] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[127\]_A_N la_oenb_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[89\] _357_/Y mprj_logic_high_inst/HI[291] vssd vssd vccd
+ vccd la_oenb_core[89] sky130_fd_sc_hd__einvp_8
XFILLER_2_934 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_411 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_455 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[67\]_A la_iena_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_614_ la_oenb_mprj[15] vssd vssd vccd vccd _614_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_545_ la_data_out_mprj[74] vssd vssd vccd vccd _545_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_315 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_18_1614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_476_ la_data_out_mprj[5] vssd vssd vccd vccd _476_/Y sky130_fd_sc_hd__inv_2
XANTENNA__407__A mprj_adr_o_core[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[58\]_A la_iena_mprj[58] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_654 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1182 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_2014 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_392 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_30_1324 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1780 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_1314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[49\]_A la_iena_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[48\] la_iena_mprj[48] mprj_logic_high_inst/HI[378] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[48\]/B sky130_fd_sc_hd__and2_1
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_65 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_330_ la_oenb_mprj[62] vssd vssd vccd vccd _330_/Y sky130_fd_sc_hd__inv_2
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_197 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_76 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_35_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[26\] la_oenb_mprj[26] la_buf_enable\[26\]/B vssd vssd vccd vccd la_buf\[26\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_35_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[28\]_TE mprj_adr_buf\[28\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1881 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[7\]_A _446_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_528_ la_data_out_mprj[57] vssd vssd vccd vccd _528_/Y sky130_fd_sc_hd__inv_2
X_459_ mprj_dat_o_core[20] vssd vssd vccd vccd _459_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1584 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__600__A la_oenb_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[60\]_TE mprj_logic_high_inst/HI[262] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_608 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_619 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_145 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_1132 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__510__A la_data_out_mprj[39] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_42 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[20\]_A user_to_mprj_in_gates\[20\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_75 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_ena_buf\[103\] la_iena_mprj[103] mprj_logic_high_inst/HI[433] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[103\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf\[123\]_A _594_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[31\] _502_/Y la_buf\[31\]/TE vssd vssd vccd vccd la_data_in_core[31] sky130_fd_sc_hd__einvp_8
XPHY_1774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_buffers\[87\]_A user_to_mprj_in_gates\[87\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_1796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_856 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[60\]_A _531_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[83\]_TE mprj_logic_high_inst/HI[285] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__420__A mprj_adr_o_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[109\] user_to_mprj_in_gates\[109\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[109] sky130_fd_sc_hd__inv_8
XFILLER_42_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[75\] user_to_mprj_in_gates\[75\]/Y vssd vssd vccd vccd la_data_in_mprj[75]
+ sky130_fd_sc_hd__inv_8
XFILLER_46_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_buffers\[11\]_A user_to_mprj_in_gates\[11\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_34_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[20\] la_data_out_core[20] user_to_mprj_in_gates\[20\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[20\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_la_buf\[114\]_A _585_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_dat_buf\[8\] _447_/Y mprj_dat_buf\[8\]/TE vssd vssd vccd vccd mprj_dat_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XANTENNA__330__A la_oenb_mprj[62] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[70\]_A_N la_oenb_mprj[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_405 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_416 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1004 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_427 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_438 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_449 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[85\]_A_N la_oenb_mprj[85] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[116\]_A user_to_mprj_in_gates\[116\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_2086 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1037 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1026 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1015 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1385 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1059 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[105\]_A _576_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1048 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__505__A la_data_out_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_22_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_1547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[23\]_A_N la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[93\] la_oenb_mprj[93] la_buf_enable\[93\]/B vssd vssd vccd vccd la_buf\[93\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[71\] _339_/Y mprj_logic_high_inst/HI[273] vssd vssd vccd
+ vccd la_oenb_core[71] sky130_fd_sc_hd__einvp_8
XFILLER_43_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[38\]_A_N la_oenb_mprj[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_74 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[79\] _550_/Y la_buf\[79\]/TE vssd vssd vccd vccd la_data_in_core[79] sky130_fd_sc_hd__einvp_8
XFILLER_21_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_421 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_972 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_961 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_950 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_buffers\[107\]_A user_to_mprj_in_gates\[107\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1403 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_1561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_994 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_983 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__415__A mprj_adr_o_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[51\]_B la_buf_enable\[51\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[68\] la_data_out_core[68] user_to_mprj_in_gates\[68\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[68\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_4_2062 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[123\]_B mprj_logic_high_inst/HI[453] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[42\]_B la_buf_enable\[42\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1261 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1169 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_527 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[114\]_B mprj_logic_high_inst/HI[444] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[30\] la_iena_mprj[30] mprj_logic_high_inst/HI[360] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[30\]/B sky130_fd_sc_hd__and2_1
XFILLER_17_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_224 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_213 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_202 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_257 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_246 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_235 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_268 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_947 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_273 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_279 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1024 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1491 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_1355 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[33\]_B la_buf_enable\[33\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1841 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[2\]_A la_iena_mprj[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_895 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[105\]_B mprj_logic_high_inst/HI[435] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_43_571 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[38\] user_to_mprj_in_gates\[38\]/Y vssd vssd vccd vccd la_data_in_mprj[38]
+ sky130_fd_sc_hd__inv_8
XPHY_780 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_1244 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_791 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[24\]_B la_buf_enable\[24\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1366 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_21_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[15\]_B la_buf_enable\[15\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[78\] la_iena_mprj[78] mprj_logic_high_inst/HI[408] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[78\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_158 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1091 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[104\] _372_/Y mprj_logic_high_inst/HI[306] vssd vssd vccd
+ vccd la_oenb_core[104] sky130_fd_sc_hd__einvp_8
XFILLER_29_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_630_ la_oenb_mprj[31] vssd vssd vccd vccd _630_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_561_ la_data_out_mprj[90] vssd vssd vccd vccd _561_/Y sky130_fd_sc_hd__inv_2
XFILLER_28_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[34\] _633_/Y mprj_logic_high_inst/HI[236] vssd vssd vccd
+ vccd la_oenb_core[34] sky130_fd_sc_hd__einvp_8
XFILLER_2_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[56\] la_oenb_mprj[56] la_buf_enable\[56\]/B vssd vssd vccd vccd la_buf\[56\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_29_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_492_ la_data_out_mprj[21] vssd vssd vccd vccd _492_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_722 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[118\]_TE mprj_logic_high_inst/HI[320] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1406 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_29_1903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1958 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_1524 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[85\]_B mprj_logic_high_inst/HI[415] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_23_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1364 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_2098 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_2103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__603__A la_oenb_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1529 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[76\]_B mprj_logic_high_inst/HI[406] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_39_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[2\]_A la_data_out_core[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[0\]_TE la_buf\[0\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__513__A la_data_out_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_423 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[67\]_B mprj_logic_high_inst/HI[397] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_613_ la_oenb_mprj[14] vssd vssd vccd vccd _613_/Y sky130_fd_sc_hd__inv_2
XFILLER_29_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[55\]_TE la_buf\[55\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_305 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[61\] _532_/Y la_buf\[61\]/TE vssd vssd vccd vccd la_data_in_core[61] sky130_fd_sc_hd__einvp_8
XFILLER_22_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_357 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_368 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_544_ la_data_out_mprj[73] vssd vssd vccd vccd _544_/Y sky130_fd_sc_hd__inv_2
X_475_ la_data_out_mprj[4] vssd vssd vccd vccd _475_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_574 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1214 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__423__A mprj_adr_o_core[16] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xmprj_adr_buf\[25\] _432_/Y mprj_adr_buf\[25\]/TE vssd vssd vccd vccd mprj_adr_o_user[25]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_283 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[50\] la_data_out_core[50] user_to_mprj_in_gates\[50\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[50\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_3_1459 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_2026 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__333__A la_oenb_mprj[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_102 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_55 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__508__A la_data_out_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_77 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[19\] la_oenb_mprj[19] la_buf_enable\[19\]/B vssd vssd vccd vccd la_buf\[19\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_10_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_13_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_irq_gates\[2\] user_irq_core[2] user_irq_gates\[2\]/B vssd vssd vccd vccd user_irq_gates\[2\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_46_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_798 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_2_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[124\] la_oenb_mprj[124] la_buf_enable\[124\]/B vssd vssd vccd vccd
+ la_buf\[124\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_18_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[27\]_TE mprj_dat_buf\[27\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_154 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_614 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_527_ la_data_out_mprj[56] vssd vssd vccd vccd _527_/Y sky130_fd_sc_hd__inv_2
XANTENNA__418__A mprj_adr_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_458_ mprj_dat_o_core[19] vssd vssd vccd vccd _458_/Y sky130_fd_sc_hd__inv_2
X_389_ la_oenb_mprj[121] vssd vssd vccd vccd _389_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_371 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_13_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[20\] user_to_mprj_in_gates\[20\]/Y vssd vssd vccd vccd la_data_in_mprj[20]
+ sky130_fd_sc_hd__inv_8
XFILLER_31_1656 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[98\] la_data_out_core[98] user_to_mprj_in_gates\[98\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[98\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_25_2128 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1613 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[111\]_A_N la_oenb_mprj[111] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_la_buf_enable\[126\]_A_N la_oenb_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_609 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[60\] la_iena_mprj[60] mprj_logic_high_inst/HI[390] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[60\]/B sky130_fd_sc_hd__and2_1
XANTENNA_mprj_sel_buf\[1\]_TE mprj_sel_buf\[1\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1972 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_463 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_42_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_606 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_19_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1776 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[24\] _495_/Y la_buf\[24\]/TE vssd vssd vccd vccd la_data_in_core[24] sky130_fd_sc_hd__einvp_8
XPHY_1797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_540 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_551 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[68\] user_to_mprj_in_gates\[68\]/Y vssd vssd vccd vccd la_data_in_mprj[68]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_989 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[13\] la_data_out_core[13] user_to_mprj_in_gates\[13\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[13\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__611__A la_oenb_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[124\] la_data_out_core[124] user_to_mprj_in_gates\[124\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[124\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_42_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_406 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_417 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1005 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_428 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_439 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1038 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1027 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1016 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1049 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[18\]_TE mprj_adr_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_mprj_adr_buf\[2\]_TE mprj_adr_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__521__A la_data_out_mprj[50] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[86\] la_oenb_mprj[86] la_buf_enable\[86\]/B vssd vssd vccd vccd la_buf\[86\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[64\] _332_/Y mprj_logic_high_inst/HI[266] vssd vssd vccd
+ vccd la_oenb_core[64] sky130_fd_sc_hd__einvp_8
XFILLER_47_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[12\] _451_/Y mprj_dat_buf\[12\]/TE vssd vssd vccd vccd mprj_dat_o_user[12]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_cyc_buf_A _400_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_227 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_86 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1699 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_962 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_951 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_940 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1573 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_995 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_984 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_973 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_oen_buffers\[50\]_TE mprj_logic_high_inst/HI[252] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1595 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__431__A mprj_adr_o_core[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[121\] user_to_mprj_in_gates\[121\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[121] sky130_fd_sc_hd__inv_8
XANTENNA_mprj_dat_buf\[6\]_TE mprj_dat_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2074 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_34_720 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__606__A la_oenb_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__341__A la_oenb_mprj[73] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1159 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_37_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_225 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_214 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_203 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[23\] la_iena_mprj[23] mprj_logic_high_inst/HI[353] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[23\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_258 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_236 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_247 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_908 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__516__A la_data_out_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_24_285 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_269 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_1036 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1312 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[2\]_B mprj_logic_high_inst/HI[332] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_47_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[91\] _562_/Y la_buf\[91\]/TE vssd vssd vccd vccd la_data_in_core[91] sky130_fd_sc_hd__einvp_8
XFILLER_47_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_222 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_200 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__426__A mprj_adr_o_core[19] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_770 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_781 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_792 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_299 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_1289 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[80\] la_data_out_core[80] user_to_mprj_in_gates\[80\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[80\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_1098 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[84\]_A_N la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[96\]_TE mprj_logic_high_inst/HI[298] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[99\]_A_N la_oenb_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[22\]_A_N la_oenb_mprj[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__336__A la_oenb_mprj[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_233 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[92\]_A la_data_out_core[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[37\]_A_N la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_1327 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_560_ la_data_out_mprj[89] vssd vssd vccd vccd _560_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_517 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_491_ la_data_out_mprj[20] vssd vssd vccd vccd _491_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[27\] _626_/Y mprj_logic_high_inst/HI[229] vssd vssd vccd
+ vccd la_oenb_core[27] sky130_fd_sc_hd__einvp_8
XFILLER_13_701 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[49\] la_oenb_mprj[49] la_buf_enable\[49\]/B vssd vssd vccd vccd la_buf\[49\]/TE
+ sky130_fd_sc_hd__and2b_1
Xuser_to_mprj_oen_buffers\[9\] _608_/Y mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd la_oenb_core[9] sky130_fd_sc_hd__einvp_8
XFILLER_44_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_734 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_gates\[83\]_A la_data_out_core[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[2\] _473_/Y la_buf\[2\]/TE vssd vssd vccd vccd la_data_in_core[2] sky130_fd_sc_hd__einvp_8
XFILLER_5_911 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1766 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_2066 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[50\] user_to_mprj_in_gates\[50\]/Y vssd vssd vccd vccd la_data_in_mprj[50]
+ sky130_fd_sc_hd__inv_8
XFILLER_16_561 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1507 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[74\]_A la_data_out_core[74] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1086 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_28_2115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[2\]_B user_to_mprj_in_gates\[2\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_41_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_39_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1153 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[65\]_A la_data_out_core[65] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_748 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1727 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[90\] la_iena_mprj[90] mprj_logic_high_inst/HI[420] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[90\]/B sky130_fd_sc_hd__and2_1
XFILLER_5_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_435 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1282 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_612_ la_oenb_mprj[13] vssd vssd vccd vccd _612_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_543_ la_data_out_mprj[72] vssd vssd vccd vccd _543_/Y sky130_fd_sc_hd__inv_2
X_474_ la_data_out_mprj[3] vssd vssd vccd vccd _474_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1053 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[126\] la_iena_mprj[126] mprj_logic_high_inst/HI[456] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[126\]/B sky130_fd_sc_hd__and2_1
Xla_buf\[54\] _525_/Y la_buf\[54\]/TE vssd vssd vccd vccd la_data_in_core[54] sky130_fd_sc_hd__einvp_8
XFILLER_13_520 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[56\]_A la_data_out_core[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[18\] _425_/Y mprj_adr_buf\[18\]/TE vssd vssd vccd vccd mprj_adr_o_user[18]
+ sky130_fd_sc_hd__einvp_8
Xla_buf\[110\] _581_/Y la_buf\[110\]/TE vssd vssd vccd vccd la_data_in_core[110] sky130_fd_sc_hd__einvp_8
XFILLER_29_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_295 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_1839 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[98\] user_to_mprj_in_gates\[98\]/Y vssd vssd vccd vccd la_data_in_mprj[98]
+ sky130_fd_sc_hd__inv_8
XFILLER_42_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[6\]_A user_to_mprj_in_gates\[6\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[43\] la_data_out_core[43] user_to_mprj_in_gates\[43\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[43\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_23_317 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_16_380 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[47\]_A la_data_out_core[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1304 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__614__A la_oenb_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[5\] la_data_out_core[5] user_to_mprj_in_gates\[5\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[5\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_41_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_56 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_34 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_89 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_648 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_78 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_67 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_22_350 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[38\]_A la_data_out_core[38] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_523 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[122\]_A la_data_out_core[122] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_6_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__524__A la_data_out_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1568 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[94\] _362_/Y mprj_logic_high_inst/HI[296] vssd vssd vccd
+ vccd la_oenb_core[94] sky130_fd_sc_hd__einvp_8
XFILLER_1_210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_711 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[22\]_TE la_buf\[22\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[7\] la_iena_mprj[7] mprj_logic_high_inst/HI[337] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[7\]/B sky130_fd_sc_hd__and2_1
XFILLER_1_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xla_buf_enable\[117\] la_oenb_mprj[117] la_buf_enable\[117\]/B vssd vssd vccd vccd
+ la_buf\[117\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_20_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1482 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_526_ la_data_out_mprj[55] vssd vssd vccd vccd _526_/Y sky130_fd_sc_hd__inv_2
XFILLER_17_199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_457_ mprj_dat_o_core[18] vssd vssd vccd vccd _457_/Y sky130_fd_sc_hd__inv_2
XFILLER_20_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_40_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[29\]_A la_data_out_core[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_388_ la_oenb_mprj[120] vssd vssd vccd vccd _388_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_gates\[113\]_A la_data_out_core[113] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__434__A mprj_adr_o_core[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[13\] user_to_mprj_in_gates\[13\]/Y vssd vssd vccd vccd la_data_in_mprj[13]
+ sky130_fd_sc_hd__inv_8
XFILLER_47_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1625 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1382 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_48_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_954 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__609__A la_oenb_mprj[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_486 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[104\]_A la_data_out_core[104] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__344__A la_oenb_mprj[76] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1230 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[53\] la_iena_mprj[53] mprj_logic_high_inst/HI[383] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[53\]/B sky130_fd_sc_hd__and2_1
XFILLER_25_1984 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_420 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__519__A la_data_out_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[5\] user_to_mprj_in_gates\[5\]/Y vssd vssd vccd vccd la_data_in_mprj[5]
+ sky130_fd_sc_hd__inv_8
Xla_buf_enable\[31\] la_oenb_mprj[31] la_buf_enable\[31\]/B vssd vssd vccd vccd la_buf\[31\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_48_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[17\] _488_/Y la_buf\[17\]/TE vssd vssd vccd vccd la_data_in_core[17] sky130_fd_sc_hd__einvp_8
XFILLER_32_1999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1387 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1759 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_762 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__429__A mprj_adr_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_509_ la_data_out_mprj[38] vssd vssd vccd vccd _509_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf\[68\]_TE la_buf\[68\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_2040 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[2\]_B la_buf_enable\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1973 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[117\] la_data_out_core[117] user_to_mprj_in_gates\[117\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[117\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA_user_to_mprj_in_ena_buf\[126\]_A la_iena_mprj[126] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_740 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__339__A la_oenb_mprj[71] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_407 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_429 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_418 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1028 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1017 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1006 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1039 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_mprj_dat_buf\[17\]_TE mprj_dat_buf\[17\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[127\] _395_/Y mprj_logic_high_inst/HI[329] vssd vssd vccd
+ vccd la_oenb_core[127] sky130_fd_sc_hd__einvp_8
XFILLER_47_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[57\] _656_/Y mprj_logic_high_inst/HI[259] vssd vssd vccd
+ vccd la_oenb_core[57] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[79\] la_oenb_mprj[79] la_buf_enable\[79\]/B vssd vssd vccd vccd la_buf\[79\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[117\]_A la_iena_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_98 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_445 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_294 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_930 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1530 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_963 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_31_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_952 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_941 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_489 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_996 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_985 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_974 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[110\]_A_N la_oenb_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1763 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_677 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[125\]_A_N la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[114\] user_to_mprj_in_gates\[114\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[114] sky130_fd_sc_hd__inv_8
XFILLER_26_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[108\]_A la_iena_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[80\] user_to_mprj_in_gates\[80\]/Y vssd vssd vccd vccd la_data_in_mprj[80]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_743 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1803 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__622__A la_oenb_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1836 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1770 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_17_57 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_215 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_204 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_259 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_237 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_248 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_226 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1794 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[16\] la_iena_mprj[16] mprj_logic_high_inst/HI[346] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[16\]/B sky130_fd_sc_hd__and2_1
XFILLER_32_1004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_419 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[30\]_A la_iena_mprj[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1048 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__532__A la_data_out_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1471 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[97\]_A la_iena_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[84\] _555_/Y la_buf\[84\]/TE vssd vssd vccd vccd la_data_in_core[84] sky130_fd_sc_hd__einvp_8
XFILLER_47_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1694 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_771 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_760 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1202 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[21\]_A la_iena_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_782 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_982 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_793 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__442__A mprj_dat_o_core[3] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[88\]_A la_iena_mprj[88] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[73\] la_data_out_core[73] user_to_mprj_in_gates\[73\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[73\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_45_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__617__A la_oenb_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[12\]_A la_iena_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__352__A la_oenb_mprj[84] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[79\]_A la_iena_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[40\]_TE mprj_logic_high_inst/HI[242] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_490_ la_data_out_mprj[19] vssd vssd vccd vccd _490_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__527__A la_data_out_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1588 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1673 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_0_694 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2078 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__437__A mprj_adr_o_core[30] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_573 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[43\] user_to_mprj_in_gates\[43\]/Y vssd vssd vccd vccd la_data_in_mprj[43]
+ sky130_fd_sc_hd__inv_8
XFILLER_34_1655 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_590 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2080 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_2127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_39_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_164 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__347__A la_oenb_mprj[79] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1739 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_11_1463 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[83\] la_iena_mprj[83] mprj_logic_high_inst/HI[413] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[83\]/B sky130_fd_sc_hd__and2_1
XFILLER_46_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_447 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_55 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1879 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_611_ la_oenb_mprj[12] vssd vssd vccd vccd _611_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_in_buffers\[50\]_A user_to_mprj_in_gates\[50\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[61\] la_oenb_mprj[61] la_buf_enable\[61\]/B vssd vssd vccd vccd la_buf\[61\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_542_ la_data_out_mprj[71] vssd vssd vccd vccd _542_/Y sky130_fd_sc_hd__inv_2
XFILLER_22_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_473_ la_data_out_mprj[2] vssd vssd vccd vccd _473_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[47\] _518_/Y la_buf\[47\]/TE vssd vssd vccd vccd la_data_in_core[47] sky130_fd_sc_hd__einvp_8
XFILLER_40_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[83\]_A_N la_oenb_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[119\] la_iena_mprj[119] mprj_logic_high_inst/HI[449] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[119\]/B sky130_fd_sc_hd__and2_1
XANTENNA_la_buf\[90\]_A _561_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[86\]_TE mprj_logic_high_inst/HI[288] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[98\]_A_N la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_797 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[103\] _574_/Y la_buf\[103\]/TE vssd vssd vccd vccd la_data_in_core[103] sky130_fd_sc_hd__einvp_8
XFILLER_42_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[21\]_A_N la_oenb_mprj[21] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[41\]_A user_to_mprj_in_gates\[41\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_657 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_A_N la_oenb_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[36\] la_data_out_core[36] user_to_mprj_in_gates\[36\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[36\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_32_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_362 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_1452 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[81\]_A _552_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__630__A la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_8_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_1434 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[32\]_A user_to_mprj_in_gates\[32\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_35 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_79 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_68 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_57 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_10_502 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_362 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_10_535 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_517 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_1672 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf\[72\]_A _543_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_539 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1260 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_1883 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__540__A la_data_out_mprj[69] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[87\] _355_/Y mprj_logic_high_inst/HI[289] vssd vssd vccd
+ vccd la_oenb_core[87] sky130_fd_sc_hd__einvp_8
XFILLER_1_222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_1632 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[23\]_A user_to_mprj_in_gates\[23\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_46_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_999 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1472 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_525_ la_data_out_mprj[54] vssd vssd vccd vccd _525_/Y sky130_fd_sc_hd__inv_2
XFILLER_33_649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[126\]_A _597_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_456_ mprj_dat_o_core[17] vssd vssd vccd vccd _456_/Y sky130_fd_sc_hd__inv_2
X_387_ la_oenb_mprj[119] vssd vssd vccd vccd _387_/Y sky130_fd_sc_hd__inv_2
XFILLER_40_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[30\] _437_/Y mprj_adr_buf\[30\]/TE vssd vssd vccd vccd mprj_adr_o_user[30]
+ sky130_fd_sc_hd__einvp_8
XFILLER_12_1013 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[63\]_A _534_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__450__A mprj_dat_o_core[11] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_29_1532 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_2108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[14\]_A user_to_mprj_in_gates\[14\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_966 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_465 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_498 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[117\]_A _588_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__625__A la_oenb_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[54\]_A _525_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__360__A la_oenb_mprj[92] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1242 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[46\] la_iena_mprj[46] mprj_logic_high_inst/HI[376] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[46\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[108\]_A _579_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_19_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__535__A la_data_out_mprj[64] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[24\] la_oenb_mprj[24] la_buf_enable\[24\]/B vssd vssd vccd vccd la_buf\[24\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[63\]_B la_buf_enable\[63\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1399 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_508_ la_data_out_mprj[37] vssd vssd vccd vccd _508_/Y sky130_fd_sc_hd__inv_2
XANTENNA__445__A mprj_dat_o_core[6] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_439_ mprj_dat_o_core[0] vssd vssd vccd vccd _439_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_1108 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_1477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[54\]_B la_buf_enable\[54\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_2052 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_391 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1401 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1985 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_82 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[126\]_B mprj_logic_high_inst/HI[456] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_28_218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_3_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_408 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[12\]_TE la_buf\[12\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_419 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1029 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1018 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1007 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__355__A la_oenb_mprj[87] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1528 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[45\]_B la_buf_enable\[45\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_47_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[117\]_B mprj_logic_high_inst/HI[447] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_19_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_284 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_920 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_43_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_953 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_942 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_931 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1542 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_997 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_986 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_975 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_964 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1775 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[101\] la_iena_mprj[101] mprj_logic_high_inst/HI[431] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[101\]/B sky130_fd_sc_hd__and2_1
XFILLER_6_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[36\]_B la_buf_enable\[36\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[5\]_A la_iena_mprj[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_26_1513 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[107\] user_to_mprj_in_gates\[107\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[107] sky130_fd_sc_hd__inv_8
XFILLER_26_1557 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_43_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[73\] user_to_mprj_in_gates\[73\]/Y vssd vssd vccd vccd la_data_in_mprj[73]
+ sky130_fd_sc_hd__inv_8
XFILLER_39_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_21_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[27\]_B la_buf_enable\[27\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1782 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[6\] _445_/Y mprj_dat_buf\[6\]/TE vssd vssd vccd vccd mprj_dat_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_42_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_216 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_205 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_40_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_238 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_249 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_227 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_16_1704 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[3\]_TE la_buf\[3\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[18\]_B la_buf_enable\[18\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[91\] la_oenb_mprj[91] la_buf_enable\[91\]/B vssd vssd vccd vccd la_buf\[91\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_ena_buf\[97\]_B mprj_logic_high_inst/HI[427] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[77\] _548_/Y la_buf\[77\]/TE vssd vssd vccd vccd la_data_in_core[77] sky130_fd_sc_hd__einvp_8
XPHY_750 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_761 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_772 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_783 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_794 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1258 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_998 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1870 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_847 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[66\] la_data_out_core[66] user_to_mprj_in_gates\[66\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[66\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_43_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1161 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1759 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1483 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__633__A la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[79\]_B mprj_logic_high_inst/HI[409] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_22_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[5\]_A la_data_out_core[5] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[124\]_A_N la_oenb_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1545 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__543__A la_data_out_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_1280 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_5_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_651 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1367 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_oen_buffers\[9\]_TE mprj_logic_high_inst/HI[211] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_buffers\[36\] user_to_mprj_in_gates\[36\]/Y vssd vssd vccd vccd la_data_in_mprj[36]
+ sky130_fd_sc_hd__inv_8
XPHY_580 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1667 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__453__A mprj_dat_o_core[14] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1509 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_591 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_795 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__628__A la_oenb_mprj[29] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_198 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_22_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__363__A la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[76\] la_iena_mprj[76] mprj_logic_high_inst/HI[406] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[76\]/B sky130_fd_sc_hd__and2_1
XFILLER_24_1814 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_oen_buffers\[102\] _370_/Y mprj_logic_high_inst/HI[304] vssd vssd vccd
+ vccd la_oenb_core[102] sky130_fd_sc_hd__einvp_8
XFILLER_44_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_610_ la_oenb_mprj[11] vssd vssd vccd vccd _610_/Y sky130_fd_sc_hd__inv_2
XANTENNA__538__A la_data_out_mprj[67] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[32\] _631_/Y mprj_logic_high_inst/HI[234] vssd vssd vccd
+ vccd la_oenb_core[32] sky130_fd_sc_hd__einvp_8
X_541_ la_data_out_mprj[70] vssd vssd vccd vccd _541_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[54\] la_oenb_mprj[54] la_buf_enable\[54\]/B vssd vssd vccd vccd la_buf\[54\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_472_ la_data_out_mprj[1] vssd vssd vccd vccd _472_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1033 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_12_1228 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_5_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__448__A mprj_dat_o_core[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_36_669 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1707 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[29\] la_data_out_core[29] user_to_mprj_in_gates\[29\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[29\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_32_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[30\]_TE mprj_logic_high_inst/HI[232] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__358__A la_oenb_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_47 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_41_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_69 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_10_547 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_17_1684 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[5\]_TE mprj_adr_buf\[5\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[28\] _467_/Y mprj_dat_buf\[28\]/TE vssd vssd vccd vccd mprj_dat_o_user[28]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1738 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_978 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_146 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_524_ la_data_out_mprj[53] vssd vssd vccd vccd _524_/Y sky130_fd_sc_hd__inv_2
X_455_ mprj_dat_o_core[16] vssd vssd vccd vccd _455_/Y sky130_fd_sc_hd__inv_2
X_386_ la_oenb_mprj[118] vssd vssd vccd vccd _386_/Y sky130_fd_sc_hd__inv_2
Xmprj_adr_buf\[23\] _430_/Y mprj_adr_buf\[23\]/TE vssd vssd vccd vccd mprj_adr_o_user[23]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[9\]_TE mprj_dat_buf\[9\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_29_1544 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1522 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1788 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[8\] la_oenb_mprj[8] la_buf_enable\[8\]/B vssd vssd vccd vccd la_buf\[8\]/TE
+ sky130_fd_sc_hd__and2b_1
XANTENNA__641__A la_oenb_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1633 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[82\]_A_N la_oenb_mprj[82] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_271 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_444 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_904 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[39\] la_iena_mprj[39] mprj_logic_high_inst/HI[369] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[39\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[97\]_A_N la_oenb_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[20\]_A_N la_oenb_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf_enable\[17\] la_oenb_mprj[17] la_buf_enable\[17\]/B vssd vssd vccd vccd la_buf\[17\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_315 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__551__A la_data_out_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_32_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[35\]_A_N la_oenb_mprj[35] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_irq_gates\[0\] user_irq_core[0] user_irq_gates\[0\]/B vssd vssd vccd vccd user_irq_gates\[0\]/Y
+ sky130_fd_sc_hd__nand2_4
XFILLER_2_521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_2_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_2142 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_2_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[122\] la_oenb_mprj[122] la_buf_enable\[122\]/B vssd vssd vccd vccd
+ la_buf\[122\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_4_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_414 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_488 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_507_ la_data_out_mprj[36] vssd vssd vccd vccd _507_/Y sky130_fd_sc_hd__inv_2
X_438_ mprj_adr_o_core[31] vssd vssd vccd vccd _438_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_369_ la_oenb_mprj[101] vssd vssd vccd vccd _369_/Y sky130_fd_sc_hd__inv_2
XANTENNA__461__A mprj_dat_o_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[96\] la_data_out_core[96] user_to_mprj_in_gates\[96\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[96\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_29_2064 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_9_1413 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1997 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_94 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[99\]_TE mprj_logic_high_inst/HI[301] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__636__A la_oenb_mprj[37] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_409 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_36_1323 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1019 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1008 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__371__A la_oenb_mprj[103] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_1349 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_56 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__546__A la_data_out_mprj[75] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_910 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_921 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_954 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_943 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_932 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_19_1554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_987 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_976 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_965 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_998 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[22\] _493_/Y la_buf\[22\]/TE vssd vssd vccd vccd la_data_in_core[22] sky130_fd_sc_hd__einvp_8
XFILLER_7_646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1787 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_156 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1175 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[5\]_B mprj_logic_high_inst/HI[335] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_3_896 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1525 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_43_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1365 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_stb_buf_TE mprj_stb_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[66\] user_to_mprj_in_gates\[66\]/Y vssd vssd vccd vccd la_data_in_mprj[66]
+ sky130_fd_sc_hd__inv_8
XFILLER_4_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_767 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__456__A mprj_dat_o_core[17] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[11\] la_data_out_core[11] user_to_mprj_in_gates\[11\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[11\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_31_1275 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_1232 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_1794 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_2061 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[122\] la_data_out_core[122] user_to_mprj_in_gates\[122\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[122\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_5_1107 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_2094 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_206 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__366__A la_oenb_mprj[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_217 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_239 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_228 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_929 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_266 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[95\]_A la_data_out_core[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1716 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1326 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[31\]_TE mprj_adr_buf\[31\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_oen_buffers\[62\] _330_/Y mprj_logic_high_inst/HI[264] vssd vssd vccd
+ vccd la_oenb_core[62] sky130_fd_sc_hd__einvp_8
XFILLER_7_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[84\] la_oenb_mprj[84] la_buf_enable\[84\]/B vssd vssd vccd vccd la_buf\[84\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_48_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[10\] _449_/Y mprj_dat_buf\[10\]/TE vssd vssd vccd vccd mprj_dat_o_user[10]
+ sky130_fd_sc_hd__einvp_8
XFILLER_0_877 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1580 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[86\]_A la_data_out_core[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_751 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_762 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_740 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_773 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_784 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_795 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_472 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[126\] _597_/Y la_buf\[126\]/TE vssd vssd vccd vccd la_data_in_core[126] sky130_fd_sc_hd__einvp_8
XFILLER_26_2001 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2067 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_user_to_mprj_in_gates\[10\]_A la_data_out_core[10] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_347 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[59\] la_data_out_core[59] user_to_mprj_in_gates\[59\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[59\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_47_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_561 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1440 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[77\]_A la_data_out_core[77] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_48_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1422 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1319 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1308 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_28_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[5\]_B user_to_mprj_in_gates\[5\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[21\] la_iena_mprj[21] mprj_logic_high_inst/HI[351] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[21\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[68\]_A la_data_out_core[68] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_247 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_16_1557 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_33_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_903 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[25\]_TE la_buf\[25\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1292 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_479 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_27_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_663 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_23_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_634 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_36_807 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_A la_data_out_core[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_570 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[29\] user_to_mprj_in_gates\[29\]/Y vssd vssd vccd vccd la_data_in_mprj[29]
+ sky130_fd_sc_hd__inv_8
XPHY_581 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_592 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1679 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_32_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_4_991 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_38_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[9\]_A user_to_mprj_in_gates\[9\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1224 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_26_339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__644__A la_oenb_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[48\]_TE la_buf\[48\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_ena_buf\[69\] la_iena_mprj[69] mprj_logic_high_inst/HI[399] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[69\]/B sky130_fd_sc_hd__and2_1
XFILLER_44_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1149 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_540_ la_data_out_mprj[69] vssd vssd vccd vccd _540_/Y sky130_fd_sc_hd__inv_2
X_471_ la_data_out_mprj[0] vssd vssd vccd vccd _471_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[7\] _606_/Y mprj_logic_high_inst/HI[209] vssd vssd vccd
+ vccd la_oenb_core[7] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[25\] _624_/Y mprj_logic_high_inst/HI[227] vssd vssd vccd
+ vccd la_oenb_core[25] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[47\] la_oenb_mprj[47] la_buf_enable\[47\]/B vssd vssd vccd vccd la_buf\[47\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_38_1056 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[125\]_A la_data_out_core[125] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XANTENNA__554__A la_data_out_mprj[83] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[0\] _471_/Y la_buf\[0\]/TE vssd vssd vccd vccd la_data_in_core[0] sky130_fd_sc_hd__einvp_8
XFILLER_5_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_431 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1959 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_40_1650 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1683 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_1719 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[116\]_A la_data_out_core[116] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_43_180 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_32_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__464__A mprj_dat_o_core[25] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[123\]_A_N la_oenb_mprj[123] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__639__A la_oenb_mprj[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_475 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_604 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_59 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_gates\[107\]_A la_data_out_core[107] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_34_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__374__A la_oenb_mprj[106] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1630 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_559 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1696 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_58 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_11_1240 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_703 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1706 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__549__A la_data_out_mprj[78] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1678 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_1441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_523_ la_data_out_mprj[52] vssd vssd vccd vccd _523_/Y sky130_fd_sc_hd__inv_2
X_454_ mprj_dat_o_core[15] vssd vssd vccd vccd _454_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_832 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_41_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[52\] _523_/Y la_buf\[52\]/TE vssd vssd vccd vccd la_data_in_core[52] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[124\] la_iena_mprj[124] mprj_logic_high_inst/HI[454] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[124\]/B sky130_fd_sc_hd__and2_1
XFILLER_9_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_385_ la_oenb_mprj[117] vssd vssd vccd vccd _385_/Y sky130_fd_sc_hd__inv_2
XFILLER_12_1015 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[16\] _423_/Y mprj_adr_buf\[16\]/TE vssd vssd vccd vccd mprj_adr_o_user[16]
+ sky130_fd_sc_hd__einvp_8
XFILLER_29_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[96\] user_to_mprj_in_gates\[96\]/Y vssd vssd vccd vccd la_data_in_mprj[96]
+ sky130_fd_sc_hd__inv_8
XFILLER_7_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__459__A mprj_dat_o_core[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_rstn_buf _396_/Y mprj_rstn_buf/TE vssd vssd vccd vccd user_resetn sky130_fd_sc_hd__einvp_8
XFILLER_7_1374 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[41\] la_data_out_core[41] user_to_mprj_in_gates\[41\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[41\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_34_1251 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_34_1284 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[5\]_B la_buf_enable\[5\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1645 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_gates\[3\] la_data_out_core[3] user_to_mprj_in_gates\[3\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[3\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_47_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__369__A la_oenb_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_283 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_23_640 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[60\]_A la_iena_mprj[60] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1713 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1702 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1724 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1735 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1746 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1757 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1768 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_367 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1779 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_327 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_13_1379 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_oen_buffers\[92\] _360_/Y mprj_logic_high_inst/HI[294] vssd vssd vccd
+ vccd la_oenb_core[92] sky130_fd_sc_hd__einvp_8
XFILLER_11_1081 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_1729 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[5\] la_iena_mprj[5] mprj_logic_high_inst/HI[335] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[5\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_1536 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1683 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[115\] la_oenb_mprj[115] la_buf_enable\[115\]/B vssd vssd vccd vccd
+ la_buf\[115\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_45_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1569 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[20\]_TE mprj_logic_high_inst/HI[222] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_938 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_33_426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_506_ la_data_out_mprj[35] vssd vssd vccd vccd _506_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1260 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_37_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[51\]_A la_iena_mprj[51] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_80 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_437_ mprj_adr_o_core[30] vssd vssd vccd vccd _437_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_109 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_2136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_368_ la_oenb_mprj[100] vssd vssd vccd vccd _368_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_in_buffers\[11\] user_to_mprj_in_gates\[11\]/Y vssd vssd vccd vccd la_data_in_mprj[11]
+ sky130_fd_sc_hd__inv_8
XFILLER_48_1910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_47_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2126 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[89\] la_data_out_core[89] user_to_mprj_in_gates\[89\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[89\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_1425 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1447 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_51 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_36_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_37_754 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_A la_iena_mprj[42] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1335 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_33_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_960 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1009 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__652__A la_oenb_mprj[53] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_22_38 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_47_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_14_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[43\]_TE mprj_logic_high_inst/HI[245] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[51\] la_iena_mprj[51] mprj_logic_high_inst/HI[381] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[51\]/B sky130_fd_sc_hd__and2_1
XFILLER_19_209 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_1615 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_41_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_220 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_cyc_buf _400_/Y mprj_cyc_buf/TE vssd vssd vccd vccd mprj_cyc_o_user sky130_fd_sc_hd__einvp_8
XFILLER_27_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_900 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[33\]_A la_iena_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_911 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_944 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_933 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[3\] user_to_mprj_in_gates\[3\]/Y vssd vssd vccd vccd la_data_in_mprj[3]
+ sky130_fd_sc_hd__inv_8
XPHY_922 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1521 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1510 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1532 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_988 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_977 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_966 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_955 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1576 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1565 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1554 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1543 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_999 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__562__A la_data_out_mprj[91] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_1598 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1587 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[15\] _486_/Y la_buf\[15\]/TE vssd vssd vccd vccd la_data_in_core[15] sky130_fd_sc_hd__einvp_8
XFILLER_6_168 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[0\]_A _439_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1187 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_adr_buf\[8\] _415_/Y mprj_adr_buf\[8\]/TE vssd vssd vccd vccd mprj_adr_o_user[8]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1300 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_2045 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_8_1480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2078 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1377 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_90 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[59\] user_to_mprj_in_gates\[59\]/Y vssd vssd vccd vccd la_data_in_mprj[59]
+ sky130_fd_sc_hd__inv_8
XANTENNA_user_to_mprj_in_ena_buf\[24\]_A la_iena_mprj[24] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1666 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_481 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__472__A la_data_out_mprj[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[81\]_A_N la_oenb_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1828 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_oen_buffers\[66\]_TE mprj_logic_high_inst/HI[268] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[96\]_A_N la_oenb_mprj[96] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1211 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_44_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1244 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_2073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1119 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[115\] la_data_out_core[115] user_to_mprj_in_gates\[115\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[115\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__647__A la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_38 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_201 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_207 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_in_ena_buf\[15\]_A la_iena_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[34\]_A_N la_oenb_mprj[34] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_40_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_218 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_229 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_24_256 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_1728 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__382__A la_oenb_mprj[114] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[49\]_A_N la_oenb_mprj[49] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_clk2_buf_TE mprj_clk2_buf/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_ena_buf\[99\] la_iena_mprj[99] mprj_logic_high_inst/HI[429] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[99\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_628 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[30\]_TE mprj_dat_buf\[30\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[125\] _393_/Y mprj_logic_high_inst/HI[327] vssd vssd vccd
+ vccd la_oenb_core[125] sky130_fd_sc_hd__einvp_8
XFILLER_27_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1918 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[55\] _654_/Y mprj_logic_high_inst/HI[257] vssd vssd vccd
+ vccd la_oenb_core[55] sky130_fd_sc_hd__einvp_8
Xla_buf_enable\[77\] la_oenb_mprj[77] la_buf_enable\[77\]/B vssd vssd vccd vccd la_buf\[77\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_1592 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_irq_ena_buf\[2\]_A user_irq_ena[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__557__A la_data_out_mprj[86] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_752 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_763 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_730 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_741 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1340 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1351 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_248 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_774 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_785 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_796 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1373 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1362 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1384 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_user_to_mprj_oen_buffers\[89\]_TE mprj_logic_high_inst/HI[291] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1395 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[119\] _590_/Y la_buf\[119\]/TE vssd vssd vccd vccd la_data_in_core[119] sky130_fd_sc_hd__einvp_8
XFILLER_48_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_26_2013 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2046 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_2118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[112\] user_to_mprj_in_gates\[112\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[112] sky130_fd_sc_hd__inv_8
XFILLER_26_2079 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[10\]_B user_to_mprj_in_gates\[10\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_38_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__467__A mprj_dat_o_core[28] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2017 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1603 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_44_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[62\]_A user_to_mprj_in_gates\[62\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_359 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__377__A la_oenb_mprj[109] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_554 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[14\] la_iena_mprj[14] mprj_logic_high_inst/HI[344] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[14\]/B sky130_fd_sc_hd__and2_1
XFILLER_40_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_208 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[100\]_A user_to_mprj_in_gates\[100\]/Y vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_buffers\[53\]_A user_to_mprj_in_gates\[53\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1665 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_27_1687 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1518 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_819 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[82\] _553_/Y la_buf\[82\]/TE vssd vssd vccd vccd la_data_in_core[82] sky130_fd_sc_hd__einvp_8
XFILLER_5_1450 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_40_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_392 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_370 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1369 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[59\]_B user_to_mprj_in_gates\[59\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_31_568 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XPHY_571 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_560 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[93\]_A _564_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_582 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_593 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1181 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1170 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1192 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_241 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_1057 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_480 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_602 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[71\] la_data_out_core[71] user_to_mprj_in_gates\[71\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[71\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_123 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[21\]_TE mprj_adr_buf\[21\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[84\]_A _555_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_22_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_30_38 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__660__A la_oenb_mprj[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1231 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_buffers\[35\]_A user_to_mprj_in_gates\[35\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_58 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1634 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_2_1623 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_17_307 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_470_ mprj_dat_o_core[31] vssd vssd vccd vccd _470_/Y sky130_fd_sc_hd__inv_2
Xuser_to_mprj_oen_buffers\[18\] _617_/Y mprj_logic_high_inst/HI[220] vssd vssd vccd
+ vccd la_oenb_core[18] sky130_fd_sc_hd__einvp_8
XFILLER_38_1068 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[75\]_A _546_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__570__A la_data_out_mprj[99] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_1705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_789 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_71 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_45_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[26\]_A user_to_mprj_in_gates\[26\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_0_494 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1695 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1662 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1166 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_170 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_599_ la_oenb_mprj[0] vssd vssd vccd vccd _599_/Y sky130_fd_sc_hd__inv_2
XFILLER_34_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_343 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_buffers\[41\] user_to_mprj_in_gates\[41\]/Y vssd vssd vccd vccd la_data_in_mprj[41]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[66\]_A _537_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1455 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_390 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_550 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__480__A la_data_out_mprj[9] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_47_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[17\]_A user_to_mprj_in_gates\[17\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1011 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1437 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_487 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_616 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[15\]_TE la_buf\[15\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_3_1987 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__655__A la_oenb_mprj[56] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_49 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_34_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[57\]_A _528_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_17_1642 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1675 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_17_1664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_398 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[75\]_B la_buf_enable\[75\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__390__A la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1886 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1875 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_46_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[81\] la_iena_mprj[81] mprj_logic_high_inst/HI[411] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[81\]/B sky130_fd_sc_hd__and2_1
XFILLER_8_1821 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1718 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_608 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_522_ la_data_out_mprj[51] vssd vssd vccd vccd _522_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_453_ mprj_dat_o_core[14] vssd vssd vccd vccd _453_/Y sky130_fd_sc_hd__inv_2
XANTENNA__565__A la_data_out_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_14_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_844 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_384_ la_oenb_mprj[116] vssd vssd vccd vccd _384_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[45\] _516_/Y la_buf\[45\]/TE vssd vssd vccd vccd la_data_in_core[45] sky130_fd_sc_hd__einvp_8
XFILLER_35_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_ena_buf\[117\] la_iena_mprj[117] mprj_logic_high_inst/HI[447] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[117\]/B sky130_fd_sc_hd__and2_1
XFILLER_12_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[101\] _572_/Y la_buf\[101\]/TE vssd vssd vccd vccd la_data_in_core[101] sky130_fd_sc_hd__einvp_8
XFILLER_7_2032 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_2065 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_291 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[89\] user_to_mprj_in_gates\[89\]/Y vssd vssd vccd vccd la_data_in_mprj[89]
+ sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_gates\[34\] la_data_out_core[34] user_to_mprj_in_gates\[34\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[34\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__475__A la_data_out_mprj[4] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_870 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[57\]_B la_buf_enable\[57\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1296 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1572 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_48 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_27_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA__385__A la_oenb_mprj[117] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1141 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_490 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[60\]_B mprj_logic_high_inst/HI[390] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_1703 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf\[6\]_TE la_buf\[6\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1714 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1725 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1736 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1747 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1758 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1769 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_10_379 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_13_1336 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_oen_buffers\[85\] _353_/Y mprj_logic_high_inst/HI[287] vssd vssd vccd
+ vccd la_oenb_core[85] sky130_fd_sc_hd__einvp_8
XFILLER_7_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1548 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[108\] la_oenb_mprj[108] la_buf_enable\[108\]/B vssd vssd vccd vccd
+ la_buf\[108\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_45_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_505_ la_data_out_mprj[34] vssd vssd vccd vccd _505_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[122\]_A_N la_oenb_mprj[122] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_436_ mprj_adr_o_core[29] vssd vssd vccd vccd _436_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_367_ la_oenb_mprj[99] vssd vssd vccd vccd _367_/Y sky130_fd_sc_hd__inv_2
XANTENNA_la_buf_enable\[39\]_B la_buf_enable\[39\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1458 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_891 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[8\]_A la_iena_mprj[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_9_2105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[106\]_A _374_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2138 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1437 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_1150 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[42\]_B mprj_logic_high_inst/HI[372] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_20_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1781 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xuser_to_mprj_in_ena_buf\[44\] la_iena_mprj[44] mprj_logic_high_inst/HI[374] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[44\]/B sky130_fd_sc_hd__and2_1
XFILLER_3_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_901 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_912 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1500 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_945 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_934 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_923 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1522 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1511 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1533 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_978 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_967 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_956 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_622 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[22\] la_oenb_mprj[22] la_buf_enable\[22\]/B vssd vssd vccd vccd la_buf\[22\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1566 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1555 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1544 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_989 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1100 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1599 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1588 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1577 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1199 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1491 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_4_1389 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_254 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_18_287 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[24\]_B mprj_logic_high_inst/HI[354] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1678 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_419_ mprj_adr_o_core[12] vssd vssd vccd vccd _419_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_953 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_14_493 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1222 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1255 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[111\]_TE mprj_logic_high_inst/HI[313] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_681 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1741 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_44_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[108\] la_data_out_core[108] user_to_mprj_in_gates\[108\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[108\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_0_1721 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1890 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[15\]_B mprj_logic_high_inst/HI[345] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1111 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_219 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_208 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_36_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_33_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_10_1339 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[10\]_TE mprj_logic_high_inst/HI[212] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[118\] _386_/Y mprj_logic_high_inst/HI[320] vssd vssd vccd
+ vccd la_oenb_core[118] sky130_fd_sc_hd__einvp_8
XFILLER_27_1858 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_868 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[8\]_A la_data_out_core[8] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_530 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[48\] _647_/Y mprj_logic_high_inst/HI[250] vssd vssd vccd
+ vccd la_oenb_core[48] sky130_fd_sc_hd__einvp_8
XFILLER_5_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_irq_ena_buf\[2\]_B user_irq_ena_buf\[2\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_720 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__573__A la_data_out_mprj[102] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_30_216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_753 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_731 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_742 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1330 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1341 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1829 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_8_913 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_764 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_775 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_786 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1374 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1363 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1352 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_797 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1396 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1385 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_485 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[105\] user_to_mprj_in_gates\[105\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[105] sky130_fd_sc_hd__inv_8
Xuser_to_mprj_in_buffers\[71\] user_to_mprj_in_gates\[71\]/Y vssd vssd vccd vccd la_data_in_mprj[71]
+ sky130_fd_sc_hd__inv_8
XFILLER_0_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2029 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__483__A la_data_out_mprj[12] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_1464 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1063 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1637 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_990 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xmprj_dat_buf\[4\] _443_/Y mprj_dat_buf\[4\]/TE vssd vssd vccd vccd mprj_dat_o_user[4]
+ sky130_fd_sc_hd__einvp_8
XFILLER_44_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__658__A la_oenb_mprj[59] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_42_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1206 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_38_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_566 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_0_1584 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__393__A la_oenb_mprj[125] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[8\]_TE mprj_adr_buf\[8\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_949 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_1611 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_0_610 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__568__A la_data_out_mprj[97] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_1699 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1833 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[80\]_A_N la_oenb_mprj[80] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_157 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_40_1866 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[71\]_TE la_buf\[71\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_1462 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_500 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[75\] _546_/Y la_buf\[75\]/TE vssd vssd vccd vccd la_data_in_core[75] sky130_fd_sc_hd__einvp_8
XFILLER_1_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[95\]_A_N la_oenb_mprj[95] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_550 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_561 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_572 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_583 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_594 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1182 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1171 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1193 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1160 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_271 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_15_1069 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_253 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[33\]_A_N la_oenb_mprj[33] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_492 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1204 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_614 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_135 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[48\]_A_N la_oenb_mprj[48] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_gates\[64\] la_data_out_core[64] user_to_mprj_in_gates\[64\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[64\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__478__A la_data_out_mprj[7] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_26_308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XANTENNA_mprj_dat_buf\[14\]_A _453_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_35_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[20\]_TE mprj_dat_buf\[20\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_10_709 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1434 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1806 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_29_113 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__388__A la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_801 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1717 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_2131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_440 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1674 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_105 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_598_ la_data_out_mprj[127] vssd vssd vccd vccd _598_/Y sky130_fd_sc_hd__inv_2
XFILLER_1_1178 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[34\] user_to_mprj_in_gates\[34\]/Y vssd vssd vccd vccd la_data_in_mprj[34]
+ sky130_fd_sc_hd__inv_8
XPHY_380 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1467 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_391 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_6_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_400 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1405 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1023 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1449 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_27_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1312 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_1_1690 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_25_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1378 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1898 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_1264 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_738 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_237 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
Xuser_to_mprj_in_ena_buf\[74\] la_iena_mprj[74] mprj_logic_high_inst/HI[404] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[74\]/B sky130_fd_sc_hd__and2_1
XFILLER_44_1073 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[100\] _368_/Y mprj_logic_high_inst/HI[302] vssd vssd vccd
+ vccd la_oenb_core[100] sky130_fd_sc_hd__einvp_8
XFILLER_45_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1410 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[30\] _629_/Y mprj_logic_high_inst/HI[232] vssd vssd vccd
+ vccd la_oenb_core[30] sky130_fd_sc_hd__einvp_8
XFILLER_45_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[52\] la_oenb_mprj[52] la_buf_enable\[52\]/B vssd vssd vccd vccd la_buf\[52\]/TE
+ sky130_fd_sc_hd__and2b_1
X_521_ la_data_out_mprj[50] vssd vssd vccd vccd _521_/Y sky130_fd_sc_hd__inv_2
X_452_ mprj_dat_o_core[13] vssd vssd vccd vccd _452_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_823 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_383_ la_oenb_mprj[115] vssd vssd vccd vccd _383_/Y sky130_fd_sc_hd__inv_2
XFILLER_14_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1743 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_41_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__581__A la_data_out_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[38\] _509_/Y la_buf\[38\]/TE vssd vssd vccd vccd la_data_in_core[38] sky130_fd_sc_hd__einvp_8
XFILLER_9_359 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_326 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[11\]_TE mprj_adr_buf\[11\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_2044 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_793 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_2077 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_irq_gates\[1\]_A user_irq_core[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_274 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_937 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[27\] la_data_out_core[27] user_to_mprj_in_gates\[27\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[27\]/Y sky130_fd_sc_hd__nand2_4
XANTENNA__491__A la_data_out_mprj[20] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1275 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_1117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_31_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1129 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_45_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_39_1120 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_adr_buf\[8\]_A _415_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1153 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1704 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1006 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1715 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_35_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1726 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1737 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1748 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1759 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[78\] _346_/Y mprj_logic_high_inst/HI[280] vssd vssd vccd
+ vccd la_oenb_core[78] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[26\] _465_/Y mprj_dat_buf\[26\]/TE vssd vssd vccd vccd mprj_dat_o_user[26]
+ sky130_fd_sc_hd__einvp_8
XFILLER_8_1652 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_1505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_41_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__576__A la_data_out_mprj[105] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_504_ la_data_out_mprj[33] vssd vssd vccd vccd _504_/Y sky130_fd_sc_hd__inv_2
XFILLER_37_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_962 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_435_ mprj_adr_o_core[28] vssd vssd vccd vccd _435_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1551 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_697 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_366_ la_oenb_mprj[98] vssd vssd vccd vccd _366_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1595 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_1426 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[21\] _428_/Y mprj_adr_buf\[21\]/TE vssd vssd vccd vccd mprj_adr_o_user[21]
+ sky130_fd_sc_hd__einvp_8
XFILLER_6_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_6_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_2117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[40\]_A la_data_out_core[40] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1162 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__486__A la_data_out_mprj[15] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_37_778 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_36_255 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_36_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_1969 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_36_2049 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[6\] la_oenb_mprj[6] la_buf_enable\[6\]/B vssd vssd vccd vccd la_buf\[6\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_47_2101 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1971 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_47_2134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[31\]_A la_data_out_core[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_47_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1786 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA__396__A caravel_rstn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_417 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[37\] la_iena_mprj[37] mprj_logic_high_inst/HI[367] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[37\]/B sky130_fd_sc_hd__and2_1
XFILLER_42_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[98\]_A la_data_out_core[98] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_902 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_3_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_935 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_913 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_924 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1523 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1512 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1501 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_979 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_968 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_957 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_946 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1567 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1556 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1545 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1534 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[15\] la_oenb_mprj[15] la_buf_enable\[15\]/B vssd vssd vccd vccd la_buf\[15\]/TE
+ sky130_fd_sc_hd__and2b_1
XPHY_1589 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1578 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_13_1112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1219 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[22\]_A la_data_out_core[22] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_2025 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[120\] la_oenb_mprj[120] la_buf_enable\[120\]/B vssd vssd vccd vccd
+ la_buf\[120\]/TE sky130_fd_sc_hd__and2b_1
XANTENNA_user_to_mprj_in_gates\[89\]_A la_data_out_core[89] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_236 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_910 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_418_ mprj_adr_o_core[11] vssd vssd vccd vccd _418_/Y sky130_fd_sc_hd__inv_2
XFILLER_41_280 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_349_ la_oenb_mprj[81] vssd vssd vccd vccd _349_/Y sky130_fd_sc_hd__inv_2
XFILLER_31_1267 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1278 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xuser_to_mprj_in_gates\[94\] la_data_out_core[94] user_to_mprj_in_gates\[94\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[94\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_6_693 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1753 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[13\]_A la_data_out_core[13] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_1279 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1396 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_1661 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1733 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_209 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_24_258 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_20_420 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_1590 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_453 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1318 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_825 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_1138 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_gates\[8\]_B user_to_mprj_in_gates\[8\]/B vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[121\]_A_N la_oenb_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_1_1519 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_710 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_743 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_754 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_921 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_721 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_732 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1331 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1320 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1342 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_30_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_765 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_776 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_787 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1375 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1364 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1353 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1532 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_7_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_798 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_23_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1397 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf\[20\] _491_/Y la_buf\[20\]/TE vssd vssd vccd vccd la_data_in_core[20] sky130_fd_sc_hd__einvp_8
XPHY_1386 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_457 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_958 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_1841 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_1852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_3_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_306 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_542 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_19_553 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_19_575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_534 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_0_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_buffers\[64\] user_to_mprj_in_gates\[64\]/Y vssd vssd vccd vccd la_data_in_mprj[64]
+ sky130_fd_sc_hd__inv_8
XFILLER_37_2144 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_34_567 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_37_1476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_15_792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_21_239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1075 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1043 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[120\] la_data_out_core[120] user_to_mprj_in_gates\[120\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[120\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_840 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1218 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_27 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_user_to_mprj_in_ena_buf\[110\]_A la_iena_mprj[110] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1830 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_294 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_4_449 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_4_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1295 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[60\] _659_/Y mprj_logic_high_inst/HI[262] vssd vssd vccd
+ vccd la_oenb_core[60] sky130_fd_sc_hd__einvp_8
XFILLER_7_1717 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf_enable\[82\] la_oenb_mprj[82] la_buf_enable\[82\]/B vssd vssd vccd vccd la_buf\[82\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_44_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_1845 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_309 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1474 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_40_1878 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_372 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[101\]_TE mprj_logic_high_inst/HI[303] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_44_876 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA__584__A la_data_out_mprj[113] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[68\] _539_/Y la_buf\[68\]/TE vssd vssd vccd vccd la_data_in_core[68] sky130_fd_sc_hd__einvp_8
XFILLER_38_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[101\]_A la_iena_mprj[101] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_34_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_540 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_551 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_562 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1150 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_573 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_584 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_595 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1026 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1183 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1172 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1161 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_755 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1194 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_265 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[124\] _595_/Y la_buf\[124\]/TE vssd vssd vccd vccd la_data_in_core[124] sky130_fd_sc_hd__einvp_8
XFILLER_7_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_972 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_626 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_1216 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1227 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[57\] la_data_out_core[57] user_to_mprj_in_gates\[57\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[57\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_46_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[119\]_A la_data_out_core[119] vssd vssd vccd vccd
+ sky130_fd_sc_hd__diode_2
XFILLER_35_876 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__494__A la_data_out_mprj[23] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1861 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_1894 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_397 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_570 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_30_581 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_11_1446 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_909 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1932 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[124\]_TE mprj_logic_high_inst/HI[326] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1531 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_ena_buf\[90\]_A la_iena_mprj[90] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_41_813 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_375 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_213 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_1729 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_27_2143 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__579__A la_data_out_mprj[108] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_7_1503 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_452 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_60 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_oen_buffers\[23\]_TE mprj_logic_high_inst/HI[225] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_489 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_35_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_180 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[81\]_A la_iena_mprj[81] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_331 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_70 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_597_ la_data_out_mprj[126] vssd vssd vccd vccd _597_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_1560 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_43_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_334 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_386 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_38_1593 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_370 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_392 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xuser_to_mprj_in_buffers\[27\] user_to_mprj_in_gates\[27\]/Y vssd vssd vccd vccd la_data_in_mprj[27]
+ sky130_fd_sc_hd__inv_8
XPHY_381 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1479 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_552 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1170 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_42 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__489__A la_data_out_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1417 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_412 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1035 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_640 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[72\]_A la_iena_mprj[72] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_26_139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_39_1324 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1508 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[8\]_B la_buf_enable\[8\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[61\]_TE la_buf\[61\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1276 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__399__A caravel_clk2 vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_oen_buffers\[46\]_TE mprj_logic_high_inst/HI[248] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf_enable\[94\]_A_N la_oenb_mprj[94] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_28_1784 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[67\] la_iena_mprj[67] mprj_logic_high_inst/HI[397] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[67\]/B sky130_fd_sc_hd__and2_1
XFILLER_41_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1085 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1422 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_2145 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_17_117 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_520_ la_data_out_mprj[49] vssd vssd vccd vccd _520_/Y sky130_fd_sc_hd__inv_2
XFILLER_18_629 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[63\]_A la_iena_mprj[63] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[23\] _622_/Y mprj_logic_high_inst/HI[225] vssd vssd vccd
+ vccd la_oenb_core[23] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_oen_buffers\[5\] _604_/Y mprj_logic_high_inst/HI[207] vssd vssd vccd
+ vccd la_oenb_core[5] sky130_fd_sc_hd__einvp_8
X_451_ mprj_dat_o_core[12] vssd vssd vccd vccd _451_/Y sky130_fd_sc_hd__inv_2
Xla_buf_enable\[45\] la_oenb_mprj[45] la_buf_enable\[45\]/B vssd vssd vccd vccd la_buf\[45\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_0_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_382_ la_oenb_mprj[114] vssd vssd vccd vccd _382_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_334 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[32\]_A_N la_oenb_mprj[32] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1711 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_356 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_14_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_338 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[47\]_A_N la_oenb_mprj[47] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_5_511 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_31_72 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[10\]_TE mprj_dat_buf\[10\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_7_1300 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_7_2089 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[54\]_A la_iena_mprj[54] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_982 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_649_ la_oenb_mprj[50] vssd vssd vccd vccd _649_/Y sky130_fd_sc_hd__inv_2
XFILLER_44_492 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_9_872 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1585 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_286 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_sel_buf\[2\]_A _405_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_3_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_ena_buf\[45\]_A la_iena_mprj[45] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_39_1132 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_621 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_1705 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1198 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1165 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1018 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_1716 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_22_131 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1727 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1738 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_827 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1749 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_46_1125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2113 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xmprj_dat_buf\[19\] _458_/Y mprj_dat_buf\[19\]/TE vssd vssd vccd vccd mprj_dat_o_user[19]
+ sky130_fd_sc_hd__einvp_8
XFILLER_41_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[36\]_A la_iena_mprj[36] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_2_1252 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_503_ la_data_out_mprj[32] vssd vssd vccd vccd _503_/Y sky130_fd_sc_hd__inv_2
X_434_ mprj_adr_o_core[27] vssd vssd vccd vccd _434_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_974 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__592__A la_data_out_mprj[121] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf\[50\] _521_/Y la_buf\[50\]/TE vssd vssd vccd vccd la_data_in_core[50] sky130_fd_sc_hd__einvp_8
Xuser_to_mprj_in_ena_buf\[122\] la_iena_mprj[122] mprj_logic_high_inst/HI[452] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[122\]/B sky130_fd_sc_hd__and2_1
X_365_ la_oenb_mprj[97] vssd vssd vccd vccd _365_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1563 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[3\]_A _442_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_31_1438 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_10_860 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[14\] _421_/Y mprj_adr_buf\[14\]/TE vssd vssd vccd vccd mprj_adr_o_user[14]
+ sky130_fd_sc_hd__einvp_8
XFILLER_48_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[94\] user_to_mprj_in_gates\[94\]/Y vssd vssd vccd vccd la_data_in_mprj[94]
+ sky130_fd_sc_hd__inv_8
XFILLER_36_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1027 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1174 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_in_ena_buf\[27\]_A la_iena_mprj[27] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1915 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_790 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_24_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_624 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_1761 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_680 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1658 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[1\] la_data_out_core[1] user_to_mprj_in_gates\[1\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[1\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_47_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_25_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1804 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_21_1618 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[18\]_A la_iena_mprj[18] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_256 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_903 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_936 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_914 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_925 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1524 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1513 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1502 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_969 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_958 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_947 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1557 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1546 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1535 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_495 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1579 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1568 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1157 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[90\] _358_/Y mprj_logic_high_inst/HI[292] vssd vssd vccd
+ vccd la_oenb_core[90] sky130_fd_sc_hd__einvp_8
XFILLER_3_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_2004 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[3\] la_iena_mprj[3] mprj_logic_high_inst/HI[333] vssd vssd
+ vccd vccd user_to_mprj_in_gates\[3\]/B sky130_fd_sc_hd__and2_1
XFILLER_4_2037 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[98\] _569_/Y la_buf\[98\]/TE vssd vssd vccd vccd la_data_in_core[98] sky130_fd_sc_hd__einvp_8
XFILLER_46_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__587__A la_data_out_mprj[116] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xla_buf_enable\[113\] la_oenb_mprj[113] la_buf_enable\[113\]/B vssd vssd vccd vccd
+ la_buf\[113\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_18_201 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_46_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_234 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_705 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_15_941 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_15_952 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_771 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_922 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_417_ mprj_adr_o_core[10] vssd vssd vccd vccd _417_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1360 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_348_ la_oenb_mprj[80] vssd vssd vccd vccd _348_/Y sky130_fd_sc_hd__inv_2
XFILLER_35_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1809 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf\[110\]_A _581_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1765 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_45_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[74\]_A user_to_mprj_in_gates\[74\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_9_1214 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[87\] la_data_out_core[87] user_to_mprj_in_gates\[87\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[87\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_42_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1269 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__497__A la_data_out_mprj[26] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_mprj_adr_buf\[24\]_TE mprj_adr_buf\[24\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_20_1673 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_20_465 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1780 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[101\]_A _572_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_43_1106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_808 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_5_1601 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_28_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_543 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1923 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_700 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_711 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_34_1809 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[1\] user_to_mprj_in_gates\[1\]/Y vssd vssd vccd vccd la_data_in_mprj[1]
+ sky130_fd_sc_hd__inv_8
XPHY_744 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_722 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_733 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1332 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1321 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1310 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_766 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_755 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_777 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_933 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_1365 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1354 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1343 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_788 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_799 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1376 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1398 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1387 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_23_95 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xla_buf\[9\] _480_/Y la_buf\[9\]/TE vssd vssd vccd vccd la_data_in_core[9] sky130_fd_sc_hd__einvp_8
Xla_buf\[13\] _484_/Y la_buf\[13\]/TE vssd vssd vccd vccd la_data_in_core[13] sky130_fd_sc_hd__einvp_8
XFILLER_7_469 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[56\]_A user_to_mprj_in_gates\[56\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_10_1864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_3_697 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_adr_buf\[6\] _413_/Y mprj_adr_buf\[6\]/TE vssd vssd vccd vccd mprj_adr_o_user[6]
+ sky130_fd_sc_hd__einvp_8
XFILLER_4_1122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_510 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_46_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1155 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2112 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_587 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_88 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[57\] user_to_mprj_in_gates\[57\]/Y vssd vssd vccd vccd la_data_in_mprj[57]
+ sky130_fd_sc_hd__inv_8
XANTENNA_la_buf\[96\]_A _567_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_34_579 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_229 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_30_796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA_user_to_mprj_in_buffers\[47\]_A user_to_mprj_in_gates\[47\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_48_1562 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_9_1055 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_in_gates\[113\] la_data_out_core[113] user_to_mprj_in_gates\[113\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[113\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_42_1161 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_852 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[18\]_TE la_buf\[18\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_38_885 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[110\]_B mprj_logic_high_inst/HI[440] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XANTENNA_la_buf\[87\]_A _558_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_33_1842 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[97\] la_iena_mprj[97] mprj_logic_high_inst/HI[427] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[97\]/B sky130_fd_sc_hd__and2_1
XANTENNA_user_to_mprj_in_buffers\[38\]_A user_to_mprj_in_gates\[38\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_oen_buffers\[123\] _391_/Y mprj_logic_high_inst/HI[325] vssd vssd vccd
+ vccd la_oenb_core[123] sky130_fd_sc_hd__einvp_8
XFILLER_5_2110 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
Xuser_to_mprj_oen_buffers\[53\] _652_/Y mprj_logic_high_inst/HI[255] vssd vssd vccd
+ vccd la_oenb_core[53] sky130_fd_sc_hd__einvp_8
XFILLER_47_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[75\] la_oenb_mprj[75] la_buf_enable\[75\]/B vssd vssd vccd vccd la_buf\[75\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_28_351 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_18_62 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_43_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_384 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_16_502 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_16_524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1731 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_505 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_38_1764 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1617 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XPHY_530 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_541 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_730 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_552 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1797 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1140 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_574 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[96\]_B la_buf_enable\[96\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_585 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_596 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_563 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1184 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1151 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1173 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1341 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1162 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1195 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_767 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_7_277 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
Xla_buf\[117\] _588_/Y la_buf\[117\]/TE vssd vssd vccd vccd la_data_in_core[117] sky130_fd_sc_hd__einvp_8
XANTENNA_user_to_mprj_in_buffers\[29\]_A user_to_mprj_in_gates\[29\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_995 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[110\] user_to_mprj_in_gates\[110\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[110] sky130_fd_sc_hd__inv_8
XFILLER_45_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[20\]_B la_buf_enable\[20\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_1239 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_340 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_35_811 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[69\]_A _540_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_1_1873 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_538 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_la_buf_enable\[120\]_A_N la_oenb_mprj[120] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_15_1550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_1458 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_48_2060 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_39 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_1944 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[11\]_B la_buf_enable\[11\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_115 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1740 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_619 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_2_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_6_1795 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_37_192 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_825 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_2095 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
Xuser_to_mprj_in_ena_buf\[12\] la_iena_mprj[12] mprj_logic_high_inst/HI[342] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[12\]/B sky130_fd_sc_hd__and2_1
XFILLER_25_387 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_9_509 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XANTENNA_la_buf_enable\[78\]_B la_buf_enable\[78\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_21_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_225 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_1_921 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_48_402 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_7_1526 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_29_50 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
Xla_buf\[80\] _551_/Y la_buf\[80\]/TE vssd vssd vccd vccd la_data_in_core[80] sky130_fd_sc_hd__einvp_8
XFILLER_29_83 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__595__A la_data_out_mprj[124] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA_user_to_mprj_in_ena_buf\[81\]_B mprj_logic_high_inst/HI[411] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_16_310 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_596_ la_data_out_mprj[125] vssd vssd vccd vccd _596_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_343 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_2137 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_360 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_la_buf_enable\[69\]_B la_buf_enable\[69\]/B vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_393 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_371 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_382 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_571 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_564 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1182 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1756 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[71\]_A _339_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_54 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_87 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_2108 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_45_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_424 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1047 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1303 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_ena_buf\[72\]_B mprj_logic_high_inst/HI[402] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_39_1336 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_652 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_22_368 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_880 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_390 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1992 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1834 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_24_1605 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1796 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1857 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1930 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_44_1097 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_1649 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1963 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1996 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_129 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_ena_buf\[63\]_B mprj_logic_high_inst/HI[393] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
X_450_ mprj_dat_o_core[11] vssd vssd vccd vccd _450_/Y sky130_fd_sc_hd__inv_2
XFILLER_25_151 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_381_ la_oenb_mprj[113] vssd vssd vccd vccd _381_/Y sky130_fd_sc_hd__inv_2
XFILLER_13_302 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[38\] la_oenb_mprj[38] la_buf_enable\[38\]/B vssd vssd vccd vccd la_buf\[38\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_25_184 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[16\] _615_/Y mprj_logic_high_inst/HI[218] vssd vssd vccd
+ vccd la_oenb_core[16] sky130_fd_sc_hd__einvp_8
XFILLER_35_1723 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1609 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_84 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_1080 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_45_961 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_600 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_648_ la_oenb_mprj[49] vssd vssd vccd vccd _648_/Y sky130_fd_sc_hd__inv_2
XFILLER_45_994 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_579_ la_data_out_mprj[108] vssd vssd vccd vccd _579_/Y sky130_fd_sc_hd__inv_2
XPHY_190 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_361 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_884 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1597 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_25_1903 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1109 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_25_1925 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_25_1947 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1732 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_298 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_23_1671 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_42_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1706 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_39_1177 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1717 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1728 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1739 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_11_839 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA_user_to_mprj_oen_buffers\[13\]_TE mprj_logic_high_inst/HI[215] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_1328 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1104 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_46_1137 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_2125 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1654 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_714 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_416 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_34_909 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_18_427 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_33_408 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_502_ la_data_out_mprj[31] vssd vssd vccd vccd _502_/Y sky130_fd_sc_hd__inv_2
X_433_ mprj_adr_o_core[26] vssd vssd vccd vccd _433_/Y sky130_fd_sc_hd__inv_2
XFILLER_42_942 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_14_644 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_986 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1531 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_364_ la_oenb_mprj[96] vssd vssd vccd vccd _364_/Y sky130_fd_sc_hd__inv_2
Xla_buf\[43\] _514_/Y la_buf\[43\]/TE vssd vssd vccd vccd la_data_in_core[43] sky130_fd_sc_hd__einvp_8
XFILLER_35_1575 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[115\] la_iena_mprj[115] mprj_logic_high_inst/HI[445] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[115\]/B sky130_fd_sc_hd__and2_1
XFILLER_35_1597 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_6_810 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_1524 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[87\] user_to_mprj_in_gates\[87\]/Y vssd vssd vccd vccd la_data_in_mprj[87]
+ sky130_fd_sc_hd__inv_8
XANTENNA_mprj_adr_buf\[22\]_A _429_/Y vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_213 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_3_1039 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[51\]_TE la_buf\[51\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_1927 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_24_408 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[32\] la_data_out_core[32] user_to_mprj_in_gates\[32\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[32\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_17_460 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_32_441 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[36\]_TE mprj_logic_high_inst/HI[238] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1339 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_la_buf_enable\[93\]_A_N la_oenb_mprj[93] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_18_1773 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_636 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_31_1951 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_34_1096 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_692 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf_enable\[31\]_A_N la_oenb_mprj[31] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_1744 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1816 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_1766 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_1849 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1540 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf_enable\[46\]_A_N la_oenb_mprj[46] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_27_268 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_904 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_915 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_926 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1514 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1503 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_959 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_948 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_937 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1525 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1558 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1547 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1536 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_607 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_11_647 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1569 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1726 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_13_1136 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_1169 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_835 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[83\] _351_/Y mprj_logic_high_inst/HI[285] vssd vssd vccd
+ vccd la_oenb_core[83] sky130_fd_sc_hd__einvp_8
Xmprj_dat_buf\[31\] _470_/Y mprj_dat_buf\[31\]/TE vssd vssd vccd vccd mprj_dat_o_user[31]
+ sky130_fd_sc_hd__einvp_8
XFILLER_3_868 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_2130 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_378 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_1451 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_2016 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_la_buf\[74\]_TE la_buf\[74\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_46_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1337 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xla_buf_enable\[106\] la_oenb_mprj[106] la_buf_enable\[106\]/B vssd vssd vccd vccd
+ la_buf\[106\]/TE sky130_fd_sc_hd__and2b_1
XFILLER_46_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_18_246 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_37_1626 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_249 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_964 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_42_783 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_416_ mprj_adr_o_core[9] vssd vssd vccd vccd _416_/Y sky130_fd_sc_hd__inv_2
X_347_ la_oenb_mprj[79] vssd vssd vccd vccd _347_/Y sky130_fd_sc_hd__inv_2
XFILLER_30_989 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_30_978 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_1670 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_172 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1799 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_9_1226 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_42_1332 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_42_1398 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_1685 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1746 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_mprj_dat_buf\[23\]_TE mprj_dat_buf\[23\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_36_1103 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_32_293 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_oen_buffers\[2\]_TE mprj_logic_high_inst/HI[204] vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
XFILLER_14_1456 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_20_488 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_20_499 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_1792 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1210 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_43_1118 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_522 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_5_1668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_28_555 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_ena_buf\[42\] la_iena_mprj[42] mprj_logic_high_inst/HI[372] vssd
+ vssd vccd vccd user_to_mprj_in_gates\[42\]/B sky130_fd_sc_hd__and2_1
XFILLER_43_514 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_1381 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1935 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1902 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XPHY_701 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_38_1968 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_745 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_712 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_723 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_734 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1300 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1333 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1322 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1311 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
Xla_buf_enable\[20\] la_oenb_mprj[20] la_buf_enable\[20\]/B vssd vssd vccd vccd la_buf\[20\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_11_433 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_767 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_756 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_778 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_956 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_23_282 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_1366 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1355 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1344 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1512 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_789 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1377 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1399 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1388 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1556 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_448 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_11_477 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1906 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_3_676 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_45_1939 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA__598__A la_data_out_mprj[127] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_4_1134 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_1167 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_46_363 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_4_1178 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_4_1189 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_19_599 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_396 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_2124 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_15_750 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_208 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_42_591 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_31_1022 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_31_1088 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_2106 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_2139 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_48_1596 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_26_1850 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1911 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_864 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_37_330 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[106\] la_data_out_core[106] user_to_mprj_in_gates\[106\]/B
+ vssd vssd vccd vccd user_to_mprj_in_gates\[106\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_38_897 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1521 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_33_1854 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_407 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_14_1264 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_429 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_1051 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[116\] _384_/Y mprj_logic_high_inst/HI[318] vssd vssd vccd
+ vccd la_oenb_core[116] sky130_fd_sc_hd__einvp_8
XFILLER_47_1084 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_668 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_5_2122 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_639 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_47_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_2008 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_oen_buffers\[46\] _645_/Y mprj_logic_high_inst/HI[248] vssd vssd vccd
+ vccd la_oenb_core[46] sky130_fd_sc_hd__einvp_8
XFILLER_18_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf_enable\[68\] la_oenb_mprj[68] la_buf_enable\[68\]/B vssd vssd vccd vccd la_buf\[68\]/TE
+ sky130_fd_sc_hd__and2b_1
XFILLER_18_85 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_43_322 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_16_536 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_43_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_38_1776 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_520 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_531 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_542 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_553 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1141 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1130 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_575 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_12_742 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_586 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_15_1028 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_564 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1152 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1174 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1320 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1163 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_7_223 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_597 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_1185 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_32_1353 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XPHY_1196 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA_mprj_adr_buf\[14\]_TE mprj_adr_buf\[14\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_1747 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_628 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_buffers\[103\] user_to_mprj_in_gates\[103\]/Y vssd vssd vccd vccd
+ la_data_in_mprj[103] sky130_fd_sc_hd__inv_8
XFILLER_35_823 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1507 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_856 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_2072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1901 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_28_1956 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_1393 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xmprj_dat_buf\[2\] _441_/Y mprj_dat_buf\[2\]/TE vssd vssd vccd vccd mprj_dat_o_user[2]
+ sky130_fd_sc_hd__einvp_8
XANTENNA_mprj_dat_buf\[2\]_TE mprj_dat_buf\[2\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_29_127 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1511 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_1752 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_22_1533 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_2_1638 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_1373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_41_837 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_la_buf\[122\]_TE la_buf\[122\]/TE vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_528 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_21_550 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_21_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_5_705 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_14_1072 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_237 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_0_476 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_7_1538 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_95 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xla_buf\[73\] _544_/Y la_buf\[73\]/TE vssd vssd vccd vccd la_data_in_core[73] sky130_fd_sc_hd__einvp_8
XFILLER_16_355 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_595_ la_data_out_mprj[124] vssd vssd vccd vccd _595_/Y sky130_fd_sc_hd__inv_2
XFILLER_16_388 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_369 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_361 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_350 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_394 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_372 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_383 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_543 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_12_583 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_8_576 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_12_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_1194 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[70\]_A la_data_out_core[70] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_6_66 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_12_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_6_99 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_4_771 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_3_270 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_1588 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_20_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_436 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
Xuser_to_mprj_in_gates\[62\] la_data_out_core[62] user_to_mprj_in_gates\[62\]/B vssd
+ vssd vccd vccd user_to_mprj_in_gates\[62\]/Y sky130_fd_sc_hd__nand2_4
XFILLER_48_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_620 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_35_664 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_1348 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_17_1646 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_31_892 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_30_1846 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XANTENNA_user_to_mprj_in_gates\[61\]_A la_data_out_core[61] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_11_1289 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_46_1308 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_1_229 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_48_1190 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_44_1010 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_1803 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_44_1054 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_24_1617 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_8_1869 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_1975 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_39_970 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_41_601 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
XFILLER_13_314 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_380_ la_oenb_mprj[112] vssd vssd vccd vccd _380_/Y sky130_fd_sc_hd__inv_2
XANTENNA_user_to_mprj_oen_buffers\[92\]_TE mprj_logic_high_inst/HI[294] vssd vssd
+ vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_25_163 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_39_1882 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_144 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_40_111 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1702 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_25_196 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_35_1735 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_35_1768 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_33_1481 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_29_1506 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_31_96 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_gates\[52\]_A la_data_out_core[52] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_0_262 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_48_233 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_647_ la_oenb_mprj[48] vssd vssd vccd vccd _647_/Y sky130_fd_sc_hd__inv_2
XFILLER_2_1980 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_32_612 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_578_ la_data_out_mprj[107] vssd vssd vccd vccd _578_/Y sky130_fd_sc_hd__inv_2
XFILLER_38_2082 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XANTENNA_user_to_mprj_in_buffers\[2\]_A user_to_mprj_in_gates\[2\]/Y vssd vssd vccd
+ vccd sky130_fd_sc_hd__diode_2
Xuser_to_mprj_in_buffers\[32\] user_to_mprj_in_gates\[32\]/Y vssd vssd vccd vccd la_data_in_mprj[32]
+ sky130_fd_sc_hd__inv_8
XPHY_180 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_191 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_8_373 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XFILLER_8_340 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
XFILLER_9_896 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_8_384 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_user_to_mprj_in_gates\[43\]_A la_data_out_core[43] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_45_2020 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
XFILLER_45_2053 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
.ends

