magic
tech sky130A
timestamp 1605923309
<< pwell >>
rect -2723 -1549 2723 1549
<< psubdiff >>
rect -2705 1514 -2657 1531
rect 2657 1514 2705 1531
rect -2705 1483 -2688 1514
rect 2688 1483 2705 1514
rect -2705 -1514 -2688 -1483
rect 2688 -1514 2705 -1483
rect -2705 -1531 -2657 -1514
rect 2657 -1531 2705 -1514
<< psubdiffcont >>
rect -2657 1514 2657 1531
rect -2705 -1483 -2688 1483
rect 2688 -1483 2705 1483
rect -2657 -1531 2657 -1514
<< xpolycontact >>
rect -2640 1250 -2571 1466
rect -2640 -1466 -2571 -1250
rect -2447 1250 -2378 1466
rect -2447 -1466 -2378 -1250
rect -2254 1250 -2185 1466
rect -2254 -1466 -2185 -1250
rect -2061 1250 -1992 1466
rect -2061 -1466 -1992 -1250
rect -1868 1250 -1799 1466
rect -1868 -1466 -1799 -1250
rect -1675 1250 -1606 1466
rect -1675 -1466 -1606 -1250
rect -1482 1250 -1413 1466
rect -1482 -1466 -1413 -1250
rect -1289 1250 -1220 1466
rect -1289 -1466 -1220 -1250
rect -1096 1250 -1027 1466
rect -1096 -1466 -1027 -1250
rect -903 1250 -834 1466
rect -903 -1466 -834 -1250
rect -710 1250 -641 1466
rect -710 -1466 -641 -1250
rect -517 1250 -448 1466
rect -517 -1466 -448 -1250
rect -324 1250 -255 1466
rect -324 -1466 -255 -1250
rect -131 1250 -62 1466
rect -131 -1466 -62 -1250
rect 62 1250 131 1466
rect 62 -1466 131 -1250
rect 255 1250 324 1466
rect 255 -1466 324 -1250
rect 448 1250 517 1466
rect 448 -1466 517 -1250
rect 641 1250 710 1466
rect 641 -1466 710 -1250
rect 834 1250 903 1466
rect 834 -1466 903 -1250
rect 1027 1250 1096 1466
rect 1027 -1466 1096 -1250
rect 1220 1250 1289 1466
rect 1220 -1466 1289 -1250
rect 1413 1250 1482 1466
rect 1413 -1466 1482 -1250
rect 1606 1250 1675 1466
rect 1606 -1466 1675 -1250
rect 1799 1250 1868 1466
rect 1799 -1466 1868 -1250
rect 1992 1250 2061 1466
rect 1992 -1466 2061 -1250
rect 2185 1250 2254 1466
rect 2185 -1466 2254 -1250
rect 2378 1250 2447 1466
rect 2378 -1466 2447 -1250
rect 2571 1250 2640 1466
rect 2571 -1466 2640 -1250
<< xpolyres >>
rect -2640 -1250 -2571 1250
rect -2447 -1250 -2378 1250
rect -2254 -1250 -2185 1250
rect -2061 -1250 -1992 1250
rect -1868 -1250 -1799 1250
rect -1675 -1250 -1606 1250
rect -1482 -1250 -1413 1250
rect -1289 -1250 -1220 1250
rect -1096 -1250 -1027 1250
rect -903 -1250 -834 1250
rect -710 -1250 -641 1250
rect -517 -1250 -448 1250
rect -324 -1250 -255 1250
rect -131 -1250 -62 1250
rect 62 -1250 131 1250
rect 255 -1250 324 1250
rect 448 -1250 517 1250
rect 641 -1250 710 1250
rect 834 -1250 903 1250
rect 1027 -1250 1096 1250
rect 1220 -1250 1289 1250
rect 1413 -1250 1482 1250
rect 1606 -1250 1675 1250
rect 1799 -1250 1868 1250
rect 1992 -1250 2061 1250
rect 2185 -1250 2254 1250
rect 2378 -1250 2447 1250
rect 2571 -1250 2640 1250
<< locali >>
rect -2705 1514 -2657 1531
rect 2657 1514 2705 1531
rect -2705 1483 -2688 1514
rect 2688 1483 2705 1514
rect -2705 -1514 -2688 -1483
rect 2688 -1514 2705 -1483
rect -2705 -1531 -2657 -1514
rect 2657 -1531 2705 -1514
<< res0p69 >>
rect -2641 -1251 -2570 1251
rect -2448 -1251 -2377 1251
rect -2255 -1251 -2184 1251
rect -2062 -1251 -1991 1251
rect -1869 -1251 -1798 1251
rect -1676 -1251 -1605 1251
rect -1483 -1251 -1412 1251
rect -1290 -1251 -1219 1251
rect -1097 -1251 -1026 1251
rect -904 -1251 -833 1251
rect -711 -1251 -640 1251
rect -518 -1251 -447 1251
rect -325 -1251 -254 1251
rect -132 -1251 -61 1251
rect 61 -1251 132 1251
rect 254 -1251 325 1251
rect 447 -1251 518 1251
rect 640 -1251 711 1251
rect 833 -1251 904 1251
rect 1026 -1251 1097 1251
rect 1219 -1251 1290 1251
rect 1412 -1251 1483 1251
rect 1605 -1251 1676 1251
rect 1798 -1251 1869 1251
rect 1991 -1251 2062 1251
rect 2184 -1251 2255 1251
rect 2377 -1251 2448 1251
rect 2570 -1251 2641 1251
<< properties >>
string gencell sky130_fd_pr__res_xhigh_po_0p69
string FIXED_BBOX -2696 -1522 2696 1522
string parameters w 0.69 l 25.0 m 1 nx 28 wmin 0.690 lmin 0.50 rho 2000 val 72.811k dummy 0 dw 0.0 term 120 sterm 0.0 caplen 0 wmax 0.690 guard 1 glc 1 grc 1 gtc 1 gbc 1 compatible {sky130_fd_pr__res_xhigh_po_0p35  sky130_fd_pr__res_xhigh_po_0p69 sky130_fd_pr__res_xhigh_po_1p41  sky130_fd_pr__res_xhigh_po_2p85 sky130_fd_pr__res_xhigh_po_5p73} full_metal 1
string library sky130
<< end >>
