magic
tech sky130A
timestamp 1618942412
<< metal2 >>
rect 4043 351760 4099 352480
rect 12139 351760 12195 352480
rect 20235 351760 20291 352480
rect 28377 351760 28433 352480
rect 36473 351760 36529 352480
rect 44569 351760 44625 352480
rect 52711 351760 52767 352480
rect 60807 351760 60863 352480
rect 68903 351760 68959 352480
rect 77045 351760 77101 352480
rect 85141 351760 85197 352480
rect 93237 351760 93293 352480
rect 101379 351760 101435 352480
rect 109475 351760 109531 352480
rect 117571 351760 117627 352480
rect 125713 351760 125769 352480
rect 133809 351760 133865 352480
rect 141905 351760 141961 352480
rect 150047 351760 150103 352480
rect 158143 351760 158199 352480
rect 166239 351760 166295 352480
rect 174381 351760 174437 352480
rect 182477 351760 182533 352480
rect 190573 351760 190629 352480
rect 198715 351760 198771 352480
rect 206811 351760 206867 352480
rect 214907 351760 214963 352480
rect 223049 351760 223105 352480
rect 231145 351760 231201 352480
rect 239241 351760 239297 352480
rect 247383 351760 247439 352480
rect 255479 351760 255535 352480
rect 263575 351760 263631 352480
rect 271717 351760 271773 352480
rect 279813 351760 279869 352480
rect 287909 351760 287965 352480
rect 271 -480 327 240
rect 823 -480 879 240
rect 1421 -480 1477 240
rect 2019 -480 2075 240
rect 2617 -480 2673 240
rect 3215 -480 3271 240
rect 3813 -480 3869 240
rect 4411 -480 4467 240
rect 5009 -480 5065 240
rect 5607 -480 5663 240
rect 6205 -480 6261 240
rect 6803 -480 6859 240
rect 7401 -480 7457 240
rect 7999 -480 8055 240
rect 8597 -480 8653 240
rect 9149 -480 9205 240
rect 9747 -480 9803 240
rect 10345 -480 10401 240
rect 10943 -480 10999 240
rect 11541 -480 11597 240
rect 12139 -480 12195 240
rect 12737 -480 12793 240
rect 13335 -480 13391 240
rect 13933 -480 13989 240
rect 14531 -480 14587 240
rect 15129 -480 15185 240
rect 15727 -480 15783 240
rect 16325 -480 16381 240
rect 16923 -480 16979 240
rect 17475 -480 17531 240
rect 18073 -480 18129 240
rect 18671 -480 18727 240
rect 19269 -480 19325 240
rect 19867 -480 19923 240
rect 20465 -480 20521 240
rect 21063 -480 21119 240
rect 21661 -480 21717 240
rect 22259 -480 22315 240
rect 22857 -480 22913 240
rect 23455 -480 23511 240
rect 24053 -480 24109 240
rect 24651 -480 24707 240
rect 25249 -480 25305 240
rect 25801 -480 25857 240
rect 26399 -480 26455 240
rect 26997 -480 27053 240
rect 27595 -480 27651 240
rect 28193 -480 28249 240
rect 28791 -480 28847 240
rect 29389 -480 29445 240
rect 29987 -480 30043 240
rect 30585 -480 30641 240
rect 31183 -480 31239 240
rect 31781 -480 31837 240
rect 32379 -480 32435 240
rect 32977 -480 33033 240
rect 33575 -480 33631 240
rect 34127 -480 34183 240
rect 34725 -480 34781 240
rect 35323 -480 35379 240
rect 35921 -480 35977 240
rect 36519 -480 36575 240
rect 37117 -480 37173 240
rect 37715 -480 37771 240
rect 38313 -480 38369 240
rect 38911 -480 38967 240
rect 39509 -480 39565 240
rect 40107 -480 40163 240
rect 40705 -480 40761 240
rect 41303 -480 41359 240
rect 41901 -480 41957 240
rect 42453 -480 42509 240
rect 43051 -480 43107 240
rect 43649 -480 43705 240
rect 44247 -480 44303 240
rect 44845 -480 44901 240
rect 45443 -480 45499 240
rect 46041 -480 46097 240
rect 46639 -480 46695 240
rect 47237 -480 47293 240
rect 47835 -480 47891 240
rect 48433 -480 48489 240
rect 49031 -480 49087 240
rect 49629 -480 49685 240
rect 50227 -480 50283 240
rect 50779 -480 50835 240
rect 51377 -480 51433 240
rect 51975 -480 52031 240
rect 52573 -480 52629 240
rect 53171 -480 53227 240
rect 53769 -480 53825 240
rect 54367 -480 54423 240
rect 54965 -480 55021 240
rect 55563 -480 55619 240
rect 56161 -480 56217 240
rect 56759 -480 56815 240
rect 57357 -480 57413 240
rect 57955 -480 58011 240
rect 58553 -480 58609 240
rect 59105 -480 59161 240
rect 59703 -480 59759 240
rect 60301 -480 60357 240
rect 60899 -480 60955 240
rect 61497 -480 61553 240
rect 62095 -480 62151 240
rect 62693 -480 62749 240
rect 63291 -480 63347 240
rect 63889 -480 63945 240
rect 64487 -480 64543 240
rect 65085 -480 65141 240
rect 65683 -480 65739 240
rect 66281 -480 66337 240
rect 66879 -480 66935 240
rect 67431 -480 67487 240
rect 68029 -480 68085 240
rect 68627 -480 68683 240
rect 69225 -480 69281 240
rect 69823 -480 69879 240
rect 70421 -480 70477 240
rect 71019 -480 71075 240
rect 71617 -480 71673 240
rect 72215 -480 72271 240
rect 72813 -480 72869 240
rect 73411 -480 73467 240
rect 74009 -480 74065 240
rect 74607 -480 74663 240
rect 75205 -480 75261 240
rect 75757 -480 75813 240
rect 76355 -480 76411 240
rect 76953 -480 77009 240
rect 77551 -480 77607 240
rect 78149 -480 78205 240
rect 78747 -480 78803 240
rect 79345 -480 79401 240
rect 79943 -480 79999 240
rect 80541 -480 80597 240
rect 81139 -480 81195 240
rect 81737 -480 81793 240
rect 82335 -480 82391 240
rect 82933 -480 82989 240
rect 83531 -480 83587 240
rect 84083 -480 84139 240
rect 84681 -480 84737 240
rect 85279 -480 85335 240
rect 85877 -480 85933 240
rect 86475 -480 86531 240
rect 87073 -480 87129 240
rect 87671 -480 87727 240
rect 88269 -480 88325 240
rect 88867 -480 88923 240
rect 89465 -480 89521 240
rect 90063 -480 90119 240
rect 90661 -480 90717 240
rect 91259 -480 91315 240
rect 91857 -480 91913 240
rect 92409 -480 92465 240
rect 93007 -480 93063 240
rect 93605 -480 93661 240
rect 94203 -480 94259 240
rect 94801 -480 94857 240
rect 95399 -480 95455 240
rect 95997 -480 96053 240
rect 96595 -480 96651 240
rect 97193 -480 97249 240
rect 97791 -480 97847 240
rect 98389 -480 98445 240
rect 98987 -480 99043 240
rect 99585 -480 99641 240
rect 100183 -480 100239 240
rect 100735 -480 100791 240
rect 101333 -480 101389 240
rect 101931 -480 101987 240
rect 102529 -480 102585 240
rect 103127 -480 103183 240
rect 103725 -480 103781 240
rect 104323 -480 104379 240
rect 104921 -480 104977 240
rect 105519 -480 105575 240
rect 106117 -480 106173 240
rect 106715 -480 106771 240
rect 107313 -480 107369 240
rect 107911 -480 107967 240
rect 108509 -480 108565 240
rect 109061 -480 109117 240
rect 109659 -480 109715 240
rect 110257 -480 110313 240
rect 110855 -480 110911 240
rect 111453 -480 111509 240
rect 112051 -480 112107 240
rect 112649 -480 112705 240
rect 113247 -480 113303 240
rect 113845 -480 113901 240
rect 114443 -480 114499 240
rect 115041 -480 115097 240
rect 115639 -480 115695 240
rect 116237 -480 116293 240
rect 116835 -480 116891 240
rect 117387 -480 117443 240
rect 117985 -480 118041 240
rect 118583 -480 118639 240
rect 119181 -480 119237 240
rect 119779 -480 119835 240
rect 120377 -480 120433 240
rect 120975 -480 121031 240
rect 121573 -480 121629 240
rect 122171 -480 122227 240
rect 122769 -480 122825 240
rect 123367 -480 123423 240
rect 123965 -480 124021 240
rect 124563 -480 124619 240
rect 125161 -480 125217 240
rect 125713 -480 125769 240
rect 126311 -480 126367 240
rect 126909 -480 126965 240
rect 127507 -480 127563 240
rect 128105 -480 128161 240
rect 128703 -480 128759 240
rect 129301 -480 129357 240
rect 129899 -480 129955 240
rect 130497 -480 130553 240
rect 131095 -480 131151 240
rect 131693 -480 131749 240
rect 132291 -480 132347 240
rect 132889 -480 132945 240
rect 133487 -480 133543 240
rect 134039 -480 134095 240
rect 134637 -480 134693 240
rect 135235 -480 135291 240
rect 135833 -480 135889 240
rect 136431 -480 136487 240
rect 137029 -480 137085 240
rect 137627 -480 137683 240
rect 138225 -480 138281 240
rect 138823 -480 138879 240
rect 139421 -480 139477 240
rect 140019 -480 140075 240
rect 140617 -480 140673 240
rect 141215 -480 141271 240
rect 141813 -480 141869 240
rect 142365 -480 142421 240
rect 142963 -480 143019 240
rect 143561 -480 143617 240
rect 144159 -480 144215 240
rect 144757 -480 144813 240
rect 145355 -480 145411 240
rect 145953 -480 146009 240
rect 146551 -480 146607 240
rect 147149 -480 147205 240
rect 147747 -480 147803 240
rect 148345 -480 148401 240
rect 148943 -480 148999 240
rect 149541 -480 149597 240
rect 150139 -480 150195 240
rect 150691 -480 150747 240
rect 151289 -480 151345 240
rect 151887 -480 151943 240
rect 152485 -480 152541 240
rect 153083 -480 153139 240
rect 153681 -480 153737 240
rect 154279 -480 154335 240
rect 154877 -480 154933 240
rect 155475 -480 155531 240
rect 156073 -480 156129 240
rect 156671 -480 156727 240
rect 157269 -480 157325 240
rect 157867 -480 157923 240
rect 158465 -480 158521 240
rect 159017 -480 159073 240
rect 159615 -480 159671 240
rect 160213 -480 160269 240
rect 160811 -480 160867 240
rect 161409 -480 161465 240
rect 162007 -480 162063 240
rect 162605 -480 162661 240
rect 163203 -480 163259 240
rect 163801 -480 163857 240
rect 164399 -480 164455 240
rect 164997 -480 165053 240
rect 165595 -480 165651 240
rect 166193 -480 166249 240
rect 166791 -480 166847 240
rect 167343 -480 167399 240
rect 167941 -480 167997 240
rect 168539 -480 168595 240
rect 169137 -480 169193 240
rect 169735 -480 169791 240
rect 170333 -480 170389 240
rect 170931 -480 170987 240
rect 171529 -480 171585 240
rect 172127 -480 172183 240
rect 172725 -480 172781 240
rect 173323 -480 173379 240
rect 173921 -480 173977 240
rect 174519 -480 174575 240
rect 175117 -480 175173 240
rect 175669 -480 175725 240
rect 176267 -480 176323 240
rect 176865 -480 176921 240
rect 177463 -480 177519 240
rect 178061 -480 178117 240
rect 178659 -480 178715 240
rect 179257 -480 179313 240
rect 179855 -480 179911 240
rect 180453 -480 180509 240
rect 181051 -480 181107 240
rect 181649 -480 181705 240
rect 182247 -480 182303 240
rect 182845 -480 182901 240
rect 183443 -480 183499 240
rect 183995 -480 184051 240
rect 184593 -480 184649 240
rect 185191 -480 185247 240
rect 185789 -480 185845 240
rect 186387 -480 186443 240
rect 186985 -480 187041 240
rect 187583 -480 187639 240
rect 188181 -480 188237 240
rect 188779 -480 188835 240
rect 189377 -480 189433 240
rect 189975 -480 190031 240
rect 190573 -480 190629 240
rect 191171 -480 191227 240
rect 191769 -480 191825 240
rect 192321 -480 192377 240
rect 192919 -480 192975 240
rect 193517 -480 193573 240
rect 194115 -480 194171 240
rect 194713 -480 194769 240
rect 195311 -480 195367 240
rect 195909 -480 195965 240
rect 196507 -480 196563 240
rect 197105 -480 197161 240
rect 197703 -480 197759 240
rect 198301 -480 198357 240
rect 198899 -480 198955 240
rect 199497 -480 199553 240
rect 200095 -480 200151 240
rect 200647 -480 200703 240
rect 201245 -480 201301 240
rect 201843 -480 201899 240
rect 202441 -480 202497 240
rect 203039 -480 203095 240
rect 203637 -480 203693 240
rect 204235 -480 204291 240
rect 204833 -480 204889 240
rect 205431 -480 205487 240
rect 206029 -480 206085 240
rect 206627 -480 206683 240
rect 207225 -480 207281 240
rect 207823 -480 207879 240
rect 208421 -480 208477 240
rect 208973 -480 209029 240
rect 209571 -480 209627 240
rect 210169 -480 210225 240
rect 210767 -480 210823 240
rect 211365 -480 211421 240
rect 211963 -480 212019 240
rect 212561 -480 212617 240
rect 213159 -480 213215 240
rect 213757 -480 213813 240
rect 214355 -480 214411 240
rect 214953 -480 215009 240
rect 215551 -480 215607 240
rect 216149 -480 216205 240
rect 216747 -480 216803 240
rect 217299 -480 217355 240
rect 217897 -480 217953 240
rect 218495 -480 218551 240
rect 219093 -480 219149 240
rect 219691 -480 219747 240
rect 220289 -480 220345 240
rect 220887 -480 220943 240
rect 221485 -480 221541 240
rect 222083 -480 222139 240
rect 222681 -480 222737 240
rect 223279 -480 223335 240
rect 223877 -480 223933 240
rect 224475 -480 224531 240
rect 225073 -480 225129 240
rect 225625 -480 225681 240
rect 226223 -480 226279 240
rect 226821 -480 226877 240
rect 227419 -480 227475 240
rect 228017 -480 228073 240
rect 228615 -480 228671 240
rect 229213 -480 229269 240
rect 229811 -480 229867 240
rect 230409 -480 230465 240
rect 231007 -480 231063 240
rect 231605 -480 231661 240
rect 232203 -480 232259 240
rect 232801 -480 232857 240
rect 233399 -480 233455 240
rect 233951 -480 234007 240
rect 234549 -480 234605 240
rect 235147 -480 235203 240
rect 235745 -480 235801 240
rect 236343 -480 236399 240
rect 236941 -480 236997 240
rect 237539 -480 237595 240
rect 238137 -480 238193 240
rect 238735 -480 238791 240
rect 239333 -480 239389 240
rect 239931 -480 239987 240
rect 240529 -480 240585 240
rect 241127 -480 241183 240
rect 241725 -480 241781 240
rect 242277 -480 242333 240
rect 242875 -480 242931 240
rect 243473 -480 243529 240
rect 244071 -480 244127 240
rect 244669 -480 244725 240
rect 245267 -480 245323 240
rect 245865 -480 245921 240
rect 246463 -480 246519 240
rect 247061 -480 247117 240
rect 247659 -480 247715 240
rect 248257 -480 248313 240
rect 248855 -480 248911 240
rect 249453 -480 249509 240
rect 250051 -480 250107 240
rect 250603 -480 250659 240
rect 251201 -480 251257 240
rect 251799 -480 251855 240
rect 252397 -480 252453 240
rect 252995 -480 253051 240
rect 253593 -480 253649 240
rect 254191 -480 254247 240
rect 254789 -480 254845 240
rect 255387 -480 255443 240
rect 255985 -480 256041 240
rect 256583 -480 256639 240
rect 257181 -480 257237 240
rect 257779 -480 257835 240
rect 258377 -480 258433 240
rect 258929 -480 258985 240
rect 259527 -480 259583 240
rect 260125 -480 260181 240
rect 260723 -480 260779 240
rect 261321 -480 261377 240
rect 261919 -480 261975 240
rect 262517 -480 262573 240
rect 263115 -480 263171 240
rect 263713 -480 263769 240
rect 264311 -480 264367 240
rect 264909 -480 264965 240
rect 265507 -480 265563 240
rect 266105 -480 266161 240
rect 266703 -480 266759 240
rect 267255 -480 267311 240
rect 267853 -480 267909 240
rect 268451 -480 268507 240
rect 269049 -480 269105 240
rect 269647 -480 269703 240
rect 270245 -480 270301 240
rect 270843 -480 270899 240
rect 271441 -480 271497 240
rect 272039 -480 272095 240
rect 272637 -480 272693 240
rect 273235 -480 273291 240
rect 273833 -480 273889 240
rect 274431 -480 274487 240
rect 275029 -480 275085 240
rect 275581 -480 275637 240
rect 276179 -480 276235 240
rect 276777 -480 276833 240
rect 277375 -480 277431 240
rect 277973 -480 278029 240
rect 278571 -480 278627 240
rect 279169 -480 279225 240
rect 279767 -480 279823 240
rect 280365 -480 280421 240
rect 280963 -480 281019 240
rect 281561 -480 281617 240
rect 282159 -480 282215 240
rect 282757 -480 282813 240
rect 283355 -480 283411 240
rect 283907 -480 283963 240
rect 284505 -480 284561 240
rect 285103 -480 285159 240
rect 285701 -480 285757 240
rect 286299 -480 286355 240
rect 286897 -480 286953 240
rect 287495 -480 287551 240
rect 288093 -480 288149 240
rect 288691 -480 288747 240
rect 289289 -480 289345 240
rect 289887 -480 289943 240
rect 290485 -480 290541 240
rect 291083 -480 291139 240
rect 291681 -480 291737 240
<< metal3 >>
rect 291760 348950 292480 349070
rect -480 348134 240 348254
rect 291760 343102 292480 343222
rect -480 340654 240 340774
rect 291760 337254 292480 337374
rect -480 333174 240 333294
rect 291760 331338 292480 331458
rect -480 325694 240 325814
rect 291760 325490 292480 325610
rect 291760 319642 292480 319762
rect -480 318214 240 318334
rect 291760 313794 292480 313914
rect -480 310734 240 310854
rect 291760 307878 292480 307998
rect -480 303254 240 303374
rect 291760 302030 292480 302150
rect 291760 296182 292480 296302
rect -480 295706 240 295826
rect 291760 290334 292480 290454
rect -480 288226 240 288346
rect 291760 284418 292480 284538
rect -480 280746 240 280866
rect 291760 278570 292480 278690
rect -480 273266 240 273386
rect 291760 272722 292480 272842
rect 291760 266874 292480 266994
rect -480 265786 240 265906
rect 291760 260958 292480 261078
rect -480 258306 240 258426
rect 291760 255110 292480 255230
rect -480 250826 240 250946
rect 291760 249262 292480 249382
rect -480 243346 240 243466
rect 291760 243346 292480 243466
rect 291760 237498 292480 237618
rect -480 235798 240 235918
rect 291760 231650 292480 231770
rect -480 228318 240 228438
rect 291760 225802 292480 225922
rect -480 220838 240 220958
rect 291760 219886 292480 220006
rect 291760 214038 292480 214158
rect -480 213358 240 213478
rect 291760 208190 292480 208310
rect -480 205878 240 205998
rect 291760 202342 292480 202462
rect -480 198398 240 198518
rect 291760 196426 292480 196546
rect -480 190918 240 191038
rect 291760 190578 292480 190698
rect 291760 184730 292480 184850
rect -480 183438 240 183558
rect 291760 178882 292480 179002
rect -480 175890 240 176010
rect 291760 172966 292480 173086
rect -480 168410 240 168530
rect 291760 167118 292480 167238
rect 291760 161270 292480 161390
rect -480 160930 240 161050
rect 291760 155354 292480 155474
rect -480 153450 240 153570
rect 291760 149506 292480 149626
rect -480 145970 240 146090
rect 291760 143658 292480 143778
rect -480 138490 240 138610
rect 291760 137810 292480 137930
rect 291760 131894 292480 132014
rect -480 131010 240 131130
rect 291760 126046 292480 126166
rect -480 123530 240 123650
rect 291760 120198 292480 120318
rect -480 115982 240 116102
rect 291760 114350 292480 114470
rect -480 108502 240 108622
rect 291760 108434 292480 108554
rect 291760 102586 292480 102706
rect -480 101022 240 101142
rect 291760 96738 292480 96858
rect -480 93542 240 93662
rect 291760 90890 292480 91010
rect -480 86062 240 86182
rect 291760 84974 292480 85094
rect 291760 79126 292480 79246
rect -480 78582 240 78702
rect 291760 73278 292480 73398
rect -480 71102 240 71222
rect 291760 67362 292480 67482
rect -480 63622 240 63742
rect 291760 61514 292480 61634
rect -480 56074 240 56194
rect 291760 55666 292480 55786
rect 291760 49818 292480 49938
rect -480 48594 240 48714
rect 291760 43902 292480 44022
rect -480 41114 240 41234
rect 291760 38054 292480 38174
rect -480 33634 240 33754
rect 291760 32206 292480 32326
rect 291760 26358 292480 26478
rect -480 26154 240 26274
rect 291760 20442 292480 20562
rect -480 18674 240 18794
rect 291760 14594 292480 14714
rect -480 11194 240 11314
rect 291760 8746 292480 8866
rect -480 3714 240 3834
rect 291760 2898 292480 3018
<< metal4 >>
rect -4288 355709 -3988 355720
rect -4288 355591 -4197 355709
rect -4079 355591 -3988 355709
rect -4288 355549 -3988 355591
rect -4288 355431 -4197 355549
rect -4079 355431 -3988 355549
rect -4288 340127 -3988 355431
rect -4288 340009 -4197 340127
rect -4079 340009 -3988 340127
rect -4288 339967 -3988 340009
rect -4288 339849 -4197 339967
rect -4079 339849 -3988 339967
rect -4288 322127 -3988 339849
rect -4288 322009 -4197 322127
rect -4079 322009 -3988 322127
rect -4288 321967 -3988 322009
rect -4288 321849 -4197 321967
rect -4079 321849 -3988 321967
rect -4288 304127 -3988 321849
rect -4288 304009 -4197 304127
rect -4079 304009 -3988 304127
rect -4288 303967 -3988 304009
rect -4288 303849 -4197 303967
rect -4079 303849 -3988 303967
rect -4288 286127 -3988 303849
rect -4288 286009 -4197 286127
rect -4079 286009 -3988 286127
rect -4288 285967 -3988 286009
rect -4288 285849 -4197 285967
rect -4079 285849 -3988 285967
rect -4288 268127 -3988 285849
rect -4288 268009 -4197 268127
rect -4079 268009 -3988 268127
rect -4288 267967 -3988 268009
rect -4288 267849 -4197 267967
rect -4079 267849 -3988 267967
rect -4288 250127 -3988 267849
rect -4288 250009 -4197 250127
rect -4079 250009 -3988 250127
rect -4288 249967 -3988 250009
rect -4288 249849 -4197 249967
rect -4079 249849 -3988 249967
rect -4288 232127 -3988 249849
rect -4288 232009 -4197 232127
rect -4079 232009 -3988 232127
rect -4288 231967 -3988 232009
rect -4288 231849 -4197 231967
rect -4079 231849 -3988 231967
rect -4288 214127 -3988 231849
rect -4288 214009 -4197 214127
rect -4079 214009 -3988 214127
rect -4288 213967 -3988 214009
rect -4288 213849 -4197 213967
rect -4079 213849 -3988 213967
rect -4288 196127 -3988 213849
rect -4288 196009 -4197 196127
rect -4079 196009 -3988 196127
rect -4288 195967 -3988 196009
rect -4288 195849 -4197 195967
rect -4079 195849 -3988 195967
rect -4288 178127 -3988 195849
rect -4288 178009 -4197 178127
rect -4079 178009 -3988 178127
rect -4288 177967 -3988 178009
rect -4288 177849 -4197 177967
rect -4079 177849 -3988 177967
rect -4288 160127 -3988 177849
rect -4288 160009 -4197 160127
rect -4079 160009 -3988 160127
rect -4288 159967 -3988 160009
rect -4288 159849 -4197 159967
rect -4079 159849 -3988 159967
rect -4288 142127 -3988 159849
rect -4288 142009 -4197 142127
rect -4079 142009 -3988 142127
rect -4288 141967 -3988 142009
rect -4288 141849 -4197 141967
rect -4079 141849 -3988 141967
rect -4288 124127 -3988 141849
rect -4288 124009 -4197 124127
rect -4079 124009 -3988 124127
rect -4288 123967 -3988 124009
rect -4288 123849 -4197 123967
rect -4079 123849 -3988 123967
rect -4288 106127 -3988 123849
rect -4288 106009 -4197 106127
rect -4079 106009 -3988 106127
rect -4288 105967 -3988 106009
rect -4288 105849 -4197 105967
rect -4079 105849 -3988 105967
rect -4288 88127 -3988 105849
rect -4288 88009 -4197 88127
rect -4079 88009 -3988 88127
rect -4288 87967 -3988 88009
rect -4288 87849 -4197 87967
rect -4079 87849 -3988 87967
rect -4288 70127 -3988 87849
rect -4288 70009 -4197 70127
rect -4079 70009 -3988 70127
rect -4288 69967 -3988 70009
rect -4288 69849 -4197 69967
rect -4079 69849 -3988 69967
rect -4288 52127 -3988 69849
rect -4288 52009 -4197 52127
rect -4079 52009 -3988 52127
rect -4288 51967 -3988 52009
rect -4288 51849 -4197 51967
rect -4079 51849 -3988 51967
rect -4288 34127 -3988 51849
rect -4288 34009 -4197 34127
rect -4079 34009 -3988 34127
rect -4288 33967 -3988 34009
rect -4288 33849 -4197 33967
rect -4079 33849 -3988 33967
rect -4288 16127 -3988 33849
rect -4288 16009 -4197 16127
rect -4079 16009 -3988 16127
rect -4288 15967 -3988 16009
rect -4288 15849 -4197 15967
rect -4079 15849 -3988 15967
rect -4288 -3463 -3988 15849
rect -3818 355239 -3518 355250
rect -3818 355121 -3727 355239
rect -3609 355121 -3518 355239
rect -3818 355079 -3518 355121
rect -3818 354961 -3727 355079
rect -3609 354961 -3518 355079
rect -3818 349127 -3518 354961
rect 6302 355239 6602 355720
rect 6302 355121 6393 355239
rect 6511 355121 6602 355239
rect 6302 355079 6602 355121
rect 6302 354961 6393 355079
rect 6511 354961 6602 355079
rect -3818 349009 -3727 349127
rect -3609 349009 -3518 349127
rect -3818 348967 -3518 349009
rect -3818 348849 -3727 348967
rect -3609 348849 -3518 348967
rect -3818 331127 -3518 348849
rect -3818 331009 -3727 331127
rect -3609 331009 -3518 331127
rect -3818 330967 -3518 331009
rect -3818 330849 -3727 330967
rect -3609 330849 -3518 330967
rect -3818 313127 -3518 330849
rect -3818 313009 -3727 313127
rect -3609 313009 -3518 313127
rect -3818 312967 -3518 313009
rect -3818 312849 -3727 312967
rect -3609 312849 -3518 312967
rect -3818 295127 -3518 312849
rect -3818 295009 -3727 295127
rect -3609 295009 -3518 295127
rect -3818 294967 -3518 295009
rect -3818 294849 -3727 294967
rect -3609 294849 -3518 294967
rect -3818 277127 -3518 294849
rect -3818 277009 -3727 277127
rect -3609 277009 -3518 277127
rect -3818 276967 -3518 277009
rect -3818 276849 -3727 276967
rect -3609 276849 -3518 276967
rect -3818 259127 -3518 276849
rect -3818 259009 -3727 259127
rect -3609 259009 -3518 259127
rect -3818 258967 -3518 259009
rect -3818 258849 -3727 258967
rect -3609 258849 -3518 258967
rect -3818 241127 -3518 258849
rect -3818 241009 -3727 241127
rect -3609 241009 -3518 241127
rect -3818 240967 -3518 241009
rect -3818 240849 -3727 240967
rect -3609 240849 -3518 240967
rect -3818 223127 -3518 240849
rect -3818 223009 -3727 223127
rect -3609 223009 -3518 223127
rect -3818 222967 -3518 223009
rect -3818 222849 -3727 222967
rect -3609 222849 -3518 222967
rect -3818 205127 -3518 222849
rect -3818 205009 -3727 205127
rect -3609 205009 -3518 205127
rect -3818 204967 -3518 205009
rect -3818 204849 -3727 204967
rect -3609 204849 -3518 204967
rect -3818 187127 -3518 204849
rect -3818 187009 -3727 187127
rect -3609 187009 -3518 187127
rect -3818 186967 -3518 187009
rect -3818 186849 -3727 186967
rect -3609 186849 -3518 186967
rect -3818 169127 -3518 186849
rect -3818 169009 -3727 169127
rect -3609 169009 -3518 169127
rect -3818 168967 -3518 169009
rect -3818 168849 -3727 168967
rect -3609 168849 -3518 168967
rect -3818 151127 -3518 168849
rect -3818 151009 -3727 151127
rect -3609 151009 -3518 151127
rect -3818 150967 -3518 151009
rect -3818 150849 -3727 150967
rect -3609 150849 -3518 150967
rect -3818 133127 -3518 150849
rect -3818 133009 -3727 133127
rect -3609 133009 -3518 133127
rect -3818 132967 -3518 133009
rect -3818 132849 -3727 132967
rect -3609 132849 -3518 132967
rect -3818 115127 -3518 132849
rect -3818 115009 -3727 115127
rect -3609 115009 -3518 115127
rect -3818 114967 -3518 115009
rect -3818 114849 -3727 114967
rect -3609 114849 -3518 114967
rect -3818 97127 -3518 114849
rect -3818 97009 -3727 97127
rect -3609 97009 -3518 97127
rect -3818 96967 -3518 97009
rect -3818 96849 -3727 96967
rect -3609 96849 -3518 96967
rect -3818 79127 -3518 96849
rect -3818 79009 -3727 79127
rect -3609 79009 -3518 79127
rect -3818 78967 -3518 79009
rect -3818 78849 -3727 78967
rect -3609 78849 -3518 78967
rect -3818 61127 -3518 78849
rect -3818 61009 -3727 61127
rect -3609 61009 -3518 61127
rect -3818 60967 -3518 61009
rect -3818 60849 -3727 60967
rect -3609 60849 -3518 60967
rect -3818 43127 -3518 60849
rect -3818 43009 -3727 43127
rect -3609 43009 -3518 43127
rect -3818 42967 -3518 43009
rect -3818 42849 -3727 42967
rect -3609 42849 -3518 42967
rect -3818 25127 -3518 42849
rect -3818 25009 -3727 25127
rect -3609 25009 -3518 25127
rect -3818 24967 -3518 25009
rect -3818 24849 -3727 24967
rect -3609 24849 -3518 24967
rect -3818 7127 -3518 24849
rect -3818 7009 -3727 7127
rect -3609 7009 -3518 7127
rect -3818 6967 -3518 7009
rect -3818 6849 -3727 6967
rect -3609 6849 -3518 6967
rect -3818 -2993 -3518 6849
rect -3348 354769 -3048 354780
rect -3348 354651 -3257 354769
rect -3139 354651 -3048 354769
rect -3348 354609 -3048 354651
rect -3348 354491 -3257 354609
rect -3139 354491 -3048 354609
rect -3348 338327 -3048 354491
rect -3348 338209 -3257 338327
rect -3139 338209 -3048 338327
rect -3348 338167 -3048 338209
rect -3348 338049 -3257 338167
rect -3139 338049 -3048 338167
rect -3348 320327 -3048 338049
rect -3348 320209 -3257 320327
rect -3139 320209 -3048 320327
rect -3348 320167 -3048 320209
rect -3348 320049 -3257 320167
rect -3139 320049 -3048 320167
rect -3348 302327 -3048 320049
rect -3348 302209 -3257 302327
rect -3139 302209 -3048 302327
rect -3348 302167 -3048 302209
rect -3348 302049 -3257 302167
rect -3139 302049 -3048 302167
rect -3348 284327 -3048 302049
rect -3348 284209 -3257 284327
rect -3139 284209 -3048 284327
rect -3348 284167 -3048 284209
rect -3348 284049 -3257 284167
rect -3139 284049 -3048 284167
rect -3348 266327 -3048 284049
rect -3348 266209 -3257 266327
rect -3139 266209 -3048 266327
rect -3348 266167 -3048 266209
rect -3348 266049 -3257 266167
rect -3139 266049 -3048 266167
rect -3348 248327 -3048 266049
rect -3348 248209 -3257 248327
rect -3139 248209 -3048 248327
rect -3348 248167 -3048 248209
rect -3348 248049 -3257 248167
rect -3139 248049 -3048 248167
rect -3348 230327 -3048 248049
rect -3348 230209 -3257 230327
rect -3139 230209 -3048 230327
rect -3348 230167 -3048 230209
rect -3348 230049 -3257 230167
rect -3139 230049 -3048 230167
rect -3348 212327 -3048 230049
rect -3348 212209 -3257 212327
rect -3139 212209 -3048 212327
rect -3348 212167 -3048 212209
rect -3348 212049 -3257 212167
rect -3139 212049 -3048 212167
rect -3348 194327 -3048 212049
rect -3348 194209 -3257 194327
rect -3139 194209 -3048 194327
rect -3348 194167 -3048 194209
rect -3348 194049 -3257 194167
rect -3139 194049 -3048 194167
rect -3348 176327 -3048 194049
rect -3348 176209 -3257 176327
rect -3139 176209 -3048 176327
rect -3348 176167 -3048 176209
rect -3348 176049 -3257 176167
rect -3139 176049 -3048 176167
rect -3348 158327 -3048 176049
rect -3348 158209 -3257 158327
rect -3139 158209 -3048 158327
rect -3348 158167 -3048 158209
rect -3348 158049 -3257 158167
rect -3139 158049 -3048 158167
rect -3348 140327 -3048 158049
rect -3348 140209 -3257 140327
rect -3139 140209 -3048 140327
rect -3348 140167 -3048 140209
rect -3348 140049 -3257 140167
rect -3139 140049 -3048 140167
rect -3348 122327 -3048 140049
rect -3348 122209 -3257 122327
rect -3139 122209 -3048 122327
rect -3348 122167 -3048 122209
rect -3348 122049 -3257 122167
rect -3139 122049 -3048 122167
rect -3348 104327 -3048 122049
rect -3348 104209 -3257 104327
rect -3139 104209 -3048 104327
rect -3348 104167 -3048 104209
rect -3348 104049 -3257 104167
rect -3139 104049 -3048 104167
rect -3348 86327 -3048 104049
rect -3348 86209 -3257 86327
rect -3139 86209 -3048 86327
rect -3348 86167 -3048 86209
rect -3348 86049 -3257 86167
rect -3139 86049 -3048 86167
rect -3348 68327 -3048 86049
rect -3348 68209 -3257 68327
rect -3139 68209 -3048 68327
rect -3348 68167 -3048 68209
rect -3348 68049 -3257 68167
rect -3139 68049 -3048 68167
rect -3348 50327 -3048 68049
rect -3348 50209 -3257 50327
rect -3139 50209 -3048 50327
rect -3348 50167 -3048 50209
rect -3348 50049 -3257 50167
rect -3139 50049 -3048 50167
rect -3348 32327 -3048 50049
rect -3348 32209 -3257 32327
rect -3139 32209 -3048 32327
rect -3348 32167 -3048 32209
rect -3348 32049 -3257 32167
rect -3139 32049 -3048 32167
rect -3348 14327 -3048 32049
rect -3348 14209 -3257 14327
rect -3139 14209 -3048 14327
rect -3348 14167 -3048 14209
rect -3348 14049 -3257 14167
rect -3139 14049 -3048 14167
rect -3348 -2523 -3048 14049
rect -2878 354299 -2578 354310
rect -2878 354181 -2787 354299
rect -2669 354181 -2578 354299
rect -2878 354139 -2578 354181
rect -2878 354021 -2787 354139
rect -2669 354021 -2578 354139
rect -2878 347327 -2578 354021
rect 4502 354299 4802 354780
rect 4502 354181 4593 354299
rect 4711 354181 4802 354299
rect 4502 354139 4802 354181
rect 4502 354021 4593 354139
rect 4711 354021 4802 354139
rect -2878 347209 -2787 347327
rect -2669 347209 -2578 347327
rect -2878 347167 -2578 347209
rect -2878 347049 -2787 347167
rect -2669 347049 -2578 347167
rect -2878 329327 -2578 347049
rect -2878 329209 -2787 329327
rect -2669 329209 -2578 329327
rect -2878 329167 -2578 329209
rect -2878 329049 -2787 329167
rect -2669 329049 -2578 329167
rect -2878 311327 -2578 329049
rect -2878 311209 -2787 311327
rect -2669 311209 -2578 311327
rect -2878 311167 -2578 311209
rect -2878 311049 -2787 311167
rect -2669 311049 -2578 311167
rect -2878 293327 -2578 311049
rect -2878 293209 -2787 293327
rect -2669 293209 -2578 293327
rect -2878 293167 -2578 293209
rect -2878 293049 -2787 293167
rect -2669 293049 -2578 293167
rect -2878 275327 -2578 293049
rect -2878 275209 -2787 275327
rect -2669 275209 -2578 275327
rect -2878 275167 -2578 275209
rect -2878 275049 -2787 275167
rect -2669 275049 -2578 275167
rect -2878 257327 -2578 275049
rect -2878 257209 -2787 257327
rect -2669 257209 -2578 257327
rect -2878 257167 -2578 257209
rect -2878 257049 -2787 257167
rect -2669 257049 -2578 257167
rect -2878 239327 -2578 257049
rect -2878 239209 -2787 239327
rect -2669 239209 -2578 239327
rect -2878 239167 -2578 239209
rect -2878 239049 -2787 239167
rect -2669 239049 -2578 239167
rect -2878 221327 -2578 239049
rect -2878 221209 -2787 221327
rect -2669 221209 -2578 221327
rect -2878 221167 -2578 221209
rect -2878 221049 -2787 221167
rect -2669 221049 -2578 221167
rect -2878 203327 -2578 221049
rect -2878 203209 -2787 203327
rect -2669 203209 -2578 203327
rect -2878 203167 -2578 203209
rect -2878 203049 -2787 203167
rect -2669 203049 -2578 203167
rect -2878 185327 -2578 203049
rect -2878 185209 -2787 185327
rect -2669 185209 -2578 185327
rect -2878 185167 -2578 185209
rect -2878 185049 -2787 185167
rect -2669 185049 -2578 185167
rect -2878 167327 -2578 185049
rect -2878 167209 -2787 167327
rect -2669 167209 -2578 167327
rect -2878 167167 -2578 167209
rect -2878 167049 -2787 167167
rect -2669 167049 -2578 167167
rect -2878 149327 -2578 167049
rect -2878 149209 -2787 149327
rect -2669 149209 -2578 149327
rect -2878 149167 -2578 149209
rect -2878 149049 -2787 149167
rect -2669 149049 -2578 149167
rect -2878 131327 -2578 149049
rect -2878 131209 -2787 131327
rect -2669 131209 -2578 131327
rect -2878 131167 -2578 131209
rect -2878 131049 -2787 131167
rect -2669 131049 -2578 131167
rect -2878 113327 -2578 131049
rect -2878 113209 -2787 113327
rect -2669 113209 -2578 113327
rect -2878 113167 -2578 113209
rect -2878 113049 -2787 113167
rect -2669 113049 -2578 113167
rect -2878 95327 -2578 113049
rect -2878 95209 -2787 95327
rect -2669 95209 -2578 95327
rect -2878 95167 -2578 95209
rect -2878 95049 -2787 95167
rect -2669 95049 -2578 95167
rect -2878 77327 -2578 95049
rect -2878 77209 -2787 77327
rect -2669 77209 -2578 77327
rect -2878 77167 -2578 77209
rect -2878 77049 -2787 77167
rect -2669 77049 -2578 77167
rect -2878 59327 -2578 77049
rect -2878 59209 -2787 59327
rect -2669 59209 -2578 59327
rect -2878 59167 -2578 59209
rect -2878 59049 -2787 59167
rect -2669 59049 -2578 59167
rect -2878 41327 -2578 59049
rect -2878 41209 -2787 41327
rect -2669 41209 -2578 41327
rect -2878 41167 -2578 41209
rect -2878 41049 -2787 41167
rect -2669 41049 -2578 41167
rect -2878 23327 -2578 41049
rect -2878 23209 -2787 23327
rect -2669 23209 -2578 23327
rect -2878 23167 -2578 23209
rect -2878 23049 -2787 23167
rect -2669 23049 -2578 23167
rect -2878 5327 -2578 23049
rect -2878 5209 -2787 5327
rect -2669 5209 -2578 5327
rect -2878 5167 -2578 5209
rect -2878 5049 -2787 5167
rect -2669 5049 -2578 5167
rect -2878 -2053 -2578 5049
rect -2408 353829 -2108 353840
rect -2408 353711 -2317 353829
rect -2199 353711 -2108 353829
rect -2408 353669 -2108 353711
rect -2408 353551 -2317 353669
rect -2199 353551 -2108 353669
rect -2408 336527 -2108 353551
rect -2408 336409 -2317 336527
rect -2199 336409 -2108 336527
rect -2408 336367 -2108 336409
rect -2408 336249 -2317 336367
rect -2199 336249 -2108 336367
rect -2408 318527 -2108 336249
rect -2408 318409 -2317 318527
rect -2199 318409 -2108 318527
rect -2408 318367 -2108 318409
rect -2408 318249 -2317 318367
rect -2199 318249 -2108 318367
rect -2408 300527 -2108 318249
rect -2408 300409 -2317 300527
rect -2199 300409 -2108 300527
rect -2408 300367 -2108 300409
rect -2408 300249 -2317 300367
rect -2199 300249 -2108 300367
rect -2408 282527 -2108 300249
rect -2408 282409 -2317 282527
rect -2199 282409 -2108 282527
rect -2408 282367 -2108 282409
rect -2408 282249 -2317 282367
rect -2199 282249 -2108 282367
rect -2408 264527 -2108 282249
rect -2408 264409 -2317 264527
rect -2199 264409 -2108 264527
rect -2408 264367 -2108 264409
rect -2408 264249 -2317 264367
rect -2199 264249 -2108 264367
rect -2408 246527 -2108 264249
rect -2408 246409 -2317 246527
rect -2199 246409 -2108 246527
rect -2408 246367 -2108 246409
rect -2408 246249 -2317 246367
rect -2199 246249 -2108 246367
rect -2408 228527 -2108 246249
rect -2408 228409 -2317 228527
rect -2199 228409 -2108 228527
rect -2408 228367 -2108 228409
rect -2408 228249 -2317 228367
rect -2199 228249 -2108 228367
rect -2408 210527 -2108 228249
rect -2408 210409 -2317 210527
rect -2199 210409 -2108 210527
rect -2408 210367 -2108 210409
rect -2408 210249 -2317 210367
rect -2199 210249 -2108 210367
rect -2408 192527 -2108 210249
rect -2408 192409 -2317 192527
rect -2199 192409 -2108 192527
rect -2408 192367 -2108 192409
rect -2408 192249 -2317 192367
rect -2199 192249 -2108 192367
rect -2408 174527 -2108 192249
rect -2408 174409 -2317 174527
rect -2199 174409 -2108 174527
rect -2408 174367 -2108 174409
rect -2408 174249 -2317 174367
rect -2199 174249 -2108 174367
rect -2408 156527 -2108 174249
rect -2408 156409 -2317 156527
rect -2199 156409 -2108 156527
rect -2408 156367 -2108 156409
rect -2408 156249 -2317 156367
rect -2199 156249 -2108 156367
rect -2408 138527 -2108 156249
rect -2408 138409 -2317 138527
rect -2199 138409 -2108 138527
rect -2408 138367 -2108 138409
rect -2408 138249 -2317 138367
rect -2199 138249 -2108 138367
rect -2408 120527 -2108 138249
rect -2408 120409 -2317 120527
rect -2199 120409 -2108 120527
rect -2408 120367 -2108 120409
rect -2408 120249 -2317 120367
rect -2199 120249 -2108 120367
rect -2408 102527 -2108 120249
rect -2408 102409 -2317 102527
rect -2199 102409 -2108 102527
rect -2408 102367 -2108 102409
rect -2408 102249 -2317 102367
rect -2199 102249 -2108 102367
rect -2408 84527 -2108 102249
rect -2408 84409 -2317 84527
rect -2199 84409 -2108 84527
rect -2408 84367 -2108 84409
rect -2408 84249 -2317 84367
rect -2199 84249 -2108 84367
rect -2408 66527 -2108 84249
rect -2408 66409 -2317 66527
rect -2199 66409 -2108 66527
rect -2408 66367 -2108 66409
rect -2408 66249 -2317 66367
rect -2199 66249 -2108 66367
rect -2408 48527 -2108 66249
rect -2408 48409 -2317 48527
rect -2199 48409 -2108 48527
rect -2408 48367 -2108 48409
rect -2408 48249 -2317 48367
rect -2199 48249 -2108 48367
rect -2408 30527 -2108 48249
rect -2408 30409 -2317 30527
rect -2199 30409 -2108 30527
rect -2408 30367 -2108 30409
rect -2408 30249 -2317 30367
rect -2199 30249 -2108 30367
rect -2408 12527 -2108 30249
rect -2408 12409 -2317 12527
rect -2199 12409 -2108 12527
rect -2408 12367 -2108 12409
rect -2408 12249 -2317 12367
rect -2199 12249 -2108 12367
rect -2408 -1583 -2108 12249
rect -1938 353359 -1638 353370
rect -1938 353241 -1847 353359
rect -1729 353241 -1638 353359
rect -1938 353199 -1638 353241
rect -1938 353081 -1847 353199
rect -1729 353081 -1638 353199
rect -1938 345527 -1638 353081
rect 2702 353359 3002 353840
rect 2702 353241 2793 353359
rect 2911 353241 3002 353359
rect 2702 353199 3002 353241
rect 2702 353081 2793 353199
rect 2911 353081 3002 353199
rect -1938 345409 -1847 345527
rect -1729 345409 -1638 345527
rect -1938 345367 -1638 345409
rect -1938 345249 -1847 345367
rect -1729 345249 -1638 345367
rect -1938 327527 -1638 345249
rect -1938 327409 -1847 327527
rect -1729 327409 -1638 327527
rect -1938 327367 -1638 327409
rect -1938 327249 -1847 327367
rect -1729 327249 -1638 327367
rect -1938 309527 -1638 327249
rect -1938 309409 -1847 309527
rect -1729 309409 -1638 309527
rect -1938 309367 -1638 309409
rect -1938 309249 -1847 309367
rect -1729 309249 -1638 309367
rect -1938 291527 -1638 309249
rect -1938 291409 -1847 291527
rect -1729 291409 -1638 291527
rect -1938 291367 -1638 291409
rect -1938 291249 -1847 291367
rect -1729 291249 -1638 291367
rect -1938 273527 -1638 291249
rect -1938 273409 -1847 273527
rect -1729 273409 -1638 273527
rect -1938 273367 -1638 273409
rect -1938 273249 -1847 273367
rect -1729 273249 -1638 273367
rect -1938 255527 -1638 273249
rect -1938 255409 -1847 255527
rect -1729 255409 -1638 255527
rect -1938 255367 -1638 255409
rect -1938 255249 -1847 255367
rect -1729 255249 -1638 255367
rect -1938 237527 -1638 255249
rect -1938 237409 -1847 237527
rect -1729 237409 -1638 237527
rect -1938 237367 -1638 237409
rect -1938 237249 -1847 237367
rect -1729 237249 -1638 237367
rect -1938 219527 -1638 237249
rect -1938 219409 -1847 219527
rect -1729 219409 -1638 219527
rect -1938 219367 -1638 219409
rect -1938 219249 -1847 219367
rect -1729 219249 -1638 219367
rect -1938 201527 -1638 219249
rect -1938 201409 -1847 201527
rect -1729 201409 -1638 201527
rect -1938 201367 -1638 201409
rect -1938 201249 -1847 201367
rect -1729 201249 -1638 201367
rect -1938 183527 -1638 201249
rect -1938 183409 -1847 183527
rect -1729 183409 -1638 183527
rect -1938 183367 -1638 183409
rect -1938 183249 -1847 183367
rect -1729 183249 -1638 183367
rect -1938 165527 -1638 183249
rect -1938 165409 -1847 165527
rect -1729 165409 -1638 165527
rect -1938 165367 -1638 165409
rect -1938 165249 -1847 165367
rect -1729 165249 -1638 165367
rect -1938 147527 -1638 165249
rect -1938 147409 -1847 147527
rect -1729 147409 -1638 147527
rect -1938 147367 -1638 147409
rect -1938 147249 -1847 147367
rect -1729 147249 -1638 147367
rect -1938 129527 -1638 147249
rect -1938 129409 -1847 129527
rect -1729 129409 -1638 129527
rect -1938 129367 -1638 129409
rect -1938 129249 -1847 129367
rect -1729 129249 -1638 129367
rect -1938 111527 -1638 129249
rect -1938 111409 -1847 111527
rect -1729 111409 -1638 111527
rect -1938 111367 -1638 111409
rect -1938 111249 -1847 111367
rect -1729 111249 -1638 111367
rect -1938 93527 -1638 111249
rect -1938 93409 -1847 93527
rect -1729 93409 -1638 93527
rect -1938 93367 -1638 93409
rect -1938 93249 -1847 93367
rect -1729 93249 -1638 93367
rect -1938 75527 -1638 93249
rect -1938 75409 -1847 75527
rect -1729 75409 -1638 75527
rect -1938 75367 -1638 75409
rect -1938 75249 -1847 75367
rect -1729 75249 -1638 75367
rect -1938 57527 -1638 75249
rect -1938 57409 -1847 57527
rect -1729 57409 -1638 57527
rect -1938 57367 -1638 57409
rect -1938 57249 -1847 57367
rect -1729 57249 -1638 57367
rect -1938 39527 -1638 57249
rect -1938 39409 -1847 39527
rect -1729 39409 -1638 39527
rect -1938 39367 -1638 39409
rect -1938 39249 -1847 39367
rect -1729 39249 -1638 39367
rect -1938 21527 -1638 39249
rect -1938 21409 -1847 21527
rect -1729 21409 -1638 21527
rect -1938 21367 -1638 21409
rect -1938 21249 -1847 21367
rect -1729 21249 -1638 21367
rect -1938 3527 -1638 21249
rect -1938 3409 -1847 3527
rect -1729 3409 -1638 3527
rect -1938 3367 -1638 3409
rect -1938 3249 -1847 3367
rect -1729 3249 -1638 3367
rect -1938 -1113 -1638 3249
rect -1468 352889 -1168 352900
rect -1468 352771 -1377 352889
rect -1259 352771 -1168 352889
rect -1468 352729 -1168 352771
rect -1468 352611 -1377 352729
rect -1259 352611 -1168 352729
rect -1468 334727 -1168 352611
rect -1468 334609 -1377 334727
rect -1259 334609 -1168 334727
rect -1468 334567 -1168 334609
rect -1468 334449 -1377 334567
rect -1259 334449 -1168 334567
rect -1468 316727 -1168 334449
rect -1468 316609 -1377 316727
rect -1259 316609 -1168 316727
rect -1468 316567 -1168 316609
rect -1468 316449 -1377 316567
rect -1259 316449 -1168 316567
rect -1468 298727 -1168 316449
rect -1468 298609 -1377 298727
rect -1259 298609 -1168 298727
rect -1468 298567 -1168 298609
rect -1468 298449 -1377 298567
rect -1259 298449 -1168 298567
rect -1468 280727 -1168 298449
rect -1468 280609 -1377 280727
rect -1259 280609 -1168 280727
rect -1468 280567 -1168 280609
rect -1468 280449 -1377 280567
rect -1259 280449 -1168 280567
rect -1468 262727 -1168 280449
rect -1468 262609 -1377 262727
rect -1259 262609 -1168 262727
rect -1468 262567 -1168 262609
rect -1468 262449 -1377 262567
rect -1259 262449 -1168 262567
rect -1468 244727 -1168 262449
rect -1468 244609 -1377 244727
rect -1259 244609 -1168 244727
rect -1468 244567 -1168 244609
rect -1468 244449 -1377 244567
rect -1259 244449 -1168 244567
rect -1468 226727 -1168 244449
rect -1468 226609 -1377 226727
rect -1259 226609 -1168 226727
rect -1468 226567 -1168 226609
rect -1468 226449 -1377 226567
rect -1259 226449 -1168 226567
rect -1468 208727 -1168 226449
rect -1468 208609 -1377 208727
rect -1259 208609 -1168 208727
rect -1468 208567 -1168 208609
rect -1468 208449 -1377 208567
rect -1259 208449 -1168 208567
rect -1468 190727 -1168 208449
rect -1468 190609 -1377 190727
rect -1259 190609 -1168 190727
rect -1468 190567 -1168 190609
rect -1468 190449 -1377 190567
rect -1259 190449 -1168 190567
rect -1468 172727 -1168 190449
rect -1468 172609 -1377 172727
rect -1259 172609 -1168 172727
rect -1468 172567 -1168 172609
rect -1468 172449 -1377 172567
rect -1259 172449 -1168 172567
rect -1468 154727 -1168 172449
rect -1468 154609 -1377 154727
rect -1259 154609 -1168 154727
rect -1468 154567 -1168 154609
rect -1468 154449 -1377 154567
rect -1259 154449 -1168 154567
rect -1468 136727 -1168 154449
rect -1468 136609 -1377 136727
rect -1259 136609 -1168 136727
rect -1468 136567 -1168 136609
rect -1468 136449 -1377 136567
rect -1259 136449 -1168 136567
rect -1468 118727 -1168 136449
rect -1468 118609 -1377 118727
rect -1259 118609 -1168 118727
rect -1468 118567 -1168 118609
rect -1468 118449 -1377 118567
rect -1259 118449 -1168 118567
rect -1468 100727 -1168 118449
rect -1468 100609 -1377 100727
rect -1259 100609 -1168 100727
rect -1468 100567 -1168 100609
rect -1468 100449 -1377 100567
rect -1259 100449 -1168 100567
rect -1468 82727 -1168 100449
rect -1468 82609 -1377 82727
rect -1259 82609 -1168 82727
rect -1468 82567 -1168 82609
rect -1468 82449 -1377 82567
rect -1259 82449 -1168 82567
rect -1468 64727 -1168 82449
rect -1468 64609 -1377 64727
rect -1259 64609 -1168 64727
rect -1468 64567 -1168 64609
rect -1468 64449 -1377 64567
rect -1259 64449 -1168 64567
rect -1468 46727 -1168 64449
rect -1468 46609 -1377 46727
rect -1259 46609 -1168 46727
rect -1468 46567 -1168 46609
rect -1468 46449 -1377 46567
rect -1259 46449 -1168 46567
rect -1468 28727 -1168 46449
rect -1468 28609 -1377 28727
rect -1259 28609 -1168 28727
rect -1468 28567 -1168 28609
rect -1468 28449 -1377 28567
rect -1259 28449 -1168 28567
rect -1468 10727 -1168 28449
rect -1468 10609 -1377 10727
rect -1259 10609 -1168 10727
rect -1468 10567 -1168 10609
rect -1468 10449 -1377 10567
rect -1259 10449 -1168 10567
rect -1468 -643 -1168 10449
rect -998 352419 -698 352430
rect -998 352301 -907 352419
rect -789 352301 -698 352419
rect -998 352259 -698 352301
rect -998 352141 -907 352259
rect -789 352141 -698 352259
rect -998 343727 -698 352141
rect -998 343609 -907 343727
rect -789 343609 -698 343727
rect -998 343567 -698 343609
rect -998 343449 -907 343567
rect -789 343449 -698 343567
rect -998 325727 -698 343449
rect -998 325609 -907 325727
rect -789 325609 -698 325727
rect -998 325567 -698 325609
rect -998 325449 -907 325567
rect -789 325449 -698 325567
rect -998 307727 -698 325449
rect -998 307609 -907 307727
rect -789 307609 -698 307727
rect -998 307567 -698 307609
rect -998 307449 -907 307567
rect -789 307449 -698 307567
rect -998 289727 -698 307449
rect -998 289609 -907 289727
rect -789 289609 -698 289727
rect -998 289567 -698 289609
rect -998 289449 -907 289567
rect -789 289449 -698 289567
rect -998 271727 -698 289449
rect -998 271609 -907 271727
rect -789 271609 -698 271727
rect -998 271567 -698 271609
rect -998 271449 -907 271567
rect -789 271449 -698 271567
rect -998 253727 -698 271449
rect -998 253609 -907 253727
rect -789 253609 -698 253727
rect -998 253567 -698 253609
rect -998 253449 -907 253567
rect -789 253449 -698 253567
rect -998 235727 -698 253449
rect -998 235609 -907 235727
rect -789 235609 -698 235727
rect -998 235567 -698 235609
rect -998 235449 -907 235567
rect -789 235449 -698 235567
rect -998 217727 -698 235449
rect -998 217609 -907 217727
rect -789 217609 -698 217727
rect -998 217567 -698 217609
rect -998 217449 -907 217567
rect -789 217449 -698 217567
rect -998 199727 -698 217449
rect -998 199609 -907 199727
rect -789 199609 -698 199727
rect -998 199567 -698 199609
rect -998 199449 -907 199567
rect -789 199449 -698 199567
rect -998 181727 -698 199449
rect -998 181609 -907 181727
rect -789 181609 -698 181727
rect -998 181567 -698 181609
rect -998 181449 -907 181567
rect -789 181449 -698 181567
rect -998 163727 -698 181449
rect -998 163609 -907 163727
rect -789 163609 -698 163727
rect -998 163567 -698 163609
rect -998 163449 -907 163567
rect -789 163449 -698 163567
rect -998 145727 -698 163449
rect -998 145609 -907 145727
rect -789 145609 -698 145727
rect -998 145567 -698 145609
rect -998 145449 -907 145567
rect -789 145449 -698 145567
rect -998 127727 -698 145449
rect -998 127609 -907 127727
rect -789 127609 -698 127727
rect -998 127567 -698 127609
rect -998 127449 -907 127567
rect -789 127449 -698 127567
rect -998 109727 -698 127449
rect -998 109609 -907 109727
rect -789 109609 -698 109727
rect -998 109567 -698 109609
rect -998 109449 -907 109567
rect -789 109449 -698 109567
rect -998 91727 -698 109449
rect -998 91609 -907 91727
rect -789 91609 -698 91727
rect -998 91567 -698 91609
rect -998 91449 -907 91567
rect -789 91449 -698 91567
rect -998 73727 -698 91449
rect -998 73609 -907 73727
rect -789 73609 -698 73727
rect -998 73567 -698 73609
rect -998 73449 -907 73567
rect -789 73449 -698 73567
rect -998 55727 -698 73449
rect -998 55609 -907 55727
rect -789 55609 -698 55727
rect -998 55567 -698 55609
rect -998 55449 -907 55567
rect -789 55449 -698 55567
rect -998 37727 -698 55449
rect -998 37609 -907 37727
rect -789 37609 -698 37727
rect -998 37567 -698 37609
rect -998 37449 -907 37567
rect -789 37449 -698 37567
rect -998 19727 -698 37449
rect -998 19609 -907 19727
rect -789 19609 -698 19727
rect -998 19567 -698 19609
rect -998 19449 -907 19567
rect -789 19449 -698 19567
rect -998 1727 -698 19449
rect -998 1609 -907 1727
rect -789 1609 -698 1727
rect -998 1567 -698 1609
rect -998 1449 -907 1567
rect -789 1449 -698 1567
rect -998 -173 -698 1449
rect -998 -291 -907 -173
rect -789 -291 -698 -173
rect -998 -333 -698 -291
rect -998 -451 -907 -333
rect -789 -451 -698 -333
rect -998 -462 -698 -451
rect 902 352419 1202 352900
rect 902 352301 993 352419
rect 1111 352301 1202 352419
rect 902 352259 1202 352301
rect 902 352141 993 352259
rect 1111 352141 1202 352259
rect 902 343727 1202 352141
rect 902 343609 993 343727
rect 1111 343609 1202 343727
rect 902 343567 1202 343609
rect 902 343449 993 343567
rect 1111 343449 1202 343567
rect 902 325727 1202 343449
rect 902 325609 993 325727
rect 1111 325609 1202 325727
rect 902 325567 1202 325609
rect 902 325449 993 325567
rect 1111 325449 1202 325567
rect 902 307727 1202 325449
rect 902 307609 993 307727
rect 1111 307609 1202 307727
rect 902 307567 1202 307609
rect 902 307449 993 307567
rect 1111 307449 1202 307567
rect 902 289727 1202 307449
rect 902 289609 993 289727
rect 1111 289609 1202 289727
rect 902 289567 1202 289609
rect 902 289449 993 289567
rect 1111 289449 1202 289567
rect 902 271727 1202 289449
rect 902 271609 993 271727
rect 1111 271609 1202 271727
rect 902 271567 1202 271609
rect 902 271449 993 271567
rect 1111 271449 1202 271567
rect 902 253727 1202 271449
rect 902 253609 993 253727
rect 1111 253609 1202 253727
rect 902 253567 1202 253609
rect 902 253449 993 253567
rect 1111 253449 1202 253567
rect 902 235727 1202 253449
rect 902 235609 993 235727
rect 1111 235609 1202 235727
rect 902 235567 1202 235609
rect 902 235449 993 235567
rect 1111 235449 1202 235567
rect 902 217727 1202 235449
rect 902 217609 993 217727
rect 1111 217609 1202 217727
rect 902 217567 1202 217609
rect 902 217449 993 217567
rect 1111 217449 1202 217567
rect 902 199727 1202 217449
rect 902 199609 993 199727
rect 1111 199609 1202 199727
rect 902 199567 1202 199609
rect 902 199449 993 199567
rect 1111 199449 1202 199567
rect 902 181727 1202 199449
rect 902 181609 993 181727
rect 1111 181609 1202 181727
rect 902 181567 1202 181609
rect 902 181449 993 181567
rect 1111 181449 1202 181567
rect 902 163727 1202 181449
rect 902 163609 993 163727
rect 1111 163609 1202 163727
rect 902 163567 1202 163609
rect 902 163449 993 163567
rect 1111 163449 1202 163567
rect 902 145727 1202 163449
rect 902 145609 993 145727
rect 1111 145609 1202 145727
rect 902 145567 1202 145609
rect 902 145449 993 145567
rect 1111 145449 1202 145567
rect 902 127727 1202 145449
rect 902 127609 993 127727
rect 1111 127609 1202 127727
rect 902 127567 1202 127609
rect 902 127449 993 127567
rect 1111 127449 1202 127567
rect 902 109727 1202 127449
rect 902 109609 993 109727
rect 1111 109609 1202 109727
rect 902 109567 1202 109609
rect 902 109449 993 109567
rect 1111 109449 1202 109567
rect 902 91727 1202 109449
rect 902 91609 993 91727
rect 1111 91609 1202 91727
rect 902 91567 1202 91609
rect 902 91449 993 91567
rect 1111 91449 1202 91567
rect 902 73727 1202 91449
rect 902 73609 993 73727
rect 1111 73609 1202 73727
rect 902 73567 1202 73609
rect 902 73449 993 73567
rect 1111 73449 1202 73567
rect 902 55727 1202 73449
rect 902 55609 993 55727
rect 1111 55609 1202 55727
rect 902 55567 1202 55609
rect 902 55449 993 55567
rect 1111 55449 1202 55567
rect 902 37727 1202 55449
rect 902 37609 993 37727
rect 1111 37609 1202 37727
rect 902 37567 1202 37609
rect 902 37449 993 37567
rect 1111 37449 1202 37567
rect 902 19727 1202 37449
rect 902 19609 993 19727
rect 1111 19609 1202 19727
rect 902 19567 1202 19609
rect 902 19449 993 19567
rect 1111 19449 1202 19567
rect 902 1727 1202 19449
rect 902 1609 993 1727
rect 1111 1609 1202 1727
rect 902 1567 1202 1609
rect 902 1449 993 1567
rect 1111 1449 1202 1567
rect 902 -173 1202 1449
rect 902 -291 993 -173
rect 1111 -291 1202 -173
rect 902 -333 1202 -291
rect 902 -451 993 -333
rect 1111 -451 1202 -333
rect -1468 -761 -1377 -643
rect -1259 -761 -1168 -643
rect -1468 -803 -1168 -761
rect -1468 -921 -1377 -803
rect -1259 -921 -1168 -803
rect -1468 -932 -1168 -921
rect 902 -932 1202 -451
rect 2702 345527 3002 353081
rect 2702 345409 2793 345527
rect 2911 345409 3002 345527
rect 2702 345367 3002 345409
rect 2702 345249 2793 345367
rect 2911 345249 3002 345367
rect 2702 327527 3002 345249
rect 2702 327409 2793 327527
rect 2911 327409 3002 327527
rect 2702 327367 3002 327409
rect 2702 327249 2793 327367
rect 2911 327249 3002 327367
rect 2702 309527 3002 327249
rect 2702 309409 2793 309527
rect 2911 309409 3002 309527
rect 2702 309367 3002 309409
rect 2702 309249 2793 309367
rect 2911 309249 3002 309367
rect 2702 291527 3002 309249
rect 2702 291409 2793 291527
rect 2911 291409 3002 291527
rect 2702 291367 3002 291409
rect 2702 291249 2793 291367
rect 2911 291249 3002 291367
rect 2702 273527 3002 291249
rect 2702 273409 2793 273527
rect 2911 273409 3002 273527
rect 2702 273367 3002 273409
rect 2702 273249 2793 273367
rect 2911 273249 3002 273367
rect 2702 255527 3002 273249
rect 2702 255409 2793 255527
rect 2911 255409 3002 255527
rect 2702 255367 3002 255409
rect 2702 255249 2793 255367
rect 2911 255249 3002 255367
rect 2702 237527 3002 255249
rect 2702 237409 2793 237527
rect 2911 237409 3002 237527
rect 2702 237367 3002 237409
rect 2702 237249 2793 237367
rect 2911 237249 3002 237367
rect 2702 219527 3002 237249
rect 2702 219409 2793 219527
rect 2911 219409 3002 219527
rect 2702 219367 3002 219409
rect 2702 219249 2793 219367
rect 2911 219249 3002 219367
rect 2702 201527 3002 219249
rect 2702 201409 2793 201527
rect 2911 201409 3002 201527
rect 2702 201367 3002 201409
rect 2702 201249 2793 201367
rect 2911 201249 3002 201367
rect 2702 183527 3002 201249
rect 2702 183409 2793 183527
rect 2911 183409 3002 183527
rect 2702 183367 3002 183409
rect 2702 183249 2793 183367
rect 2911 183249 3002 183367
rect 2702 165527 3002 183249
rect 2702 165409 2793 165527
rect 2911 165409 3002 165527
rect 2702 165367 3002 165409
rect 2702 165249 2793 165367
rect 2911 165249 3002 165367
rect 2702 147527 3002 165249
rect 2702 147409 2793 147527
rect 2911 147409 3002 147527
rect 2702 147367 3002 147409
rect 2702 147249 2793 147367
rect 2911 147249 3002 147367
rect 2702 129527 3002 147249
rect 2702 129409 2793 129527
rect 2911 129409 3002 129527
rect 2702 129367 3002 129409
rect 2702 129249 2793 129367
rect 2911 129249 3002 129367
rect 2702 111527 3002 129249
rect 2702 111409 2793 111527
rect 2911 111409 3002 111527
rect 2702 111367 3002 111409
rect 2702 111249 2793 111367
rect 2911 111249 3002 111367
rect 2702 93527 3002 111249
rect 2702 93409 2793 93527
rect 2911 93409 3002 93527
rect 2702 93367 3002 93409
rect 2702 93249 2793 93367
rect 2911 93249 3002 93367
rect 2702 75527 3002 93249
rect 2702 75409 2793 75527
rect 2911 75409 3002 75527
rect 2702 75367 3002 75409
rect 2702 75249 2793 75367
rect 2911 75249 3002 75367
rect 2702 57527 3002 75249
rect 2702 57409 2793 57527
rect 2911 57409 3002 57527
rect 2702 57367 3002 57409
rect 2702 57249 2793 57367
rect 2911 57249 3002 57367
rect 2702 39527 3002 57249
rect 2702 39409 2793 39527
rect 2911 39409 3002 39527
rect 2702 39367 3002 39409
rect 2702 39249 2793 39367
rect 2911 39249 3002 39367
rect 2702 21527 3002 39249
rect 2702 21409 2793 21527
rect 2911 21409 3002 21527
rect 2702 21367 3002 21409
rect 2702 21249 2793 21367
rect 2911 21249 3002 21367
rect 2702 3527 3002 21249
rect 2702 3409 2793 3527
rect 2911 3409 3002 3527
rect 2702 3367 3002 3409
rect 2702 3249 2793 3367
rect 2911 3249 3002 3367
rect -1938 -1231 -1847 -1113
rect -1729 -1231 -1638 -1113
rect -1938 -1273 -1638 -1231
rect -1938 -1391 -1847 -1273
rect -1729 -1391 -1638 -1273
rect -1938 -1402 -1638 -1391
rect 2702 -1113 3002 3249
rect 2702 -1231 2793 -1113
rect 2911 -1231 3002 -1113
rect 2702 -1273 3002 -1231
rect 2702 -1391 2793 -1273
rect 2911 -1391 3002 -1273
rect -2408 -1701 -2317 -1583
rect -2199 -1701 -2108 -1583
rect -2408 -1743 -2108 -1701
rect -2408 -1861 -2317 -1743
rect -2199 -1861 -2108 -1743
rect -2408 -1872 -2108 -1861
rect 2702 -1872 3002 -1391
rect 4502 347327 4802 354021
rect 4502 347209 4593 347327
rect 4711 347209 4802 347327
rect 4502 347167 4802 347209
rect 4502 347049 4593 347167
rect 4711 347049 4802 347167
rect 4502 329327 4802 347049
rect 4502 329209 4593 329327
rect 4711 329209 4802 329327
rect 4502 329167 4802 329209
rect 4502 329049 4593 329167
rect 4711 329049 4802 329167
rect 4502 311327 4802 329049
rect 4502 311209 4593 311327
rect 4711 311209 4802 311327
rect 4502 311167 4802 311209
rect 4502 311049 4593 311167
rect 4711 311049 4802 311167
rect 4502 293327 4802 311049
rect 4502 293209 4593 293327
rect 4711 293209 4802 293327
rect 4502 293167 4802 293209
rect 4502 293049 4593 293167
rect 4711 293049 4802 293167
rect 4502 275327 4802 293049
rect 4502 275209 4593 275327
rect 4711 275209 4802 275327
rect 4502 275167 4802 275209
rect 4502 275049 4593 275167
rect 4711 275049 4802 275167
rect 4502 257327 4802 275049
rect 4502 257209 4593 257327
rect 4711 257209 4802 257327
rect 4502 257167 4802 257209
rect 4502 257049 4593 257167
rect 4711 257049 4802 257167
rect 4502 239327 4802 257049
rect 4502 239209 4593 239327
rect 4711 239209 4802 239327
rect 4502 239167 4802 239209
rect 4502 239049 4593 239167
rect 4711 239049 4802 239167
rect 4502 221327 4802 239049
rect 4502 221209 4593 221327
rect 4711 221209 4802 221327
rect 4502 221167 4802 221209
rect 4502 221049 4593 221167
rect 4711 221049 4802 221167
rect 4502 203327 4802 221049
rect 4502 203209 4593 203327
rect 4711 203209 4802 203327
rect 4502 203167 4802 203209
rect 4502 203049 4593 203167
rect 4711 203049 4802 203167
rect 4502 185327 4802 203049
rect 4502 185209 4593 185327
rect 4711 185209 4802 185327
rect 4502 185167 4802 185209
rect 4502 185049 4593 185167
rect 4711 185049 4802 185167
rect 4502 167327 4802 185049
rect 4502 167209 4593 167327
rect 4711 167209 4802 167327
rect 4502 167167 4802 167209
rect 4502 167049 4593 167167
rect 4711 167049 4802 167167
rect 4502 149327 4802 167049
rect 4502 149209 4593 149327
rect 4711 149209 4802 149327
rect 4502 149167 4802 149209
rect 4502 149049 4593 149167
rect 4711 149049 4802 149167
rect 4502 131327 4802 149049
rect 4502 131209 4593 131327
rect 4711 131209 4802 131327
rect 4502 131167 4802 131209
rect 4502 131049 4593 131167
rect 4711 131049 4802 131167
rect 4502 113327 4802 131049
rect 4502 113209 4593 113327
rect 4711 113209 4802 113327
rect 4502 113167 4802 113209
rect 4502 113049 4593 113167
rect 4711 113049 4802 113167
rect 4502 95327 4802 113049
rect 4502 95209 4593 95327
rect 4711 95209 4802 95327
rect 4502 95167 4802 95209
rect 4502 95049 4593 95167
rect 4711 95049 4802 95167
rect 4502 77327 4802 95049
rect 4502 77209 4593 77327
rect 4711 77209 4802 77327
rect 4502 77167 4802 77209
rect 4502 77049 4593 77167
rect 4711 77049 4802 77167
rect 4502 59327 4802 77049
rect 4502 59209 4593 59327
rect 4711 59209 4802 59327
rect 4502 59167 4802 59209
rect 4502 59049 4593 59167
rect 4711 59049 4802 59167
rect 4502 41327 4802 59049
rect 4502 41209 4593 41327
rect 4711 41209 4802 41327
rect 4502 41167 4802 41209
rect 4502 41049 4593 41167
rect 4711 41049 4802 41167
rect 4502 23327 4802 41049
rect 4502 23209 4593 23327
rect 4711 23209 4802 23327
rect 4502 23167 4802 23209
rect 4502 23049 4593 23167
rect 4711 23049 4802 23167
rect 4502 5327 4802 23049
rect 4502 5209 4593 5327
rect 4711 5209 4802 5327
rect 4502 5167 4802 5209
rect 4502 5049 4593 5167
rect 4711 5049 4802 5167
rect -2878 -2171 -2787 -2053
rect -2669 -2171 -2578 -2053
rect -2878 -2213 -2578 -2171
rect -2878 -2331 -2787 -2213
rect -2669 -2331 -2578 -2213
rect -2878 -2342 -2578 -2331
rect 4502 -2053 4802 5049
rect 4502 -2171 4593 -2053
rect 4711 -2171 4802 -2053
rect 4502 -2213 4802 -2171
rect 4502 -2331 4593 -2213
rect 4711 -2331 4802 -2213
rect -3348 -2641 -3257 -2523
rect -3139 -2641 -3048 -2523
rect -3348 -2683 -3048 -2641
rect -3348 -2801 -3257 -2683
rect -3139 -2801 -3048 -2683
rect -3348 -2812 -3048 -2801
rect 4502 -2812 4802 -2331
rect 6302 349127 6602 354961
rect 15302 355709 15602 355720
rect 15302 355591 15393 355709
rect 15511 355591 15602 355709
rect 15302 355549 15602 355591
rect 15302 355431 15393 355549
rect 15511 355431 15602 355549
rect 13502 354769 13802 354780
rect 13502 354651 13593 354769
rect 13711 354651 13802 354769
rect 13502 354609 13802 354651
rect 13502 354491 13593 354609
rect 13711 354491 13802 354609
rect 11702 353829 12002 353840
rect 11702 353711 11793 353829
rect 11911 353711 12002 353829
rect 11702 353669 12002 353711
rect 11702 353551 11793 353669
rect 11911 353551 12002 353669
rect 6302 349009 6393 349127
rect 6511 349009 6602 349127
rect 6302 348967 6602 349009
rect 6302 348849 6393 348967
rect 6511 348849 6602 348967
rect 6302 331127 6602 348849
rect 6302 331009 6393 331127
rect 6511 331009 6602 331127
rect 6302 330967 6602 331009
rect 6302 330849 6393 330967
rect 6511 330849 6602 330967
rect 6302 313127 6602 330849
rect 6302 313009 6393 313127
rect 6511 313009 6602 313127
rect 6302 312967 6602 313009
rect 6302 312849 6393 312967
rect 6511 312849 6602 312967
rect 6302 295127 6602 312849
rect 6302 295009 6393 295127
rect 6511 295009 6602 295127
rect 6302 294967 6602 295009
rect 6302 294849 6393 294967
rect 6511 294849 6602 294967
rect 6302 277127 6602 294849
rect 6302 277009 6393 277127
rect 6511 277009 6602 277127
rect 6302 276967 6602 277009
rect 6302 276849 6393 276967
rect 6511 276849 6602 276967
rect 6302 259127 6602 276849
rect 6302 259009 6393 259127
rect 6511 259009 6602 259127
rect 6302 258967 6602 259009
rect 6302 258849 6393 258967
rect 6511 258849 6602 258967
rect 6302 241127 6602 258849
rect 6302 241009 6393 241127
rect 6511 241009 6602 241127
rect 6302 240967 6602 241009
rect 6302 240849 6393 240967
rect 6511 240849 6602 240967
rect 6302 223127 6602 240849
rect 6302 223009 6393 223127
rect 6511 223009 6602 223127
rect 6302 222967 6602 223009
rect 6302 222849 6393 222967
rect 6511 222849 6602 222967
rect 6302 205127 6602 222849
rect 6302 205009 6393 205127
rect 6511 205009 6602 205127
rect 6302 204967 6602 205009
rect 6302 204849 6393 204967
rect 6511 204849 6602 204967
rect 6302 187127 6602 204849
rect 6302 187009 6393 187127
rect 6511 187009 6602 187127
rect 6302 186967 6602 187009
rect 6302 186849 6393 186967
rect 6511 186849 6602 186967
rect 6302 169127 6602 186849
rect 6302 169009 6393 169127
rect 6511 169009 6602 169127
rect 6302 168967 6602 169009
rect 6302 168849 6393 168967
rect 6511 168849 6602 168967
rect 6302 151127 6602 168849
rect 6302 151009 6393 151127
rect 6511 151009 6602 151127
rect 6302 150967 6602 151009
rect 6302 150849 6393 150967
rect 6511 150849 6602 150967
rect 6302 133127 6602 150849
rect 6302 133009 6393 133127
rect 6511 133009 6602 133127
rect 6302 132967 6602 133009
rect 6302 132849 6393 132967
rect 6511 132849 6602 132967
rect 6302 115127 6602 132849
rect 6302 115009 6393 115127
rect 6511 115009 6602 115127
rect 6302 114967 6602 115009
rect 6302 114849 6393 114967
rect 6511 114849 6602 114967
rect 6302 97127 6602 114849
rect 6302 97009 6393 97127
rect 6511 97009 6602 97127
rect 6302 96967 6602 97009
rect 6302 96849 6393 96967
rect 6511 96849 6602 96967
rect 6302 79127 6602 96849
rect 6302 79009 6393 79127
rect 6511 79009 6602 79127
rect 6302 78967 6602 79009
rect 6302 78849 6393 78967
rect 6511 78849 6602 78967
rect 6302 61127 6602 78849
rect 6302 61009 6393 61127
rect 6511 61009 6602 61127
rect 6302 60967 6602 61009
rect 6302 60849 6393 60967
rect 6511 60849 6602 60967
rect 6302 43127 6602 60849
rect 6302 43009 6393 43127
rect 6511 43009 6602 43127
rect 6302 42967 6602 43009
rect 6302 42849 6393 42967
rect 6511 42849 6602 42967
rect 6302 25127 6602 42849
rect 6302 25009 6393 25127
rect 6511 25009 6602 25127
rect 6302 24967 6602 25009
rect 6302 24849 6393 24967
rect 6511 24849 6602 24967
rect 6302 7127 6602 24849
rect 6302 7009 6393 7127
rect 6511 7009 6602 7127
rect 6302 6967 6602 7009
rect 6302 6849 6393 6967
rect 6511 6849 6602 6967
rect -3818 -3111 -3727 -2993
rect -3609 -3111 -3518 -2993
rect -3818 -3153 -3518 -3111
rect -3818 -3271 -3727 -3153
rect -3609 -3271 -3518 -3153
rect -3818 -3282 -3518 -3271
rect 6302 -2993 6602 6849
rect 9902 352889 10202 352900
rect 9902 352771 9993 352889
rect 10111 352771 10202 352889
rect 9902 352729 10202 352771
rect 9902 352611 9993 352729
rect 10111 352611 10202 352729
rect 9902 334727 10202 352611
rect 9902 334609 9993 334727
rect 10111 334609 10202 334727
rect 9902 334567 10202 334609
rect 9902 334449 9993 334567
rect 10111 334449 10202 334567
rect 9902 316727 10202 334449
rect 9902 316609 9993 316727
rect 10111 316609 10202 316727
rect 9902 316567 10202 316609
rect 9902 316449 9993 316567
rect 10111 316449 10202 316567
rect 9902 298727 10202 316449
rect 9902 298609 9993 298727
rect 10111 298609 10202 298727
rect 9902 298567 10202 298609
rect 9902 298449 9993 298567
rect 10111 298449 10202 298567
rect 9902 280727 10202 298449
rect 9902 280609 9993 280727
rect 10111 280609 10202 280727
rect 9902 280567 10202 280609
rect 9902 280449 9993 280567
rect 10111 280449 10202 280567
rect 9902 262727 10202 280449
rect 9902 262609 9993 262727
rect 10111 262609 10202 262727
rect 9902 262567 10202 262609
rect 9902 262449 9993 262567
rect 10111 262449 10202 262567
rect 9902 244727 10202 262449
rect 9902 244609 9993 244727
rect 10111 244609 10202 244727
rect 9902 244567 10202 244609
rect 9902 244449 9993 244567
rect 10111 244449 10202 244567
rect 9902 226727 10202 244449
rect 9902 226609 9993 226727
rect 10111 226609 10202 226727
rect 9902 226567 10202 226609
rect 9902 226449 9993 226567
rect 10111 226449 10202 226567
rect 9902 208727 10202 226449
rect 9902 208609 9993 208727
rect 10111 208609 10202 208727
rect 9902 208567 10202 208609
rect 9902 208449 9993 208567
rect 10111 208449 10202 208567
rect 9902 190727 10202 208449
rect 9902 190609 9993 190727
rect 10111 190609 10202 190727
rect 9902 190567 10202 190609
rect 9902 190449 9993 190567
rect 10111 190449 10202 190567
rect 9902 172727 10202 190449
rect 9902 172609 9993 172727
rect 10111 172609 10202 172727
rect 9902 172567 10202 172609
rect 9902 172449 9993 172567
rect 10111 172449 10202 172567
rect 9902 154727 10202 172449
rect 9902 154609 9993 154727
rect 10111 154609 10202 154727
rect 9902 154567 10202 154609
rect 9902 154449 9993 154567
rect 10111 154449 10202 154567
rect 9902 136727 10202 154449
rect 9902 136609 9993 136727
rect 10111 136609 10202 136727
rect 9902 136567 10202 136609
rect 9902 136449 9993 136567
rect 10111 136449 10202 136567
rect 9902 118727 10202 136449
rect 9902 118609 9993 118727
rect 10111 118609 10202 118727
rect 9902 118567 10202 118609
rect 9902 118449 9993 118567
rect 10111 118449 10202 118567
rect 9902 100727 10202 118449
rect 9902 100609 9993 100727
rect 10111 100609 10202 100727
rect 9902 100567 10202 100609
rect 9902 100449 9993 100567
rect 10111 100449 10202 100567
rect 9902 82727 10202 100449
rect 9902 82609 9993 82727
rect 10111 82609 10202 82727
rect 9902 82567 10202 82609
rect 9902 82449 9993 82567
rect 10111 82449 10202 82567
rect 9902 64727 10202 82449
rect 9902 64609 9993 64727
rect 10111 64609 10202 64727
rect 9902 64567 10202 64609
rect 9902 64449 9993 64567
rect 10111 64449 10202 64567
rect 9902 46727 10202 64449
rect 9902 46609 9993 46727
rect 10111 46609 10202 46727
rect 9902 46567 10202 46609
rect 9902 46449 9993 46567
rect 10111 46449 10202 46567
rect 9902 28727 10202 46449
rect 9902 28609 9993 28727
rect 10111 28609 10202 28727
rect 9902 28567 10202 28609
rect 9902 28449 9993 28567
rect 10111 28449 10202 28567
rect 9902 10727 10202 28449
rect 9902 10609 9993 10727
rect 10111 10609 10202 10727
rect 9902 10567 10202 10609
rect 9902 10449 9993 10567
rect 10111 10449 10202 10567
rect 9902 -643 10202 10449
rect 9902 -761 9993 -643
rect 10111 -761 10202 -643
rect 9902 -803 10202 -761
rect 9902 -921 9993 -803
rect 10111 -921 10202 -803
rect 9902 -932 10202 -921
rect 11702 336527 12002 353551
rect 11702 336409 11793 336527
rect 11911 336409 12002 336527
rect 11702 336367 12002 336409
rect 11702 336249 11793 336367
rect 11911 336249 12002 336367
rect 11702 318527 12002 336249
rect 11702 318409 11793 318527
rect 11911 318409 12002 318527
rect 11702 318367 12002 318409
rect 11702 318249 11793 318367
rect 11911 318249 12002 318367
rect 11702 300527 12002 318249
rect 11702 300409 11793 300527
rect 11911 300409 12002 300527
rect 11702 300367 12002 300409
rect 11702 300249 11793 300367
rect 11911 300249 12002 300367
rect 11702 282527 12002 300249
rect 11702 282409 11793 282527
rect 11911 282409 12002 282527
rect 11702 282367 12002 282409
rect 11702 282249 11793 282367
rect 11911 282249 12002 282367
rect 11702 264527 12002 282249
rect 11702 264409 11793 264527
rect 11911 264409 12002 264527
rect 11702 264367 12002 264409
rect 11702 264249 11793 264367
rect 11911 264249 12002 264367
rect 11702 246527 12002 264249
rect 11702 246409 11793 246527
rect 11911 246409 12002 246527
rect 11702 246367 12002 246409
rect 11702 246249 11793 246367
rect 11911 246249 12002 246367
rect 11702 228527 12002 246249
rect 11702 228409 11793 228527
rect 11911 228409 12002 228527
rect 11702 228367 12002 228409
rect 11702 228249 11793 228367
rect 11911 228249 12002 228367
rect 11702 210527 12002 228249
rect 11702 210409 11793 210527
rect 11911 210409 12002 210527
rect 11702 210367 12002 210409
rect 11702 210249 11793 210367
rect 11911 210249 12002 210367
rect 11702 192527 12002 210249
rect 11702 192409 11793 192527
rect 11911 192409 12002 192527
rect 11702 192367 12002 192409
rect 11702 192249 11793 192367
rect 11911 192249 12002 192367
rect 11702 174527 12002 192249
rect 11702 174409 11793 174527
rect 11911 174409 12002 174527
rect 11702 174367 12002 174409
rect 11702 174249 11793 174367
rect 11911 174249 12002 174367
rect 11702 156527 12002 174249
rect 11702 156409 11793 156527
rect 11911 156409 12002 156527
rect 11702 156367 12002 156409
rect 11702 156249 11793 156367
rect 11911 156249 12002 156367
rect 11702 138527 12002 156249
rect 11702 138409 11793 138527
rect 11911 138409 12002 138527
rect 11702 138367 12002 138409
rect 11702 138249 11793 138367
rect 11911 138249 12002 138367
rect 11702 120527 12002 138249
rect 11702 120409 11793 120527
rect 11911 120409 12002 120527
rect 11702 120367 12002 120409
rect 11702 120249 11793 120367
rect 11911 120249 12002 120367
rect 11702 102527 12002 120249
rect 11702 102409 11793 102527
rect 11911 102409 12002 102527
rect 11702 102367 12002 102409
rect 11702 102249 11793 102367
rect 11911 102249 12002 102367
rect 11702 84527 12002 102249
rect 11702 84409 11793 84527
rect 11911 84409 12002 84527
rect 11702 84367 12002 84409
rect 11702 84249 11793 84367
rect 11911 84249 12002 84367
rect 11702 66527 12002 84249
rect 11702 66409 11793 66527
rect 11911 66409 12002 66527
rect 11702 66367 12002 66409
rect 11702 66249 11793 66367
rect 11911 66249 12002 66367
rect 11702 48527 12002 66249
rect 11702 48409 11793 48527
rect 11911 48409 12002 48527
rect 11702 48367 12002 48409
rect 11702 48249 11793 48367
rect 11911 48249 12002 48367
rect 11702 30527 12002 48249
rect 11702 30409 11793 30527
rect 11911 30409 12002 30527
rect 11702 30367 12002 30409
rect 11702 30249 11793 30367
rect 11911 30249 12002 30367
rect 11702 12527 12002 30249
rect 11702 12409 11793 12527
rect 11911 12409 12002 12527
rect 11702 12367 12002 12409
rect 11702 12249 11793 12367
rect 11911 12249 12002 12367
rect 11702 -1583 12002 12249
rect 11702 -1701 11793 -1583
rect 11911 -1701 12002 -1583
rect 11702 -1743 12002 -1701
rect 11702 -1861 11793 -1743
rect 11911 -1861 12002 -1743
rect 11702 -1872 12002 -1861
rect 13502 338327 13802 354491
rect 13502 338209 13593 338327
rect 13711 338209 13802 338327
rect 13502 338167 13802 338209
rect 13502 338049 13593 338167
rect 13711 338049 13802 338167
rect 13502 320327 13802 338049
rect 13502 320209 13593 320327
rect 13711 320209 13802 320327
rect 13502 320167 13802 320209
rect 13502 320049 13593 320167
rect 13711 320049 13802 320167
rect 13502 302327 13802 320049
rect 13502 302209 13593 302327
rect 13711 302209 13802 302327
rect 13502 302167 13802 302209
rect 13502 302049 13593 302167
rect 13711 302049 13802 302167
rect 13502 284327 13802 302049
rect 13502 284209 13593 284327
rect 13711 284209 13802 284327
rect 13502 284167 13802 284209
rect 13502 284049 13593 284167
rect 13711 284049 13802 284167
rect 13502 266327 13802 284049
rect 13502 266209 13593 266327
rect 13711 266209 13802 266327
rect 13502 266167 13802 266209
rect 13502 266049 13593 266167
rect 13711 266049 13802 266167
rect 13502 248327 13802 266049
rect 13502 248209 13593 248327
rect 13711 248209 13802 248327
rect 13502 248167 13802 248209
rect 13502 248049 13593 248167
rect 13711 248049 13802 248167
rect 13502 230327 13802 248049
rect 13502 230209 13593 230327
rect 13711 230209 13802 230327
rect 13502 230167 13802 230209
rect 13502 230049 13593 230167
rect 13711 230049 13802 230167
rect 13502 212327 13802 230049
rect 13502 212209 13593 212327
rect 13711 212209 13802 212327
rect 13502 212167 13802 212209
rect 13502 212049 13593 212167
rect 13711 212049 13802 212167
rect 13502 194327 13802 212049
rect 13502 194209 13593 194327
rect 13711 194209 13802 194327
rect 13502 194167 13802 194209
rect 13502 194049 13593 194167
rect 13711 194049 13802 194167
rect 13502 176327 13802 194049
rect 13502 176209 13593 176327
rect 13711 176209 13802 176327
rect 13502 176167 13802 176209
rect 13502 176049 13593 176167
rect 13711 176049 13802 176167
rect 13502 158327 13802 176049
rect 13502 158209 13593 158327
rect 13711 158209 13802 158327
rect 13502 158167 13802 158209
rect 13502 158049 13593 158167
rect 13711 158049 13802 158167
rect 13502 140327 13802 158049
rect 13502 140209 13593 140327
rect 13711 140209 13802 140327
rect 13502 140167 13802 140209
rect 13502 140049 13593 140167
rect 13711 140049 13802 140167
rect 13502 122327 13802 140049
rect 13502 122209 13593 122327
rect 13711 122209 13802 122327
rect 13502 122167 13802 122209
rect 13502 122049 13593 122167
rect 13711 122049 13802 122167
rect 13502 104327 13802 122049
rect 13502 104209 13593 104327
rect 13711 104209 13802 104327
rect 13502 104167 13802 104209
rect 13502 104049 13593 104167
rect 13711 104049 13802 104167
rect 13502 86327 13802 104049
rect 13502 86209 13593 86327
rect 13711 86209 13802 86327
rect 13502 86167 13802 86209
rect 13502 86049 13593 86167
rect 13711 86049 13802 86167
rect 13502 68327 13802 86049
rect 13502 68209 13593 68327
rect 13711 68209 13802 68327
rect 13502 68167 13802 68209
rect 13502 68049 13593 68167
rect 13711 68049 13802 68167
rect 13502 50327 13802 68049
rect 13502 50209 13593 50327
rect 13711 50209 13802 50327
rect 13502 50167 13802 50209
rect 13502 50049 13593 50167
rect 13711 50049 13802 50167
rect 13502 32327 13802 50049
rect 13502 32209 13593 32327
rect 13711 32209 13802 32327
rect 13502 32167 13802 32209
rect 13502 32049 13593 32167
rect 13711 32049 13802 32167
rect 13502 14327 13802 32049
rect 13502 14209 13593 14327
rect 13711 14209 13802 14327
rect 13502 14167 13802 14209
rect 13502 14049 13593 14167
rect 13711 14049 13802 14167
rect 13502 -2523 13802 14049
rect 13502 -2641 13593 -2523
rect 13711 -2641 13802 -2523
rect 13502 -2683 13802 -2641
rect 13502 -2801 13593 -2683
rect 13711 -2801 13802 -2683
rect 13502 -2812 13802 -2801
rect 15302 340127 15602 355431
rect 24302 355239 24602 355720
rect 24302 355121 24393 355239
rect 24511 355121 24602 355239
rect 24302 355079 24602 355121
rect 24302 354961 24393 355079
rect 24511 354961 24602 355079
rect 22502 354299 22802 354780
rect 22502 354181 22593 354299
rect 22711 354181 22802 354299
rect 22502 354139 22802 354181
rect 22502 354021 22593 354139
rect 22711 354021 22802 354139
rect 20702 353359 21002 353840
rect 20702 353241 20793 353359
rect 20911 353241 21002 353359
rect 20702 353199 21002 353241
rect 20702 353081 20793 353199
rect 20911 353081 21002 353199
rect 15302 340009 15393 340127
rect 15511 340009 15602 340127
rect 15302 339967 15602 340009
rect 15302 339849 15393 339967
rect 15511 339849 15602 339967
rect 15302 322127 15602 339849
rect 15302 322009 15393 322127
rect 15511 322009 15602 322127
rect 15302 321967 15602 322009
rect 15302 321849 15393 321967
rect 15511 321849 15602 321967
rect 15302 304127 15602 321849
rect 15302 304009 15393 304127
rect 15511 304009 15602 304127
rect 15302 303967 15602 304009
rect 15302 303849 15393 303967
rect 15511 303849 15602 303967
rect 15302 286127 15602 303849
rect 15302 286009 15393 286127
rect 15511 286009 15602 286127
rect 15302 285967 15602 286009
rect 15302 285849 15393 285967
rect 15511 285849 15602 285967
rect 15302 268127 15602 285849
rect 15302 268009 15393 268127
rect 15511 268009 15602 268127
rect 15302 267967 15602 268009
rect 15302 267849 15393 267967
rect 15511 267849 15602 267967
rect 15302 250127 15602 267849
rect 15302 250009 15393 250127
rect 15511 250009 15602 250127
rect 15302 249967 15602 250009
rect 15302 249849 15393 249967
rect 15511 249849 15602 249967
rect 15302 232127 15602 249849
rect 15302 232009 15393 232127
rect 15511 232009 15602 232127
rect 15302 231967 15602 232009
rect 15302 231849 15393 231967
rect 15511 231849 15602 231967
rect 15302 214127 15602 231849
rect 15302 214009 15393 214127
rect 15511 214009 15602 214127
rect 15302 213967 15602 214009
rect 15302 213849 15393 213967
rect 15511 213849 15602 213967
rect 15302 196127 15602 213849
rect 15302 196009 15393 196127
rect 15511 196009 15602 196127
rect 15302 195967 15602 196009
rect 15302 195849 15393 195967
rect 15511 195849 15602 195967
rect 15302 178127 15602 195849
rect 15302 178009 15393 178127
rect 15511 178009 15602 178127
rect 15302 177967 15602 178009
rect 15302 177849 15393 177967
rect 15511 177849 15602 177967
rect 15302 160127 15602 177849
rect 15302 160009 15393 160127
rect 15511 160009 15602 160127
rect 15302 159967 15602 160009
rect 15302 159849 15393 159967
rect 15511 159849 15602 159967
rect 15302 142127 15602 159849
rect 15302 142009 15393 142127
rect 15511 142009 15602 142127
rect 15302 141967 15602 142009
rect 15302 141849 15393 141967
rect 15511 141849 15602 141967
rect 15302 124127 15602 141849
rect 15302 124009 15393 124127
rect 15511 124009 15602 124127
rect 15302 123967 15602 124009
rect 15302 123849 15393 123967
rect 15511 123849 15602 123967
rect 15302 106127 15602 123849
rect 15302 106009 15393 106127
rect 15511 106009 15602 106127
rect 15302 105967 15602 106009
rect 15302 105849 15393 105967
rect 15511 105849 15602 105967
rect 15302 88127 15602 105849
rect 15302 88009 15393 88127
rect 15511 88009 15602 88127
rect 15302 87967 15602 88009
rect 15302 87849 15393 87967
rect 15511 87849 15602 87967
rect 15302 70127 15602 87849
rect 15302 70009 15393 70127
rect 15511 70009 15602 70127
rect 15302 69967 15602 70009
rect 15302 69849 15393 69967
rect 15511 69849 15602 69967
rect 15302 52127 15602 69849
rect 15302 52009 15393 52127
rect 15511 52009 15602 52127
rect 15302 51967 15602 52009
rect 15302 51849 15393 51967
rect 15511 51849 15602 51967
rect 15302 34127 15602 51849
rect 15302 34009 15393 34127
rect 15511 34009 15602 34127
rect 15302 33967 15602 34009
rect 15302 33849 15393 33967
rect 15511 33849 15602 33967
rect 15302 16127 15602 33849
rect 15302 16009 15393 16127
rect 15511 16009 15602 16127
rect 15302 15967 15602 16009
rect 15302 15849 15393 15967
rect 15511 15849 15602 15967
rect 6302 -3111 6393 -2993
rect 6511 -3111 6602 -2993
rect 6302 -3153 6602 -3111
rect 6302 -3271 6393 -3153
rect 6511 -3271 6602 -3153
rect -4288 -3581 -4197 -3463
rect -4079 -3581 -3988 -3463
rect -4288 -3623 -3988 -3581
rect -4288 -3741 -4197 -3623
rect -4079 -3741 -3988 -3623
rect -4288 -3752 -3988 -3741
rect 6302 -3752 6602 -3271
rect 15302 -3463 15602 15849
rect 18902 352419 19202 352900
rect 18902 352301 18993 352419
rect 19111 352301 19202 352419
rect 18902 352259 19202 352301
rect 18902 352141 18993 352259
rect 19111 352141 19202 352259
rect 18902 343727 19202 352141
rect 18902 343609 18993 343727
rect 19111 343609 19202 343727
rect 18902 343567 19202 343609
rect 18902 343449 18993 343567
rect 19111 343449 19202 343567
rect 18902 325727 19202 343449
rect 18902 325609 18993 325727
rect 19111 325609 19202 325727
rect 18902 325567 19202 325609
rect 18902 325449 18993 325567
rect 19111 325449 19202 325567
rect 18902 307727 19202 325449
rect 18902 307609 18993 307727
rect 19111 307609 19202 307727
rect 18902 307567 19202 307609
rect 18902 307449 18993 307567
rect 19111 307449 19202 307567
rect 18902 289727 19202 307449
rect 18902 289609 18993 289727
rect 19111 289609 19202 289727
rect 18902 289567 19202 289609
rect 18902 289449 18993 289567
rect 19111 289449 19202 289567
rect 18902 271727 19202 289449
rect 18902 271609 18993 271727
rect 19111 271609 19202 271727
rect 18902 271567 19202 271609
rect 18902 271449 18993 271567
rect 19111 271449 19202 271567
rect 18902 253727 19202 271449
rect 18902 253609 18993 253727
rect 19111 253609 19202 253727
rect 18902 253567 19202 253609
rect 18902 253449 18993 253567
rect 19111 253449 19202 253567
rect 18902 235727 19202 253449
rect 18902 235609 18993 235727
rect 19111 235609 19202 235727
rect 18902 235567 19202 235609
rect 18902 235449 18993 235567
rect 19111 235449 19202 235567
rect 18902 217727 19202 235449
rect 18902 217609 18993 217727
rect 19111 217609 19202 217727
rect 18902 217567 19202 217609
rect 18902 217449 18993 217567
rect 19111 217449 19202 217567
rect 18902 199727 19202 217449
rect 18902 199609 18993 199727
rect 19111 199609 19202 199727
rect 18902 199567 19202 199609
rect 18902 199449 18993 199567
rect 19111 199449 19202 199567
rect 18902 181727 19202 199449
rect 18902 181609 18993 181727
rect 19111 181609 19202 181727
rect 18902 181567 19202 181609
rect 18902 181449 18993 181567
rect 19111 181449 19202 181567
rect 18902 163727 19202 181449
rect 18902 163609 18993 163727
rect 19111 163609 19202 163727
rect 18902 163567 19202 163609
rect 18902 163449 18993 163567
rect 19111 163449 19202 163567
rect 18902 145727 19202 163449
rect 18902 145609 18993 145727
rect 19111 145609 19202 145727
rect 18902 145567 19202 145609
rect 18902 145449 18993 145567
rect 19111 145449 19202 145567
rect 18902 127727 19202 145449
rect 18902 127609 18993 127727
rect 19111 127609 19202 127727
rect 18902 127567 19202 127609
rect 18902 127449 18993 127567
rect 19111 127449 19202 127567
rect 18902 109727 19202 127449
rect 18902 109609 18993 109727
rect 19111 109609 19202 109727
rect 18902 109567 19202 109609
rect 18902 109449 18993 109567
rect 19111 109449 19202 109567
rect 18902 91727 19202 109449
rect 18902 91609 18993 91727
rect 19111 91609 19202 91727
rect 18902 91567 19202 91609
rect 18902 91449 18993 91567
rect 19111 91449 19202 91567
rect 18902 73727 19202 91449
rect 18902 73609 18993 73727
rect 19111 73609 19202 73727
rect 18902 73567 19202 73609
rect 18902 73449 18993 73567
rect 19111 73449 19202 73567
rect 18902 55727 19202 73449
rect 18902 55609 18993 55727
rect 19111 55609 19202 55727
rect 18902 55567 19202 55609
rect 18902 55449 18993 55567
rect 19111 55449 19202 55567
rect 18902 37727 19202 55449
rect 18902 37609 18993 37727
rect 19111 37609 19202 37727
rect 18902 37567 19202 37609
rect 18902 37449 18993 37567
rect 19111 37449 19202 37567
rect 18902 19727 19202 37449
rect 18902 19609 18993 19727
rect 19111 19609 19202 19727
rect 18902 19567 19202 19609
rect 18902 19449 18993 19567
rect 19111 19449 19202 19567
rect 18902 1727 19202 19449
rect 18902 1609 18993 1727
rect 19111 1609 19202 1727
rect 18902 1567 19202 1609
rect 18902 1449 18993 1567
rect 19111 1449 19202 1567
rect 18902 -173 19202 1449
rect 18902 -291 18993 -173
rect 19111 -291 19202 -173
rect 18902 -333 19202 -291
rect 18902 -451 18993 -333
rect 19111 -451 19202 -333
rect 18902 -932 19202 -451
rect 20702 345527 21002 353081
rect 20702 345409 20793 345527
rect 20911 345409 21002 345527
rect 20702 345367 21002 345409
rect 20702 345249 20793 345367
rect 20911 345249 21002 345367
rect 20702 327527 21002 345249
rect 20702 327409 20793 327527
rect 20911 327409 21002 327527
rect 20702 327367 21002 327409
rect 20702 327249 20793 327367
rect 20911 327249 21002 327367
rect 20702 309527 21002 327249
rect 20702 309409 20793 309527
rect 20911 309409 21002 309527
rect 20702 309367 21002 309409
rect 20702 309249 20793 309367
rect 20911 309249 21002 309367
rect 20702 291527 21002 309249
rect 20702 291409 20793 291527
rect 20911 291409 21002 291527
rect 20702 291367 21002 291409
rect 20702 291249 20793 291367
rect 20911 291249 21002 291367
rect 20702 273527 21002 291249
rect 20702 273409 20793 273527
rect 20911 273409 21002 273527
rect 20702 273367 21002 273409
rect 20702 273249 20793 273367
rect 20911 273249 21002 273367
rect 20702 255527 21002 273249
rect 20702 255409 20793 255527
rect 20911 255409 21002 255527
rect 20702 255367 21002 255409
rect 20702 255249 20793 255367
rect 20911 255249 21002 255367
rect 20702 237527 21002 255249
rect 20702 237409 20793 237527
rect 20911 237409 21002 237527
rect 20702 237367 21002 237409
rect 20702 237249 20793 237367
rect 20911 237249 21002 237367
rect 20702 219527 21002 237249
rect 20702 219409 20793 219527
rect 20911 219409 21002 219527
rect 20702 219367 21002 219409
rect 20702 219249 20793 219367
rect 20911 219249 21002 219367
rect 20702 201527 21002 219249
rect 20702 201409 20793 201527
rect 20911 201409 21002 201527
rect 20702 201367 21002 201409
rect 20702 201249 20793 201367
rect 20911 201249 21002 201367
rect 20702 183527 21002 201249
rect 20702 183409 20793 183527
rect 20911 183409 21002 183527
rect 20702 183367 21002 183409
rect 20702 183249 20793 183367
rect 20911 183249 21002 183367
rect 20702 165527 21002 183249
rect 20702 165409 20793 165527
rect 20911 165409 21002 165527
rect 20702 165367 21002 165409
rect 20702 165249 20793 165367
rect 20911 165249 21002 165367
rect 20702 147527 21002 165249
rect 20702 147409 20793 147527
rect 20911 147409 21002 147527
rect 20702 147367 21002 147409
rect 20702 147249 20793 147367
rect 20911 147249 21002 147367
rect 20702 129527 21002 147249
rect 20702 129409 20793 129527
rect 20911 129409 21002 129527
rect 20702 129367 21002 129409
rect 20702 129249 20793 129367
rect 20911 129249 21002 129367
rect 20702 111527 21002 129249
rect 20702 111409 20793 111527
rect 20911 111409 21002 111527
rect 20702 111367 21002 111409
rect 20702 111249 20793 111367
rect 20911 111249 21002 111367
rect 20702 93527 21002 111249
rect 20702 93409 20793 93527
rect 20911 93409 21002 93527
rect 20702 93367 21002 93409
rect 20702 93249 20793 93367
rect 20911 93249 21002 93367
rect 20702 75527 21002 93249
rect 20702 75409 20793 75527
rect 20911 75409 21002 75527
rect 20702 75367 21002 75409
rect 20702 75249 20793 75367
rect 20911 75249 21002 75367
rect 20702 57527 21002 75249
rect 20702 57409 20793 57527
rect 20911 57409 21002 57527
rect 20702 57367 21002 57409
rect 20702 57249 20793 57367
rect 20911 57249 21002 57367
rect 20702 39527 21002 57249
rect 20702 39409 20793 39527
rect 20911 39409 21002 39527
rect 20702 39367 21002 39409
rect 20702 39249 20793 39367
rect 20911 39249 21002 39367
rect 20702 21527 21002 39249
rect 20702 21409 20793 21527
rect 20911 21409 21002 21527
rect 20702 21367 21002 21409
rect 20702 21249 20793 21367
rect 20911 21249 21002 21367
rect 20702 3527 21002 21249
rect 20702 3409 20793 3527
rect 20911 3409 21002 3527
rect 20702 3367 21002 3409
rect 20702 3249 20793 3367
rect 20911 3249 21002 3367
rect 20702 -1113 21002 3249
rect 20702 -1231 20793 -1113
rect 20911 -1231 21002 -1113
rect 20702 -1273 21002 -1231
rect 20702 -1391 20793 -1273
rect 20911 -1391 21002 -1273
rect 20702 -1872 21002 -1391
rect 22502 347327 22802 354021
rect 22502 347209 22593 347327
rect 22711 347209 22802 347327
rect 22502 347167 22802 347209
rect 22502 347049 22593 347167
rect 22711 347049 22802 347167
rect 22502 329327 22802 347049
rect 22502 329209 22593 329327
rect 22711 329209 22802 329327
rect 22502 329167 22802 329209
rect 22502 329049 22593 329167
rect 22711 329049 22802 329167
rect 22502 311327 22802 329049
rect 22502 311209 22593 311327
rect 22711 311209 22802 311327
rect 22502 311167 22802 311209
rect 22502 311049 22593 311167
rect 22711 311049 22802 311167
rect 22502 293327 22802 311049
rect 22502 293209 22593 293327
rect 22711 293209 22802 293327
rect 22502 293167 22802 293209
rect 22502 293049 22593 293167
rect 22711 293049 22802 293167
rect 22502 275327 22802 293049
rect 22502 275209 22593 275327
rect 22711 275209 22802 275327
rect 22502 275167 22802 275209
rect 22502 275049 22593 275167
rect 22711 275049 22802 275167
rect 22502 257327 22802 275049
rect 22502 257209 22593 257327
rect 22711 257209 22802 257327
rect 22502 257167 22802 257209
rect 22502 257049 22593 257167
rect 22711 257049 22802 257167
rect 22502 239327 22802 257049
rect 22502 239209 22593 239327
rect 22711 239209 22802 239327
rect 22502 239167 22802 239209
rect 22502 239049 22593 239167
rect 22711 239049 22802 239167
rect 22502 221327 22802 239049
rect 22502 221209 22593 221327
rect 22711 221209 22802 221327
rect 22502 221167 22802 221209
rect 22502 221049 22593 221167
rect 22711 221049 22802 221167
rect 22502 203327 22802 221049
rect 22502 203209 22593 203327
rect 22711 203209 22802 203327
rect 22502 203167 22802 203209
rect 22502 203049 22593 203167
rect 22711 203049 22802 203167
rect 22502 185327 22802 203049
rect 22502 185209 22593 185327
rect 22711 185209 22802 185327
rect 22502 185167 22802 185209
rect 22502 185049 22593 185167
rect 22711 185049 22802 185167
rect 22502 167327 22802 185049
rect 22502 167209 22593 167327
rect 22711 167209 22802 167327
rect 22502 167167 22802 167209
rect 22502 167049 22593 167167
rect 22711 167049 22802 167167
rect 22502 149327 22802 167049
rect 22502 149209 22593 149327
rect 22711 149209 22802 149327
rect 22502 149167 22802 149209
rect 22502 149049 22593 149167
rect 22711 149049 22802 149167
rect 22502 131327 22802 149049
rect 22502 131209 22593 131327
rect 22711 131209 22802 131327
rect 22502 131167 22802 131209
rect 22502 131049 22593 131167
rect 22711 131049 22802 131167
rect 22502 113327 22802 131049
rect 22502 113209 22593 113327
rect 22711 113209 22802 113327
rect 22502 113167 22802 113209
rect 22502 113049 22593 113167
rect 22711 113049 22802 113167
rect 22502 95327 22802 113049
rect 22502 95209 22593 95327
rect 22711 95209 22802 95327
rect 22502 95167 22802 95209
rect 22502 95049 22593 95167
rect 22711 95049 22802 95167
rect 22502 77327 22802 95049
rect 22502 77209 22593 77327
rect 22711 77209 22802 77327
rect 22502 77167 22802 77209
rect 22502 77049 22593 77167
rect 22711 77049 22802 77167
rect 22502 59327 22802 77049
rect 22502 59209 22593 59327
rect 22711 59209 22802 59327
rect 22502 59167 22802 59209
rect 22502 59049 22593 59167
rect 22711 59049 22802 59167
rect 22502 41327 22802 59049
rect 22502 41209 22593 41327
rect 22711 41209 22802 41327
rect 22502 41167 22802 41209
rect 22502 41049 22593 41167
rect 22711 41049 22802 41167
rect 22502 23327 22802 41049
rect 22502 23209 22593 23327
rect 22711 23209 22802 23327
rect 22502 23167 22802 23209
rect 22502 23049 22593 23167
rect 22711 23049 22802 23167
rect 22502 5327 22802 23049
rect 22502 5209 22593 5327
rect 22711 5209 22802 5327
rect 22502 5167 22802 5209
rect 22502 5049 22593 5167
rect 22711 5049 22802 5167
rect 22502 -2053 22802 5049
rect 22502 -2171 22593 -2053
rect 22711 -2171 22802 -2053
rect 22502 -2213 22802 -2171
rect 22502 -2331 22593 -2213
rect 22711 -2331 22802 -2213
rect 22502 -2812 22802 -2331
rect 24302 349127 24602 354961
rect 33302 355709 33602 355720
rect 33302 355591 33393 355709
rect 33511 355591 33602 355709
rect 33302 355549 33602 355591
rect 33302 355431 33393 355549
rect 33511 355431 33602 355549
rect 31502 354769 31802 354780
rect 31502 354651 31593 354769
rect 31711 354651 31802 354769
rect 31502 354609 31802 354651
rect 31502 354491 31593 354609
rect 31711 354491 31802 354609
rect 29702 353829 30002 353840
rect 29702 353711 29793 353829
rect 29911 353711 30002 353829
rect 29702 353669 30002 353711
rect 29702 353551 29793 353669
rect 29911 353551 30002 353669
rect 24302 349009 24393 349127
rect 24511 349009 24602 349127
rect 24302 348967 24602 349009
rect 24302 348849 24393 348967
rect 24511 348849 24602 348967
rect 24302 331127 24602 348849
rect 24302 331009 24393 331127
rect 24511 331009 24602 331127
rect 24302 330967 24602 331009
rect 24302 330849 24393 330967
rect 24511 330849 24602 330967
rect 24302 313127 24602 330849
rect 24302 313009 24393 313127
rect 24511 313009 24602 313127
rect 24302 312967 24602 313009
rect 24302 312849 24393 312967
rect 24511 312849 24602 312967
rect 24302 295127 24602 312849
rect 24302 295009 24393 295127
rect 24511 295009 24602 295127
rect 24302 294967 24602 295009
rect 24302 294849 24393 294967
rect 24511 294849 24602 294967
rect 24302 277127 24602 294849
rect 24302 277009 24393 277127
rect 24511 277009 24602 277127
rect 24302 276967 24602 277009
rect 24302 276849 24393 276967
rect 24511 276849 24602 276967
rect 24302 259127 24602 276849
rect 24302 259009 24393 259127
rect 24511 259009 24602 259127
rect 24302 258967 24602 259009
rect 24302 258849 24393 258967
rect 24511 258849 24602 258967
rect 24302 241127 24602 258849
rect 24302 241009 24393 241127
rect 24511 241009 24602 241127
rect 24302 240967 24602 241009
rect 24302 240849 24393 240967
rect 24511 240849 24602 240967
rect 24302 223127 24602 240849
rect 24302 223009 24393 223127
rect 24511 223009 24602 223127
rect 24302 222967 24602 223009
rect 24302 222849 24393 222967
rect 24511 222849 24602 222967
rect 24302 205127 24602 222849
rect 24302 205009 24393 205127
rect 24511 205009 24602 205127
rect 24302 204967 24602 205009
rect 24302 204849 24393 204967
rect 24511 204849 24602 204967
rect 24302 187127 24602 204849
rect 24302 187009 24393 187127
rect 24511 187009 24602 187127
rect 24302 186967 24602 187009
rect 24302 186849 24393 186967
rect 24511 186849 24602 186967
rect 24302 169127 24602 186849
rect 24302 169009 24393 169127
rect 24511 169009 24602 169127
rect 24302 168967 24602 169009
rect 24302 168849 24393 168967
rect 24511 168849 24602 168967
rect 24302 151127 24602 168849
rect 24302 151009 24393 151127
rect 24511 151009 24602 151127
rect 24302 150967 24602 151009
rect 24302 150849 24393 150967
rect 24511 150849 24602 150967
rect 24302 133127 24602 150849
rect 24302 133009 24393 133127
rect 24511 133009 24602 133127
rect 24302 132967 24602 133009
rect 24302 132849 24393 132967
rect 24511 132849 24602 132967
rect 24302 115127 24602 132849
rect 24302 115009 24393 115127
rect 24511 115009 24602 115127
rect 24302 114967 24602 115009
rect 24302 114849 24393 114967
rect 24511 114849 24602 114967
rect 24302 97127 24602 114849
rect 24302 97009 24393 97127
rect 24511 97009 24602 97127
rect 24302 96967 24602 97009
rect 24302 96849 24393 96967
rect 24511 96849 24602 96967
rect 24302 79127 24602 96849
rect 24302 79009 24393 79127
rect 24511 79009 24602 79127
rect 24302 78967 24602 79009
rect 24302 78849 24393 78967
rect 24511 78849 24602 78967
rect 24302 61127 24602 78849
rect 24302 61009 24393 61127
rect 24511 61009 24602 61127
rect 24302 60967 24602 61009
rect 24302 60849 24393 60967
rect 24511 60849 24602 60967
rect 24302 43127 24602 60849
rect 24302 43009 24393 43127
rect 24511 43009 24602 43127
rect 24302 42967 24602 43009
rect 24302 42849 24393 42967
rect 24511 42849 24602 42967
rect 24302 25127 24602 42849
rect 24302 25009 24393 25127
rect 24511 25009 24602 25127
rect 24302 24967 24602 25009
rect 24302 24849 24393 24967
rect 24511 24849 24602 24967
rect 24302 7127 24602 24849
rect 24302 7009 24393 7127
rect 24511 7009 24602 7127
rect 24302 6967 24602 7009
rect 24302 6849 24393 6967
rect 24511 6849 24602 6967
rect 15302 -3581 15393 -3463
rect 15511 -3581 15602 -3463
rect 15302 -3623 15602 -3581
rect 15302 -3741 15393 -3623
rect 15511 -3741 15602 -3623
rect 15302 -3752 15602 -3741
rect 24302 -2993 24602 6849
rect 27902 352889 28202 352900
rect 27902 352771 27993 352889
rect 28111 352771 28202 352889
rect 27902 352729 28202 352771
rect 27902 352611 27993 352729
rect 28111 352611 28202 352729
rect 27902 334727 28202 352611
rect 27902 334609 27993 334727
rect 28111 334609 28202 334727
rect 27902 334567 28202 334609
rect 27902 334449 27993 334567
rect 28111 334449 28202 334567
rect 27902 316727 28202 334449
rect 27902 316609 27993 316727
rect 28111 316609 28202 316727
rect 27902 316567 28202 316609
rect 27902 316449 27993 316567
rect 28111 316449 28202 316567
rect 27902 298727 28202 316449
rect 27902 298609 27993 298727
rect 28111 298609 28202 298727
rect 27902 298567 28202 298609
rect 27902 298449 27993 298567
rect 28111 298449 28202 298567
rect 27902 280727 28202 298449
rect 27902 280609 27993 280727
rect 28111 280609 28202 280727
rect 27902 280567 28202 280609
rect 27902 280449 27993 280567
rect 28111 280449 28202 280567
rect 27902 262727 28202 280449
rect 27902 262609 27993 262727
rect 28111 262609 28202 262727
rect 27902 262567 28202 262609
rect 27902 262449 27993 262567
rect 28111 262449 28202 262567
rect 27902 244727 28202 262449
rect 27902 244609 27993 244727
rect 28111 244609 28202 244727
rect 27902 244567 28202 244609
rect 27902 244449 27993 244567
rect 28111 244449 28202 244567
rect 27902 226727 28202 244449
rect 27902 226609 27993 226727
rect 28111 226609 28202 226727
rect 27902 226567 28202 226609
rect 27902 226449 27993 226567
rect 28111 226449 28202 226567
rect 27902 208727 28202 226449
rect 27902 208609 27993 208727
rect 28111 208609 28202 208727
rect 27902 208567 28202 208609
rect 27902 208449 27993 208567
rect 28111 208449 28202 208567
rect 27902 190727 28202 208449
rect 27902 190609 27993 190727
rect 28111 190609 28202 190727
rect 27902 190567 28202 190609
rect 27902 190449 27993 190567
rect 28111 190449 28202 190567
rect 27902 172727 28202 190449
rect 27902 172609 27993 172727
rect 28111 172609 28202 172727
rect 27902 172567 28202 172609
rect 27902 172449 27993 172567
rect 28111 172449 28202 172567
rect 27902 154727 28202 172449
rect 27902 154609 27993 154727
rect 28111 154609 28202 154727
rect 27902 154567 28202 154609
rect 27902 154449 27993 154567
rect 28111 154449 28202 154567
rect 27902 136727 28202 154449
rect 27902 136609 27993 136727
rect 28111 136609 28202 136727
rect 27902 136567 28202 136609
rect 27902 136449 27993 136567
rect 28111 136449 28202 136567
rect 27902 118727 28202 136449
rect 27902 118609 27993 118727
rect 28111 118609 28202 118727
rect 27902 118567 28202 118609
rect 27902 118449 27993 118567
rect 28111 118449 28202 118567
rect 27902 100727 28202 118449
rect 27902 100609 27993 100727
rect 28111 100609 28202 100727
rect 27902 100567 28202 100609
rect 27902 100449 27993 100567
rect 28111 100449 28202 100567
rect 27902 82727 28202 100449
rect 27902 82609 27993 82727
rect 28111 82609 28202 82727
rect 27902 82567 28202 82609
rect 27902 82449 27993 82567
rect 28111 82449 28202 82567
rect 27902 64727 28202 82449
rect 27902 64609 27993 64727
rect 28111 64609 28202 64727
rect 27902 64567 28202 64609
rect 27902 64449 27993 64567
rect 28111 64449 28202 64567
rect 27902 46727 28202 64449
rect 27902 46609 27993 46727
rect 28111 46609 28202 46727
rect 27902 46567 28202 46609
rect 27902 46449 27993 46567
rect 28111 46449 28202 46567
rect 27902 28727 28202 46449
rect 27902 28609 27993 28727
rect 28111 28609 28202 28727
rect 27902 28567 28202 28609
rect 27902 28449 27993 28567
rect 28111 28449 28202 28567
rect 27902 10727 28202 28449
rect 27902 10609 27993 10727
rect 28111 10609 28202 10727
rect 27902 10567 28202 10609
rect 27902 10449 27993 10567
rect 28111 10449 28202 10567
rect 27902 -643 28202 10449
rect 27902 -761 27993 -643
rect 28111 -761 28202 -643
rect 27902 -803 28202 -761
rect 27902 -921 27993 -803
rect 28111 -921 28202 -803
rect 27902 -932 28202 -921
rect 29702 336527 30002 353551
rect 29702 336409 29793 336527
rect 29911 336409 30002 336527
rect 29702 336367 30002 336409
rect 29702 336249 29793 336367
rect 29911 336249 30002 336367
rect 29702 318527 30002 336249
rect 29702 318409 29793 318527
rect 29911 318409 30002 318527
rect 29702 318367 30002 318409
rect 29702 318249 29793 318367
rect 29911 318249 30002 318367
rect 29702 300527 30002 318249
rect 29702 300409 29793 300527
rect 29911 300409 30002 300527
rect 29702 300367 30002 300409
rect 29702 300249 29793 300367
rect 29911 300249 30002 300367
rect 29702 282527 30002 300249
rect 29702 282409 29793 282527
rect 29911 282409 30002 282527
rect 29702 282367 30002 282409
rect 29702 282249 29793 282367
rect 29911 282249 30002 282367
rect 29702 264527 30002 282249
rect 29702 264409 29793 264527
rect 29911 264409 30002 264527
rect 29702 264367 30002 264409
rect 29702 264249 29793 264367
rect 29911 264249 30002 264367
rect 29702 246527 30002 264249
rect 29702 246409 29793 246527
rect 29911 246409 30002 246527
rect 29702 246367 30002 246409
rect 29702 246249 29793 246367
rect 29911 246249 30002 246367
rect 29702 228527 30002 246249
rect 29702 228409 29793 228527
rect 29911 228409 30002 228527
rect 29702 228367 30002 228409
rect 29702 228249 29793 228367
rect 29911 228249 30002 228367
rect 29702 210527 30002 228249
rect 29702 210409 29793 210527
rect 29911 210409 30002 210527
rect 29702 210367 30002 210409
rect 29702 210249 29793 210367
rect 29911 210249 30002 210367
rect 29702 192527 30002 210249
rect 29702 192409 29793 192527
rect 29911 192409 30002 192527
rect 29702 192367 30002 192409
rect 29702 192249 29793 192367
rect 29911 192249 30002 192367
rect 29702 174527 30002 192249
rect 29702 174409 29793 174527
rect 29911 174409 30002 174527
rect 29702 174367 30002 174409
rect 29702 174249 29793 174367
rect 29911 174249 30002 174367
rect 29702 156527 30002 174249
rect 29702 156409 29793 156527
rect 29911 156409 30002 156527
rect 29702 156367 30002 156409
rect 29702 156249 29793 156367
rect 29911 156249 30002 156367
rect 29702 138527 30002 156249
rect 29702 138409 29793 138527
rect 29911 138409 30002 138527
rect 29702 138367 30002 138409
rect 29702 138249 29793 138367
rect 29911 138249 30002 138367
rect 29702 120527 30002 138249
rect 29702 120409 29793 120527
rect 29911 120409 30002 120527
rect 29702 120367 30002 120409
rect 29702 120249 29793 120367
rect 29911 120249 30002 120367
rect 29702 102527 30002 120249
rect 29702 102409 29793 102527
rect 29911 102409 30002 102527
rect 29702 102367 30002 102409
rect 29702 102249 29793 102367
rect 29911 102249 30002 102367
rect 29702 84527 30002 102249
rect 29702 84409 29793 84527
rect 29911 84409 30002 84527
rect 29702 84367 30002 84409
rect 29702 84249 29793 84367
rect 29911 84249 30002 84367
rect 29702 66527 30002 84249
rect 29702 66409 29793 66527
rect 29911 66409 30002 66527
rect 29702 66367 30002 66409
rect 29702 66249 29793 66367
rect 29911 66249 30002 66367
rect 29702 48527 30002 66249
rect 29702 48409 29793 48527
rect 29911 48409 30002 48527
rect 29702 48367 30002 48409
rect 29702 48249 29793 48367
rect 29911 48249 30002 48367
rect 29702 30527 30002 48249
rect 29702 30409 29793 30527
rect 29911 30409 30002 30527
rect 29702 30367 30002 30409
rect 29702 30249 29793 30367
rect 29911 30249 30002 30367
rect 29702 12527 30002 30249
rect 29702 12409 29793 12527
rect 29911 12409 30002 12527
rect 29702 12367 30002 12409
rect 29702 12249 29793 12367
rect 29911 12249 30002 12367
rect 29702 -1583 30002 12249
rect 29702 -1701 29793 -1583
rect 29911 -1701 30002 -1583
rect 29702 -1743 30002 -1701
rect 29702 -1861 29793 -1743
rect 29911 -1861 30002 -1743
rect 29702 -1872 30002 -1861
rect 31502 338327 31802 354491
rect 31502 338209 31593 338327
rect 31711 338209 31802 338327
rect 31502 338167 31802 338209
rect 31502 338049 31593 338167
rect 31711 338049 31802 338167
rect 31502 320327 31802 338049
rect 31502 320209 31593 320327
rect 31711 320209 31802 320327
rect 31502 320167 31802 320209
rect 31502 320049 31593 320167
rect 31711 320049 31802 320167
rect 31502 302327 31802 320049
rect 31502 302209 31593 302327
rect 31711 302209 31802 302327
rect 31502 302167 31802 302209
rect 31502 302049 31593 302167
rect 31711 302049 31802 302167
rect 31502 284327 31802 302049
rect 31502 284209 31593 284327
rect 31711 284209 31802 284327
rect 31502 284167 31802 284209
rect 31502 284049 31593 284167
rect 31711 284049 31802 284167
rect 31502 266327 31802 284049
rect 31502 266209 31593 266327
rect 31711 266209 31802 266327
rect 31502 266167 31802 266209
rect 31502 266049 31593 266167
rect 31711 266049 31802 266167
rect 31502 248327 31802 266049
rect 31502 248209 31593 248327
rect 31711 248209 31802 248327
rect 31502 248167 31802 248209
rect 31502 248049 31593 248167
rect 31711 248049 31802 248167
rect 31502 230327 31802 248049
rect 31502 230209 31593 230327
rect 31711 230209 31802 230327
rect 31502 230167 31802 230209
rect 31502 230049 31593 230167
rect 31711 230049 31802 230167
rect 31502 212327 31802 230049
rect 31502 212209 31593 212327
rect 31711 212209 31802 212327
rect 31502 212167 31802 212209
rect 31502 212049 31593 212167
rect 31711 212049 31802 212167
rect 31502 194327 31802 212049
rect 31502 194209 31593 194327
rect 31711 194209 31802 194327
rect 31502 194167 31802 194209
rect 31502 194049 31593 194167
rect 31711 194049 31802 194167
rect 31502 176327 31802 194049
rect 31502 176209 31593 176327
rect 31711 176209 31802 176327
rect 31502 176167 31802 176209
rect 31502 176049 31593 176167
rect 31711 176049 31802 176167
rect 31502 158327 31802 176049
rect 31502 158209 31593 158327
rect 31711 158209 31802 158327
rect 31502 158167 31802 158209
rect 31502 158049 31593 158167
rect 31711 158049 31802 158167
rect 31502 140327 31802 158049
rect 31502 140209 31593 140327
rect 31711 140209 31802 140327
rect 31502 140167 31802 140209
rect 31502 140049 31593 140167
rect 31711 140049 31802 140167
rect 31502 122327 31802 140049
rect 31502 122209 31593 122327
rect 31711 122209 31802 122327
rect 31502 122167 31802 122209
rect 31502 122049 31593 122167
rect 31711 122049 31802 122167
rect 31502 104327 31802 122049
rect 31502 104209 31593 104327
rect 31711 104209 31802 104327
rect 31502 104167 31802 104209
rect 31502 104049 31593 104167
rect 31711 104049 31802 104167
rect 31502 86327 31802 104049
rect 31502 86209 31593 86327
rect 31711 86209 31802 86327
rect 31502 86167 31802 86209
rect 31502 86049 31593 86167
rect 31711 86049 31802 86167
rect 31502 68327 31802 86049
rect 31502 68209 31593 68327
rect 31711 68209 31802 68327
rect 31502 68167 31802 68209
rect 31502 68049 31593 68167
rect 31711 68049 31802 68167
rect 31502 50327 31802 68049
rect 31502 50209 31593 50327
rect 31711 50209 31802 50327
rect 31502 50167 31802 50209
rect 31502 50049 31593 50167
rect 31711 50049 31802 50167
rect 31502 32327 31802 50049
rect 31502 32209 31593 32327
rect 31711 32209 31802 32327
rect 31502 32167 31802 32209
rect 31502 32049 31593 32167
rect 31711 32049 31802 32167
rect 31502 14327 31802 32049
rect 31502 14209 31593 14327
rect 31711 14209 31802 14327
rect 31502 14167 31802 14209
rect 31502 14049 31593 14167
rect 31711 14049 31802 14167
rect 31502 -2523 31802 14049
rect 31502 -2641 31593 -2523
rect 31711 -2641 31802 -2523
rect 31502 -2683 31802 -2641
rect 31502 -2801 31593 -2683
rect 31711 -2801 31802 -2683
rect 31502 -2812 31802 -2801
rect 33302 340127 33602 355431
rect 42302 355239 42602 355720
rect 42302 355121 42393 355239
rect 42511 355121 42602 355239
rect 42302 355079 42602 355121
rect 42302 354961 42393 355079
rect 42511 354961 42602 355079
rect 40502 354299 40802 354780
rect 40502 354181 40593 354299
rect 40711 354181 40802 354299
rect 40502 354139 40802 354181
rect 40502 354021 40593 354139
rect 40711 354021 40802 354139
rect 38702 353359 39002 353840
rect 38702 353241 38793 353359
rect 38911 353241 39002 353359
rect 38702 353199 39002 353241
rect 38702 353081 38793 353199
rect 38911 353081 39002 353199
rect 33302 340009 33393 340127
rect 33511 340009 33602 340127
rect 33302 339967 33602 340009
rect 33302 339849 33393 339967
rect 33511 339849 33602 339967
rect 33302 322127 33602 339849
rect 33302 322009 33393 322127
rect 33511 322009 33602 322127
rect 33302 321967 33602 322009
rect 33302 321849 33393 321967
rect 33511 321849 33602 321967
rect 33302 304127 33602 321849
rect 33302 304009 33393 304127
rect 33511 304009 33602 304127
rect 33302 303967 33602 304009
rect 33302 303849 33393 303967
rect 33511 303849 33602 303967
rect 33302 286127 33602 303849
rect 33302 286009 33393 286127
rect 33511 286009 33602 286127
rect 33302 285967 33602 286009
rect 33302 285849 33393 285967
rect 33511 285849 33602 285967
rect 33302 268127 33602 285849
rect 33302 268009 33393 268127
rect 33511 268009 33602 268127
rect 33302 267967 33602 268009
rect 33302 267849 33393 267967
rect 33511 267849 33602 267967
rect 33302 250127 33602 267849
rect 33302 250009 33393 250127
rect 33511 250009 33602 250127
rect 33302 249967 33602 250009
rect 33302 249849 33393 249967
rect 33511 249849 33602 249967
rect 33302 232127 33602 249849
rect 33302 232009 33393 232127
rect 33511 232009 33602 232127
rect 33302 231967 33602 232009
rect 33302 231849 33393 231967
rect 33511 231849 33602 231967
rect 33302 214127 33602 231849
rect 33302 214009 33393 214127
rect 33511 214009 33602 214127
rect 33302 213967 33602 214009
rect 33302 213849 33393 213967
rect 33511 213849 33602 213967
rect 33302 196127 33602 213849
rect 33302 196009 33393 196127
rect 33511 196009 33602 196127
rect 33302 195967 33602 196009
rect 33302 195849 33393 195967
rect 33511 195849 33602 195967
rect 33302 178127 33602 195849
rect 33302 178009 33393 178127
rect 33511 178009 33602 178127
rect 33302 177967 33602 178009
rect 33302 177849 33393 177967
rect 33511 177849 33602 177967
rect 33302 160127 33602 177849
rect 33302 160009 33393 160127
rect 33511 160009 33602 160127
rect 33302 159967 33602 160009
rect 33302 159849 33393 159967
rect 33511 159849 33602 159967
rect 33302 142127 33602 159849
rect 33302 142009 33393 142127
rect 33511 142009 33602 142127
rect 33302 141967 33602 142009
rect 33302 141849 33393 141967
rect 33511 141849 33602 141967
rect 33302 124127 33602 141849
rect 33302 124009 33393 124127
rect 33511 124009 33602 124127
rect 33302 123967 33602 124009
rect 33302 123849 33393 123967
rect 33511 123849 33602 123967
rect 33302 106127 33602 123849
rect 33302 106009 33393 106127
rect 33511 106009 33602 106127
rect 33302 105967 33602 106009
rect 33302 105849 33393 105967
rect 33511 105849 33602 105967
rect 33302 88127 33602 105849
rect 33302 88009 33393 88127
rect 33511 88009 33602 88127
rect 33302 87967 33602 88009
rect 33302 87849 33393 87967
rect 33511 87849 33602 87967
rect 33302 70127 33602 87849
rect 33302 70009 33393 70127
rect 33511 70009 33602 70127
rect 33302 69967 33602 70009
rect 33302 69849 33393 69967
rect 33511 69849 33602 69967
rect 33302 52127 33602 69849
rect 33302 52009 33393 52127
rect 33511 52009 33602 52127
rect 33302 51967 33602 52009
rect 33302 51849 33393 51967
rect 33511 51849 33602 51967
rect 33302 34127 33602 51849
rect 33302 34009 33393 34127
rect 33511 34009 33602 34127
rect 33302 33967 33602 34009
rect 33302 33849 33393 33967
rect 33511 33849 33602 33967
rect 33302 16127 33602 33849
rect 33302 16009 33393 16127
rect 33511 16009 33602 16127
rect 33302 15967 33602 16009
rect 33302 15849 33393 15967
rect 33511 15849 33602 15967
rect 24302 -3111 24393 -2993
rect 24511 -3111 24602 -2993
rect 24302 -3153 24602 -3111
rect 24302 -3271 24393 -3153
rect 24511 -3271 24602 -3153
rect 24302 -3752 24602 -3271
rect 33302 -3463 33602 15849
rect 36902 352419 37202 352900
rect 36902 352301 36993 352419
rect 37111 352301 37202 352419
rect 36902 352259 37202 352301
rect 36902 352141 36993 352259
rect 37111 352141 37202 352259
rect 36902 343727 37202 352141
rect 36902 343609 36993 343727
rect 37111 343609 37202 343727
rect 36902 343567 37202 343609
rect 36902 343449 36993 343567
rect 37111 343449 37202 343567
rect 36902 325727 37202 343449
rect 36902 325609 36993 325727
rect 37111 325609 37202 325727
rect 36902 325567 37202 325609
rect 36902 325449 36993 325567
rect 37111 325449 37202 325567
rect 36902 307727 37202 325449
rect 36902 307609 36993 307727
rect 37111 307609 37202 307727
rect 36902 307567 37202 307609
rect 36902 307449 36993 307567
rect 37111 307449 37202 307567
rect 36902 289727 37202 307449
rect 36902 289609 36993 289727
rect 37111 289609 37202 289727
rect 36902 289567 37202 289609
rect 36902 289449 36993 289567
rect 37111 289449 37202 289567
rect 36902 271727 37202 289449
rect 36902 271609 36993 271727
rect 37111 271609 37202 271727
rect 36902 271567 37202 271609
rect 36902 271449 36993 271567
rect 37111 271449 37202 271567
rect 36902 253727 37202 271449
rect 36902 253609 36993 253727
rect 37111 253609 37202 253727
rect 36902 253567 37202 253609
rect 36902 253449 36993 253567
rect 37111 253449 37202 253567
rect 36902 235727 37202 253449
rect 36902 235609 36993 235727
rect 37111 235609 37202 235727
rect 36902 235567 37202 235609
rect 36902 235449 36993 235567
rect 37111 235449 37202 235567
rect 36902 217727 37202 235449
rect 36902 217609 36993 217727
rect 37111 217609 37202 217727
rect 36902 217567 37202 217609
rect 36902 217449 36993 217567
rect 37111 217449 37202 217567
rect 36902 199727 37202 217449
rect 36902 199609 36993 199727
rect 37111 199609 37202 199727
rect 36902 199567 37202 199609
rect 36902 199449 36993 199567
rect 37111 199449 37202 199567
rect 36902 181727 37202 199449
rect 36902 181609 36993 181727
rect 37111 181609 37202 181727
rect 36902 181567 37202 181609
rect 36902 181449 36993 181567
rect 37111 181449 37202 181567
rect 36902 163727 37202 181449
rect 36902 163609 36993 163727
rect 37111 163609 37202 163727
rect 36902 163567 37202 163609
rect 36902 163449 36993 163567
rect 37111 163449 37202 163567
rect 36902 145727 37202 163449
rect 36902 145609 36993 145727
rect 37111 145609 37202 145727
rect 36902 145567 37202 145609
rect 36902 145449 36993 145567
rect 37111 145449 37202 145567
rect 36902 127727 37202 145449
rect 36902 127609 36993 127727
rect 37111 127609 37202 127727
rect 36902 127567 37202 127609
rect 36902 127449 36993 127567
rect 37111 127449 37202 127567
rect 36902 109727 37202 127449
rect 36902 109609 36993 109727
rect 37111 109609 37202 109727
rect 36902 109567 37202 109609
rect 36902 109449 36993 109567
rect 37111 109449 37202 109567
rect 36902 91727 37202 109449
rect 36902 91609 36993 91727
rect 37111 91609 37202 91727
rect 36902 91567 37202 91609
rect 36902 91449 36993 91567
rect 37111 91449 37202 91567
rect 36902 73727 37202 91449
rect 36902 73609 36993 73727
rect 37111 73609 37202 73727
rect 36902 73567 37202 73609
rect 36902 73449 36993 73567
rect 37111 73449 37202 73567
rect 36902 55727 37202 73449
rect 36902 55609 36993 55727
rect 37111 55609 37202 55727
rect 36902 55567 37202 55609
rect 36902 55449 36993 55567
rect 37111 55449 37202 55567
rect 36902 37727 37202 55449
rect 36902 37609 36993 37727
rect 37111 37609 37202 37727
rect 36902 37567 37202 37609
rect 36902 37449 36993 37567
rect 37111 37449 37202 37567
rect 36902 19727 37202 37449
rect 36902 19609 36993 19727
rect 37111 19609 37202 19727
rect 36902 19567 37202 19609
rect 36902 19449 36993 19567
rect 37111 19449 37202 19567
rect 36902 1727 37202 19449
rect 36902 1609 36993 1727
rect 37111 1609 37202 1727
rect 36902 1567 37202 1609
rect 36902 1449 36993 1567
rect 37111 1449 37202 1567
rect 36902 -173 37202 1449
rect 36902 -291 36993 -173
rect 37111 -291 37202 -173
rect 36902 -333 37202 -291
rect 36902 -451 36993 -333
rect 37111 -451 37202 -333
rect 36902 -932 37202 -451
rect 38702 345527 39002 353081
rect 38702 345409 38793 345527
rect 38911 345409 39002 345527
rect 38702 345367 39002 345409
rect 38702 345249 38793 345367
rect 38911 345249 39002 345367
rect 38702 327527 39002 345249
rect 38702 327409 38793 327527
rect 38911 327409 39002 327527
rect 38702 327367 39002 327409
rect 38702 327249 38793 327367
rect 38911 327249 39002 327367
rect 38702 309527 39002 327249
rect 38702 309409 38793 309527
rect 38911 309409 39002 309527
rect 38702 309367 39002 309409
rect 38702 309249 38793 309367
rect 38911 309249 39002 309367
rect 38702 291527 39002 309249
rect 38702 291409 38793 291527
rect 38911 291409 39002 291527
rect 38702 291367 39002 291409
rect 38702 291249 38793 291367
rect 38911 291249 39002 291367
rect 38702 273527 39002 291249
rect 38702 273409 38793 273527
rect 38911 273409 39002 273527
rect 38702 273367 39002 273409
rect 38702 273249 38793 273367
rect 38911 273249 39002 273367
rect 38702 255527 39002 273249
rect 38702 255409 38793 255527
rect 38911 255409 39002 255527
rect 38702 255367 39002 255409
rect 38702 255249 38793 255367
rect 38911 255249 39002 255367
rect 38702 237527 39002 255249
rect 38702 237409 38793 237527
rect 38911 237409 39002 237527
rect 38702 237367 39002 237409
rect 38702 237249 38793 237367
rect 38911 237249 39002 237367
rect 38702 219527 39002 237249
rect 38702 219409 38793 219527
rect 38911 219409 39002 219527
rect 38702 219367 39002 219409
rect 38702 219249 38793 219367
rect 38911 219249 39002 219367
rect 38702 201527 39002 219249
rect 38702 201409 38793 201527
rect 38911 201409 39002 201527
rect 38702 201367 39002 201409
rect 38702 201249 38793 201367
rect 38911 201249 39002 201367
rect 38702 183527 39002 201249
rect 38702 183409 38793 183527
rect 38911 183409 39002 183527
rect 38702 183367 39002 183409
rect 38702 183249 38793 183367
rect 38911 183249 39002 183367
rect 38702 165527 39002 183249
rect 38702 165409 38793 165527
rect 38911 165409 39002 165527
rect 38702 165367 39002 165409
rect 38702 165249 38793 165367
rect 38911 165249 39002 165367
rect 38702 147527 39002 165249
rect 38702 147409 38793 147527
rect 38911 147409 39002 147527
rect 38702 147367 39002 147409
rect 38702 147249 38793 147367
rect 38911 147249 39002 147367
rect 38702 129527 39002 147249
rect 38702 129409 38793 129527
rect 38911 129409 39002 129527
rect 38702 129367 39002 129409
rect 38702 129249 38793 129367
rect 38911 129249 39002 129367
rect 38702 111527 39002 129249
rect 38702 111409 38793 111527
rect 38911 111409 39002 111527
rect 38702 111367 39002 111409
rect 38702 111249 38793 111367
rect 38911 111249 39002 111367
rect 38702 93527 39002 111249
rect 38702 93409 38793 93527
rect 38911 93409 39002 93527
rect 38702 93367 39002 93409
rect 38702 93249 38793 93367
rect 38911 93249 39002 93367
rect 38702 75527 39002 93249
rect 38702 75409 38793 75527
rect 38911 75409 39002 75527
rect 38702 75367 39002 75409
rect 38702 75249 38793 75367
rect 38911 75249 39002 75367
rect 38702 57527 39002 75249
rect 38702 57409 38793 57527
rect 38911 57409 39002 57527
rect 38702 57367 39002 57409
rect 38702 57249 38793 57367
rect 38911 57249 39002 57367
rect 38702 39527 39002 57249
rect 38702 39409 38793 39527
rect 38911 39409 39002 39527
rect 38702 39367 39002 39409
rect 38702 39249 38793 39367
rect 38911 39249 39002 39367
rect 38702 21527 39002 39249
rect 38702 21409 38793 21527
rect 38911 21409 39002 21527
rect 38702 21367 39002 21409
rect 38702 21249 38793 21367
rect 38911 21249 39002 21367
rect 38702 3527 39002 21249
rect 38702 3409 38793 3527
rect 38911 3409 39002 3527
rect 38702 3367 39002 3409
rect 38702 3249 38793 3367
rect 38911 3249 39002 3367
rect 38702 -1113 39002 3249
rect 38702 -1231 38793 -1113
rect 38911 -1231 39002 -1113
rect 38702 -1273 39002 -1231
rect 38702 -1391 38793 -1273
rect 38911 -1391 39002 -1273
rect 38702 -1872 39002 -1391
rect 40502 347327 40802 354021
rect 40502 347209 40593 347327
rect 40711 347209 40802 347327
rect 40502 347167 40802 347209
rect 40502 347049 40593 347167
rect 40711 347049 40802 347167
rect 40502 329327 40802 347049
rect 40502 329209 40593 329327
rect 40711 329209 40802 329327
rect 40502 329167 40802 329209
rect 40502 329049 40593 329167
rect 40711 329049 40802 329167
rect 40502 311327 40802 329049
rect 40502 311209 40593 311327
rect 40711 311209 40802 311327
rect 40502 311167 40802 311209
rect 40502 311049 40593 311167
rect 40711 311049 40802 311167
rect 40502 293327 40802 311049
rect 40502 293209 40593 293327
rect 40711 293209 40802 293327
rect 40502 293167 40802 293209
rect 40502 293049 40593 293167
rect 40711 293049 40802 293167
rect 40502 275327 40802 293049
rect 40502 275209 40593 275327
rect 40711 275209 40802 275327
rect 40502 275167 40802 275209
rect 40502 275049 40593 275167
rect 40711 275049 40802 275167
rect 40502 257327 40802 275049
rect 40502 257209 40593 257327
rect 40711 257209 40802 257327
rect 40502 257167 40802 257209
rect 40502 257049 40593 257167
rect 40711 257049 40802 257167
rect 40502 239327 40802 257049
rect 40502 239209 40593 239327
rect 40711 239209 40802 239327
rect 40502 239167 40802 239209
rect 40502 239049 40593 239167
rect 40711 239049 40802 239167
rect 40502 221327 40802 239049
rect 40502 221209 40593 221327
rect 40711 221209 40802 221327
rect 40502 221167 40802 221209
rect 40502 221049 40593 221167
rect 40711 221049 40802 221167
rect 40502 203327 40802 221049
rect 40502 203209 40593 203327
rect 40711 203209 40802 203327
rect 40502 203167 40802 203209
rect 40502 203049 40593 203167
rect 40711 203049 40802 203167
rect 40502 185327 40802 203049
rect 40502 185209 40593 185327
rect 40711 185209 40802 185327
rect 40502 185167 40802 185209
rect 40502 185049 40593 185167
rect 40711 185049 40802 185167
rect 40502 167327 40802 185049
rect 40502 167209 40593 167327
rect 40711 167209 40802 167327
rect 40502 167167 40802 167209
rect 40502 167049 40593 167167
rect 40711 167049 40802 167167
rect 40502 149327 40802 167049
rect 40502 149209 40593 149327
rect 40711 149209 40802 149327
rect 40502 149167 40802 149209
rect 40502 149049 40593 149167
rect 40711 149049 40802 149167
rect 40502 131327 40802 149049
rect 40502 131209 40593 131327
rect 40711 131209 40802 131327
rect 40502 131167 40802 131209
rect 40502 131049 40593 131167
rect 40711 131049 40802 131167
rect 40502 113327 40802 131049
rect 40502 113209 40593 113327
rect 40711 113209 40802 113327
rect 40502 113167 40802 113209
rect 40502 113049 40593 113167
rect 40711 113049 40802 113167
rect 40502 95327 40802 113049
rect 40502 95209 40593 95327
rect 40711 95209 40802 95327
rect 40502 95167 40802 95209
rect 40502 95049 40593 95167
rect 40711 95049 40802 95167
rect 40502 77327 40802 95049
rect 40502 77209 40593 77327
rect 40711 77209 40802 77327
rect 40502 77167 40802 77209
rect 40502 77049 40593 77167
rect 40711 77049 40802 77167
rect 40502 59327 40802 77049
rect 40502 59209 40593 59327
rect 40711 59209 40802 59327
rect 40502 59167 40802 59209
rect 40502 59049 40593 59167
rect 40711 59049 40802 59167
rect 40502 41327 40802 59049
rect 40502 41209 40593 41327
rect 40711 41209 40802 41327
rect 40502 41167 40802 41209
rect 40502 41049 40593 41167
rect 40711 41049 40802 41167
rect 40502 23327 40802 41049
rect 40502 23209 40593 23327
rect 40711 23209 40802 23327
rect 40502 23167 40802 23209
rect 40502 23049 40593 23167
rect 40711 23049 40802 23167
rect 40502 5327 40802 23049
rect 40502 5209 40593 5327
rect 40711 5209 40802 5327
rect 40502 5167 40802 5209
rect 40502 5049 40593 5167
rect 40711 5049 40802 5167
rect 40502 -2053 40802 5049
rect 40502 -2171 40593 -2053
rect 40711 -2171 40802 -2053
rect 40502 -2213 40802 -2171
rect 40502 -2331 40593 -2213
rect 40711 -2331 40802 -2213
rect 40502 -2812 40802 -2331
rect 42302 349127 42602 354961
rect 51302 355709 51602 355720
rect 51302 355591 51393 355709
rect 51511 355591 51602 355709
rect 51302 355549 51602 355591
rect 51302 355431 51393 355549
rect 51511 355431 51602 355549
rect 49502 354769 49802 354780
rect 49502 354651 49593 354769
rect 49711 354651 49802 354769
rect 49502 354609 49802 354651
rect 49502 354491 49593 354609
rect 49711 354491 49802 354609
rect 47702 353829 48002 353840
rect 47702 353711 47793 353829
rect 47911 353711 48002 353829
rect 47702 353669 48002 353711
rect 47702 353551 47793 353669
rect 47911 353551 48002 353669
rect 42302 349009 42393 349127
rect 42511 349009 42602 349127
rect 42302 348967 42602 349009
rect 42302 348849 42393 348967
rect 42511 348849 42602 348967
rect 42302 331127 42602 348849
rect 42302 331009 42393 331127
rect 42511 331009 42602 331127
rect 42302 330967 42602 331009
rect 42302 330849 42393 330967
rect 42511 330849 42602 330967
rect 42302 313127 42602 330849
rect 42302 313009 42393 313127
rect 42511 313009 42602 313127
rect 42302 312967 42602 313009
rect 42302 312849 42393 312967
rect 42511 312849 42602 312967
rect 42302 295127 42602 312849
rect 42302 295009 42393 295127
rect 42511 295009 42602 295127
rect 42302 294967 42602 295009
rect 42302 294849 42393 294967
rect 42511 294849 42602 294967
rect 42302 277127 42602 294849
rect 42302 277009 42393 277127
rect 42511 277009 42602 277127
rect 42302 276967 42602 277009
rect 42302 276849 42393 276967
rect 42511 276849 42602 276967
rect 42302 259127 42602 276849
rect 42302 259009 42393 259127
rect 42511 259009 42602 259127
rect 42302 258967 42602 259009
rect 42302 258849 42393 258967
rect 42511 258849 42602 258967
rect 42302 241127 42602 258849
rect 42302 241009 42393 241127
rect 42511 241009 42602 241127
rect 42302 240967 42602 241009
rect 42302 240849 42393 240967
rect 42511 240849 42602 240967
rect 42302 223127 42602 240849
rect 42302 223009 42393 223127
rect 42511 223009 42602 223127
rect 42302 222967 42602 223009
rect 42302 222849 42393 222967
rect 42511 222849 42602 222967
rect 42302 205127 42602 222849
rect 42302 205009 42393 205127
rect 42511 205009 42602 205127
rect 42302 204967 42602 205009
rect 42302 204849 42393 204967
rect 42511 204849 42602 204967
rect 42302 187127 42602 204849
rect 42302 187009 42393 187127
rect 42511 187009 42602 187127
rect 42302 186967 42602 187009
rect 42302 186849 42393 186967
rect 42511 186849 42602 186967
rect 42302 169127 42602 186849
rect 42302 169009 42393 169127
rect 42511 169009 42602 169127
rect 42302 168967 42602 169009
rect 42302 168849 42393 168967
rect 42511 168849 42602 168967
rect 42302 151127 42602 168849
rect 42302 151009 42393 151127
rect 42511 151009 42602 151127
rect 42302 150967 42602 151009
rect 42302 150849 42393 150967
rect 42511 150849 42602 150967
rect 42302 133127 42602 150849
rect 42302 133009 42393 133127
rect 42511 133009 42602 133127
rect 42302 132967 42602 133009
rect 42302 132849 42393 132967
rect 42511 132849 42602 132967
rect 42302 115127 42602 132849
rect 42302 115009 42393 115127
rect 42511 115009 42602 115127
rect 42302 114967 42602 115009
rect 42302 114849 42393 114967
rect 42511 114849 42602 114967
rect 42302 97127 42602 114849
rect 42302 97009 42393 97127
rect 42511 97009 42602 97127
rect 42302 96967 42602 97009
rect 42302 96849 42393 96967
rect 42511 96849 42602 96967
rect 42302 79127 42602 96849
rect 42302 79009 42393 79127
rect 42511 79009 42602 79127
rect 42302 78967 42602 79009
rect 42302 78849 42393 78967
rect 42511 78849 42602 78967
rect 42302 61127 42602 78849
rect 42302 61009 42393 61127
rect 42511 61009 42602 61127
rect 42302 60967 42602 61009
rect 42302 60849 42393 60967
rect 42511 60849 42602 60967
rect 42302 43127 42602 60849
rect 42302 43009 42393 43127
rect 42511 43009 42602 43127
rect 42302 42967 42602 43009
rect 42302 42849 42393 42967
rect 42511 42849 42602 42967
rect 42302 25127 42602 42849
rect 42302 25009 42393 25127
rect 42511 25009 42602 25127
rect 42302 24967 42602 25009
rect 42302 24849 42393 24967
rect 42511 24849 42602 24967
rect 42302 7127 42602 24849
rect 42302 7009 42393 7127
rect 42511 7009 42602 7127
rect 42302 6967 42602 7009
rect 42302 6849 42393 6967
rect 42511 6849 42602 6967
rect 33302 -3581 33393 -3463
rect 33511 -3581 33602 -3463
rect 33302 -3623 33602 -3581
rect 33302 -3741 33393 -3623
rect 33511 -3741 33602 -3623
rect 33302 -3752 33602 -3741
rect 42302 -2993 42602 6849
rect 45902 352889 46202 352900
rect 45902 352771 45993 352889
rect 46111 352771 46202 352889
rect 45902 352729 46202 352771
rect 45902 352611 45993 352729
rect 46111 352611 46202 352729
rect 45902 334727 46202 352611
rect 45902 334609 45993 334727
rect 46111 334609 46202 334727
rect 45902 334567 46202 334609
rect 45902 334449 45993 334567
rect 46111 334449 46202 334567
rect 45902 316727 46202 334449
rect 45902 316609 45993 316727
rect 46111 316609 46202 316727
rect 45902 316567 46202 316609
rect 45902 316449 45993 316567
rect 46111 316449 46202 316567
rect 45902 298727 46202 316449
rect 45902 298609 45993 298727
rect 46111 298609 46202 298727
rect 45902 298567 46202 298609
rect 45902 298449 45993 298567
rect 46111 298449 46202 298567
rect 45902 280727 46202 298449
rect 45902 280609 45993 280727
rect 46111 280609 46202 280727
rect 45902 280567 46202 280609
rect 45902 280449 45993 280567
rect 46111 280449 46202 280567
rect 45902 262727 46202 280449
rect 45902 262609 45993 262727
rect 46111 262609 46202 262727
rect 45902 262567 46202 262609
rect 45902 262449 45993 262567
rect 46111 262449 46202 262567
rect 45902 244727 46202 262449
rect 45902 244609 45993 244727
rect 46111 244609 46202 244727
rect 45902 244567 46202 244609
rect 45902 244449 45993 244567
rect 46111 244449 46202 244567
rect 45902 226727 46202 244449
rect 45902 226609 45993 226727
rect 46111 226609 46202 226727
rect 45902 226567 46202 226609
rect 45902 226449 45993 226567
rect 46111 226449 46202 226567
rect 45902 208727 46202 226449
rect 45902 208609 45993 208727
rect 46111 208609 46202 208727
rect 45902 208567 46202 208609
rect 45902 208449 45993 208567
rect 46111 208449 46202 208567
rect 45902 190727 46202 208449
rect 45902 190609 45993 190727
rect 46111 190609 46202 190727
rect 45902 190567 46202 190609
rect 45902 190449 45993 190567
rect 46111 190449 46202 190567
rect 45902 172727 46202 190449
rect 45902 172609 45993 172727
rect 46111 172609 46202 172727
rect 45902 172567 46202 172609
rect 45902 172449 45993 172567
rect 46111 172449 46202 172567
rect 45902 154727 46202 172449
rect 45902 154609 45993 154727
rect 46111 154609 46202 154727
rect 45902 154567 46202 154609
rect 45902 154449 45993 154567
rect 46111 154449 46202 154567
rect 45902 136727 46202 154449
rect 45902 136609 45993 136727
rect 46111 136609 46202 136727
rect 45902 136567 46202 136609
rect 45902 136449 45993 136567
rect 46111 136449 46202 136567
rect 45902 118727 46202 136449
rect 45902 118609 45993 118727
rect 46111 118609 46202 118727
rect 45902 118567 46202 118609
rect 45902 118449 45993 118567
rect 46111 118449 46202 118567
rect 45902 100727 46202 118449
rect 45902 100609 45993 100727
rect 46111 100609 46202 100727
rect 45902 100567 46202 100609
rect 45902 100449 45993 100567
rect 46111 100449 46202 100567
rect 45902 82727 46202 100449
rect 45902 82609 45993 82727
rect 46111 82609 46202 82727
rect 45902 82567 46202 82609
rect 45902 82449 45993 82567
rect 46111 82449 46202 82567
rect 45902 64727 46202 82449
rect 45902 64609 45993 64727
rect 46111 64609 46202 64727
rect 45902 64567 46202 64609
rect 45902 64449 45993 64567
rect 46111 64449 46202 64567
rect 45902 46727 46202 64449
rect 45902 46609 45993 46727
rect 46111 46609 46202 46727
rect 45902 46567 46202 46609
rect 45902 46449 45993 46567
rect 46111 46449 46202 46567
rect 45902 28727 46202 46449
rect 45902 28609 45993 28727
rect 46111 28609 46202 28727
rect 45902 28567 46202 28609
rect 45902 28449 45993 28567
rect 46111 28449 46202 28567
rect 45902 10727 46202 28449
rect 45902 10609 45993 10727
rect 46111 10609 46202 10727
rect 45902 10567 46202 10609
rect 45902 10449 45993 10567
rect 46111 10449 46202 10567
rect 45902 -643 46202 10449
rect 45902 -761 45993 -643
rect 46111 -761 46202 -643
rect 45902 -803 46202 -761
rect 45902 -921 45993 -803
rect 46111 -921 46202 -803
rect 45902 -932 46202 -921
rect 47702 336527 48002 353551
rect 47702 336409 47793 336527
rect 47911 336409 48002 336527
rect 47702 336367 48002 336409
rect 47702 336249 47793 336367
rect 47911 336249 48002 336367
rect 47702 318527 48002 336249
rect 47702 318409 47793 318527
rect 47911 318409 48002 318527
rect 47702 318367 48002 318409
rect 47702 318249 47793 318367
rect 47911 318249 48002 318367
rect 47702 300527 48002 318249
rect 47702 300409 47793 300527
rect 47911 300409 48002 300527
rect 47702 300367 48002 300409
rect 47702 300249 47793 300367
rect 47911 300249 48002 300367
rect 47702 282527 48002 300249
rect 47702 282409 47793 282527
rect 47911 282409 48002 282527
rect 47702 282367 48002 282409
rect 47702 282249 47793 282367
rect 47911 282249 48002 282367
rect 47702 264527 48002 282249
rect 47702 264409 47793 264527
rect 47911 264409 48002 264527
rect 47702 264367 48002 264409
rect 47702 264249 47793 264367
rect 47911 264249 48002 264367
rect 47702 246527 48002 264249
rect 47702 246409 47793 246527
rect 47911 246409 48002 246527
rect 47702 246367 48002 246409
rect 47702 246249 47793 246367
rect 47911 246249 48002 246367
rect 47702 228527 48002 246249
rect 47702 228409 47793 228527
rect 47911 228409 48002 228527
rect 47702 228367 48002 228409
rect 47702 228249 47793 228367
rect 47911 228249 48002 228367
rect 47702 210527 48002 228249
rect 47702 210409 47793 210527
rect 47911 210409 48002 210527
rect 47702 210367 48002 210409
rect 47702 210249 47793 210367
rect 47911 210249 48002 210367
rect 47702 192527 48002 210249
rect 47702 192409 47793 192527
rect 47911 192409 48002 192527
rect 47702 192367 48002 192409
rect 47702 192249 47793 192367
rect 47911 192249 48002 192367
rect 47702 174527 48002 192249
rect 47702 174409 47793 174527
rect 47911 174409 48002 174527
rect 47702 174367 48002 174409
rect 47702 174249 47793 174367
rect 47911 174249 48002 174367
rect 47702 156527 48002 174249
rect 47702 156409 47793 156527
rect 47911 156409 48002 156527
rect 47702 156367 48002 156409
rect 47702 156249 47793 156367
rect 47911 156249 48002 156367
rect 47702 138527 48002 156249
rect 47702 138409 47793 138527
rect 47911 138409 48002 138527
rect 47702 138367 48002 138409
rect 47702 138249 47793 138367
rect 47911 138249 48002 138367
rect 47702 120527 48002 138249
rect 47702 120409 47793 120527
rect 47911 120409 48002 120527
rect 47702 120367 48002 120409
rect 47702 120249 47793 120367
rect 47911 120249 48002 120367
rect 47702 102527 48002 120249
rect 47702 102409 47793 102527
rect 47911 102409 48002 102527
rect 47702 102367 48002 102409
rect 47702 102249 47793 102367
rect 47911 102249 48002 102367
rect 47702 84527 48002 102249
rect 47702 84409 47793 84527
rect 47911 84409 48002 84527
rect 47702 84367 48002 84409
rect 47702 84249 47793 84367
rect 47911 84249 48002 84367
rect 47702 66527 48002 84249
rect 47702 66409 47793 66527
rect 47911 66409 48002 66527
rect 47702 66367 48002 66409
rect 47702 66249 47793 66367
rect 47911 66249 48002 66367
rect 47702 48527 48002 66249
rect 47702 48409 47793 48527
rect 47911 48409 48002 48527
rect 47702 48367 48002 48409
rect 47702 48249 47793 48367
rect 47911 48249 48002 48367
rect 47702 30527 48002 48249
rect 47702 30409 47793 30527
rect 47911 30409 48002 30527
rect 47702 30367 48002 30409
rect 47702 30249 47793 30367
rect 47911 30249 48002 30367
rect 47702 12527 48002 30249
rect 47702 12409 47793 12527
rect 47911 12409 48002 12527
rect 47702 12367 48002 12409
rect 47702 12249 47793 12367
rect 47911 12249 48002 12367
rect 47702 -1583 48002 12249
rect 47702 -1701 47793 -1583
rect 47911 -1701 48002 -1583
rect 47702 -1743 48002 -1701
rect 47702 -1861 47793 -1743
rect 47911 -1861 48002 -1743
rect 47702 -1872 48002 -1861
rect 49502 338327 49802 354491
rect 49502 338209 49593 338327
rect 49711 338209 49802 338327
rect 49502 338167 49802 338209
rect 49502 338049 49593 338167
rect 49711 338049 49802 338167
rect 49502 320327 49802 338049
rect 49502 320209 49593 320327
rect 49711 320209 49802 320327
rect 49502 320167 49802 320209
rect 49502 320049 49593 320167
rect 49711 320049 49802 320167
rect 49502 302327 49802 320049
rect 49502 302209 49593 302327
rect 49711 302209 49802 302327
rect 49502 302167 49802 302209
rect 49502 302049 49593 302167
rect 49711 302049 49802 302167
rect 49502 284327 49802 302049
rect 49502 284209 49593 284327
rect 49711 284209 49802 284327
rect 49502 284167 49802 284209
rect 49502 284049 49593 284167
rect 49711 284049 49802 284167
rect 49502 266327 49802 284049
rect 49502 266209 49593 266327
rect 49711 266209 49802 266327
rect 49502 266167 49802 266209
rect 49502 266049 49593 266167
rect 49711 266049 49802 266167
rect 49502 248327 49802 266049
rect 49502 248209 49593 248327
rect 49711 248209 49802 248327
rect 49502 248167 49802 248209
rect 49502 248049 49593 248167
rect 49711 248049 49802 248167
rect 49502 230327 49802 248049
rect 49502 230209 49593 230327
rect 49711 230209 49802 230327
rect 49502 230167 49802 230209
rect 49502 230049 49593 230167
rect 49711 230049 49802 230167
rect 49502 212327 49802 230049
rect 49502 212209 49593 212327
rect 49711 212209 49802 212327
rect 49502 212167 49802 212209
rect 49502 212049 49593 212167
rect 49711 212049 49802 212167
rect 49502 194327 49802 212049
rect 49502 194209 49593 194327
rect 49711 194209 49802 194327
rect 49502 194167 49802 194209
rect 49502 194049 49593 194167
rect 49711 194049 49802 194167
rect 49502 176327 49802 194049
rect 49502 176209 49593 176327
rect 49711 176209 49802 176327
rect 49502 176167 49802 176209
rect 49502 176049 49593 176167
rect 49711 176049 49802 176167
rect 49502 158327 49802 176049
rect 49502 158209 49593 158327
rect 49711 158209 49802 158327
rect 49502 158167 49802 158209
rect 49502 158049 49593 158167
rect 49711 158049 49802 158167
rect 49502 140327 49802 158049
rect 49502 140209 49593 140327
rect 49711 140209 49802 140327
rect 49502 140167 49802 140209
rect 49502 140049 49593 140167
rect 49711 140049 49802 140167
rect 49502 122327 49802 140049
rect 49502 122209 49593 122327
rect 49711 122209 49802 122327
rect 49502 122167 49802 122209
rect 49502 122049 49593 122167
rect 49711 122049 49802 122167
rect 49502 104327 49802 122049
rect 49502 104209 49593 104327
rect 49711 104209 49802 104327
rect 49502 104167 49802 104209
rect 49502 104049 49593 104167
rect 49711 104049 49802 104167
rect 49502 86327 49802 104049
rect 49502 86209 49593 86327
rect 49711 86209 49802 86327
rect 49502 86167 49802 86209
rect 49502 86049 49593 86167
rect 49711 86049 49802 86167
rect 49502 68327 49802 86049
rect 49502 68209 49593 68327
rect 49711 68209 49802 68327
rect 49502 68167 49802 68209
rect 49502 68049 49593 68167
rect 49711 68049 49802 68167
rect 49502 50327 49802 68049
rect 49502 50209 49593 50327
rect 49711 50209 49802 50327
rect 49502 50167 49802 50209
rect 49502 50049 49593 50167
rect 49711 50049 49802 50167
rect 49502 32327 49802 50049
rect 49502 32209 49593 32327
rect 49711 32209 49802 32327
rect 49502 32167 49802 32209
rect 49502 32049 49593 32167
rect 49711 32049 49802 32167
rect 49502 14327 49802 32049
rect 49502 14209 49593 14327
rect 49711 14209 49802 14327
rect 49502 14167 49802 14209
rect 49502 14049 49593 14167
rect 49711 14049 49802 14167
rect 49502 -2523 49802 14049
rect 49502 -2641 49593 -2523
rect 49711 -2641 49802 -2523
rect 49502 -2683 49802 -2641
rect 49502 -2801 49593 -2683
rect 49711 -2801 49802 -2683
rect 49502 -2812 49802 -2801
rect 51302 340127 51602 355431
rect 60302 355239 60602 355720
rect 60302 355121 60393 355239
rect 60511 355121 60602 355239
rect 60302 355079 60602 355121
rect 60302 354961 60393 355079
rect 60511 354961 60602 355079
rect 58502 354299 58802 354780
rect 58502 354181 58593 354299
rect 58711 354181 58802 354299
rect 58502 354139 58802 354181
rect 58502 354021 58593 354139
rect 58711 354021 58802 354139
rect 56702 353359 57002 353840
rect 56702 353241 56793 353359
rect 56911 353241 57002 353359
rect 56702 353199 57002 353241
rect 56702 353081 56793 353199
rect 56911 353081 57002 353199
rect 51302 340009 51393 340127
rect 51511 340009 51602 340127
rect 51302 339967 51602 340009
rect 51302 339849 51393 339967
rect 51511 339849 51602 339967
rect 51302 322127 51602 339849
rect 51302 322009 51393 322127
rect 51511 322009 51602 322127
rect 51302 321967 51602 322009
rect 51302 321849 51393 321967
rect 51511 321849 51602 321967
rect 51302 304127 51602 321849
rect 51302 304009 51393 304127
rect 51511 304009 51602 304127
rect 51302 303967 51602 304009
rect 51302 303849 51393 303967
rect 51511 303849 51602 303967
rect 51302 286127 51602 303849
rect 51302 286009 51393 286127
rect 51511 286009 51602 286127
rect 51302 285967 51602 286009
rect 51302 285849 51393 285967
rect 51511 285849 51602 285967
rect 51302 268127 51602 285849
rect 51302 268009 51393 268127
rect 51511 268009 51602 268127
rect 51302 267967 51602 268009
rect 51302 267849 51393 267967
rect 51511 267849 51602 267967
rect 51302 250127 51602 267849
rect 51302 250009 51393 250127
rect 51511 250009 51602 250127
rect 51302 249967 51602 250009
rect 51302 249849 51393 249967
rect 51511 249849 51602 249967
rect 51302 232127 51602 249849
rect 51302 232009 51393 232127
rect 51511 232009 51602 232127
rect 51302 231967 51602 232009
rect 51302 231849 51393 231967
rect 51511 231849 51602 231967
rect 51302 214127 51602 231849
rect 51302 214009 51393 214127
rect 51511 214009 51602 214127
rect 51302 213967 51602 214009
rect 51302 213849 51393 213967
rect 51511 213849 51602 213967
rect 51302 196127 51602 213849
rect 51302 196009 51393 196127
rect 51511 196009 51602 196127
rect 51302 195967 51602 196009
rect 51302 195849 51393 195967
rect 51511 195849 51602 195967
rect 51302 178127 51602 195849
rect 51302 178009 51393 178127
rect 51511 178009 51602 178127
rect 51302 177967 51602 178009
rect 51302 177849 51393 177967
rect 51511 177849 51602 177967
rect 51302 160127 51602 177849
rect 51302 160009 51393 160127
rect 51511 160009 51602 160127
rect 51302 159967 51602 160009
rect 51302 159849 51393 159967
rect 51511 159849 51602 159967
rect 51302 142127 51602 159849
rect 51302 142009 51393 142127
rect 51511 142009 51602 142127
rect 51302 141967 51602 142009
rect 51302 141849 51393 141967
rect 51511 141849 51602 141967
rect 51302 124127 51602 141849
rect 51302 124009 51393 124127
rect 51511 124009 51602 124127
rect 51302 123967 51602 124009
rect 51302 123849 51393 123967
rect 51511 123849 51602 123967
rect 51302 106127 51602 123849
rect 51302 106009 51393 106127
rect 51511 106009 51602 106127
rect 51302 105967 51602 106009
rect 51302 105849 51393 105967
rect 51511 105849 51602 105967
rect 51302 88127 51602 105849
rect 51302 88009 51393 88127
rect 51511 88009 51602 88127
rect 51302 87967 51602 88009
rect 51302 87849 51393 87967
rect 51511 87849 51602 87967
rect 51302 70127 51602 87849
rect 51302 70009 51393 70127
rect 51511 70009 51602 70127
rect 51302 69967 51602 70009
rect 51302 69849 51393 69967
rect 51511 69849 51602 69967
rect 51302 52127 51602 69849
rect 51302 52009 51393 52127
rect 51511 52009 51602 52127
rect 51302 51967 51602 52009
rect 51302 51849 51393 51967
rect 51511 51849 51602 51967
rect 51302 34127 51602 51849
rect 51302 34009 51393 34127
rect 51511 34009 51602 34127
rect 51302 33967 51602 34009
rect 51302 33849 51393 33967
rect 51511 33849 51602 33967
rect 51302 16127 51602 33849
rect 51302 16009 51393 16127
rect 51511 16009 51602 16127
rect 51302 15967 51602 16009
rect 51302 15849 51393 15967
rect 51511 15849 51602 15967
rect 42302 -3111 42393 -2993
rect 42511 -3111 42602 -2993
rect 42302 -3153 42602 -3111
rect 42302 -3271 42393 -3153
rect 42511 -3271 42602 -3153
rect 42302 -3752 42602 -3271
rect 51302 -3463 51602 15849
rect 54902 352419 55202 352900
rect 54902 352301 54993 352419
rect 55111 352301 55202 352419
rect 54902 352259 55202 352301
rect 54902 352141 54993 352259
rect 55111 352141 55202 352259
rect 54902 343727 55202 352141
rect 54902 343609 54993 343727
rect 55111 343609 55202 343727
rect 54902 343567 55202 343609
rect 54902 343449 54993 343567
rect 55111 343449 55202 343567
rect 54902 325727 55202 343449
rect 54902 325609 54993 325727
rect 55111 325609 55202 325727
rect 54902 325567 55202 325609
rect 54902 325449 54993 325567
rect 55111 325449 55202 325567
rect 54902 307727 55202 325449
rect 54902 307609 54993 307727
rect 55111 307609 55202 307727
rect 54902 307567 55202 307609
rect 54902 307449 54993 307567
rect 55111 307449 55202 307567
rect 54902 289727 55202 307449
rect 54902 289609 54993 289727
rect 55111 289609 55202 289727
rect 54902 289567 55202 289609
rect 54902 289449 54993 289567
rect 55111 289449 55202 289567
rect 54902 271727 55202 289449
rect 54902 271609 54993 271727
rect 55111 271609 55202 271727
rect 54902 271567 55202 271609
rect 54902 271449 54993 271567
rect 55111 271449 55202 271567
rect 54902 253727 55202 271449
rect 54902 253609 54993 253727
rect 55111 253609 55202 253727
rect 54902 253567 55202 253609
rect 54902 253449 54993 253567
rect 55111 253449 55202 253567
rect 54902 235727 55202 253449
rect 54902 235609 54993 235727
rect 55111 235609 55202 235727
rect 54902 235567 55202 235609
rect 54902 235449 54993 235567
rect 55111 235449 55202 235567
rect 54902 217727 55202 235449
rect 54902 217609 54993 217727
rect 55111 217609 55202 217727
rect 54902 217567 55202 217609
rect 54902 217449 54993 217567
rect 55111 217449 55202 217567
rect 54902 199727 55202 217449
rect 54902 199609 54993 199727
rect 55111 199609 55202 199727
rect 54902 199567 55202 199609
rect 54902 199449 54993 199567
rect 55111 199449 55202 199567
rect 54902 181727 55202 199449
rect 54902 181609 54993 181727
rect 55111 181609 55202 181727
rect 54902 181567 55202 181609
rect 54902 181449 54993 181567
rect 55111 181449 55202 181567
rect 54902 163727 55202 181449
rect 54902 163609 54993 163727
rect 55111 163609 55202 163727
rect 54902 163567 55202 163609
rect 54902 163449 54993 163567
rect 55111 163449 55202 163567
rect 54902 145727 55202 163449
rect 54902 145609 54993 145727
rect 55111 145609 55202 145727
rect 54902 145567 55202 145609
rect 54902 145449 54993 145567
rect 55111 145449 55202 145567
rect 54902 127727 55202 145449
rect 54902 127609 54993 127727
rect 55111 127609 55202 127727
rect 54902 127567 55202 127609
rect 54902 127449 54993 127567
rect 55111 127449 55202 127567
rect 54902 109727 55202 127449
rect 54902 109609 54993 109727
rect 55111 109609 55202 109727
rect 54902 109567 55202 109609
rect 54902 109449 54993 109567
rect 55111 109449 55202 109567
rect 54902 91727 55202 109449
rect 54902 91609 54993 91727
rect 55111 91609 55202 91727
rect 54902 91567 55202 91609
rect 54902 91449 54993 91567
rect 55111 91449 55202 91567
rect 54902 73727 55202 91449
rect 54902 73609 54993 73727
rect 55111 73609 55202 73727
rect 54902 73567 55202 73609
rect 54902 73449 54993 73567
rect 55111 73449 55202 73567
rect 54902 55727 55202 73449
rect 54902 55609 54993 55727
rect 55111 55609 55202 55727
rect 54902 55567 55202 55609
rect 54902 55449 54993 55567
rect 55111 55449 55202 55567
rect 54902 37727 55202 55449
rect 54902 37609 54993 37727
rect 55111 37609 55202 37727
rect 54902 37567 55202 37609
rect 54902 37449 54993 37567
rect 55111 37449 55202 37567
rect 54902 19727 55202 37449
rect 54902 19609 54993 19727
rect 55111 19609 55202 19727
rect 54902 19567 55202 19609
rect 54902 19449 54993 19567
rect 55111 19449 55202 19567
rect 54902 1727 55202 19449
rect 54902 1609 54993 1727
rect 55111 1609 55202 1727
rect 54902 1567 55202 1609
rect 54902 1449 54993 1567
rect 55111 1449 55202 1567
rect 54902 -173 55202 1449
rect 54902 -291 54993 -173
rect 55111 -291 55202 -173
rect 54902 -333 55202 -291
rect 54902 -451 54993 -333
rect 55111 -451 55202 -333
rect 54902 -932 55202 -451
rect 56702 345527 57002 353081
rect 56702 345409 56793 345527
rect 56911 345409 57002 345527
rect 56702 345367 57002 345409
rect 56702 345249 56793 345367
rect 56911 345249 57002 345367
rect 56702 327527 57002 345249
rect 56702 327409 56793 327527
rect 56911 327409 57002 327527
rect 56702 327367 57002 327409
rect 56702 327249 56793 327367
rect 56911 327249 57002 327367
rect 56702 309527 57002 327249
rect 56702 309409 56793 309527
rect 56911 309409 57002 309527
rect 56702 309367 57002 309409
rect 56702 309249 56793 309367
rect 56911 309249 57002 309367
rect 56702 291527 57002 309249
rect 56702 291409 56793 291527
rect 56911 291409 57002 291527
rect 56702 291367 57002 291409
rect 56702 291249 56793 291367
rect 56911 291249 57002 291367
rect 56702 273527 57002 291249
rect 56702 273409 56793 273527
rect 56911 273409 57002 273527
rect 56702 273367 57002 273409
rect 56702 273249 56793 273367
rect 56911 273249 57002 273367
rect 56702 255527 57002 273249
rect 56702 255409 56793 255527
rect 56911 255409 57002 255527
rect 56702 255367 57002 255409
rect 56702 255249 56793 255367
rect 56911 255249 57002 255367
rect 56702 237527 57002 255249
rect 56702 237409 56793 237527
rect 56911 237409 57002 237527
rect 56702 237367 57002 237409
rect 56702 237249 56793 237367
rect 56911 237249 57002 237367
rect 56702 219527 57002 237249
rect 56702 219409 56793 219527
rect 56911 219409 57002 219527
rect 56702 219367 57002 219409
rect 56702 219249 56793 219367
rect 56911 219249 57002 219367
rect 56702 201527 57002 219249
rect 56702 201409 56793 201527
rect 56911 201409 57002 201527
rect 56702 201367 57002 201409
rect 56702 201249 56793 201367
rect 56911 201249 57002 201367
rect 56702 183527 57002 201249
rect 56702 183409 56793 183527
rect 56911 183409 57002 183527
rect 56702 183367 57002 183409
rect 56702 183249 56793 183367
rect 56911 183249 57002 183367
rect 56702 165527 57002 183249
rect 56702 165409 56793 165527
rect 56911 165409 57002 165527
rect 56702 165367 57002 165409
rect 56702 165249 56793 165367
rect 56911 165249 57002 165367
rect 56702 147527 57002 165249
rect 56702 147409 56793 147527
rect 56911 147409 57002 147527
rect 56702 147367 57002 147409
rect 56702 147249 56793 147367
rect 56911 147249 57002 147367
rect 56702 129527 57002 147249
rect 56702 129409 56793 129527
rect 56911 129409 57002 129527
rect 56702 129367 57002 129409
rect 56702 129249 56793 129367
rect 56911 129249 57002 129367
rect 56702 111527 57002 129249
rect 56702 111409 56793 111527
rect 56911 111409 57002 111527
rect 56702 111367 57002 111409
rect 56702 111249 56793 111367
rect 56911 111249 57002 111367
rect 56702 93527 57002 111249
rect 56702 93409 56793 93527
rect 56911 93409 57002 93527
rect 56702 93367 57002 93409
rect 56702 93249 56793 93367
rect 56911 93249 57002 93367
rect 56702 75527 57002 93249
rect 56702 75409 56793 75527
rect 56911 75409 57002 75527
rect 56702 75367 57002 75409
rect 56702 75249 56793 75367
rect 56911 75249 57002 75367
rect 56702 57527 57002 75249
rect 56702 57409 56793 57527
rect 56911 57409 57002 57527
rect 56702 57367 57002 57409
rect 56702 57249 56793 57367
rect 56911 57249 57002 57367
rect 56702 39527 57002 57249
rect 56702 39409 56793 39527
rect 56911 39409 57002 39527
rect 56702 39367 57002 39409
rect 56702 39249 56793 39367
rect 56911 39249 57002 39367
rect 56702 21527 57002 39249
rect 56702 21409 56793 21527
rect 56911 21409 57002 21527
rect 56702 21367 57002 21409
rect 56702 21249 56793 21367
rect 56911 21249 57002 21367
rect 56702 3527 57002 21249
rect 56702 3409 56793 3527
rect 56911 3409 57002 3527
rect 56702 3367 57002 3409
rect 56702 3249 56793 3367
rect 56911 3249 57002 3367
rect 56702 -1113 57002 3249
rect 56702 -1231 56793 -1113
rect 56911 -1231 57002 -1113
rect 56702 -1273 57002 -1231
rect 56702 -1391 56793 -1273
rect 56911 -1391 57002 -1273
rect 56702 -1872 57002 -1391
rect 58502 347327 58802 354021
rect 58502 347209 58593 347327
rect 58711 347209 58802 347327
rect 58502 347167 58802 347209
rect 58502 347049 58593 347167
rect 58711 347049 58802 347167
rect 58502 329327 58802 347049
rect 58502 329209 58593 329327
rect 58711 329209 58802 329327
rect 58502 329167 58802 329209
rect 58502 329049 58593 329167
rect 58711 329049 58802 329167
rect 58502 311327 58802 329049
rect 58502 311209 58593 311327
rect 58711 311209 58802 311327
rect 58502 311167 58802 311209
rect 58502 311049 58593 311167
rect 58711 311049 58802 311167
rect 58502 293327 58802 311049
rect 58502 293209 58593 293327
rect 58711 293209 58802 293327
rect 58502 293167 58802 293209
rect 58502 293049 58593 293167
rect 58711 293049 58802 293167
rect 58502 275327 58802 293049
rect 58502 275209 58593 275327
rect 58711 275209 58802 275327
rect 58502 275167 58802 275209
rect 58502 275049 58593 275167
rect 58711 275049 58802 275167
rect 58502 257327 58802 275049
rect 58502 257209 58593 257327
rect 58711 257209 58802 257327
rect 58502 257167 58802 257209
rect 58502 257049 58593 257167
rect 58711 257049 58802 257167
rect 58502 239327 58802 257049
rect 58502 239209 58593 239327
rect 58711 239209 58802 239327
rect 58502 239167 58802 239209
rect 58502 239049 58593 239167
rect 58711 239049 58802 239167
rect 58502 221327 58802 239049
rect 58502 221209 58593 221327
rect 58711 221209 58802 221327
rect 58502 221167 58802 221209
rect 58502 221049 58593 221167
rect 58711 221049 58802 221167
rect 58502 203327 58802 221049
rect 58502 203209 58593 203327
rect 58711 203209 58802 203327
rect 58502 203167 58802 203209
rect 58502 203049 58593 203167
rect 58711 203049 58802 203167
rect 58502 185327 58802 203049
rect 58502 185209 58593 185327
rect 58711 185209 58802 185327
rect 58502 185167 58802 185209
rect 58502 185049 58593 185167
rect 58711 185049 58802 185167
rect 58502 167327 58802 185049
rect 58502 167209 58593 167327
rect 58711 167209 58802 167327
rect 58502 167167 58802 167209
rect 58502 167049 58593 167167
rect 58711 167049 58802 167167
rect 58502 149327 58802 167049
rect 58502 149209 58593 149327
rect 58711 149209 58802 149327
rect 58502 149167 58802 149209
rect 58502 149049 58593 149167
rect 58711 149049 58802 149167
rect 58502 131327 58802 149049
rect 58502 131209 58593 131327
rect 58711 131209 58802 131327
rect 58502 131167 58802 131209
rect 58502 131049 58593 131167
rect 58711 131049 58802 131167
rect 58502 113327 58802 131049
rect 58502 113209 58593 113327
rect 58711 113209 58802 113327
rect 58502 113167 58802 113209
rect 58502 113049 58593 113167
rect 58711 113049 58802 113167
rect 58502 95327 58802 113049
rect 58502 95209 58593 95327
rect 58711 95209 58802 95327
rect 58502 95167 58802 95209
rect 58502 95049 58593 95167
rect 58711 95049 58802 95167
rect 58502 77327 58802 95049
rect 58502 77209 58593 77327
rect 58711 77209 58802 77327
rect 58502 77167 58802 77209
rect 58502 77049 58593 77167
rect 58711 77049 58802 77167
rect 58502 59327 58802 77049
rect 58502 59209 58593 59327
rect 58711 59209 58802 59327
rect 58502 59167 58802 59209
rect 58502 59049 58593 59167
rect 58711 59049 58802 59167
rect 58502 41327 58802 59049
rect 58502 41209 58593 41327
rect 58711 41209 58802 41327
rect 58502 41167 58802 41209
rect 58502 41049 58593 41167
rect 58711 41049 58802 41167
rect 58502 23327 58802 41049
rect 58502 23209 58593 23327
rect 58711 23209 58802 23327
rect 58502 23167 58802 23209
rect 58502 23049 58593 23167
rect 58711 23049 58802 23167
rect 58502 5327 58802 23049
rect 58502 5209 58593 5327
rect 58711 5209 58802 5327
rect 58502 5167 58802 5209
rect 58502 5049 58593 5167
rect 58711 5049 58802 5167
rect 58502 -2053 58802 5049
rect 58502 -2171 58593 -2053
rect 58711 -2171 58802 -2053
rect 58502 -2213 58802 -2171
rect 58502 -2331 58593 -2213
rect 58711 -2331 58802 -2213
rect 58502 -2812 58802 -2331
rect 60302 349127 60602 354961
rect 69302 355709 69602 355720
rect 69302 355591 69393 355709
rect 69511 355591 69602 355709
rect 69302 355549 69602 355591
rect 69302 355431 69393 355549
rect 69511 355431 69602 355549
rect 67502 354769 67802 354780
rect 67502 354651 67593 354769
rect 67711 354651 67802 354769
rect 67502 354609 67802 354651
rect 67502 354491 67593 354609
rect 67711 354491 67802 354609
rect 65702 353829 66002 353840
rect 65702 353711 65793 353829
rect 65911 353711 66002 353829
rect 65702 353669 66002 353711
rect 65702 353551 65793 353669
rect 65911 353551 66002 353669
rect 60302 349009 60393 349127
rect 60511 349009 60602 349127
rect 60302 348967 60602 349009
rect 60302 348849 60393 348967
rect 60511 348849 60602 348967
rect 60302 331127 60602 348849
rect 60302 331009 60393 331127
rect 60511 331009 60602 331127
rect 60302 330967 60602 331009
rect 60302 330849 60393 330967
rect 60511 330849 60602 330967
rect 60302 313127 60602 330849
rect 60302 313009 60393 313127
rect 60511 313009 60602 313127
rect 60302 312967 60602 313009
rect 60302 312849 60393 312967
rect 60511 312849 60602 312967
rect 60302 295127 60602 312849
rect 60302 295009 60393 295127
rect 60511 295009 60602 295127
rect 60302 294967 60602 295009
rect 60302 294849 60393 294967
rect 60511 294849 60602 294967
rect 60302 277127 60602 294849
rect 60302 277009 60393 277127
rect 60511 277009 60602 277127
rect 60302 276967 60602 277009
rect 60302 276849 60393 276967
rect 60511 276849 60602 276967
rect 60302 259127 60602 276849
rect 60302 259009 60393 259127
rect 60511 259009 60602 259127
rect 60302 258967 60602 259009
rect 60302 258849 60393 258967
rect 60511 258849 60602 258967
rect 60302 241127 60602 258849
rect 60302 241009 60393 241127
rect 60511 241009 60602 241127
rect 60302 240967 60602 241009
rect 60302 240849 60393 240967
rect 60511 240849 60602 240967
rect 60302 223127 60602 240849
rect 60302 223009 60393 223127
rect 60511 223009 60602 223127
rect 60302 222967 60602 223009
rect 60302 222849 60393 222967
rect 60511 222849 60602 222967
rect 60302 205127 60602 222849
rect 60302 205009 60393 205127
rect 60511 205009 60602 205127
rect 60302 204967 60602 205009
rect 60302 204849 60393 204967
rect 60511 204849 60602 204967
rect 60302 187127 60602 204849
rect 60302 187009 60393 187127
rect 60511 187009 60602 187127
rect 60302 186967 60602 187009
rect 60302 186849 60393 186967
rect 60511 186849 60602 186967
rect 60302 169127 60602 186849
rect 60302 169009 60393 169127
rect 60511 169009 60602 169127
rect 60302 168967 60602 169009
rect 60302 168849 60393 168967
rect 60511 168849 60602 168967
rect 60302 151127 60602 168849
rect 60302 151009 60393 151127
rect 60511 151009 60602 151127
rect 60302 150967 60602 151009
rect 60302 150849 60393 150967
rect 60511 150849 60602 150967
rect 60302 133127 60602 150849
rect 60302 133009 60393 133127
rect 60511 133009 60602 133127
rect 60302 132967 60602 133009
rect 60302 132849 60393 132967
rect 60511 132849 60602 132967
rect 60302 115127 60602 132849
rect 60302 115009 60393 115127
rect 60511 115009 60602 115127
rect 60302 114967 60602 115009
rect 60302 114849 60393 114967
rect 60511 114849 60602 114967
rect 60302 97127 60602 114849
rect 60302 97009 60393 97127
rect 60511 97009 60602 97127
rect 60302 96967 60602 97009
rect 60302 96849 60393 96967
rect 60511 96849 60602 96967
rect 60302 79127 60602 96849
rect 60302 79009 60393 79127
rect 60511 79009 60602 79127
rect 60302 78967 60602 79009
rect 60302 78849 60393 78967
rect 60511 78849 60602 78967
rect 60302 61127 60602 78849
rect 60302 61009 60393 61127
rect 60511 61009 60602 61127
rect 60302 60967 60602 61009
rect 60302 60849 60393 60967
rect 60511 60849 60602 60967
rect 60302 43127 60602 60849
rect 60302 43009 60393 43127
rect 60511 43009 60602 43127
rect 60302 42967 60602 43009
rect 60302 42849 60393 42967
rect 60511 42849 60602 42967
rect 60302 25127 60602 42849
rect 60302 25009 60393 25127
rect 60511 25009 60602 25127
rect 60302 24967 60602 25009
rect 60302 24849 60393 24967
rect 60511 24849 60602 24967
rect 60302 7127 60602 24849
rect 60302 7009 60393 7127
rect 60511 7009 60602 7127
rect 60302 6967 60602 7009
rect 60302 6849 60393 6967
rect 60511 6849 60602 6967
rect 51302 -3581 51393 -3463
rect 51511 -3581 51602 -3463
rect 51302 -3623 51602 -3581
rect 51302 -3741 51393 -3623
rect 51511 -3741 51602 -3623
rect 51302 -3752 51602 -3741
rect 60302 -2993 60602 6849
rect 63902 352889 64202 352900
rect 63902 352771 63993 352889
rect 64111 352771 64202 352889
rect 63902 352729 64202 352771
rect 63902 352611 63993 352729
rect 64111 352611 64202 352729
rect 63902 334727 64202 352611
rect 63902 334609 63993 334727
rect 64111 334609 64202 334727
rect 63902 334567 64202 334609
rect 63902 334449 63993 334567
rect 64111 334449 64202 334567
rect 63902 316727 64202 334449
rect 63902 316609 63993 316727
rect 64111 316609 64202 316727
rect 63902 316567 64202 316609
rect 63902 316449 63993 316567
rect 64111 316449 64202 316567
rect 63902 298727 64202 316449
rect 63902 298609 63993 298727
rect 64111 298609 64202 298727
rect 63902 298567 64202 298609
rect 63902 298449 63993 298567
rect 64111 298449 64202 298567
rect 63902 280727 64202 298449
rect 63902 280609 63993 280727
rect 64111 280609 64202 280727
rect 63902 280567 64202 280609
rect 63902 280449 63993 280567
rect 64111 280449 64202 280567
rect 63902 262727 64202 280449
rect 63902 262609 63993 262727
rect 64111 262609 64202 262727
rect 63902 262567 64202 262609
rect 63902 262449 63993 262567
rect 64111 262449 64202 262567
rect 63902 244727 64202 262449
rect 63902 244609 63993 244727
rect 64111 244609 64202 244727
rect 63902 244567 64202 244609
rect 63902 244449 63993 244567
rect 64111 244449 64202 244567
rect 63902 226727 64202 244449
rect 63902 226609 63993 226727
rect 64111 226609 64202 226727
rect 63902 226567 64202 226609
rect 63902 226449 63993 226567
rect 64111 226449 64202 226567
rect 63902 208727 64202 226449
rect 63902 208609 63993 208727
rect 64111 208609 64202 208727
rect 63902 208567 64202 208609
rect 63902 208449 63993 208567
rect 64111 208449 64202 208567
rect 63902 190727 64202 208449
rect 63902 190609 63993 190727
rect 64111 190609 64202 190727
rect 63902 190567 64202 190609
rect 63902 190449 63993 190567
rect 64111 190449 64202 190567
rect 63902 172727 64202 190449
rect 63902 172609 63993 172727
rect 64111 172609 64202 172727
rect 63902 172567 64202 172609
rect 63902 172449 63993 172567
rect 64111 172449 64202 172567
rect 63902 154727 64202 172449
rect 63902 154609 63993 154727
rect 64111 154609 64202 154727
rect 63902 154567 64202 154609
rect 63902 154449 63993 154567
rect 64111 154449 64202 154567
rect 63902 136727 64202 154449
rect 63902 136609 63993 136727
rect 64111 136609 64202 136727
rect 63902 136567 64202 136609
rect 63902 136449 63993 136567
rect 64111 136449 64202 136567
rect 63902 118727 64202 136449
rect 63902 118609 63993 118727
rect 64111 118609 64202 118727
rect 63902 118567 64202 118609
rect 63902 118449 63993 118567
rect 64111 118449 64202 118567
rect 63902 100727 64202 118449
rect 63902 100609 63993 100727
rect 64111 100609 64202 100727
rect 63902 100567 64202 100609
rect 63902 100449 63993 100567
rect 64111 100449 64202 100567
rect 63902 82727 64202 100449
rect 63902 82609 63993 82727
rect 64111 82609 64202 82727
rect 63902 82567 64202 82609
rect 63902 82449 63993 82567
rect 64111 82449 64202 82567
rect 63902 64727 64202 82449
rect 63902 64609 63993 64727
rect 64111 64609 64202 64727
rect 63902 64567 64202 64609
rect 63902 64449 63993 64567
rect 64111 64449 64202 64567
rect 63902 46727 64202 64449
rect 63902 46609 63993 46727
rect 64111 46609 64202 46727
rect 63902 46567 64202 46609
rect 63902 46449 63993 46567
rect 64111 46449 64202 46567
rect 63902 28727 64202 46449
rect 63902 28609 63993 28727
rect 64111 28609 64202 28727
rect 63902 28567 64202 28609
rect 63902 28449 63993 28567
rect 64111 28449 64202 28567
rect 63902 10727 64202 28449
rect 63902 10609 63993 10727
rect 64111 10609 64202 10727
rect 63902 10567 64202 10609
rect 63902 10449 63993 10567
rect 64111 10449 64202 10567
rect 63902 -643 64202 10449
rect 63902 -761 63993 -643
rect 64111 -761 64202 -643
rect 63902 -803 64202 -761
rect 63902 -921 63993 -803
rect 64111 -921 64202 -803
rect 63902 -932 64202 -921
rect 65702 336527 66002 353551
rect 65702 336409 65793 336527
rect 65911 336409 66002 336527
rect 65702 336367 66002 336409
rect 65702 336249 65793 336367
rect 65911 336249 66002 336367
rect 65702 318527 66002 336249
rect 65702 318409 65793 318527
rect 65911 318409 66002 318527
rect 65702 318367 66002 318409
rect 65702 318249 65793 318367
rect 65911 318249 66002 318367
rect 65702 300527 66002 318249
rect 65702 300409 65793 300527
rect 65911 300409 66002 300527
rect 65702 300367 66002 300409
rect 65702 300249 65793 300367
rect 65911 300249 66002 300367
rect 65702 282527 66002 300249
rect 65702 282409 65793 282527
rect 65911 282409 66002 282527
rect 65702 282367 66002 282409
rect 65702 282249 65793 282367
rect 65911 282249 66002 282367
rect 65702 264527 66002 282249
rect 65702 264409 65793 264527
rect 65911 264409 66002 264527
rect 65702 264367 66002 264409
rect 65702 264249 65793 264367
rect 65911 264249 66002 264367
rect 65702 246527 66002 264249
rect 65702 246409 65793 246527
rect 65911 246409 66002 246527
rect 65702 246367 66002 246409
rect 65702 246249 65793 246367
rect 65911 246249 66002 246367
rect 65702 228527 66002 246249
rect 65702 228409 65793 228527
rect 65911 228409 66002 228527
rect 65702 228367 66002 228409
rect 65702 228249 65793 228367
rect 65911 228249 66002 228367
rect 65702 210527 66002 228249
rect 65702 210409 65793 210527
rect 65911 210409 66002 210527
rect 65702 210367 66002 210409
rect 65702 210249 65793 210367
rect 65911 210249 66002 210367
rect 65702 192527 66002 210249
rect 65702 192409 65793 192527
rect 65911 192409 66002 192527
rect 65702 192367 66002 192409
rect 65702 192249 65793 192367
rect 65911 192249 66002 192367
rect 65702 174527 66002 192249
rect 65702 174409 65793 174527
rect 65911 174409 66002 174527
rect 65702 174367 66002 174409
rect 65702 174249 65793 174367
rect 65911 174249 66002 174367
rect 65702 156527 66002 174249
rect 65702 156409 65793 156527
rect 65911 156409 66002 156527
rect 65702 156367 66002 156409
rect 65702 156249 65793 156367
rect 65911 156249 66002 156367
rect 65702 138527 66002 156249
rect 65702 138409 65793 138527
rect 65911 138409 66002 138527
rect 65702 138367 66002 138409
rect 65702 138249 65793 138367
rect 65911 138249 66002 138367
rect 65702 120527 66002 138249
rect 65702 120409 65793 120527
rect 65911 120409 66002 120527
rect 65702 120367 66002 120409
rect 65702 120249 65793 120367
rect 65911 120249 66002 120367
rect 65702 102527 66002 120249
rect 65702 102409 65793 102527
rect 65911 102409 66002 102527
rect 65702 102367 66002 102409
rect 65702 102249 65793 102367
rect 65911 102249 66002 102367
rect 65702 84527 66002 102249
rect 65702 84409 65793 84527
rect 65911 84409 66002 84527
rect 65702 84367 66002 84409
rect 65702 84249 65793 84367
rect 65911 84249 66002 84367
rect 65702 66527 66002 84249
rect 65702 66409 65793 66527
rect 65911 66409 66002 66527
rect 65702 66367 66002 66409
rect 65702 66249 65793 66367
rect 65911 66249 66002 66367
rect 65702 48527 66002 66249
rect 65702 48409 65793 48527
rect 65911 48409 66002 48527
rect 65702 48367 66002 48409
rect 65702 48249 65793 48367
rect 65911 48249 66002 48367
rect 65702 30527 66002 48249
rect 65702 30409 65793 30527
rect 65911 30409 66002 30527
rect 65702 30367 66002 30409
rect 65702 30249 65793 30367
rect 65911 30249 66002 30367
rect 65702 12527 66002 30249
rect 65702 12409 65793 12527
rect 65911 12409 66002 12527
rect 65702 12367 66002 12409
rect 65702 12249 65793 12367
rect 65911 12249 66002 12367
rect 65702 -1583 66002 12249
rect 65702 -1701 65793 -1583
rect 65911 -1701 66002 -1583
rect 65702 -1743 66002 -1701
rect 65702 -1861 65793 -1743
rect 65911 -1861 66002 -1743
rect 65702 -1872 66002 -1861
rect 67502 338327 67802 354491
rect 67502 338209 67593 338327
rect 67711 338209 67802 338327
rect 67502 338167 67802 338209
rect 67502 338049 67593 338167
rect 67711 338049 67802 338167
rect 67502 320327 67802 338049
rect 67502 320209 67593 320327
rect 67711 320209 67802 320327
rect 67502 320167 67802 320209
rect 67502 320049 67593 320167
rect 67711 320049 67802 320167
rect 67502 302327 67802 320049
rect 67502 302209 67593 302327
rect 67711 302209 67802 302327
rect 67502 302167 67802 302209
rect 67502 302049 67593 302167
rect 67711 302049 67802 302167
rect 67502 284327 67802 302049
rect 67502 284209 67593 284327
rect 67711 284209 67802 284327
rect 67502 284167 67802 284209
rect 67502 284049 67593 284167
rect 67711 284049 67802 284167
rect 67502 266327 67802 284049
rect 67502 266209 67593 266327
rect 67711 266209 67802 266327
rect 67502 266167 67802 266209
rect 67502 266049 67593 266167
rect 67711 266049 67802 266167
rect 67502 248327 67802 266049
rect 67502 248209 67593 248327
rect 67711 248209 67802 248327
rect 67502 248167 67802 248209
rect 67502 248049 67593 248167
rect 67711 248049 67802 248167
rect 67502 230327 67802 248049
rect 67502 230209 67593 230327
rect 67711 230209 67802 230327
rect 67502 230167 67802 230209
rect 67502 230049 67593 230167
rect 67711 230049 67802 230167
rect 67502 212327 67802 230049
rect 67502 212209 67593 212327
rect 67711 212209 67802 212327
rect 67502 212167 67802 212209
rect 67502 212049 67593 212167
rect 67711 212049 67802 212167
rect 67502 194327 67802 212049
rect 67502 194209 67593 194327
rect 67711 194209 67802 194327
rect 67502 194167 67802 194209
rect 67502 194049 67593 194167
rect 67711 194049 67802 194167
rect 67502 176327 67802 194049
rect 67502 176209 67593 176327
rect 67711 176209 67802 176327
rect 67502 176167 67802 176209
rect 67502 176049 67593 176167
rect 67711 176049 67802 176167
rect 67502 158327 67802 176049
rect 67502 158209 67593 158327
rect 67711 158209 67802 158327
rect 67502 158167 67802 158209
rect 67502 158049 67593 158167
rect 67711 158049 67802 158167
rect 67502 140327 67802 158049
rect 67502 140209 67593 140327
rect 67711 140209 67802 140327
rect 67502 140167 67802 140209
rect 67502 140049 67593 140167
rect 67711 140049 67802 140167
rect 67502 122327 67802 140049
rect 67502 122209 67593 122327
rect 67711 122209 67802 122327
rect 67502 122167 67802 122209
rect 67502 122049 67593 122167
rect 67711 122049 67802 122167
rect 67502 104327 67802 122049
rect 67502 104209 67593 104327
rect 67711 104209 67802 104327
rect 67502 104167 67802 104209
rect 67502 104049 67593 104167
rect 67711 104049 67802 104167
rect 67502 86327 67802 104049
rect 67502 86209 67593 86327
rect 67711 86209 67802 86327
rect 67502 86167 67802 86209
rect 67502 86049 67593 86167
rect 67711 86049 67802 86167
rect 67502 68327 67802 86049
rect 67502 68209 67593 68327
rect 67711 68209 67802 68327
rect 67502 68167 67802 68209
rect 67502 68049 67593 68167
rect 67711 68049 67802 68167
rect 67502 50327 67802 68049
rect 67502 50209 67593 50327
rect 67711 50209 67802 50327
rect 67502 50167 67802 50209
rect 67502 50049 67593 50167
rect 67711 50049 67802 50167
rect 67502 32327 67802 50049
rect 67502 32209 67593 32327
rect 67711 32209 67802 32327
rect 67502 32167 67802 32209
rect 67502 32049 67593 32167
rect 67711 32049 67802 32167
rect 67502 14327 67802 32049
rect 67502 14209 67593 14327
rect 67711 14209 67802 14327
rect 67502 14167 67802 14209
rect 67502 14049 67593 14167
rect 67711 14049 67802 14167
rect 67502 -2523 67802 14049
rect 67502 -2641 67593 -2523
rect 67711 -2641 67802 -2523
rect 67502 -2683 67802 -2641
rect 67502 -2801 67593 -2683
rect 67711 -2801 67802 -2683
rect 67502 -2812 67802 -2801
rect 69302 340127 69602 355431
rect 78302 355239 78602 355720
rect 78302 355121 78393 355239
rect 78511 355121 78602 355239
rect 78302 355079 78602 355121
rect 78302 354961 78393 355079
rect 78511 354961 78602 355079
rect 76502 354299 76802 354780
rect 76502 354181 76593 354299
rect 76711 354181 76802 354299
rect 76502 354139 76802 354181
rect 76502 354021 76593 354139
rect 76711 354021 76802 354139
rect 74702 353359 75002 353840
rect 74702 353241 74793 353359
rect 74911 353241 75002 353359
rect 74702 353199 75002 353241
rect 74702 353081 74793 353199
rect 74911 353081 75002 353199
rect 69302 340009 69393 340127
rect 69511 340009 69602 340127
rect 69302 339967 69602 340009
rect 69302 339849 69393 339967
rect 69511 339849 69602 339967
rect 69302 322127 69602 339849
rect 69302 322009 69393 322127
rect 69511 322009 69602 322127
rect 69302 321967 69602 322009
rect 69302 321849 69393 321967
rect 69511 321849 69602 321967
rect 69302 304127 69602 321849
rect 69302 304009 69393 304127
rect 69511 304009 69602 304127
rect 69302 303967 69602 304009
rect 69302 303849 69393 303967
rect 69511 303849 69602 303967
rect 69302 286127 69602 303849
rect 69302 286009 69393 286127
rect 69511 286009 69602 286127
rect 69302 285967 69602 286009
rect 69302 285849 69393 285967
rect 69511 285849 69602 285967
rect 69302 268127 69602 285849
rect 69302 268009 69393 268127
rect 69511 268009 69602 268127
rect 69302 267967 69602 268009
rect 69302 267849 69393 267967
rect 69511 267849 69602 267967
rect 69302 250127 69602 267849
rect 69302 250009 69393 250127
rect 69511 250009 69602 250127
rect 69302 249967 69602 250009
rect 69302 249849 69393 249967
rect 69511 249849 69602 249967
rect 69302 232127 69602 249849
rect 69302 232009 69393 232127
rect 69511 232009 69602 232127
rect 69302 231967 69602 232009
rect 69302 231849 69393 231967
rect 69511 231849 69602 231967
rect 69302 214127 69602 231849
rect 69302 214009 69393 214127
rect 69511 214009 69602 214127
rect 69302 213967 69602 214009
rect 69302 213849 69393 213967
rect 69511 213849 69602 213967
rect 69302 196127 69602 213849
rect 69302 196009 69393 196127
rect 69511 196009 69602 196127
rect 69302 195967 69602 196009
rect 69302 195849 69393 195967
rect 69511 195849 69602 195967
rect 69302 178127 69602 195849
rect 69302 178009 69393 178127
rect 69511 178009 69602 178127
rect 69302 177967 69602 178009
rect 69302 177849 69393 177967
rect 69511 177849 69602 177967
rect 69302 160127 69602 177849
rect 69302 160009 69393 160127
rect 69511 160009 69602 160127
rect 69302 159967 69602 160009
rect 69302 159849 69393 159967
rect 69511 159849 69602 159967
rect 69302 142127 69602 159849
rect 69302 142009 69393 142127
rect 69511 142009 69602 142127
rect 69302 141967 69602 142009
rect 69302 141849 69393 141967
rect 69511 141849 69602 141967
rect 69302 124127 69602 141849
rect 69302 124009 69393 124127
rect 69511 124009 69602 124127
rect 69302 123967 69602 124009
rect 69302 123849 69393 123967
rect 69511 123849 69602 123967
rect 69302 106127 69602 123849
rect 69302 106009 69393 106127
rect 69511 106009 69602 106127
rect 69302 105967 69602 106009
rect 69302 105849 69393 105967
rect 69511 105849 69602 105967
rect 69302 88127 69602 105849
rect 69302 88009 69393 88127
rect 69511 88009 69602 88127
rect 69302 87967 69602 88009
rect 69302 87849 69393 87967
rect 69511 87849 69602 87967
rect 69302 70127 69602 87849
rect 69302 70009 69393 70127
rect 69511 70009 69602 70127
rect 69302 69967 69602 70009
rect 69302 69849 69393 69967
rect 69511 69849 69602 69967
rect 69302 52127 69602 69849
rect 69302 52009 69393 52127
rect 69511 52009 69602 52127
rect 69302 51967 69602 52009
rect 69302 51849 69393 51967
rect 69511 51849 69602 51967
rect 69302 34127 69602 51849
rect 69302 34009 69393 34127
rect 69511 34009 69602 34127
rect 69302 33967 69602 34009
rect 69302 33849 69393 33967
rect 69511 33849 69602 33967
rect 69302 16127 69602 33849
rect 69302 16009 69393 16127
rect 69511 16009 69602 16127
rect 69302 15967 69602 16009
rect 69302 15849 69393 15967
rect 69511 15849 69602 15967
rect 60302 -3111 60393 -2993
rect 60511 -3111 60602 -2993
rect 60302 -3153 60602 -3111
rect 60302 -3271 60393 -3153
rect 60511 -3271 60602 -3153
rect 60302 -3752 60602 -3271
rect 69302 -3463 69602 15849
rect 72902 352419 73202 352900
rect 72902 352301 72993 352419
rect 73111 352301 73202 352419
rect 72902 352259 73202 352301
rect 72902 352141 72993 352259
rect 73111 352141 73202 352259
rect 72902 343727 73202 352141
rect 72902 343609 72993 343727
rect 73111 343609 73202 343727
rect 72902 343567 73202 343609
rect 72902 343449 72993 343567
rect 73111 343449 73202 343567
rect 72902 325727 73202 343449
rect 72902 325609 72993 325727
rect 73111 325609 73202 325727
rect 72902 325567 73202 325609
rect 72902 325449 72993 325567
rect 73111 325449 73202 325567
rect 72902 307727 73202 325449
rect 72902 307609 72993 307727
rect 73111 307609 73202 307727
rect 72902 307567 73202 307609
rect 72902 307449 72993 307567
rect 73111 307449 73202 307567
rect 72902 289727 73202 307449
rect 72902 289609 72993 289727
rect 73111 289609 73202 289727
rect 72902 289567 73202 289609
rect 72902 289449 72993 289567
rect 73111 289449 73202 289567
rect 72902 271727 73202 289449
rect 72902 271609 72993 271727
rect 73111 271609 73202 271727
rect 72902 271567 73202 271609
rect 72902 271449 72993 271567
rect 73111 271449 73202 271567
rect 72902 253727 73202 271449
rect 72902 253609 72993 253727
rect 73111 253609 73202 253727
rect 72902 253567 73202 253609
rect 72902 253449 72993 253567
rect 73111 253449 73202 253567
rect 72902 235727 73202 253449
rect 72902 235609 72993 235727
rect 73111 235609 73202 235727
rect 72902 235567 73202 235609
rect 72902 235449 72993 235567
rect 73111 235449 73202 235567
rect 72902 217727 73202 235449
rect 72902 217609 72993 217727
rect 73111 217609 73202 217727
rect 72902 217567 73202 217609
rect 72902 217449 72993 217567
rect 73111 217449 73202 217567
rect 72902 199727 73202 217449
rect 72902 199609 72993 199727
rect 73111 199609 73202 199727
rect 72902 199567 73202 199609
rect 72902 199449 72993 199567
rect 73111 199449 73202 199567
rect 72902 181727 73202 199449
rect 72902 181609 72993 181727
rect 73111 181609 73202 181727
rect 72902 181567 73202 181609
rect 72902 181449 72993 181567
rect 73111 181449 73202 181567
rect 72902 163727 73202 181449
rect 72902 163609 72993 163727
rect 73111 163609 73202 163727
rect 72902 163567 73202 163609
rect 72902 163449 72993 163567
rect 73111 163449 73202 163567
rect 72902 145727 73202 163449
rect 72902 145609 72993 145727
rect 73111 145609 73202 145727
rect 72902 145567 73202 145609
rect 72902 145449 72993 145567
rect 73111 145449 73202 145567
rect 72902 127727 73202 145449
rect 72902 127609 72993 127727
rect 73111 127609 73202 127727
rect 72902 127567 73202 127609
rect 72902 127449 72993 127567
rect 73111 127449 73202 127567
rect 72902 109727 73202 127449
rect 72902 109609 72993 109727
rect 73111 109609 73202 109727
rect 72902 109567 73202 109609
rect 72902 109449 72993 109567
rect 73111 109449 73202 109567
rect 72902 91727 73202 109449
rect 72902 91609 72993 91727
rect 73111 91609 73202 91727
rect 72902 91567 73202 91609
rect 72902 91449 72993 91567
rect 73111 91449 73202 91567
rect 72902 73727 73202 91449
rect 72902 73609 72993 73727
rect 73111 73609 73202 73727
rect 72902 73567 73202 73609
rect 72902 73449 72993 73567
rect 73111 73449 73202 73567
rect 72902 55727 73202 73449
rect 72902 55609 72993 55727
rect 73111 55609 73202 55727
rect 72902 55567 73202 55609
rect 72902 55449 72993 55567
rect 73111 55449 73202 55567
rect 72902 37727 73202 55449
rect 72902 37609 72993 37727
rect 73111 37609 73202 37727
rect 72902 37567 73202 37609
rect 72902 37449 72993 37567
rect 73111 37449 73202 37567
rect 72902 19727 73202 37449
rect 72902 19609 72993 19727
rect 73111 19609 73202 19727
rect 72902 19567 73202 19609
rect 72902 19449 72993 19567
rect 73111 19449 73202 19567
rect 72902 1727 73202 19449
rect 72902 1609 72993 1727
rect 73111 1609 73202 1727
rect 72902 1567 73202 1609
rect 72902 1449 72993 1567
rect 73111 1449 73202 1567
rect 72902 -173 73202 1449
rect 72902 -291 72993 -173
rect 73111 -291 73202 -173
rect 72902 -333 73202 -291
rect 72902 -451 72993 -333
rect 73111 -451 73202 -333
rect 72902 -932 73202 -451
rect 74702 345527 75002 353081
rect 74702 345409 74793 345527
rect 74911 345409 75002 345527
rect 74702 345367 75002 345409
rect 74702 345249 74793 345367
rect 74911 345249 75002 345367
rect 74702 327527 75002 345249
rect 74702 327409 74793 327527
rect 74911 327409 75002 327527
rect 74702 327367 75002 327409
rect 74702 327249 74793 327367
rect 74911 327249 75002 327367
rect 74702 309527 75002 327249
rect 74702 309409 74793 309527
rect 74911 309409 75002 309527
rect 74702 309367 75002 309409
rect 74702 309249 74793 309367
rect 74911 309249 75002 309367
rect 74702 291527 75002 309249
rect 74702 291409 74793 291527
rect 74911 291409 75002 291527
rect 74702 291367 75002 291409
rect 74702 291249 74793 291367
rect 74911 291249 75002 291367
rect 74702 273527 75002 291249
rect 74702 273409 74793 273527
rect 74911 273409 75002 273527
rect 74702 273367 75002 273409
rect 74702 273249 74793 273367
rect 74911 273249 75002 273367
rect 74702 255527 75002 273249
rect 74702 255409 74793 255527
rect 74911 255409 75002 255527
rect 74702 255367 75002 255409
rect 74702 255249 74793 255367
rect 74911 255249 75002 255367
rect 74702 237527 75002 255249
rect 74702 237409 74793 237527
rect 74911 237409 75002 237527
rect 74702 237367 75002 237409
rect 74702 237249 74793 237367
rect 74911 237249 75002 237367
rect 74702 219527 75002 237249
rect 74702 219409 74793 219527
rect 74911 219409 75002 219527
rect 74702 219367 75002 219409
rect 74702 219249 74793 219367
rect 74911 219249 75002 219367
rect 74702 201527 75002 219249
rect 74702 201409 74793 201527
rect 74911 201409 75002 201527
rect 74702 201367 75002 201409
rect 74702 201249 74793 201367
rect 74911 201249 75002 201367
rect 74702 183527 75002 201249
rect 74702 183409 74793 183527
rect 74911 183409 75002 183527
rect 74702 183367 75002 183409
rect 74702 183249 74793 183367
rect 74911 183249 75002 183367
rect 74702 165527 75002 183249
rect 74702 165409 74793 165527
rect 74911 165409 75002 165527
rect 74702 165367 75002 165409
rect 74702 165249 74793 165367
rect 74911 165249 75002 165367
rect 74702 147527 75002 165249
rect 74702 147409 74793 147527
rect 74911 147409 75002 147527
rect 74702 147367 75002 147409
rect 74702 147249 74793 147367
rect 74911 147249 75002 147367
rect 74702 129527 75002 147249
rect 74702 129409 74793 129527
rect 74911 129409 75002 129527
rect 74702 129367 75002 129409
rect 74702 129249 74793 129367
rect 74911 129249 75002 129367
rect 74702 111527 75002 129249
rect 74702 111409 74793 111527
rect 74911 111409 75002 111527
rect 74702 111367 75002 111409
rect 74702 111249 74793 111367
rect 74911 111249 75002 111367
rect 74702 93527 75002 111249
rect 74702 93409 74793 93527
rect 74911 93409 75002 93527
rect 74702 93367 75002 93409
rect 74702 93249 74793 93367
rect 74911 93249 75002 93367
rect 74702 75527 75002 93249
rect 74702 75409 74793 75527
rect 74911 75409 75002 75527
rect 74702 75367 75002 75409
rect 74702 75249 74793 75367
rect 74911 75249 75002 75367
rect 74702 57527 75002 75249
rect 74702 57409 74793 57527
rect 74911 57409 75002 57527
rect 74702 57367 75002 57409
rect 74702 57249 74793 57367
rect 74911 57249 75002 57367
rect 74702 39527 75002 57249
rect 74702 39409 74793 39527
rect 74911 39409 75002 39527
rect 74702 39367 75002 39409
rect 74702 39249 74793 39367
rect 74911 39249 75002 39367
rect 74702 21527 75002 39249
rect 74702 21409 74793 21527
rect 74911 21409 75002 21527
rect 74702 21367 75002 21409
rect 74702 21249 74793 21367
rect 74911 21249 75002 21367
rect 74702 3527 75002 21249
rect 74702 3409 74793 3527
rect 74911 3409 75002 3527
rect 74702 3367 75002 3409
rect 74702 3249 74793 3367
rect 74911 3249 75002 3367
rect 74702 -1113 75002 3249
rect 74702 -1231 74793 -1113
rect 74911 -1231 75002 -1113
rect 74702 -1273 75002 -1231
rect 74702 -1391 74793 -1273
rect 74911 -1391 75002 -1273
rect 74702 -1872 75002 -1391
rect 76502 347327 76802 354021
rect 76502 347209 76593 347327
rect 76711 347209 76802 347327
rect 76502 347167 76802 347209
rect 76502 347049 76593 347167
rect 76711 347049 76802 347167
rect 76502 329327 76802 347049
rect 76502 329209 76593 329327
rect 76711 329209 76802 329327
rect 76502 329167 76802 329209
rect 76502 329049 76593 329167
rect 76711 329049 76802 329167
rect 76502 311327 76802 329049
rect 76502 311209 76593 311327
rect 76711 311209 76802 311327
rect 76502 311167 76802 311209
rect 76502 311049 76593 311167
rect 76711 311049 76802 311167
rect 76502 293327 76802 311049
rect 76502 293209 76593 293327
rect 76711 293209 76802 293327
rect 76502 293167 76802 293209
rect 76502 293049 76593 293167
rect 76711 293049 76802 293167
rect 76502 275327 76802 293049
rect 76502 275209 76593 275327
rect 76711 275209 76802 275327
rect 76502 275167 76802 275209
rect 76502 275049 76593 275167
rect 76711 275049 76802 275167
rect 76502 257327 76802 275049
rect 76502 257209 76593 257327
rect 76711 257209 76802 257327
rect 76502 257167 76802 257209
rect 76502 257049 76593 257167
rect 76711 257049 76802 257167
rect 76502 239327 76802 257049
rect 76502 239209 76593 239327
rect 76711 239209 76802 239327
rect 76502 239167 76802 239209
rect 76502 239049 76593 239167
rect 76711 239049 76802 239167
rect 76502 221327 76802 239049
rect 76502 221209 76593 221327
rect 76711 221209 76802 221327
rect 76502 221167 76802 221209
rect 76502 221049 76593 221167
rect 76711 221049 76802 221167
rect 76502 203327 76802 221049
rect 76502 203209 76593 203327
rect 76711 203209 76802 203327
rect 76502 203167 76802 203209
rect 76502 203049 76593 203167
rect 76711 203049 76802 203167
rect 76502 185327 76802 203049
rect 76502 185209 76593 185327
rect 76711 185209 76802 185327
rect 76502 185167 76802 185209
rect 76502 185049 76593 185167
rect 76711 185049 76802 185167
rect 76502 167327 76802 185049
rect 76502 167209 76593 167327
rect 76711 167209 76802 167327
rect 76502 167167 76802 167209
rect 76502 167049 76593 167167
rect 76711 167049 76802 167167
rect 76502 149327 76802 167049
rect 76502 149209 76593 149327
rect 76711 149209 76802 149327
rect 76502 149167 76802 149209
rect 76502 149049 76593 149167
rect 76711 149049 76802 149167
rect 76502 131327 76802 149049
rect 76502 131209 76593 131327
rect 76711 131209 76802 131327
rect 76502 131167 76802 131209
rect 76502 131049 76593 131167
rect 76711 131049 76802 131167
rect 76502 113327 76802 131049
rect 76502 113209 76593 113327
rect 76711 113209 76802 113327
rect 76502 113167 76802 113209
rect 76502 113049 76593 113167
rect 76711 113049 76802 113167
rect 76502 95327 76802 113049
rect 76502 95209 76593 95327
rect 76711 95209 76802 95327
rect 76502 95167 76802 95209
rect 76502 95049 76593 95167
rect 76711 95049 76802 95167
rect 76502 77327 76802 95049
rect 76502 77209 76593 77327
rect 76711 77209 76802 77327
rect 76502 77167 76802 77209
rect 76502 77049 76593 77167
rect 76711 77049 76802 77167
rect 76502 59327 76802 77049
rect 76502 59209 76593 59327
rect 76711 59209 76802 59327
rect 76502 59167 76802 59209
rect 76502 59049 76593 59167
rect 76711 59049 76802 59167
rect 76502 41327 76802 59049
rect 76502 41209 76593 41327
rect 76711 41209 76802 41327
rect 76502 41167 76802 41209
rect 76502 41049 76593 41167
rect 76711 41049 76802 41167
rect 76502 23327 76802 41049
rect 76502 23209 76593 23327
rect 76711 23209 76802 23327
rect 76502 23167 76802 23209
rect 76502 23049 76593 23167
rect 76711 23049 76802 23167
rect 76502 5327 76802 23049
rect 76502 5209 76593 5327
rect 76711 5209 76802 5327
rect 76502 5167 76802 5209
rect 76502 5049 76593 5167
rect 76711 5049 76802 5167
rect 76502 -2053 76802 5049
rect 76502 -2171 76593 -2053
rect 76711 -2171 76802 -2053
rect 76502 -2213 76802 -2171
rect 76502 -2331 76593 -2213
rect 76711 -2331 76802 -2213
rect 76502 -2812 76802 -2331
rect 78302 349127 78602 354961
rect 87302 355709 87602 355720
rect 87302 355591 87393 355709
rect 87511 355591 87602 355709
rect 87302 355549 87602 355591
rect 87302 355431 87393 355549
rect 87511 355431 87602 355549
rect 85502 354769 85802 354780
rect 85502 354651 85593 354769
rect 85711 354651 85802 354769
rect 85502 354609 85802 354651
rect 85502 354491 85593 354609
rect 85711 354491 85802 354609
rect 83702 353829 84002 353840
rect 83702 353711 83793 353829
rect 83911 353711 84002 353829
rect 83702 353669 84002 353711
rect 83702 353551 83793 353669
rect 83911 353551 84002 353669
rect 78302 349009 78393 349127
rect 78511 349009 78602 349127
rect 78302 348967 78602 349009
rect 78302 348849 78393 348967
rect 78511 348849 78602 348967
rect 78302 331127 78602 348849
rect 78302 331009 78393 331127
rect 78511 331009 78602 331127
rect 78302 330967 78602 331009
rect 78302 330849 78393 330967
rect 78511 330849 78602 330967
rect 78302 313127 78602 330849
rect 78302 313009 78393 313127
rect 78511 313009 78602 313127
rect 78302 312967 78602 313009
rect 78302 312849 78393 312967
rect 78511 312849 78602 312967
rect 78302 295127 78602 312849
rect 78302 295009 78393 295127
rect 78511 295009 78602 295127
rect 78302 294967 78602 295009
rect 78302 294849 78393 294967
rect 78511 294849 78602 294967
rect 78302 277127 78602 294849
rect 78302 277009 78393 277127
rect 78511 277009 78602 277127
rect 78302 276967 78602 277009
rect 78302 276849 78393 276967
rect 78511 276849 78602 276967
rect 78302 259127 78602 276849
rect 78302 259009 78393 259127
rect 78511 259009 78602 259127
rect 78302 258967 78602 259009
rect 78302 258849 78393 258967
rect 78511 258849 78602 258967
rect 78302 241127 78602 258849
rect 78302 241009 78393 241127
rect 78511 241009 78602 241127
rect 78302 240967 78602 241009
rect 78302 240849 78393 240967
rect 78511 240849 78602 240967
rect 78302 223127 78602 240849
rect 78302 223009 78393 223127
rect 78511 223009 78602 223127
rect 78302 222967 78602 223009
rect 78302 222849 78393 222967
rect 78511 222849 78602 222967
rect 78302 205127 78602 222849
rect 78302 205009 78393 205127
rect 78511 205009 78602 205127
rect 78302 204967 78602 205009
rect 78302 204849 78393 204967
rect 78511 204849 78602 204967
rect 78302 187127 78602 204849
rect 78302 187009 78393 187127
rect 78511 187009 78602 187127
rect 78302 186967 78602 187009
rect 78302 186849 78393 186967
rect 78511 186849 78602 186967
rect 78302 169127 78602 186849
rect 78302 169009 78393 169127
rect 78511 169009 78602 169127
rect 78302 168967 78602 169009
rect 78302 168849 78393 168967
rect 78511 168849 78602 168967
rect 78302 151127 78602 168849
rect 78302 151009 78393 151127
rect 78511 151009 78602 151127
rect 78302 150967 78602 151009
rect 78302 150849 78393 150967
rect 78511 150849 78602 150967
rect 78302 133127 78602 150849
rect 78302 133009 78393 133127
rect 78511 133009 78602 133127
rect 78302 132967 78602 133009
rect 78302 132849 78393 132967
rect 78511 132849 78602 132967
rect 78302 115127 78602 132849
rect 78302 115009 78393 115127
rect 78511 115009 78602 115127
rect 78302 114967 78602 115009
rect 78302 114849 78393 114967
rect 78511 114849 78602 114967
rect 78302 97127 78602 114849
rect 78302 97009 78393 97127
rect 78511 97009 78602 97127
rect 78302 96967 78602 97009
rect 78302 96849 78393 96967
rect 78511 96849 78602 96967
rect 78302 79127 78602 96849
rect 78302 79009 78393 79127
rect 78511 79009 78602 79127
rect 78302 78967 78602 79009
rect 78302 78849 78393 78967
rect 78511 78849 78602 78967
rect 78302 61127 78602 78849
rect 78302 61009 78393 61127
rect 78511 61009 78602 61127
rect 78302 60967 78602 61009
rect 78302 60849 78393 60967
rect 78511 60849 78602 60967
rect 78302 43127 78602 60849
rect 78302 43009 78393 43127
rect 78511 43009 78602 43127
rect 78302 42967 78602 43009
rect 78302 42849 78393 42967
rect 78511 42849 78602 42967
rect 78302 25127 78602 42849
rect 78302 25009 78393 25127
rect 78511 25009 78602 25127
rect 78302 24967 78602 25009
rect 78302 24849 78393 24967
rect 78511 24849 78602 24967
rect 78302 7127 78602 24849
rect 78302 7009 78393 7127
rect 78511 7009 78602 7127
rect 78302 6967 78602 7009
rect 78302 6849 78393 6967
rect 78511 6849 78602 6967
rect 69302 -3581 69393 -3463
rect 69511 -3581 69602 -3463
rect 69302 -3623 69602 -3581
rect 69302 -3741 69393 -3623
rect 69511 -3741 69602 -3623
rect 69302 -3752 69602 -3741
rect 78302 -2993 78602 6849
rect 81902 352889 82202 352900
rect 81902 352771 81993 352889
rect 82111 352771 82202 352889
rect 81902 352729 82202 352771
rect 81902 352611 81993 352729
rect 82111 352611 82202 352729
rect 81902 334727 82202 352611
rect 81902 334609 81993 334727
rect 82111 334609 82202 334727
rect 81902 334567 82202 334609
rect 81902 334449 81993 334567
rect 82111 334449 82202 334567
rect 81902 316727 82202 334449
rect 81902 316609 81993 316727
rect 82111 316609 82202 316727
rect 81902 316567 82202 316609
rect 81902 316449 81993 316567
rect 82111 316449 82202 316567
rect 81902 298727 82202 316449
rect 81902 298609 81993 298727
rect 82111 298609 82202 298727
rect 81902 298567 82202 298609
rect 81902 298449 81993 298567
rect 82111 298449 82202 298567
rect 81902 280727 82202 298449
rect 81902 280609 81993 280727
rect 82111 280609 82202 280727
rect 81902 280567 82202 280609
rect 81902 280449 81993 280567
rect 82111 280449 82202 280567
rect 81902 262727 82202 280449
rect 81902 262609 81993 262727
rect 82111 262609 82202 262727
rect 81902 262567 82202 262609
rect 81902 262449 81993 262567
rect 82111 262449 82202 262567
rect 81902 244727 82202 262449
rect 81902 244609 81993 244727
rect 82111 244609 82202 244727
rect 81902 244567 82202 244609
rect 81902 244449 81993 244567
rect 82111 244449 82202 244567
rect 81902 226727 82202 244449
rect 81902 226609 81993 226727
rect 82111 226609 82202 226727
rect 81902 226567 82202 226609
rect 81902 226449 81993 226567
rect 82111 226449 82202 226567
rect 81902 208727 82202 226449
rect 81902 208609 81993 208727
rect 82111 208609 82202 208727
rect 81902 208567 82202 208609
rect 81902 208449 81993 208567
rect 82111 208449 82202 208567
rect 81902 190727 82202 208449
rect 81902 190609 81993 190727
rect 82111 190609 82202 190727
rect 81902 190567 82202 190609
rect 81902 190449 81993 190567
rect 82111 190449 82202 190567
rect 81902 172727 82202 190449
rect 81902 172609 81993 172727
rect 82111 172609 82202 172727
rect 81902 172567 82202 172609
rect 81902 172449 81993 172567
rect 82111 172449 82202 172567
rect 81902 154727 82202 172449
rect 81902 154609 81993 154727
rect 82111 154609 82202 154727
rect 81902 154567 82202 154609
rect 81902 154449 81993 154567
rect 82111 154449 82202 154567
rect 81902 136727 82202 154449
rect 81902 136609 81993 136727
rect 82111 136609 82202 136727
rect 81902 136567 82202 136609
rect 81902 136449 81993 136567
rect 82111 136449 82202 136567
rect 81902 118727 82202 136449
rect 81902 118609 81993 118727
rect 82111 118609 82202 118727
rect 81902 118567 82202 118609
rect 81902 118449 81993 118567
rect 82111 118449 82202 118567
rect 81902 100727 82202 118449
rect 81902 100609 81993 100727
rect 82111 100609 82202 100727
rect 81902 100567 82202 100609
rect 81902 100449 81993 100567
rect 82111 100449 82202 100567
rect 81902 82727 82202 100449
rect 81902 82609 81993 82727
rect 82111 82609 82202 82727
rect 81902 82567 82202 82609
rect 81902 82449 81993 82567
rect 82111 82449 82202 82567
rect 81902 64727 82202 82449
rect 81902 64609 81993 64727
rect 82111 64609 82202 64727
rect 81902 64567 82202 64609
rect 81902 64449 81993 64567
rect 82111 64449 82202 64567
rect 81902 46727 82202 64449
rect 81902 46609 81993 46727
rect 82111 46609 82202 46727
rect 81902 46567 82202 46609
rect 81902 46449 81993 46567
rect 82111 46449 82202 46567
rect 81902 28727 82202 46449
rect 81902 28609 81993 28727
rect 82111 28609 82202 28727
rect 81902 28567 82202 28609
rect 81902 28449 81993 28567
rect 82111 28449 82202 28567
rect 81902 10727 82202 28449
rect 81902 10609 81993 10727
rect 82111 10609 82202 10727
rect 81902 10567 82202 10609
rect 81902 10449 81993 10567
rect 82111 10449 82202 10567
rect 81902 -643 82202 10449
rect 81902 -761 81993 -643
rect 82111 -761 82202 -643
rect 81902 -803 82202 -761
rect 81902 -921 81993 -803
rect 82111 -921 82202 -803
rect 81902 -932 82202 -921
rect 83702 336527 84002 353551
rect 83702 336409 83793 336527
rect 83911 336409 84002 336527
rect 83702 336367 84002 336409
rect 83702 336249 83793 336367
rect 83911 336249 84002 336367
rect 83702 318527 84002 336249
rect 83702 318409 83793 318527
rect 83911 318409 84002 318527
rect 83702 318367 84002 318409
rect 83702 318249 83793 318367
rect 83911 318249 84002 318367
rect 83702 300527 84002 318249
rect 83702 300409 83793 300527
rect 83911 300409 84002 300527
rect 83702 300367 84002 300409
rect 83702 300249 83793 300367
rect 83911 300249 84002 300367
rect 83702 282527 84002 300249
rect 83702 282409 83793 282527
rect 83911 282409 84002 282527
rect 83702 282367 84002 282409
rect 83702 282249 83793 282367
rect 83911 282249 84002 282367
rect 83702 264527 84002 282249
rect 83702 264409 83793 264527
rect 83911 264409 84002 264527
rect 83702 264367 84002 264409
rect 83702 264249 83793 264367
rect 83911 264249 84002 264367
rect 83702 246527 84002 264249
rect 83702 246409 83793 246527
rect 83911 246409 84002 246527
rect 83702 246367 84002 246409
rect 83702 246249 83793 246367
rect 83911 246249 84002 246367
rect 83702 228527 84002 246249
rect 83702 228409 83793 228527
rect 83911 228409 84002 228527
rect 83702 228367 84002 228409
rect 83702 228249 83793 228367
rect 83911 228249 84002 228367
rect 83702 210527 84002 228249
rect 83702 210409 83793 210527
rect 83911 210409 84002 210527
rect 83702 210367 84002 210409
rect 83702 210249 83793 210367
rect 83911 210249 84002 210367
rect 83702 192527 84002 210249
rect 83702 192409 83793 192527
rect 83911 192409 84002 192527
rect 83702 192367 84002 192409
rect 83702 192249 83793 192367
rect 83911 192249 84002 192367
rect 83702 174527 84002 192249
rect 83702 174409 83793 174527
rect 83911 174409 84002 174527
rect 83702 174367 84002 174409
rect 83702 174249 83793 174367
rect 83911 174249 84002 174367
rect 83702 156527 84002 174249
rect 83702 156409 83793 156527
rect 83911 156409 84002 156527
rect 83702 156367 84002 156409
rect 83702 156249 83793 156367
rect 83911 156249 84002 156367
rect 83702 138527 84002 156249
rect 83702 138409 83793 138527
rect 83911 138409 84002 138527
rect 83702 138367 84002 138409
rect 83702 138249 83793 138367
rect 83911 138249 84002 138367
rect 83702 120527 84002 138249
rect 83702 120409 83793 120527
rect 83911 120409 84002 120527
rect 83702 120367 84002 120409
rect 83702 120249 83793 120367
rect 83911 120249 84002 120367
rect 83702 102527 84002 120249
rect 83702 102409 83793 102527
rect 83911 102409 84002 102527
rect 83702 102367 84002 102409
rect 83702 102249 83793 102367
rect 83911 102249 84002 102367
rect 83702 84527 84002 102249
rect 83702 84409 83793 84527
rect 83911 84409 84002 84527
rect 83702 84367 84002 84409
rect 83702 84249 83793 84367
rect 83911 84249 84002 84367
rect 83702 66527 84002 84249
rect 83702 66409 83793 66527
rect 83911 66409 84002 66527
rect 83702 66367 84002 66409
rect 83702 66249 83793 66367
rect 83911 66249 84002 66367
rect 83702 48527 84002 66249
rect 83702 48409 83793 48527
rect 83911 48409 84002 48527
rect 83702 48367 84002 48409
rect 83702 48249 83793 48367
rect 83911 48249 84002 48367
rect 83702 30527 84002 48249
rect 83702 30409 83793 30527
rect 83911 30409 84002 30527
rect 83702 30367 84002 30409
rect 83702 30249 83793 30367
rect 83911 30249 84002 30367
rect 83702 12527 84002 30249
rect 83702 12409 83793 12527
rect 83911 12409 84002 12527
rect 83702 12367 84002 12409
rect 83702 12249 83793 12367
rect 83911 12249 84002 12367
rect 83702 -1583 84002 12249
rect 83702 -1701 83793 -1583
rect 83911 -1701 84002 -1583
rect 83702 -1743 84002 -1701
rect 83702 -1861 83793 -1743
rect 83911 -1861 84002 -1743
rect 83702 -1872 84002 -1861
rect 85502 338327 85802 354491
rect 85502 338209 85593 338327
rect 85711 338209 85802 338327
rect 85502 338167 85802 338209
rect 85502 338049 85593 338167
rect 85711 338049 85802 338167
rect 85502 320327 85802 338049
rect 85502 320209 85593 320327
rect 85711 320209 85802 320327
rect 85502 320167 85802 320209
rect 85502 320049 85593 320167
rect 85711 320049 85802 320167
rect 85502 302327 85802 320049
rect 85502 302209 85593 302327
rect 85711 302209 85802 302327
rect 85502 302167 85802 302209
rect 85502 302049 85593 302167
rect 85711 302049 85802 302167
rect 85502 284327 85802 302049
rect 85502 284209 85593 284327
rect 85711 284209 85802 284327
rect 85502 284167 85802 284209
rect 85502 284049 85593 284167
rect 85711 284049 85802 284167
rect 85502 266327 85802 284049
rect 85502 266209 85593 266327
rect 85711 266209 85802 266327
rect 85502 266167 85802 266209
rect 85502 266049 85593 266167
rect 85711 266049 85802 266167
rect 85502 248327 85802 266049
rect 85502 248209 85593 248327
rect 85711 248209 85802 248327
rect 85502 248167 85802 248209
rect 85502 248049 85593 248167
rect 85711 248049 85802 248167
rect 85502 230327 85802 248049
rect 85502 230209 85593 230327
rect 85711 230209 85802 230327
rect 85502 230167 85802 230209
rect 85502 230049 85593 230167
rect 85711 230049 85802 230167
rect 85502 212327 85802 230049
rect 85502 212209 85593 212327
rect 85711 212209 85802 212327
rect 85502 212167 85802 212209
rect 85502 212049 85593 212167
rect 85711 212049 85802 212167
rect 85502 194327 85802 212049
rect 85502 194209 85593 194327
rect 85711 194209 85802 194327
rect 85502 194167 85802 194209
rect 85502 194049 85593 194167
rect 85711 194049 85802 194167
rect 85502 176327 85802 194049
rect 85502 176209 85593 176327
rect 85711 176209 85802 176327
rect 85502 176167 85802 176209
rect 85502 176049 85593 176167
rect 85711 176049 85802 176167
rect 85502 158327 85802 176049
rect 85502 158209 85593 158327
rect 85711 158209 85802 158327
rect 85502 158167 85802 158209
rect 85502 158049 85593 158167
rect 85711 158049 85802 158167
rect 85502 140327 85802 158049
rect 85502 140209 85593 140327
rect 85711 140209 85802 140327
rect 85502 140167 85802 140209
rect 85502 140049 85593 140167
rect 85711 140049 85802 140167
rect 85502 122327 85802 140049
rect 85502 122209 85593 122327
rect 85711 122209 85802 122327
rect 85502 122167 85802 122209
rect 85502 122049 85593 122167
rect 85711 122049 85802 122167
rect 85502 104327 85802 122049
rect 85502 104209 85593 104327
rect 85711 104209 85802 104327
rect 85502 104167 85802 104209
rect 85502 104049 85593 104167
rect 85711 104049 85802 104167
rect 85502 86327 85802 104049
rect 85502 86209 85593 86327
rect 85711 86209 85802 86327
rect 85502 86167 85802 86209
rect 85502 86049 85593 86167
rect 85711 86049 85802 86167
rect 85502 68327 85802 86049
rect 85502 68209 85593 68327
rect 85711 68209 85802 68327
rect 85502 68167 85802 68209
rect 85502 68049 85593 68167
rect 85711 68049 85802 68167
rect 85502 50327 85802 68049
rect 85502 50209 85593 50327
rect 85711 50209 85802 50327
rect 85502 50167 85802 50209
rect 85502 50049 85593 50167
rect 85711 50049 85802 50167
rect 85502 32327 85802 50049
rect 85502 32209 85593 32327
rect 85711 32209 85802 32327
rect 85502 32167 85802 32209
rect 85502 32049 85593 32167
rect 85711 32049 85802 32167
rect 85502 14327 85802 32049
rect 85502 14209 85593 14327
rect 85711 14209 85802 14327
rect 85502 14167 85802 14209
rect 85502 14049 85593 14167
rect 85711 14049 85802 14167
rect 85502 -2523 85802 14049
rect 85502 -2641 85593 -2523
rect 85711 -2641 85802 -2523
rect 85502 -2683 85802 -2641
rect 85502 -2801 85593 -2683
rect 85711 -2801 85802 -2683
rect 85502 -2812 85802 -2801
rect 87302 340127 87602 355431
rect 96302 355239 96602 355720
rect 96302 355121 96393 355239
rect 96511 355121 96602 355239
rect 96302 355079 96602 355121
rect 96302 354961 96393 355079
rect 96511 354961 96602 355079
rect 94502 354299 94802 354780
rect 94502 354181 94593 354299
rect 94711 354181 94802 354299
rect 94502 354139 94802 354181
rect 94502 354021 94593 354139
rect 94711 354021 94802 354139
rect 92702 353359 93002 353840
rect 92702 353241 92793 353359
rect 92911 353241 93002 353359
rect 92702 353199 93002 353241
rect 92702 353081 92793 353199
rect 92911 353081 93002 353199
rect 87302 340009 87393 340127
rect 87511 340009 87602 340127
rect 87302 339967 87602 340009
rect 87302 339849 87393 339967
rect 87511 339849 87602 339967
rect 87302 322127 87602 339849
rect 87302 322009 87393 322127
rect 87511 322009 87602 322127
rect 87302 321967 87602 322009
rect 87302 321849 87393 321967
rect 87511 321849 87602 321967
rect 87302 304127 87602 321849
rect 87302 304009 87393 304127
rect 87511 304009 87602 304127
rect 87302 303967 87602 304009
rect 87302 303849 87393 303967
rect 87511 303849 87602 303967
rect 87302 286127 87602 303849
rect 87302 286009 87393 286127
rect 87511 286009 87602 286127
rect 87302 285967 87602 286009
rect 87302 285849 87393 285967
rect 87511 285849 87602 285967
rect 87302 268127 87602 285849
rect 87302 268009 87393 268127
rect 87511 268009 87602 268127
rect 87302 267967 87602 268009
rect 87302 267849 87393 267967
rect 87511 267849 87602 267967
rect 87302 250127 87602 267849
rect 87302 250009 87393 250127
rect 87511 250009 87602 250127
rect 87302 249967 87602 250009
rect 87302 249849 87393 249967
rect 87511 249849 87602 249967
rect 87302 232127 87602 249849
rect 87302 232009 87393 232127
rect 87511 232009 87602 232127
rect 87302 231967 87602 232009
rect 87302 231849 87393 231967
rect 87511 231849 87602 231967
rect 87302 214127 87602 231849
rect 87302 214009 87393 214127
rect 87511 214009 87602 214127
rect 87302 213967 87602 214009
rect 87302 213849 87393 213967
rect 87511 213849 87602 213967
rect 87302 196127 87602 213849
rect 87302 196009 87393 196127
rect 87511 196009 87602 196127
rect 87302 195967 87602 196009
rect 87302 195849 87393 195967
rect 87511 195849 87602 195967
rect 87302 178127 87602 195849
rect 87302 178009 87393 178127
rect 87511 178009 87602 178127
rect 87302 177967 87602 178009
rect 87302 177849 87393 177967
rect 87511 177849 87602 177967
rect 87302 160127 87602 177849
rect 87302 160009 87393 160127
rect 87511 160009 87602 160127
rect 87302 159967 87602 160009
rect 87302 159849 87393 159967
rect 87511 159849 87602 159967
rect 87302 142127 87602 159849
rect 87302 142009 87393 142127
rect 87511 142009 87602 142127
rect 87302 141967 87602 142009
rect 87302 141849 87393 141967
rect 87511 141849 87602 141967
rect 87302 124127 87602 141849
rect 87302 124009 87393 124127
rect 87511 124009 87602 124127
rect 87302 123967 87602 124009
rect 87302 123849 87393 123967
rect 87511 123849 87602 123967
rect 87302 106127 87602 123849
rect 87302 106009 87393 106127
rect 87511 106009 87602 106127
rect 87302 105967 87602 106009
rect 87302 105849 87393 105967
rect 87511 105849 87602 105967
rect 87302 88127 87602 105849
rect 87302 88009 87393 88127
rect 87511 88009 87602 88127
rect 87302 87967 87602 88009
rect 87302 87849 87393 87967
rect 87511 87849 87602 87967
rect 87302 70127 87602 87849
rect 87302 70009 87393 70127
rect 87511 70009 87602 70127
rect 87302 69967 87602 70009
rect 87302 69849 87393 69967
rect 87511 69849 87602 69967
rect 87302 52127 87602 69849
rect 87302 52009 87393 52127
rect 87511 52009 87602 52127
rect 87302 51967 87602 52009
rect 87302 51849 87393 51967
rect 87511 51849 87602 51967
rect 87302 34127 87602 51849
rect 87302 34009 87393 34127
rect 87511 34009 87602 34127
rect 87302 33967 87602 34009
rect 87302 33849 87393 33967
rect 87511 33849 87602 33967
rect 87302 16127 87602 33849
rect 87302 16009 87393 16127
rect 87511 16009 87602 16127
rect 87302 15967 87602 16009
rect 87302 15849 87393 15967
rect 87511 15849 87602 15967
rect 78302 -3111 78393 -2993
rect 78511 -3111 78602 -2993
rect 78302 -3153 78602 -3111
rect 78302 -3271 78393 -3153
rect 78511 -3271 78602 -3153
rect 78302 -3752 78602 -3271
rect 87302 -3463 87602 15849
rect 90902 352419 91202 352900
rect 90902 352301 90993 352419
rect 91111 352301 91202 352419
rect 90902 352259 91202 352301
rect 90902 352141 90993 352259
rect 91111 352141 91202 352259
rect 90902 343727 91202 352141
rect 90902 343609 90993 343727
rect 91111 343609 91202 343727
rect 90902 343567 91202 343609
rect 90902 343449 90993 343567
rect 91111 343449 91202 343567
rect 90902 325727 91202 343449
rect 90902 325609 90993 325727
rect 91111 325609 91202 325727
rect 90902 325567 91202 325609
rect 90902 325449 90993 325567
rect 91111 325449 91202 325567
rect 90902 307727 91202 325449
rect 90902 307609 90993 307727
rect 91111 307609 91202 307727
rect 90902 307567 91202 307609
rect 90902 307449 90993 307567
rect 91111 307449 91202 307567
rect 90902 289727 91202 307449
rect 90902 289609 90993 289727
rect 91111 289609 91202 289727
rect 90902 289567 91202 289609
rect 90902 289449 90993 289567
rect 91111 289449 91202 289567
rect 90902 271727 91202 289449
rect 90902 271609 90993 271727
rect 91111 271609 91202 271727
rect 90902 271567 91202 271609
rect 90902 271449 90993 271567
rect 91111 271449 91202 271567
rect 90902 253727 91202 271449
rect 90902 253609 90993 253727
rect 91111 253609 91202 253727
rect 90902 253567 91202 253609
rect 90902 253449 90993 253567
rect 91111 253449 91202 253567
rect 90902 235727 91202 253449
rect 90902 235609 90993 235727
rect 91111 235609 91202 235727
rect 90902 235567 91202 235609
rect 90902 235449 90993 235567
rect 91111 235449 91202 235567
rect 90902 217727 91202 235449
rect 90902 217609 90993 217727
rect 91111 217609 91202 217727
rect 90902 217567 91202 217609
rect 90902 217449 90993 217567
rect 91111 217449 91202 217567
rect 90902 199727 91202 217449
rect 90902 199609 90993 199727
rect 91111 199609 91202 199727
rect 90902 199567 91202 199609
rect 90902 199449 90993 199567
rect 91111 199449 91202 199567
rect 90902 181727 91202 199449
rect 90902 181609 90993 181727
rect 91111 181609 91202 181727
rect 90902 181567 91202 181609
rect 90902 181449 90993 181567
rect 91111 181449 91202 181567
rect 90902 163727 91202 181449
rect 90902 163609 90993 163727
rect 91111 163609 91202 163727
rect 90902 163567 91202 163609
rect 90902 163449 90993 163567
rect 91111 163449 91202 163567
rect 90902 145727 91202 163449
rect 90902 145609 90993 145727
rect 91111 145609 91202 145727
rect 90902 145567 91202 145609
rect 90902 145449 90993 145567
rect 91111 145449 91202 145567
rect 90902 127727 91202 145449
rect 90902 127609 90993 127727
rect 91111 127609 91202 127727
rect 90902 127567 91202 127609
rect 90902 127449 90993 127567
rect 91111 127449 91202 127567
rect 90902 109727 91202 127449
rect 90902 109609 90993 109727
rect 91111 109609 91202 109727
rect 90902 109567 91202 109609
rect 90902 109449 90993 109567
rect 91111 109449 91202 109567
rect 90902 91727 91202 109449
rect 90902 91609 90993 91727
rect 91111 91609 91202 91727
rect 90902 91567 91202 91609
rect 90902 91449 90993 91567
rect 91111 91449 91202 91567
rect 90902 73727 91202 91449
rect 90902 73609 90993 73727
rect 91111 73609 91202 73727
rect 90902 73567 91202 73609
rect 90902 73449 90993 73567
rect 91111 73449 91202 73567
rect 90902 55727 91202 73449
rect 90902 55609 90993 55727
rect 91111 55609 91202 55727
rect 90902 55567 91202 55609
rect 90902 55449 90993 55567
rect 91111 55449 91202 55567
rect 90902 37727 91202 55449
rect 90902 37609 90993 37727
rect 91111 37609 91202 37727
rect 90902 37567 91202 37609
rect 90902 37449 90993 37567
rect 91111 37449 91202 37567
rect 90902 19727 91202 37449
rect 90902 19609 90993 19727
rect 91111 19609 91202 19727
rect 90902 19567 91202 19609
rect 90902 19449 90993 19567
rect 91111 19449 91202 19567
rect 90902 1727 91202 19449
rect 90902 1609 90993 1727
rect 91111 1609 91202 1727
rect 90902 1567 91202 1609
rect 90902 1449 90993 1567
rect 91111 1449 91202 1567
rect 90902 -173 91202 1449
rect 90902 -291 90993 -173
rect 91111 -291 91202 -173
rect 90902 -333 91202 -291
rect 90902 -451 90993 -333
rect 91111 -451 91202 -333
rect 90902 -932 91202 -451
rect 92702 345527 93002 353081
rect 92702 345409 92793 345527
rect 92911 345409 93002 345527
rect 92702 345367 93002 345409
rect 92702 345249 92793 345367
rect 92911 345249 93002 345367
rect 92702 327527 93002 345249
rect 92702 327409 92793 327527
rect 92911 327409 93002 327527
rect 92702 327367 93002 327409
rect 92702 327249 92793 327367
rect 92911 327249 93002 327367
rect 92702 309527 93002 327249
rect 92702 309409 92793 309527
rect 92911 309409 93002 309527
rect 92702 309367 93002 309409
rect 92702 309249 92793 309367
rect 92911 309249 93002 309367
rect 92702 291527 93002 309249
rect 92702 291409 92793 291527
rect 92911 291409 93002 291527
rect 92702 291367 93002 291409
rect 92702 291249 92793 291367
rect 92911 291249 93002 291367
rect 92702 273527 93002 291249
rect 92702 273409 92793 273527
rect 92911 273409 93002 273527
rect 92702 273367 93002 273409
rect 92702 273249 92793 273367
rect 92911 273249 93002 273367
rect 92702 255527 93002 273249
rect 92702 255409 92793 255527
rect 92911 255409 93002 255527
rect 92702 255367 93002 255409
rect 92702 255249 92793 255367
rect 92911 255249 93002 255367
rect 92702 237527 93002 255249
rect 92702 237409 92793 237527
rect 92911 237409 93002 237527
rect 92702 237367 93002 237409
rect 92702 237249 92793 237367
rect 92911 237249 93002 237367
rect 92702 219527 93002 237249
rect 92702 219409 92793 219527
rect 92911 219409 93002 219527
rect 92702 219367 93002 219409
rect 92702 219249 92793 219367
rect 92911 219249 93002 219367
rect 92702 201527 93002 219249
rect 92702 201409 92793 201527
rect 92911 201409 93002 201527
rect 92702 201367 93002 201409
rect 92702 201249 92793 201367
rect 92911 201249 93002 201367
rect 92702 183527 93002 201249
rect 92702 183409 92793 183527
rect 92911 183409 93002 183527
rect 92702 183367 93002 183409
rect 92702 183249 92793 183367
rect 92911 183249 93002 183367
rect 92702 165527 93002 183249
rect 92702 165409 92793 165527
rect 92911 165409 93002 165527
rect 92702 165367 93002 165409
rect 92702 165249 92793 165367
rect 92911 165249 93002 165367
rect 92702 147527 93002 165249
rect 92702 147409 92793 147527
rect 92911 147409 93002 147527
rect 92702 147367 93002 147409
rect 92702 147249 92793 147367
rect 92911 147249 93002 147367
rect 92702 129527 93002 147249
rect 92702 129409 92793 129527
rect 92911 129409 93002 129527
rect 92702 129367 93002 129409
rect 92702 129249 92793 129367
rect 92911 129249 93002 129367
rect 92702 111527 93002 129249
rect 92702 111409 92793 111527
rect 92911 111409 93002 111527
rect 92702 111367 93002 111409
rect 92702 111249 92793 111367
rect 92911 111249 93002 111367
rect 92702 93527 93002 111249
rect 92702 93409 92793 93527
rect 92911 93409 93002 93527
rect 92702 93367 93002 93409
rect 92702 93249 92793 93367
rect 92911 93249 93002 93367
rect 92702 75527 93002 93249
rect 92702 75409 92793 75527
rect 92911 75409 93002 75527
rect 92702 75367 93002 75409
rect 92702 75249 92793 75367
rect 92911 75249 93002 75367
rect 92702 57527 93002 75249
rect 92702 57409 92793 57527
rect 92911 57409 93002 57527
rect 92702 57367 93002 57409
rect 92702 57249 92793 57367
rect 92911 57249 93002 57367
rect 92702 39527 93002 57249
rect 92702 39409 92793 39527
rect 92911 39409 93002 39527
rect 92702 39367 93002 39409
rect 92702 39249 92793 39367
rect 92911 39249 93002 39367
rect 92702 21527 93002 39249
rect 92702 21409 92793 21527
rect 92911 21409 93002 21527
rect 92702 21367 93002 21409
rect 92702 21249 92793 21367
rect 92911 21249 93002 21367
rect 92702 3527 93002 21249
rect 92702 3409 92793 3527
rect 92911 3409 93002 3527
rect 92702 3367 93002 3409
rect 92702 3249 92793 3367
rect 92911 3249 93002 3367
rect 92702 -1113 93002 3249
rect 92702 -1231 92793 -1113
rect 92911 -1231 93002 -1113
rect 92702 -1273 93002 -1231
rect 92702 -1391 92793 -1273
rect 92911 -1391 93002 -1273
rect 92702 -1872 93002 -1391
rect 94502 347327 94802 354021
rect 94502 347209 94593 347327
rect 94711 347209 94802 347327
rect 94502 347167 94802 347209
rect 94502 347049 94593 347167
rect 94711 347049 94802 347167
rect 94502 329327 94802 347049
rect 94502 329209 94593 329327
rect 94711 329209 94802 329327
rect 94502 329167 94802 329209
rect 94502 329049 94593 329167
rect 94711 329049 94802 329167
rect 94502 311327 94802 329049
rect 94502 311209 94593 311327
rect 94711 311209 94802 311327
rect 94502 311167 94802 311209
rect 94502 311049 94593 311167
rect 94711 311049 94802 311167
rect 94502 293327 94802 311049
rect 94502 293209 94593 293327
rect 94711 293209 94802 293327
rect 94502 293167 94802 293209
rect 94502 293049 94593 293167
rect 94711 293049 94802 293167
rect 94502 275327 94802 293049
rect 94502 275209 94593 275327
rect 94711 275209 94802 275327
rect 94502 275167 94802 275209
rect 94502 275049 94593 275167
rect 94711 275049 94802 275167
rect 94502 257327 94802 275049
rect 94502 257209 94593 257327
rect 94711 257209 94802 257327
rect 94502 257167 94802 257209
rect 94502 257049 94593 257167
rect 94711 257049 94802 257167
rect 94502 239327 94802 257049
rect 94502 239209 94593 239327
rect 94711 239209 94802 239327
rect 94502 239167 94802 239209
rect 94502 239049 94593 239167
rect 94711 239049 94802 239167
rect 94502 221327 94802 239049
rect 94502 221209 94593 221327
rect 94711 221209 94802 221327
rect 94502 221167 94802 221209
rect 94502 221049 94593 221167
rect 94711 221049 94802 221167
rect 94502 203327 94802 221049
rect 94502 203209 94593 203327
rect 94711 203209 94802 203327
rect 94502 203167 94802 203209
rect 94502 203049 94593 203167
rect 94711 203049 94802 203167
rect 94502 185327 94802 203049
rect 94502 185209 94593 185327
rect 94711 185209 94802 185327
rect 94502 185167 94802 185209
rect 94502 185049 94593 185167
rect 94711 185049 94802 185167
rect 94502 167327 94802 185049
rect 94502 167209 94593 167327
rect 94711 167209 94802 167327
rect 94502 167167 94802 167209
rect 94502 167049 94593 167167
rect 94711 167049 94802 167167
rect 94502 149327 94802 167049
rect 94502 149209 94593 149327
rect 94711 149209 94802 149327
rect 94502 149167 94802 149209
rect 94502 149049 94593 149167
rect 94711 149049 94802 149167
rect 94502 131327 94802 149049
rect 94502 131209 94593 131327
rect 94711 131209 94802 131327
rect 94502 131167 94802 131209
rect 94502 131049 94593 131167
rect 94711 131049 94802 131167
rect 94502 113327 94802 131049
rect 94502 113209 94593 113327
rect 94711 113209 94802 113327
rect 94502 113167 94802 113209
rect 94502 113049 94593 113167
rect 94711 113049 94802 113167
rect 94502 95327 94802 113049
rect 94502 95209 94593 95327
rect 94711 95209 94802 95327
rect 94502 95167 94802 95209
rect 94502 95049 94593 95167
rect 94711 95049 94802 95167
rect 94502 77327 94802 95049
rect 94502 77209 94593 77327
rect 94711 77209 94802 77327
rect 94502 77167 94802 77209
rect 94502 77049 94593 77167
rect 94711 77049 94802 77167
rect 94502 59327 94802 77049
rect 94502 59209 94593 59327
rect 94711 59209 94802 59327
rect 94502 59167 94802 59209
rect 94502 59049 94593 59167
rect 94711 59049 94802 59167
rect 94502 41327 94802 59049
rect 94502 41209 94593 41327
rect 94711 41209 94802 41327
rect 94502 41167 94802 41209
rect 94502 41049 94593 41167
rect 94711 41049 94802 41167
rect 94502 23327 94802 41049
rect 94502 23209 94593 23327
rect 94711 23209 94802 23327
rect 94502 23167 94802 23209
rect 94502 23049 94593 23167
rect 94711 23049 94802 23167
rect 94502 5327 94802 23049
rect 94502 5209 94593 5327
rect 94711 5209 94802 5327
rect 94502 5167 94802 5209
rect 94502 5049 94593 5167
rect 94711 5049 94802 5167
rect 94502 -2053 94802 5049
rect 94502 -2171 94593 -2053
rect 94711 -2171 94802 -2053
rect 94502 -2213 94802 -2171
rect 94502 -2331 94593 -2213
rect 94711 -2331 94802 -2213
rect 94502 -2812 94802 -2331
rect 96302 349127 96602 354961
rect 105302 355709 105602 355720
rect 105302 355591 105393 355709
rect 105511 355591 105602 355709
rect 105302 355549 105602 355591
rect 105302 355431 105393 355549
rect 105511 355431 105602 355549
rect 103502 354769 103802 354780
rect 103502 354651 103593 354769
rect 103711 354651 103802 354769
rect 103502 354609 103802 354651
rect 103502 354491 103593 354609
rect 103711 354491 103802 354609
rect 101702 353829 102002 353840
rect 101702 353711 101793 353829
rect 101911 353711 102002 353829
rect 101702 353669 102002 353711
rect 101702 353551 101793 353669
rect 101911 353551 102002 353669
rect 96302 349009 96393 349127
rect 96511 349009 96602 349127
rect 96302 348967 96602 349009
rect 96302 348849 96393 348967
rect 96511 348849 96602 348967
rect 96302 331127 96602 348849
rect 96302 331009 96393 331127
rect 96511 331009 96602 331127
rect 96302 330967 96602 331009
rect 96302 330849 96393 330967
rect 96511 330849 96602 330967
rect 96302 313127 96602 330849
rect 96302 313009 96393 313127
rect 96511 313009 96602 313127
rect 96302 312967 96602 313009
rect 96302 312849 96393 312967
rect 96511 312849 96602 312967
rect 96302 295127 96602 312849
rect 96302 295009 96393 295127
rect 96511 295009 96602 295127
rect 96302 294967 96602 295009
rect 96302 294849 96393 294967
rect 96511 294849 96602 294967
rect 96302 277127 96602 294849
rect 96302 277009 96393 277127
rect 96511 277009 96602 277127
rect 96302 276967 96602 277009
rect 96302 276849 96393 276967
rect 96511 276849 96602 276967
rect 96302 259127 96602 276849
rect 96302 259009 96393 259127
rect 96511 259009 96602 259127
rect 96302 258967 96602 259009
rect 96302 258849 96393 258967
rect 96511 258849 96602 258967
rect 96302 241127 96602 258849
rect 96302 241009 96393 241127
rect 96511 241009 96602 241127
rect 96302 240967 96602 241009
rect 96302 240849 96393 240967
rect 96511 240849 96602 240967
rect 96302 223127 96602 240849
rect 96302 223009 96393 223127
rect 96511 223009 96602 223127
rect 96302 222967 96602 223009
rect 96302 222849 96393 222967
rect 96511 222849 96602 222967
rect 96302 205127 96602 222849
rect 96302 205009 96393 205127
rect 96511 205009 96602 205127
rect 96302 204967 96602 205009
rect 96302 204849 96393 204967
rect 96511 204849 96602 204967
rect 96302 187127 96602 204849
rect 96302 187009 96393 187127
rect 96511 187009 96602 187127
rect 96302 186967 96602 187009
rect 96302 186849 96393 186967
rect 96511 186849 96602 186967
rect 96302 169127 96602 186849
rect 96302 169009 96393 169127
rect 96511 169009 96602 169127
rect 96302 168967 96602 169009
rect 96302 168849 96393 168967
rect 96511 168849 96602 168967
rect 96302 151127 96602 168849
rect 96302 151009 96393 151127
rect 96511 151009 96602 151127
rect 96302 150967 96602 151009
rect 96302 150849 96393 150967
rect 96511 150849 96602 150967
rect 96302 133127 96602 150849
rect 96302 133009 96393 133127
rect 96511 133009 96602 133127
rect 96302 132967 96602 133009
rect 96302 132849 96393 132967
rect 96511 132849 96602 132967
rect 96302 115127 96602 132849
rect 96302 115009 96393 115127
rect 96511 115009 96602 115127
rect 96302 114967 96602 115009
rect 96302 114849 96393 114967
rect 96511 114849 96602 114967
rect 96302 97127 96602 114849
rect 96302 97009 96393 97127
rect 96511 97009 96602 97127
rect 96302 96967 96602 97009
rect 96302 96849 96393 96967
rect 96511 96849 96602 96967
rect 96302 79127 96602 96849
rect 96302 79009 96393 79127
rect 96511 79009 96602 79127
rect 96302 78967 96602 79009
rect 96302 78849 96393 78967
rect 96511 78849 96602 78967
rect 96302 61127 96602 78849
rect 96302 61009 96393 61127
rect 96511 61009 96602 61127
rect 96302 60967 96602 61009
rect 96302 60849 96393 60967
rect 96511 60849 96602 60967
rect 96302 43127 96602 60849
rect 96302 43009 96393 43127
rect 96511 43009 96602 43127
rect 96302 42967 96602 43009
rect 96302 42849 96393 42967
rect 96511 42849 96602 42967
rect 96302 25127 96602 42849
rect 96302 25009 96393 25127
rect 96511 25009 96602 25127
rect 96302 24967 96602 25009
rect 96302 24849 96393 24967
rect 96511 24849 96602 24967
rect 96302 7127 96602 24849
rect 96302 7009 96393 7127
rect 96511 7009 96602 7127
rect 96302 6967 96602 7009
rect 96302 6849 96393 6967
rect 96511 6849 96602 6967
rect 87302 -3581 87393 -3463
rect 87511 -3581 87602 -3463
rect 87302 -3623 87602 -3581
rect 87302 -3741 87393 -3623
rect 87511 -3741 87602 -3623
rect 87302 -3752 87602 -3741
rect 96302 -2993 96602 6849
rect 99902 352889 100202 352900
rect 99902 352771 99993 352889
rect 100111 352771 100202 352889
rect 99902 352729 100202 352771
rect 99902 352611 99993 352729
rect 100111 352611 100202 352729
rect 99902 334727 100202 352611
rect 99902 334609 99993 334727
rect 100111 334609 100202 334727
rect 99902 334567 100202 334609
rect 99902 334449 99993 334567
rect 100111 334449 100202 334567
rect 99902 316727 100202 334449
rect 99902 316609 99993 316727
rect 100111 316609 100202 316727
rect 99902 316567 100202 316609
rect 99902 316449 99993 316567
rect 100111 316449 100202 316567
rect 99902 298727 100202 316449
rect 99902 298609 99993 298727
rect 100111 298609 100202 298727
rect 99902 298567 100202 298609
rect 99902 298449 99993 298567
rect 100111 298449 100202 298567
rect 99902 280727 100202 298449
rect 99902 280609 99993 280727
rect 100111 280609 100202 280727
rect 99902 280567 100202 280609
rect 99902 280449 99993 280567
rect 100111 280449 100202 280567
rect 99902 262727 100202 280449
rect 99902 262609 99993 262727
rect 100111 262609 100202 262727
rect 99902 262567 100202 262609
rect 99902 262449 99993 262567
rect 100111 262449 100202 262567
rect 99902 244727 100202 262449
rect 99902 244609 99993 244727
rect 100111 244609 100202 244727
rect 99902 244567 100202 244609
rect 99902 244449 99993 244567
rect 100111 244449 100202 244567
rect 99902 226727 100202 244449
rect 99902 226609 99993 226727
rect 100111 226609 100202 226727
rect 99902 226567 100202 226609
rect 99902 226449 99993 226567
rect 100111 226449 100202 226567
rect 99902 208727 100202 226449
rect 99902 208609 99993 208727
rect 100111 208609 100202 208727
rect 99902 208567 100202 208609
rect 99902 208449 99993 208567
rect 100111 208449 100202 208567
rect 99902 190727 100202 208449
rect 99902 190609 99993 190727
rect 100111 190609 100202 190727
rect 99902 190567 100202 190609
rect 99902 190449 99993 190567
rect 100111 190449 100202 190567
rect 99902 172727 100202 190449
rect 99902 172609 99993 172727
rect 100111 172609 100202 172727
rect 99902 172567 100202 172609
rect 99902 172449 99993 172567
rect 100111 172449 100202 172567
rect 99902 154727 100202 172449
rect 99902 154609 99993 154727
rect 100111 154609 100202 154727
rect 99902 154567 100202 154609
rect 99902 154449 99993 154567
rect 100111 154449 100202 154567
rect 99902 136727 100202 154449
rect 99902 136609 99993 136727
rect 100111 136609 100202 136727
rect 99902 136567 100202 136609
rect 99902 136449 99993 136567
rect 100111 136449 100202 136567
rect 99902 118727 100202 136449
rect 99902 118609 99993 118727
rect 100111 118609 100202 118727
rect 99902 118567 100202 118609
rect 99902 118449 99993 118567
rect 100111 118449 100202 118567
rect 99902 100727 100202 118449
rect 99902 100609 99993 100727
rect 100111 100609 100202 100727
rect 99902 100567 100202 100609
rect 99902 100449 99993 100567
rect 100111 100449 100202 100567
rect 99902 82727 100202 100449
rect 99902 82609 99993 82727
rect 100111 82609 100202 82727
rect 99902 82567 100202 82609
rect 99902 82449 99993 82567
rect 100111 82449 100202 82567
rect 99902 64727 100202 82449
rect 99902 64609 99993 64727
rect 100111 64609 100202 64727
rect 99902 64567 100202 64609
rect 99902 64449 99993 64567
rect 100111 64449 100202 64567
rect 99902 46727 100202 64449
rect 99902 46609 99993 46727
rect 100111 46609 100202 46727
rect 99902 46567 100202 46609
rect 99902 46449 99993 46567
rect 100111 46449 100202 46567
rect 99902 28727 100202 46449
rect 99902 28609 99993 28727
rect 100111 28609 100202 28727
rect 99902 28567 100202 28609
rect 99902 28449 99993 28567
rect 100111 28449 100202 28567
rect 99902 10727 100202 28449
rect 99902 10609 99993 10727
rect 100111 10609 100202 10727
rect 99902 10567 100202 10609
rect 99902 10449 99993 10567
rect 100111 10449 100202 10567
rect 99902 -643 100202 10449
rect 99902 -761 99993 -643
rect 100111 -761 100202 -643
rect 99902 -803 100202 -761
rect 99902 -921 99993 -803
rect 100111 -921 100202 -803
rect 99902 -932 100202 -921
rect 101702 336527 102002 353551
rect 101702 336409 101793 336527
rect 101911 336409 102002 336527
rect 101702 336367 102002 336409
rect 101702 336249 101793 336367
rect 101911 336249 102002 336367
rect 101702 318527 102002 336249
rect 101702 318409 101793 318527
rect 101911 318409 102002 318527
rect 101702 318367 102002 318409
rect 101702 318249 101793 318367
rect 101911 318249 102002 318367
rect 101702 300527 102002 318249
rect 101702 300409 101793 300527
rect 101911 300409 102002 300527
rect 101702 300367 102002 300409
rect 101702 300249 101793 300367
rect 101911 300249 102002 300367
rect 101702 282527 102002 300249
rect 101702 282409 101793 282527
rect 101911 282409 102002 282527
rect 101702 282367 102002 282409
rect 101702 282249 101793 282367
rect 101911 282249 102002 282367
rect 101702 264527 102002 282249
rect 101702 264409 101793 264527
rect 101911 264409 102002 264527
rect 101702 264367 102002 264409
rect 101702 264249 101793 264367
rect 101911 264249 102002 264367
rect 101702 246527 102002 264249
rect 101702 246409 101793 246527
rect 101911 246409 102002 246527
rect 101702 246367 102002 246409
rect 101702 246249 101793 246367
rect 101911 246249 102002 246367
rect 101702 228527 102002 246249
rect 101702 228409 101793 228527
rect 101911 228409 102002 228527
rect 101702 228367 102002 228409
rect 101702 228249 101793 228367
rect 101911 228249 102002 228367
rect 101702 210527 102002 228249
rect 101702 210409 101793 210527
rect 101911 210409 102002 210527
rect 101702 210367 102002 210409
rect 101702 210249 101793 210367
rect 101911 210249 102002 210367
rect 101702 192527 102002 210249
rect 101702 192409 101793 192527
rect 101911 192409 102002 192527
rect 101702 192367 102002 192409
rect 101702 192249 101793 192367
rect 101911 192249 102002 192367
rect 101702 174527 102002 192249
rect 101702 174409 101793 174527
rect 101911 174409 102002 174527
rect 101702 174367 102002 174409
rect 101702 174249 101793 174367
rect 101911 174249 102002 174367
rect 101702 156527 102002 174249
rect 101702 156409 101793 156527
rect 101911 156409 102002 156527
rect 101702 156367 102002 156409
rect 101702 156249 101793 156367
rect 101911 156249 102002 156367
rect 101702 138527 102002 156249
rect 101702 138409 101793 138527
rect 101911 138409 102002 138527
rect 101702 138367 102002 138409
rect 101702 138249 101793 138367
rect 101911 138249 102002 138367
rect 101702 120527 102002 138249
rect 101702 120409 101793 120527
rect 101911 120409 102002 120527
rect 101702 120367 102002 120409
rect 101702 120249 101793 120367
rect 101911 120249 102002 120367
rect 101702 102527 102002 120249
rect 101702 102409 101793 102527
rect 101911 102409 102002 102527
rect 101702 102367 102002 102409
rect 101702 102249 101793 102367
rect 101911 102249 102002 102367
rect 101702 84527 102002 102249
rect 101702 84409 101793 84527
rect 101911 84409 102002 84527
rect 101702 84367 102002 84409
rect 101702 84249 101793 84367
rect 101911 84249 102002 84367
rect 101702 66527 102002 84249
rect 101702 66409 101793 66527
rect 101911 66409 102002 66527
rect 101702 66367 102002 66409
rect 101702 66249 101793 66367
rect 101911 66249 102002 66367
rect 101702 48527 102002 66249
rect 101702 48409 101793 48527
rect 101911 48409 102002 48527
rect 101702 48367 102002 48409
rect 101702 48249 101793 48367
rect 101911 48249 102002 48367
rect 101702 30527 102002 48249
rect 101702 30409 101793 30527
rect 101911 30409 102002 30527
rect 101702 30367 102002 30409
rect 101702 30249 101793 30367
rect 101911 30249 102002 30367
rect 101702 12527 102002 30249
rect 101702 12409 101793 12527
rect 101911 12409 102002 12527
rect 101702 12367 102002 12409
rect 101702 12249 101793 12367
rect 101911 12249 102002 12367
rect 101702 -1583 102002 12249
rect 101702 -1701 101793 -1583
rect 101911 -1701 102002 -1583
rect 101702 -1743 102002 -1701
rect 101702 -1861 101793 -1743
rect 101911 -1861 102002 -1743
rect 101702 -1872 102002 -1861
rect 103502 338327 103802 354491
rect 103502 338209 103593 338327
rect 103711 338209 103802 338327
rect 103502 338167 103802 338209
rect 103502 338049 103593 338167
rect 103711 338049 103802 338167
rect 103502 320327 103802 338049
rect 103502 320209 103593 320327
rect 103711 320209 103802 320327
rect 103502 320167 103802 320209
rect 103502 320049 103593 320167
rect 103711 320049 103802 320167
rect 103502 302327 103802 320049
rect 103502 302209 103593 302327
rect 103711 302209 103802 302327
rect 103502 302167 103802 302209
rect 103502 302049 103593 302167
rect 103711 302049 103802 302167
rect 103502 284327 103802 302049
rect 103502 284209 103593 284327
rect 103711 284209 103802 284327
rect 103502 284167 103802 284209
rect 103502 284049 103593 284167
rect 103711 284049 103802 284167
rect 103502 266327 103802 284049
rect 103502 266209 103593 266327
rect 103711 266209 103802 266327
rect 103502 266167 103802 266209
rect 103502 266049 103593 266167
rect 103711 266049 103802 266167
rect 103502 248327 103802 266049
rect 103502 248209 103593 248327
rect 103711 248209 103802 248327
rect 103502 248167 103802 248209
rect 103502 248049 103593 248167
rect 103711 248049 103802 248167
rect 103502 230327 103802 248049
rect 103502 230209 103593 230327
rect 103711 230209 103802 230327
rect 103502 230167 103802 230209
rect 103502 230049 103593 230167
rect 103711 230049 103802 230167
rect 103502 212327 103802 230049
rect 103502 212209 103593 212327
rect 103711 212209 103802 212327
rect 103502 212167 103802 212209
rect 103502 212049 103593 212167
rect 103711 212049 103802 212167
rect 103502 194327 103802 212049
rect 103502 194209 103593 194327
rect 103711 194209 103802 194327
rect 103502 194167 103802 194209
rect 103502 194049 103593 194167
rect 103711 194049 103802 194167
rect 103502 176327 103802 194049
rect 103502 176209 103593 176327
rect 103711 176209 103802 176327
rect 103502 176167 103802 176209
rect 103502 176049 103593 176167
rect 103711 176049 103802 176167
rect 103502 158327 103802 176049
rect 103502 158209 103593 158327
rect 103711 158209 103802 158327
rect 103502 158167 103802 158209
rect 103502 158049 103593 158167
rect 103711 158049 103802 158167
rect 103502 140327 103802 158049
rect 103502 140209 103593 140327
rect 103711 140209 103802 140327
rect 103502 140167 103802 140209
rect 103502 140049 103593 140167
rect 103711 140049 103802 140167
rect 103502 122327 103802 140049
rect 103502 122209 103593 122327
rect 103711 122209 103802 122327
rect 103502 122167 103802 122209
rect 103502 122049 103593 122167
rect 103711 122049 103802 122167
rect 103502 104327 103802 122049
rect 103502 104209 103593 104327
rect 103711 104209 103802 104327
rect 103502 104167 103802 104209
rect 103502 104049 103593 104167
rect 103711 104049 103802 104167
rect 103502 86327 103802 104049
rect 103502 86209 103593 86327
rect 103711 86209 103802 86327
rect 103502 86167 103802 86209
rect 103502 86049 103593 86167
rect 103711 86049 103802 86167
rect 103502 68327 103802 86049
rect 103502 68209 103593 68327
rect 103711 68209 103802 68327
rect 103502 68167 103802 68209
rect 103502 68049 103593 68167
rect 103711 68049 103802 68167
rect 103502 50327 103802 68049
rect 103502 50209 103593 50327
rect 103711 50209 103802 50327
rect 103502 50167 103802 50209
rect 103502 50049 103593 50167
rect 103711 50049 103802 50167
rect 103502 32327 103802 50049
rect 103502 32209 103593 32327
rect 103711 32209 103802 32327
rect 103502 32167 103802 32209
rect 103502 32049 103593 32167
rect 103711 32049 103802 32167
rect 103502 14327 103802 32049
rect 103502 14209 103593 14327
rect 103711 14209 103802 14327
rect 103502 14167 103802 14209
rect 103502 14049 103593 14167
rect 103711 14049 103802 14167
rect 103502 -2523 103802 14049
rect 103502 -2641 103593 -2523
rect 103711 -2641 103802 -2523
rect 103502 -2683 103802 -2641
rect 103502 -2801 103593 -2683
rect 103711 -2801 103802 -2683
rect 103502 -2812 103802 -2801
rect 105302 340127 105602 355431
rect 114302 355239 114602 355720
rect 114302 355121 114393 355239
rect 114511 355121 114602 355239
rect 114302 355079 114602 355121
rect 114302 354961 114393 355079
rect 114511 354961 114602 355079
rect 112502 354299 112802 354780
rect 112502 354181 112593 354299
rect 112711 354181 112802 354299
rect 112502 354139 112802 354181
rect 112502 354021 112593 354139
rect 112711 354021 112802 354139
rect 110702 353359 111002 353840
rect 110702 353241 110793 353359
rect 110911 353241 111002 353359
rect 110702 353199 111002 353241
rect 110702 353081 110793 353199
rect 110911 353081 111002 353199
rect 105302 340009 105393 340127
rect 105511 340009 105602 340127
rect 105302 339967 105602 340009
rect 105302 339849 105393 339967
rect 105511 339849 105602 339967
rect 105302 322127 105602 339849
rect 105302 322009 105393 322127
rect 105511 322009 105602 322127
rect 105302 321967 105602 322009
rect 105302 321849 105393 321967
rect 105511 321849 105602 321967
rect 105302 304127 105602 321849
rect 105302 304009 105393 304127
rect 105511 304009 105602 304127
rect 105302 303967 105602 304009
rect 105302 303849 105393 303967
rect 105511 303849 105602 303967
rect 105302 286127 105602 303849
rect 105302 286009 105393 286127
rect 105511 286009 105602 286127
rect 105302 285967 105602 286009
rect 105302 285849 105393 285967
rect 105511 285849 105602 285967
rect 105302 268127 105602 285849
rect 105302 268009 105393 268127
rect 105511 268009 105602 268127
rect 105302 267967 105602 268009
rect 105302 267849 105393 267967
rect 105511 267849 105602 267967
rect 105302 250127 105602 267849
rect 105302 250009 105393 250127
rect 105511 250009 105602 250127
rect 105302 249967 105602 250009
rect 105302 249849 105393 249967
rect 105511 249849 105602 249967
rect 105302 232127 105602 249849
rect 105302 232009 105393 232127
rect 105511 232009 105602 232127
rect 105302 231967 105602 232009
rect 105302 231849 105393 231967
rect 105511 231849 105602 231967
rect 105302 214127 105602 231849
rect 105302 214009 105393 214127
rect 105511 214009 105602 214127
rect 105302 213967 105602 214009
rect 105302 213849 105393 213967
rect 105511 213849 105602 213967
rect 105302 196127 105602 213849
rect 105302 196009 105393 196127
rect 105511 196009 105602 196127
rect 105302 195967 105602 196009
rect 105302 195849 105393 195967
rect 105511 195849 105602 195967
rect 105302 178127 105602 195849
rect 105302 178009 105393 178127
rect 105511 178009 105602 178127
rect 105302 177967 105602 178009
rect 105302 177849 105393 177967
rect 105511 177849 105602 177967
rect 105302 160127 105602 177849
rect 105302 160009 105393 160127
rect 105511 160009 105602 160127
rect 105302 159967 105602 160009
rect 105302 159849 105393 159967
rect 105511 159849 105602 159967
rect 105302 142127 105602 159849
rect 105302 142009 105393 142127
rect 105511 142009 105602 142127
rect 105302 141967 105602 142009
rect 105302 141849 105393 141967
rect 105511 141849 105602 141967
rect 105302 124127 105602 141849
rect 105302 124009 105393 124127
rect 105511 124009 105602 124127
rect 105302 123967 105602 124009
rect 105302 123849 105393 123967
rect 105511 123849 105602 123967
rect 105302 106127 105602 123849
rect 105302 106009 105393 106127
rect 105511 106009 105602 106127
rect 105302 105967 105602 106009
rect 105302 105849 105393 105967
rect 105511 105849 105602 105967
rect 105302 88127 105602 105849
rect 105302 88009 105393 88127
rect 105511 88009 105602 88127
rect 105302 87967 105602 88009
rect 105302 87849 105393 87967
rect 105511 87849 105602 87967
rect 105302 70127 105602 87849
rect 105302 70009 105393 70127
rect 105511 70009 105602 70127
rect 105302 69967 105602 70009
rect 105302 69849 105393 69967
rect 105511 69849 105602 69967
rect 105302 52127 105602 69849
rect 105302 52009 105393 52127
rect 105511 52009 105602 52127
rect 105302 51967 105602 52009
rect 105302 51849 105393 51967
rect 105511 51849 105602 51967
rect 105302 34127 105602 51849
rect 105302 34009 105393 34127
rect 105511 34009 105602 34127
rect 105302 33967 105602 34009
rect 105302 33849 105393 33967
rect 105511 33849 105602 33967
rect 105302 16127 105602 33849
rect 105302 16009 105393 16127
rect 105511 16009 105602 16127
rect 105302 15967 105602 16009
rect 105302 15849 105393 15967
rect 105511 15849 105602 15967
rect 96302 -3111 96393 -2993
rect 96511 -3111 96602 -2993
rect 96302 -3153 96602 -3111
rect 96302 -3271 96393 -3153
rect 96511 -3271 96602 -3153
rect 96302 -3752 96602 -3271
rect 105302 -3463 105602 15849
rect 108902 352419 109202 352900
rect 108902 352301 108993 352419
rect 109111 352301 109202 352419
rect 108902 352259 109202 352301
rect 108902 352141 108993 352259
rect 109111 352141 109202 352259
rect 108902 343727 109202 352141
rect 108902 343609 108993 343727
rect 109111 343609 109202 343727
rect 108902 343567 109202 343609
rect 108902 343449 108993 343567
rect 109111 343449 109202 343567
rect 108902 325727 109202 343449
rect 108902 325609 108993 325727
rect 109111 325609 109202 325727
rect 108902 325567 109202 325609
rect 108902 325449 108993 325567
rect 109111 325449 109202 325567
rect 108902 307727 109202 325449
rect 108902 307609 108993 307727
rect 109111 307609 109202 307727
rect 108902 307567 109202 307609
rect 108902 307449 108993 307567
rect 109111 307449 109202 307567
rect 108902 289727 109202 307449
rect 108902 289609 108993 289727
rect 109111 289609 109202 289727
rect 108902 289567 109202 289609
rect 108902 289449 108993 289567
rect 109111 289449 109202 289567
rect 108902 271727 109202 289449
rect 108902 271609 108993 271727
rect 109111 271609 109202 271727
rect 108902 271567 109202 271609
rect 108902 271449 108993 271567
rect 109111 271449 109202 271567
rect 108902 253727 109202 271449
rect 108902 253609 108993 253727
rect 109111 253609 109202 253727
rect 108902 253567 109202 253609
rect 108902 253449 108993 253567
rect 109111 253449 109202 253567
rect 108902 235727 109202 253449
rect 108902 235609 108993 235727
rect 109111 235609 109202 235727
rect 108902 235567 109202 235609
rect 108902 235449 108993 235567
rect 109111 235449 109202 235567
rect 108902 217727 109202 235449
rect 108902 217609 108993 217727
rect 109111 217609 109202 217727
rect 108902 217567 109202 217609
rect 108902 217449 108993 217567
rect 109111 217449 109202 217567
rect 108902 199727 109202 217449
rect 108902 199609 108993 199727
rect 109111 199609 109202 199727
rect 108902 199567 109202 199609
rect 108902 199449 108993 199567
rect 109111 199449 109202 199567
rect 108902 181727 109202 199449
rect 108902 181609 108993 181727
rect 109111 181609 109202 181727
rect 108902 181567 109202 181609
rect 108902 181449 108993 181567
rect 109111 181449 109202 181567
rect 108902 163727 109202 181449
rect 108902 163609 108993 163727
rect 109111 163609 109202 163727
rect 108902 163567 109202 163609
rect 108902 163449 108993 163567
rect 109111 163449 109202 163567
rect 108902 145727 109202 163449
rect 108902 145609 108993 145727
rect 109111 145609 109202 145727
rect 108902 145567 109202 145609
rect 108902 145449 108993 145567
rect 109111 145449 109202 145567
rect 108902 127727 109202 145449
rect 108902 127609 108993 127727
rect 109111 127609 109202 127727
rect 108902 127567 109202 127609
rect 108902 127449 108993 127567
rect 109111 127449 109202 127567
rect 108902 109727 109202 127449
rect 108902 109609 108993 109727
rect 109111 109609 109202 109727
rect 108902 109567 109202 109609
rect 108902 109449 108993 109567
rect 109111 109449 109202 109567
rect 108902 91727 109202 109449
rect 108902 91609 108993 91727
rect 109111 91609 109202 91727
rect 108902 91567 109202 91609
rect 108902 91449 108993 91567
rect 109111 91449 109202 91567
rect 108902 73727 109202 91449
rect 108902 73609 108993 73727
rect 109111 73609 109202 73727
rect 108902 73567 109202 73609
rect 108902 73449 108993 73567
rect 109111 73449 109202 73567
rect 108902 55727 109202 73449
rect 108902 55609 108993 55727
rect 109111 55609 109202 55727
rect 108902 55567 109202 55609
rect 108902 55449 108993 55567
rect 109111 55449 109202 55567
rect 108902 37727 109202 55449
rect 108902 37609 108993 37727
rect 109111 37609 109202 37727
rect 108902 37567 109202 37609
rect 108902 37449 108993 37567
rect 109111 37449 109202 37567
rect 108902 19727 109202 37449
rect 108902 19609 108993 19727
rect 109111 19609 109202 19727
rect 108902 19567 109202 19609
rect 108902 19449 108993 19567
rect 109111 19449 109202 19567
rect 108902 1727 109202 19449
rect 108902 1609 108993 1727
rect 109111 1609 109202 1727
rect 108902 1567 109202 1609
rect 108902 1449 108993 1567
rect 109111 1449 109202 1567
rect 108902 -173 109202 1449
rect 108902 -291 108993 -173
rect 109111 -291 109202 -173
rect 108902 -333 109202 -291
rect 108902 -451 108993 -333
rect 109111 -451 109202 -333
rect 108902 -932 109202 -451
rect 110702 345527 111002 353081
rect 110702 345409 110793 345527
rect 110911 345409 111002 345527
rect 110702 345367 111002 345409
rect 110702 345249 110793 345367
rect 110911 345249 111002 345367
rect 110702 327527 111002 345249
rect 110702 327409 110793 327527
rect 110911 327409 111002 327527
rect 110702 327367 111002 327409
rect 110702 327249 110793 327367
rect 110911 327249 111002 327367
rect 110702 309527 111002 327249
rect 110702 309409 110793 309527
rect 110911 309409 111002 309527
rect 110702 309367 111002 309409
rect 110702 309249 110793 309367
rect 110911 309249 111002 309367
rect 110702 291527 111002 309249
rect 110702 291409 110793 291527
rect 110911 291409 111002 291527
rect 110702 291367 111002 291409
rect 110702 291249 110793 291367
rect 110911 291249 111002 291367
rect 110702 273527 111002 291249
rect 110702 273409 110793 273527
rect 110911 273409 111002 273527
rect 110702 273367 111002 273409
rect 110702 273249 110793 273367
rect 110911 273249 111002 273367
rect 110702 255527 111002 273249
rect 110702 255409 110793 255527
rect 110911 255409 111002 255527
rect 110702 255367 111002 255409
rect 110702 255249 110793 255367
rect 110911 255249 111002 255367
rect 110702 237527 111002 255249
rect 110702 237409 110793 237527
rect 110911 237409 111002 237527
rect 110702 237367 111002 237409
rect 110702 237249 110793 237367
rect 110911 237249 111002 237367
rect 110702 219527 111002 237249
rect 110702 219409 110793 219527
rect 110911 219409 111002 219527
rect 110702 219367 111002 219409
rect 110702 219249 110793 219367
rect 110911 219249 111002 219367
rect 110702 201527 111002 219249
rect 110702 201409 110793 201527
rect 110911 201409 111002 201527
rect 110702 201367 111002 201409
rect 110702 201249 110793 201367
rect 110911 201249 111002 201367
rect 110702 183527 111002 201249
rect 110702 183409 110793 183527
rect 110911 183409 111002 183527
rect 110702 183367 111002 183409
rect 110702 183249 110793 183367
rect 110911 183249 111002 183367
rect 110702 165527 111002 183249
rect 110702 165409 110793 165527
rect 110911 165409 111002 165527
rect 110702 165367 111002 165409
rect 110702 165249 110793 165367
rect 110911 165249 111002 165367
rect 110702 147527 111002 165249
rect 110702 147409 110793 147527
rect 110911 147409 111002 147527
rect 110702 147367 111002 147409
rect 110702 147249 110793 147367
rect 110911 147249 111002 147367
rect 110702 129527 111002 147249
rect 110702 129409 110793 129527
rect 110911 129409 111002 129527
rect 110702 129367 111002 129409
rect 110702 129249 110793 129367
rect 110911 129249 111002 129367
rect 110702 111527 111002 129249
rect 110702 111409 110793 111527
rect 110911 111409 111002 111527
rect 110702 111367 111002 111409
rect 110702 111249 110793 111367
rect 110911 111249 111002 111367
rect 110702 93527 111002 111249
rect 110702 93409 110793 93527
rect 110911 93409 111002 93527
rect 110702 93367 111002 93409
rect 110702 93249 110793 93367
rect 110911 93249 111002 93367
rect 110702 75527 111002 93249
rect 110702 75409 110793 75527
rect 110911 75409 111002 75527
rect 110702 75367 111002 75409
rect 110702 75249 110793 75367
rect 110911 75249 111002 75367
rect 110702 57527 111002 75249
rect 110702 57409 110793 57527
rect 110911 57409 111002 57527
rect 110702 57367 111002 57409
rect 110702 57249 110793 57367
rect 110911 57249 111002 57367
rect 110702 39527 111002 57249
rect 110702 39409 110793 39527
rect 110911 39409 111002 39527
rect 110702 39367 111002 39409
rect 110702 39249 110793 39367
rect 110911 39249 111002 39367
rect 110702 21527 111002 39249
rect 110702 21409 110793 21527
rect 110911 21409 111002 21527
rect 110702 21367 111002 21409
rect 110702 21249 110793 21367
rect 110911 21249 111002 21367
rect 110702 3527 111002 21249
rect 110702 3409 110793 3527
rect 110911 3409 111002 3527
rect 110702 3367 111002 3409
rect 110702 3249 110793 3367
rect 110911 3249 111002 3367
rect 110702 -1113 111002 3249
rect 110702 -1231 110793 -1113
rect 110911 -1231 111002 -1113
rect 110702 -1273 111002 -1231
rect 110702 -1391 110793 -1273
rect 110911 -1391 111002 -1273
rect 110702 -1872 111002 -1391
rect 112502 347327 112802 354021
rect 112502 347209 112593 347327
rect 112711 347209 112802 347327
rect 112502 347167 112802 347209
rect 112502 347049 112593 347167
rect 112711 347049 112802 347167
rect 112502 329327 112802 347049
rect 112502 329209 112593 329327
rect 112711 329209 112802 329327
rect 112502 329167 112802 329209
rect 112502 329049 112593 329167
rect 112711 329049 112802 329167
rect 112502 311327 112802 329049
rect 112502 311209 112593 311327
rect 112711 311209 112802 311327
rect 112502 311167 112802 311209
rect 112502 311049 112593 311167
rect 112711 311049 112802 311167
rect 112502 293327 112802 311049
rect 112502 293209 112593 293327
rect 112711 293209 112802 293327
rect 112502 293167 112802 293209
rect 112502 293049 112593 293167
rect 112711 293049 112802 293167
rect 112502 275327 112802 293049
rect 112502 275209 112593 275327
rect 112711 275209 112802 275327
rect 112502 275167 112802 275209
rect 112502 275049 112593 275167
rect 112711 275049 112802 275167
rect 112502 257327 112802 275049
rect 112502 257209 112593 257327
rect 112711 257209 112802 257327
rect 112502 257167 112802 257209
rect 112502 257049 112593 257167
rect 112711 257049 112802 257167
rect 112502 239327 112802 257049
rect 112502 239209 112593 239327
rect 112711 239209 112802 239327
rect 112502 239167 112802 239209
rect 112502 239049 112593 239167
rect 112711 239049 112802 239167
rect 112502 221327 112802 239049
rect 112502 221209 112593 221327
rect 112711 221209 112802 221327
rect 112502 221167 112802 221209
rect 112502 221049 112593 221167
rect 112711 221049 112802 221167
rect 112502 203327 112802 221049
rect 112502 203209 112593 203327
rect 112711 203209 112802 203327
rect 112502 203167 112802 203209
rect 112502 203049 112593 203167
rect 112711 203049 112802 203167
rect 112502 185327 112802 203049
rect 112502 185209 112593 185327
rect 112711 185209 112802 185327
rect 112502 185167 112802 185209
rect 112502 185049 112593 185167
rect 112711 185049 112802 185167
rect 112502 167327 112802 185049
rect 112502 167209 112593 167327
rect 112711 167209 112802 167327
rect 112502 167167 112802 167209
rect 112502 167049 112593 167167
rect 112711 167049 112802 167167
rect 112502 149327 112802 167049
rect 112502 149209 112593 149327
rect 112711 149209 112802 149327
rect 112502 149167 112802 149209
rect 112502 149049 112593 149167
rect 112711 149049 112802 149167
rect 112502 131327 112802 149049
rect 112502 131209 112593 131327
rect 112711 131209 112802 131327
rect 112502 131167 112802 131209
rect 112502 131049 112593 131167
rect 112711 131049 112802 131167
rect 112502 113327 112802 131049
rect 112502 113209 112593 113327
rect 112711 113209 112802 113327
rect 112502 113167 112802 113209
rect 112502 113049 112593 113167
rect 112711 113049 112802 113167
rect 112502 95327 112802 113049
rect 112502 95209 112593 95327
rect 112711 95209 112802 95327
rect 112502 95167 112802 95209
rect 112502 95049 112593 95167
rect 112711 95049 112802 95167
rect 112502 77327 112802 95049
rect 112502 77209 112593 77327
rect 112711 77209 112802 77327
rect 112502 77167 112802 77209
rect 112502 77049 112593 77167
rect 112711 77049 112802 77167
rect 112502 59327 112802 77049
rect 112502 59209 112593 59327
rect 112711 59209 112802 59327
rect 112502 59167 112802 59209
rect 112502 59049 112593 59167
rect 112711 59049 112802 59167
rect 112502 41327 112802 59049
rect 112502 41209 112593 41327
rect 112711 41209 112802 41327
rect 112502 41167 112802 41209
rect 112502 41049 112593 41167
rect 112711 41049 112802 41167
rect 112502 23327 112802 41049
rect 112502 23209 112593 23327
rect 112711 23209 112802 23327
rect 112502 23167 112802 23209
rect 112502 23049 112593 23167
rect 112711 23049 112802 23167
rect 112502 5327 112802 23049
rect 112502 5209 112593 5327
rect 112711 5209 112802 5327
rect 112502 5167 112802 5209
rect 112502 5049 112593 5167
rect 112711 5049 112802 5167
rect 112502 -2053 112802 5049
rect 112502 -2171 112593 -2053
rect 112711 -2171 112802 -2053
rect 112502 -2213 112802 -2171
rect 112502 -2331 112593 -2213
rect 112711 -2331 112802 -2213
rect 112502 -2812 112802 -2331
rect 114302 349127 114602 354961
rect 123302 355709 123602 355720
rect 123302 355591 123393 355709
rect 123511 355591 123602 355709
rect 123302 355549 123602 355591
rect 123302 355431 123393 355549
rect 123511 355431 123602 355549
rect 121502 354769 121802 354780
rect 121502 354651 121593 354769
rect 121711 354651 121802 354769
rect 121502 354609 121802 354651
rect 121502 354491 121593 354609
rect 121711 354491 121802 354609
rect 119702 353829 120002 353840
rect 119702 353711 119793 353829
rect 119911 353711 120002 353829
rect 119702 353669 120002 353711
rect 119702 353551 119793 353669
rect 119911 353551 120002 353669
rect 114302 349009 114393 349127
rect 114511 349009 114602 349127
rect 114302 348967 114602 349009
rect 114302 348849 114393 348967
rect 114511 348849 114602 348967
rect 114302 331127 114602 348849
rect 114302 331009 114393 331127
rect 114511 331009 114602 331127
rect 114302 330967 114602 331009
rect 114302 330849 114393 330967
rect 114511 330849 114602 330967
rect 114302 313127 114602 330849
rect 114302 313009 114393 313127
rect 114511 313009 114602 313127
rect 114302 312967 114602 313009
rect 114302 312849 114393 312967
rect 114511 312849 114602 312967
rect 114302 295127 114602 312849
rect 114302 295009 114393 295127
rect 114511 295009 114602 295127
rect 114302 294967 114602 295009
rect 114302 294849 114393 294967
rect 114511 294849 114602 294967
rect 114302 277127 114602 294849
rect 114302 277009 114393 277127
rect 114511 277009 114602 277127
rect 114302 276967 114602 277009
rect 114302 276849 114393 276967
rect 114511 276849 114602 276967
rect 114302 259127 114602 276849
rect 114302 259009 114393 259127
rect 114511 259009 114602 259127
rect 114302 258967 114602 259009
rect 114302 258849 114393 258967
rect 114511 258849 114602 258967
rect 114302 241127 114602 258849
rect 114302 241009 114393 241127
rect 114511 241009 114602 241127
rect 114302 240967 114602 241009
rect 114302 240849 114393 240967
rect 114511 240849 114602 240967
rect 114302 223127 114602 240849
rect 114302 223009 114393 223127
rect 114511 223009 114602 223127
rect 114302 222967 114602 223009
rect 114302 222849 114393 222967
rect 114511 222849 114602 222967
rect 114302 205127 114602 222849
rect 114302 205009 114393 205127
rect 114511 205009 114602 205127
rect 114302 204967 114602 205009
rect 114302 204849 114393 204967
rect 114511 204849 114602 204967
rect 114302 187127 114602 204849
rect 114302 187009 114393 187127
rect 114511 187009 114602 187127
rect 114302 186967 114602 187009
rect 114302 186849 114393 186967
rect 114511 186849 114602 186967
rect 114302 169127 114602 186849
rect 114302 169009 114393 169127
rect 114511 169009 114602 169127
rect 114302 168967 114602 169009
rect 114302 168849 114393 168967
rect 114511 168849 114602 168967
rect 114302 151127 114602 168849
rect 114302 151009 114393 151127
rect 114511 151009 114602 151127
rect 114302 150967 114602 151009
rect 114302 150849 114393 150967
rect 114511 150849 114602 150967
rect 114302 133127 114602 150849
rect 114302 133009 114393 133127
rect 114511 133009 114602 133127
rect 114302 132967 114602 133009
rect 114302 132849 114393 132967
rect 114511 132849 114602 132967
rect 114302 115127 114602 132849
rect 114302 115009 114393 115127
rect 114511 115009 114602 115127
rect 114302 114967 114602 115009
rect 114302 114849 114393 114967
rect 114511 114849 114602 114967
rect 114302 97127 114602 114849
rect 114302 97009 114393 97127
rect 114511 97009 114602 97127
rect 114302 96967 114602 97009
rect 114302 96849 114393 96967
rect 114511 96849 114602 96967
rect 114302 79127 114602 96849
rect 114302 79009 114393 79127
rect 114511 79009 114602 79127
rect 114302 78967 114602 79009
rect 114302 78849 114393 78967
rect 114511 78849 114602 78967
rect 114302 61127 114602 78849
rect 114302 61009 114393 61127
rect 114511 61009 114602 61127
rect 114302 60967 114602 61009
rect 114302 60849 114393 60967
rect 114511 60849 114602 60967
rect 114302 43127 114602 60849
rect 114302 43009 114393 43127
rect 114511 43009 114602 43127
rect 114302 42967 114602 43009
rect 114302 42849 114393 42967
rect 114511 42849 114602 42967
rect 114302 25127 114602 42849
rect 114302 25009 114393 25127
rect 114511 25009 114602 25127
rect 114302 24967 114602 25009
rect 114302 24849 114393 24967
rect 114511 24849 114602 24967
rect 114302 7127 114602 24849
rect 114302 7009 114393 7127
rect 114511 7009 114602 7127
rect 114302 6967 114602 7009
rect 114302 6849 114393 6967
rect 114511 6849 114602 6967
rect 105302 -3581 105393 -3463
rect 105511 -3581 105602 -3463
rect 105302 -3623 105602 -3581
rect 105302 -3741 105393 -3623
rect 105511 -3741 105602 -3623
rect 105302 -3752 105602 -3741
rect 114302 -2993 114602 6849
rect 117902 352889 118202 352900
rect 117902 352771 117993 352889
rect 118111 352771 118202 352889
rect 117902 352729 118202 352771
rect 117902 352611 117993 352729
rect 118111 352611 118202 352729
rect 117902 334727 118202 352611
rect 117902 334609 117993 334727
rect 118111 334609 118202 334727
rect 117902 334567 118202 334609
rect 117902 334449 117993 334567
rect 118111 334449 118202 334567
rect 117902 316727 118202 334449
rect 117902 316609 117993 316727
rect 118111 316609 118202 316727
rect 117902 316567 118202 316609
rect 117902 316449 117993 316567
rect 118111 316449 118202 316567
rect 117902 298727 118202 316449
rect 117902 298609 117993 298727
rect 118111 298609 118202 298727
rect 117902 298567 118202 298609
rect 117902 298449 117993 298567
rect 118111 298449 118202 298567
rect 117902 280727 118202 298449
rect 117902 280609 117993 280727
rect 118111 280609 118202 280727
rect 117902 280567 118202 280609
rect 117902 280449 117993 280567
rect 118111 280449 118202 280567
rect 117902 262727 118202 280449
rect 117902 262609 117993 262727
rect 118111 262609 118202 262727
rect 117902 262567 118202 262609
rect 117902 262449 117993 262567
rect 118111 262449 118202 262567
rect 117902 244727 118202 262449
rect 117902 244609 117993 244727
rect 118111 244609 118202 244727
rect 117902 244567 118202 244609
rect 117902 244449 117993 244567
rect 118111 244449 118202 244567
rect 117902 226727 118202 244449
rect 117902 226609 117993 226727
rect 118111 226609 118202 226727
rect 117902 226567 118202 226609
rect 117902 226449 117993 226567
rect 118111 226449 118202 226567
rect 117902 208727 118202 226449
rect 117902 208609 117993 208727
rect 118111 208609 118202 208727
rect 117902 208567 118202 208609
rect 117902 208449 117993 208567
rect 118111 208449 118202 208567
rect 117902 190727 118202 208449
rect 117902 190609 117993 190727
rect 118111 190609 118202 190727
rect 117902 190567 118202 190609
rect 117902 190449 117993 190567
rect 118111 190449 118202 190567
rect 117902 172727 118202 190449
rect 117902 172609 117993 172727
rect 118111 172609 118202 172727
rect 117902 172567 118202 172609
rect 117902 172449 117993 172567
rect 118111 172449 118202 172567
rect 117902 154727 118202 172449
rect 117902 154609 117993 154727
rect 118111 154609 118202 154727
rect 117902 154567 118202 154609
rect 117902 154449 117993 154567
rect 118111 154449 118202 154567
rect 117902 136727 118202 154449
rect 117902 136609 117993 136727
rect 118111 136609 118202 136727
rect 117902 136567 118202 136609
rect 117902 136449 117993 136567
rect 118111 136449 118202 136567
rect 117902 118727 118202 136449
rect 117902 118609 117993 118727
rect 118111 118609 118202 118727
rect 117902 118567 118202 118609
rect 117902 118449 117993 118567
rect 118111 118449 118202 118567
rect 117902 100727 118202 118449
rect 117902 100609 117993 100727
rect 118111 100609 118202 100727
rect 117902 100567 118202 100609
rect 117902 100449 117993 100567
rect 118111 100449 118202 100567
rect 117902 82727 118202 100449
rect 117902 82609 117993 82727
rect 118111 82609 118202 82727
rect 117902 82567 118202 82609
rect 117902 82449 117993 82567
rect 118111 82449 118202 82567
rect 117902 64727 118202 82449
rect 117902 64609 117993 64727
rect 118111 64609 118202 64727
rect 117902 64567 118202 64609
rect 117902 64449 117993 64567
rect 118111 64449 118202 64567
rect 117902 46727 118202 64449
rect 117902 46609 117993 46727
rect 118111 46609 118202 46727
rect 117902 46567 118202 46609
rect 117902 46449 117993 46567
rect 118111 46449 118202 46567
rect 117902 28727 118202 46449
rect 117902 28609 117993 28727
rect 118111 28609 118202 28727
rect 117902 28567 118202 28609
rect 117902 28449 117993 28567
rect 118111 28449 118202 28567
rect 117902 10727 118202 28449
rect 117902 10609 117993 10727
rect 118111 10609 118202 10727
rect 117902 10567 118202 10609
rect 117902 10449 117993 10567
rect 118111 10449 118202 10567
rect 117902 -643 118202 10449
rect 117902 -761 117993 -643
rect 118111 -761 118202 -643
rect 117902 -803 118202 -761
rect 117902 -921 117993 -803
rect 118111 -921 118202 -803
rect 117902 -932 118202 -921
rect 119702 336527 120002 353551
rect 119702 336409 119793 336527
rect 119911 336409 120002 336527
rect 119702 336367 120002 336409
rect 119702 336249 119793 336367
rect 119911 336249 120002 336367
rect 119702 318527 120002 336249
rect 119702 318409 119793 318527
rect 119911 318409 120002 318527
rect 119702 318367 120002 318409
rect 119702 318249 119793 318367
rect 119911 318249 120002 318367
rect 119702 300527 120002 318249
rect 119702 300409 119793 300527
rect 119911 300409 120002 300527
rect 119702 300367 120002 300409
rect 119702 300249 119793 300367
rect 119911 300249 120002 300367
rect 119702 282527 120002 300249
rect 119702 282409 119793 282527
rect 119911 282409 120002 282527
rect 119702 282367 120002 282409
rect 119702 282249 119793 282367
rect 119911 282249 120002 282367
rect 119702 264527 120002 282249
rect 119702 264409 119793 264527
rect 119911 264409 120002 264527
rect 119702 264367 120002 264409
rect 119702 264249 119793 264367
rect 119911 264249 120002 264367
rect 119702 246527 120002 264249
rect 119702 246409 119793 246527
rect 119911 246409 120002 246527
rect 119702 246367 120002 246409
rect 119702 246249 119793 246367
rect 119911 246249 120002 246367
rect 119702 228527 120002 246249
rect 119702 228409 119793 228527
rect 119911 228409 120002 228527
rect 119702 228367 120002 228409
rect 119702 228249 119793 228367
rect 119911 228249 120002 228367
rect 119702 210527 120002 228249
rect 119702 210409 119793 210527
rect 119911 210409 120002 210527
rect 119702 210367 120002 210409
rect 119702 210249 119793 210367
rect 119911 210249 120002 210367
rect 119702 192527 120002 210249
rect 119702 192409 119793 192527
rect 119911 192409 120002 192527
rect 119702 192367 120002 192409
rect 119702 192249 119793 192367
rect 119911 192249 120002 192367
rect 119702 174527 120002 192249
rect 119702 174409 119793 174527
rect 119911 174409 120002 174527
rect 119702 174367 120002 174409
rect 119702 174249 119793 174367
rect 119911 174249 120002 174367
rect 119702 156527 120002 174249
rect 119702 156409 119793 156527
rect 119911 156409 120002 156527
rect 119702 156367 120002 156409
rect 119702 156249 119793 156367
rect 119911 156249 120002 156367
rect 119702 138527 120002 156249
rect 119702 138409 119793 138527
rect 119911 138409 120002 138527
rect 119702 138367 120002 138409
rect 119702 138249 119793 138367
rect 119911 138249 120002 138367
rect 119702 120527 120002 138249
rect 119702 120409 119793 120527
rect 119911 120409 120002 120527
rect 119702 120367 120002 120409
rect 119702 120249 119793 120367
rect 119911 120249 120002 120367
rect 119702 102527 120002 120249
rect 119702 102409 119793 102527
rect 119911 102409 120002 102527
rect 119702 102367 120002 102409
rect 119702 102249 119793 102367
rect 119911 102249 120002 102367
rect 119702 84527 120002 102249
rect 119702 84409 119793 84527
rect 119911 84409 120002 84527
rect 119702 84367 120002 84409
rect 119702 84249 119793 84367
rect 119911 84249 120002 84367
rect 119702 66527 120002 84249
rect 119702 66409 119793 66527
rect 119911 66409 120002 66527
rect 119702 66367 120002 66409
rect 119702 66249 119793 66367
rect 119911 66249 120002 66367
rect 119702 48527 120002 66249
rect 119702 48409 119793 48527
rect 119911 48409 120002 48527
rect 119702 48367 120002 48409
rect 119702 48249 119793 48367
rect 119911 48249 120002 48367
rect 119702 30527 120002 48249
rect 119702 30409 119793 30527
rect 119911 30409 120002 30527
rect 119702 30367 120002 30409
rect 119702 30249 119793 30367
rect 119911 30249 120002 30367
rect 119702 12527 120002 30249
rect 119702 12409 119793 12527
rect 119911 12409 120002 12527
rect 119702 12367 120002 12409
rect 119702 12249 119793 12367
rect 119911 12249 120002 12367
rect 119702 -1583 120002 12249
rect 119702 -1701 119793 -1583
rect 119911 -1701 120002 -1583
rect 119702 -1743 120002 -1701
rect 119702 -1861 119793 -1743
rect 119911 -1861 120002 -1743
rect 119702 -1872 120002 -1861
rect 121502 338327 121802 354491
rect 121502 338209 121593 338327
rect 121711 338209 121802 338327
rect 121502 338167 121802 338209
rect 121502 338049 121593 338167
rect 121711 338049 121802 338167
rect 121502 320327 121802 338049
rect 121502 320209 121593 320327
rect 121711 320209 121802 320327
rect 121502 320167 121802 320209
rect 121502 320049 121593 320167
rect 121711 320049 121802 320167
rect 121502 302327 121802 320049
rect 121502 302209 121593 302327
rect 121711 302209 121802 302327
rect 121502 302167 121802 302209
rect 121502 302049 121593 302167
rect 121711 302049 121802 302167
rect 121502 284327 121802 302049
rect 121502 284209 121593 284327
rect 121711 284209 121802 284327
rect 121502 284167 121802 284209
rect 121502 284049 121593 284167
rect 121711 284049 121802 284167
rect 121502 266327 121802 284049
rect 121502 266209 121593 266327
rect 121711 266209 121802 266327
rect 121502 266167 121802 266209
rect 121502 266049 121593 266167
rect 121711 266049 121802 266167
rect 121502 248327 121802 266049
rect 121502 248209 121593 248327
rect 121711 248209 121802 248327
rect 121502 248167 121802 248209
rect 121502 248049 121593 248167
rect 121711 248049 121802 248167
rect 121502 230327 121802 248049
rect 121502 230209 121593 230327
rect 121711 230209 121802 230327
rect 121502 230167 121802 230209
rect 121502 230049 121593 230167
rect 121711 230049 121802 230167
rect 121502 212327 121802 230049
rect 121502 212209 121593 212327
rect 121711 212209 121802 212327
rect 121502 212167 121802 212209
rect 121502 212049 121593 212167
rect 121711 212049 121802 212167
rect 121502 194327 121802 212049
rect 121502 194209 121593 194327
rect 121711 194209 121802 194327
rect 121502 194167 121802 194209
rect 121502 194049 121593 194167
rect 121711 194049 121802 194167
rect 121502 176327 121802 194049
rect 121502 176209 121593 176327
rect 121711 176209 121802 176327
rect 121502 176167 121802 176209
rect 121502 176049 121593 176167
rect 121711 176049 121802 176167
rect 121502 158327 121802 176049
rect 121502 158209 121593 158327
rect 121711 158209 121802 158327
rect 121502 158167 121802 158209
rect 121502 158049 121593 158167
rect 121711 158049 121802 158167
rect 121502 140327 121802 158049
rect 121502 140209 121593 140327
rect 121711 140209 121802 140327
rect 121502 140167 121802 140209
rect 121502 140049 121593 140167
rect 121711 140049 121802 140167
rect 121502 122327 121802 140049
rect 121502 122209 121593 122327
rect 121711 122209 121802 122327
rect 121502 122167 121802 122209
rect 121502 122049 121593 122167
rect 121711 122049 121802 122167
rect 121502 104327 121802 122049
rect 121502 104209 121593 104327
rect 121711 104209 121802 104327
rect 121502 104167 121802 104209
rect 121502 104049 121593 104167
rect 121711 104049 121802 104167
rect 121502 86327 121802 104049
rect 121502 86209 121593 86327
rect 121711 86209 121802 86327
rect 121502 86167 121802 86209
rect 121502 86049 121593 86167
rect 121711 86049 121802 86167
rect 121502 68327 121802 86049
rect 121502 68209 121593 68327
rect 121711 68209 121802 68327
rect 121502 68167 121802 68209
rect 121502 68049 121593 68167
rect 121711 68049 121802 68167
rect 121502 50327 121802 68049
rect 121502 50209 121593 50327
rect 121711 50209 121802 50327
rect 121502 50167 121802 50209
rect 121502 50049 121593 50167
rect 121711 50049 121802 50167
rect 121502 32327 121802 50049
rect 121502 32209 121593 32327
rect 121711 32209 121802 32327
rect 121502 32167 121802 32209
rect 121502 32049 121593 32167
rect 121711 32049 121802 32167
rect 121502 14327 121802 32049
rect 121502 14209 121593 14327
rect 121711 14209 121802 14327
rect 121502 14167 121802 14209
rect 121502 14049 121593 14167
rect 121711 14049 121802 14167
rect 121502 -2523 121802 14049
rect 121502 -2641 121593 -2523
rect 121711 -2641 121802 -2523
rect 121502 -2683 121802 -2641
rect 121502 -2801 121593 -2683
rect 121711 -2801 121802 -2683
rect 121502 -2812 121802 -2801
rect 123302 340127 123602 355431
rect 132302 355239 132602 355720
rect 132302 355121 132393 355239
rect 132511 355121 132602 355239
rect 132302 355079 132602 355121
rect 132302 354961 132393 355079
rect 132511 354961 132602 355079
rect 130502 354299 130802 354780
rect 130502 354181 130593 354299
rect 130711 354181 130802 354299
rect 130502 354139 130802 354181
rect 130502 354021 130593 354139
rect 130711 354021 130802 354139
rect 128702 353359 129002 353840
rect 128702 353241 128793 353359
rect 128911 353241 129002 353359
rect 128702 353199 129002 353241
rect 128702 353081 128793 353199
rect 128911 353081 129002 353199
rect 123302 340009 123393 340127
rect 123511 340009 123602 340127
rect 123302 339967 123602 340009
rect 123302 339849 123393 339967
rect 123511 339849 123602 339967
rect 123302 322127 123602 339849
rect 123302 322009 123393 322127
rect 123511 322009 123602 322127
rect 123302 321967 123602 322009
rect 123302 321849 123393 321967
rect 123511 321849 123602 321967
rect 123302 304127 123602 321849
rect 123302 304009 123393 304127
rect 123511 304009 123602 304127
rect 123302 303967 123602 304009
rect 123302 303849 123393 303967
rect 123511 303849 123602 303967
rect 123302 286127 123602 303849
rect 123302 286009 123393 286127
rect 123511 286009 123602 286127
rect 123302 285967 123602 286009
rect 123302 285849 123393 285967
rect 123511 285849 123602 285967
rect 123302 268127 123602 285849
rect 123302 268009 123393 268127
rect 123511 268009 123602 268127
rect 123302 267967 123602 268009
rect 123302 267849 123393 267967
rect 123511 267849 123602 267967
rect 123302 250127 123602 267849
rect 123302 250009 123393 250127
rect 123511 250009 123602 250127
rect 123302 249967 123602 250009
rect 123302 249849 123393 249967
rect 123511 249849 123602 249967
rect 123302 232127 123602 249849
rect 123302 232009 123393 232127
rect 123511 232009 123602 232127
rect 123302 231967 123602 232009
rect 123302 231849 123393 231967
rect 123511 231849 123602 231967
rect 123302 214127 123602 231849
rect 123302 214009 123393 214127
rect 123511 214009 123602 214127
rect 123302 213967 123602 214009
rect 123302 213849 123393 213967
rect 123511 213849 123602 213967
rect 123302 196127 123602 213849
rect 123302 196009 123393 196127
rect 123511 196009 123602 196127
rect 123302 195967 123602 196009
rect 123302 195849 123393 195967
rect 123511 195849 123602 195967
rect 123302 178127 123602 195849
rect 123302 178009 123393 178127
rect 123511 178009 123602 178127
rect 123302 177967 123602 178009
rect 123302 177849 123393 177967
rect 123511 177849 123602 177967
rect 123302 160127 123602 177849
rect 123302 160009 123393 160127
rect 123511 160009 123602 160127
rect 123302 159967 123602 160009
rect 123302 159849 123393 159967
rect 123511 159849 123602 159967
rect 123302 142127 123602 159849
rect 123302 142009 123393 142127
rect 123511 142009 123602 142127
rect 123302 141967 123602 142009
rect 123302 141849 123393 141967
rect 123511 141849 123602 141967
rect 123302 124127 123602 141849
rect 123302 124009 123393 124127
rect 123511 124009 123602 124127
rect 123302 123967 123602 124009
rect 123302 123849 123393 123967
rect 123511 123849 123602 123967
rect 123302 106127 123602 123849
rect 123302 106009 123393 106127
rect 123511 106009 123602 106127
rect 123302 105967 123602 106009
rect 123302 105849 123393 105967
rect 123511 105849 123602 105967
rect 123302 88127 123602 105849
rect 123302 88009 123393 88127
rect 123511 88009 123602 88127
rect 123302 87967 123602 88009
rect 123302 87849 123393 87967
rect 123511 87849 123602 87967
rect 123302 70127 123602 87849
rect 123302 70009 123393 70127
rect 123511 70009 123602 70127
rect 123302 69967 123602 70009
rect 123302 69849 123393 69967
rect 123511 69849 123602 69967
rect 123302 52127 123602 69849
rect 123302 52009 123393 52127
rect 123511 52009 123602 52127
rect 123302 51967 123602 52009
rect 123302 51849 123393 51967
rect 123511 51849 123602 51967
rect 123302 34127 123602 51849
rect 123302 34009 123393 34127
rect 123511 34009 123602 34127
rect 123302 33967 123602 34009
rect 123302 33849 123393 33967
rect 123511 33849 123602 33967
rect 123302 16127 123602 33849
rect 123302 16009 123393 16127
rect 123511 16009 123602 16127
rect 123302 15967 123602 16009
rect 123302 15849 123393 15967
rect 123511 15849 123602 15967
rect 114302 -3111 114393 -2993
rect 114511 -3111 114602 -2993
rect 114302 -3153 114602 -3111
rect 114302 -3271 114393 -3153
rect 114511 -3271 114602 -3153
rect 114302 -3752 114602 -3271
rect 123302 -3463 123602 15849
rect 126902 352419 127202 352900
rect 126902 352301 126993 352419
rect 127111 352301 127202 352419
rect 126902 352259 127202 352301
rect 126902 352141 126993 352259
rect 127111 352141 127202 352259
rect 126902 343727 127202 352141
rect 126902 343609 126993 343727
rect 127111 343609 127202 343727
rect 126902 343567 127202 343609
rect 126902 343449 126993 343567
rect 127111 343449 127202 343567
rect 126902 325727 127202 343449
rect 126902 325609 126993 325727
rect 127111 325609 127202 325727
rect 126902 325567 127202 325609
rect 126902 325449 126993 325567
rect 127111 325449 127202 325567
rect 126902 307727 127202 325449
rect 126902 307609 126993 307727
rect 127111 307609 127202 307727
rect 126902 307567 127202 307609
rect 126902 307449 126993 307567
rect 127111 307449 127202 307567
rect 126902 289727 127202 307449
rect 126902 289609 126993 289727
rect 127111 289609 127202 289727
rect 126902 289567 127202 289609
rect 126902 289449 126993 289567
rect 127111 289449 127202 289567
rect 126902 271727 127202 289449
rect 126902 271609 126993 271727
rect 127111 271609 127202 271727
rect 126902 271567 127202 271609
rect 126902 271449 126993 271567
rect 127111 271449 127202 271567
rect 126902 253727 127202 271449
rect 126902 253609 126993 253727
rect 127111 253609 127202 253727
rect 126902 253567 127202 253609
rect 126902 253449 126993 253567
rect 127111 253449 127202 253567
rect 126902 235727 127202 253449
rect 126902 235609 126993 235727
rect 127111 235609 127202 235727
rect 126902 235567 127202 235609
rect 126902 235449 126993 235567
rect 127111 235449 127202 235567
rect 126902 217727 127202 235449
rect 126902 217609 126993 217727
rect 127111 217609 127202 217727
rect 126902 217567 127202 217609
rect 126902 217449 126993 217567
rect 127111 217449 127202 217567
rect 126902 199727 127202 217449
rect 126902 199609 126993 199727
rect 127111 199609 127202 199727
rect 126902 199567 127202 199609
rect 126902 199449 126993 199567
rect 127111 199449 127202 199567
rect 126902 181727 127202 199449
rect 126902 181609 126993 181727
rect 127111 181609 127202 181727
rect 126902 181567 127202 181609
rect 126902 181449 126993 181567
rect 127111 181449 127202 181567
rect 126902 163727 127202 181449
rect 126902 163609 126993 163727
rect 127111 163609 127202 163727
rect 126902 163567 127202 163609
rect 126902 163449 126993 163567
rect 127111 163449 127202 163567
rect 126902 145727 127202 163449
rect 126902 145609 126993 145727
rect 127111 145609 127202 145727
rect 126902 145567 127202 145609
rect 126902 145449 126993 145567
rect 127111 145449 127202 145567
rect 126902 127727 127202 145449
rect 126902 127609 126993 127727
rect 127111 127609 127202 127727
rect 126902 127567 127202 127609
rect 126902 127449 126993 127567
rect 127111 127449 127202 127567
rect 126902 109727 127202 127449
rect 126902 109609 126993 109727
rect 127111 109609 127202 109727
rect 126902 109567 127202 109609
rect 126902 109449 126993 109567
rect 127111 109449 127202 109567
rect 126902 91727 127202 109449
rect 126902 91609 126993 91727
rect 127111 91609 127202 91727
rect 126902 91567 127202 91609
rect 126902 91449 126993 91567
rect 127111 91449 127202 91567
rect 126902 73727 127202 91449
rect 126902 73609 126993 73727
rect 127111 73609 127202 73727
rect 126902 73567 127202 73609
rect 126902 73449 126993 73567
rect 127111 73449 127202 73567
rect 126902 55727 127202 73449
rect 126902 55609 126993 55727
rect 127111 55609 127202 55727
rect 126902 55567 127202 55609
rect 126902 55449 126993 55567
rect 127111 55449 127202 55567
rect 126902 37727 127202 55449
rect 126902 37609 126993 37727
rect 127111 37609 127202 37727
rect 126902 37567 127202 37609
rect 126902 37449 126993 37567
rect 127111 37449 127202 37567
rect 126902 19727 127202 37449
rect 126902 19609 126993 19727
rect 127111 19609 127202 19727
rect 126902 19567 127202 19609
rect 126902 19449 126993 19567
rect 127111 19449 127202 19567
rect 126902 1727 127202 19449
rect 126902 1609 126993 1727
rect 127111 1609 127202 1727
rect 126902 1567 127202 1609
rect 126902 1449 126993 1567
rect 127111 1449 127202 1567
rect 126902 -173 127202 1449
rect 126902 -291 126993 -173
rect 127111 -291 127202 -173
rect 126902 -333 127202 -291
rect 126902 -451 126993 -333
rect 127111 -451 127202 -333
rect 126902 -932 127202 -451
rect 128702 345527 129002 353081
rect 128702 345409 128793 345527
rect 128911 345409 129002 345527
rect 128702 345367 129002 345409
rect 128702 345249 128793 345367
rect 128911 345249 129002 345367
rect 128702 327527 129002 345249
rect 128702 327409 128793 327527
rect 128911 327409 129002 327527
rect 128702 327367 129002 327409
rect 128702 327249 128793 327367
rect 128911 327249 129002 327367
rect 128702 309527 129002 327249
rect 128702 309409 128793 309527
rect 128911 309409 129002 309527
rect 128702 309367 129002 309409
rect 128702 309249 128793 309367
rect 128911 309249 129002 309367
rect 128702 291527 129002 309249
rect 128702 291409 128793 291527
rect 128911 291409 129002 291527
rect 128702 291367 129002 291409
rect 128702 291249 128793 291367
rect 128911 291249 129002 291367
rect 128702 273527 129002 291249
rect 128702 273409 128793 273527
rect 128911 273409 129002 273527
rect 128702 273367 129002 273409
rect 128702 273249 128793 273367
rect 128911 273249 129002 273367
rect 128702 255527 129002 273249
rect 128702 255409 128793 255527
rect 128911 255409 129002 255527
rect 128702 255367 129002 255409
rect 128702 255249 128793 255367
rect 128911 255249 129002 255367
rect 128702 237527 129002 255249
rect 128702 237409 128793 237527
rect 128911 237409 129002 237527
rect 128702 237367 129002 237409
rect 128702 237249 128793 237367
rect 128911 237249 129002 237367
rect 128702 219527 129002 237249
rect 128702 219409 128793 219527
rect 128911 219409 129002 219527
rect 128702 219367 129002 219409
rect 128702 219249 128793 219367
rect 128911 219249 129002 219367
rect 128702 201527 129002 219249
rect 128702 201409 128793 201527
rect 128911 201409 129002 201527
rect 128702 201367 129002 201409
rect 128702 201249 128793 201367
rect 128911 201249 129002 201367
rect 128702 183527 129002 201249
rect 128702 183409 128793 183527
rect 128911 183409 129002 183527
rect 128702 183367 129002 183409
rect 128702 183249 128793 183367
rect 128911 183249 129002 183367
rect 128702 165527 129002 183249
rect 128702 165409 128793 165527
rect 128911 165409 129002 165527
rect 128702 165367 129002 165409
rect 128702 165249 128793 165367
rect 128911 165249 129002 165367
rect 128702 147527 129002 165249
rect 128702 147409 128793 147527
rect 128911 147409 129002 147527
rect 128702 147367 129002 147409
rect 128702 147249 128793 147367
rect 128911 147249 129002 147367
rect 128702 129527 129002 147249
rect 128702 129409 128793 129527
rect 128911 129409 129002 129527
rect 128702 129367 129002 129409
rect 128702 129249 128793 129367
rect 128911 129249 129002 129367
rect 128702 111527 129002 129249
rect 128702 111409 128793 111527
rect 128911 111409 129002 111527
rect 128702 111367 129002 111409
rect 128702 111249 128793 111367
rect 128911 111249 129002 111367
rect 128702 93527 129002 111249
rect 128702 93409 128793 93527
rect 128911 93409 129002 93527
rect 128702 93367 129002 93409
rect 128702 93249 128793 93367
rect 128911 93249 129002 93367
rect 128702 75527 129002 93249
rect 128702 75409 128793 75527
rect 128911 75409 129002 75527
rect 128702 75367 129002 75409
rect 128702 75249 128793 75367
rect 128911 75249 129002 75367
rect 128702 57527 129002 75249
rect 128702 57409 128793 57527
rect 128911 57409 129002 57527
rect 128702 57367 129002 57409
rect 128702 57249 128793 57367
rect 128911 57249 129002 57367
rect 128702 39527 129002 57249
rect 128702 39409 128793 39527
rect 128911 39409 129002 39527
rect 128702 39367 129002 39409
rect 128702 39249 128793 39367
rect 128911 39249 129002 39367
rect 128702 21527 129002 39249
rect 128702 21409 128793 21527
rect 128911 21409 129002 21527
rect 128702 21367 129002 21409
rect 128702 21249 128793 21367
rect 128911 21249 129002 21367
rect 128702 3527 129002 21249
rect 128702 3409 128793 3527
rect 128911 3409 129002 3527
rect 128702 3367 129002 3409
rect 128702 3249 128793 3367
rect 128911 3249 129002 3367
rect 128702 -1113 129002 3249
rect 128702 -1231 128793 -1113
rect 128911 -1231 129002 -1113
rect 128702 -1273 129002 -1231
rect 128702 -1391 128793 -1273
rect 128911 -1391 129002 -1273
rect 128702 -1872 129002 -1391
rect 130502 347327 130802 354021
rect 130502 347209 130593 347327
rect 130711 347209 130802 347327
rect 130502 347167 130802 347209
rect 130502 347049 130593 347167
rect 130711 347049 130802 347167
rect 130502 329327 130802 347049
rect 130502 329209 130593 329327
rect 130711 329209 130802 329327
rect 130502 329167 130802 329209
rect 130502 329049 130593 329167
rect 130711 329049 130802 329167
rect 130502 311327 130802 329049
rect 130502 311209 130593 311327
rect 130711 311209 130802 311327
rect 130502 311167 130802 311209
rect 130502 311049 130593 311167
rect 130711 311049 130802 311167
rect 130502 293327 130802 311049
rect 130502 293209 130593 293327
rect 130711 293209 130802 293327
rect 130502 293167 130802 293209
rect 130502 293049 130593 293167
rect 130711 293049 130802 293167
rect 130502 275327 130802 293049
rect 130502 275209 130593 275327
rect 130711 275209 130802 275327
rect 130502 275167 130802 275209
rect 130502 275049 130593 275167
rect 130711 275049 130802 275167
rect 130502 257327 130802 275049
rect 130502 257209 130593 257327
rect 130711 257209 130802 257327
rect 130502 257167 130802 257209
rect 130502 257049 130593 257167
rect 130711 257049 130802 257167
rect 130502 239327 130802 257049
rect 130502 239209 130593 239327
rect 130711 239209 130802 239327
rect 130502 239167 130802 239209
rect 130502 239049 130593 239167
rect 130711 239049 130802 239167
rect 130502 221327 130802 239049
rect 130502 221209 130593 221327
rect 130711 221209 130802 221327
rect 130502 221167 130802 221209
rect 130502 221049 130593 221167
rect 130711 221049 130802 221167
rect 130502 203327 130802 221049
rect 130502 203209 130593 203327
rect 130711 203209 130802 203327
rect 130502 203167 130802 203209
rect 130502 203049 130593 203167
rect 130711 203049 130802 203167
rect 130502 185327 130802 203049
rect 130502 185209 130593 185327
rect 130711 185209 130802 185327
rect 130502 185167 130802 185209
rect 130502 185049 130593 185167
rect 130711 185049 130802 185167
rect 130502 167327 130802 185049
rect 130502 167209 130593 167327
rect 130711 167209 130802 167327
rect 130502 167167 130802 167209
rect 130502 167049 130593 167167
rect 130711 167049 130802 167167
rect 130502 149327 130802 167049
rect 130502 149209 130593 149327
rect 130711 149209 130802 149327
rect 130502 149167 130802 149209
rect 130502 149049 130593 149167
rect 130711 149049 130802 149167
rect 130502 131327 130802 149049
rect 130502 131209 130593 131327
rect 130711 131209 130802 131327
rect 130502 131167 130802 131209
rect 130502 131049 130593 131167
rect 130711 131049 130802 131167
rect 130502 113327 130802 131049
rect 130502 113209 130593 113327
rect 130711 113209 130802 113327
rect 130502 113167 130802 113209
rect 130502 113049 130593 113167
rect 130711 113049 130802 113167
rect 130502 95327 130802 113049
rect 130502 95209 130593 95327
rect 130711 95209 130802 95327
rect 130502 95167 130802 95209
rect 130502 95049 130593 95167
rect 130711 95049 130802 95167
rect 130502 77327 130802 95049
rect 130502 77209 130593 77327
rect 130711 77209 130802 77327
rect 130502 77167 130802 77209
rect 130502 77049 130593 77167
rect 130711 77049 130802 77167
rect 130502 59327 130802 77049
rect 130502 59209 130593 59327
rect 130711 59209 130802 59327
rect 130502 59167 130802 59209
rect 130502 59049 130593 59167
rect 130711 59049 130802 59167
rect 130502 41327 130802 59049
rect 130502 41209 130593 41327
rect 130711 41209 130802 41327
rect 130502 41167 130802 41209
rect 130502 41049 130593 41167
rect 130711 41049 130802 41167
rect 130502 23327 130802 41049
rect 130502 23209 130593 23327
rect 130711 23209 130802 23327
rect 130502 23167 130802 23209
rect 130502 23049 130593 23167
rect 130711 23049 130802 23167
rect 130502 5327 130802 23049
rect 130502 5209 130593 5327
rect 130711 5209 130802 5327
rect 130502 5167 130802 5209
rect 130502 5049 130593 5167
rect 130711 5049 130802 5167
rect 130502 -2053 130802 5049
rect 130502 -2171 130593 -2053
rect 130711 -2171 130802 -2053
rect 130502 -2213 130802 -2171
rect 130502 -2331 130593 -2213
rect 130711 -2331 130802 -2213
rect 130502 -2812 130802 -2331
rect 132302 349127 132602 354961
rect 141302 355709 141602 355720
rect 141302 355591 141393 355709
rect 141511 355591 141602 355709
rect 141302 355549 141602 355591
rect 141302 355431 141393 355549
rect 141511 355431 141602 355549
rect 139502 354769 139802 354780
rect 139502 354651 139593 354769
rect 139711 354651 139802 354769
rect 139502 354609 139802 354651
rect 139502 354491 139593 354609
rect 139711 354491 139802 354609
rect 137702 353829 138002 353840
rect 137702 353711 137793 353829
rect 137911 353711 138002 353829
rect 137702 353669 138002 353711
rect 137702 353551 137793 353669
rect 137911 353551 138002 353669
rect 132302 349009 132393 349127
rect 132511 349009 132602 349127
rect 132302 348967 132602 349009
rect 132302 348849 132393 348967
rect 132511 348849 132602 348967
rect 132302 331127 132602 348849
rect 132302 331009 132393 331127
rect 132511 331009 132602 331127
rect 132302 330967 132602 331009
rect 132302 330849 132393 330967
rect 132511 330849 132602 330967
rect 132302 313127 132602 330849
rect 132302 313009 132393 313127
rect 132511 313009 132602 313127
rect 132302 312967 132602 313009
rect 132302 312849 132393 312967
rect 132511 312849 132602 312967
rect 132302 295127 132602 312849
rect 132302 295009 132393 295127
rect 132511 295009 132602 295127
rect 132302 294967 132602 295009
rect 132302 294849 132393 294967
rect 132511 294849 132602 294967
rect 132302 277127 132602 294849
rect 132302 277009 132393 277127
rect 132511 277009 132602 277127
rect 132302 276967 132602 277009
rect 132302 276849 132393 276967
rect 132511 276849 132602 276967
rect 132302 259127 132602 276849
rect 132302 259009 132393 259127
rect 132511 259009 132602 259127
rect 132302 258967 132602 259009
rect 132302 258849 132393 258967
rect 132511 258849 132602 258967
rect 132302 241127 132602 258849
rect 132302 241009 132393 241127
rect 132511 241009 132602 241127
rect 132302 240967 132602 241009
rect 132302 240849 132393 240967
rect 132511 240849 132602 240967
rect 132302 223127 132602 240849
rect 132302 223009 132393 223127
rect 132511 223009 132602 223127
rect 132302 222967 132602 223009
rect 132302 222849 132393 222967
rect 132511 222849 132602 222967
rect 132302 205127 132602 222849
rect 132302 205009 132393 205127
rect 132511 205009 132602 205127
rect 132302 204967 132602 205009
rect 132302 204849 132393 204967
rect 132511 204849 132602 204967
rect 132302 187127 132602 204849
rect 132302 187009 132393 187127
rect 132511 187009 132602 187127
rect 132302 186967 132602 187009
rect 132302 186849 132393 186967
rect 132511 186849 132602 186967
rect 132302 169127 132602 186849
rect 132302 169009 132393 169127
rect 132511 169009 132602 169127
rect 132302 168967 132602 169009
rect 132302 168849 132393 168967
rect 132511 168849 132602 168967
rect 132302 151127 132602 168849
rect 132302 151009 132393 151127
rect 132511 151009 132602 151127
rect 132302 150967 132602 151009
rect 132302 150849 132393 150967
rect 132511 150849 132602 150967
rect 132302 133127 132602 150849
rect 132302 133009 132393 133127
rect 132511 133009 132602 133127
rect 132302 132967 132602 133009
rect 132302 132849 132393 132967
rect 132511 132849 132602 132967
rect 132302 115127 132602 132849
rect 132302 115009 132393 115127
rect 132511 115009 132602 115127
rect 132302 114967 132602 115009
rect 132302 114849 132393 114967
rect 132511 114849 132602 114967
rect 132302 97127 132602 114849
rect 132302 97009 132393 97127
rect 132511 97009 132602 97127
rect 132302 96967 132602 97009
rect 132302 96849 132393 96967
rect 132511 96849 132602 96967
rect 132302 79127 132602 96849
rect 132302 79009 132393 79127
rect 132511 79009 132602 79127
rect 132302 78967 132602 79009
rect 132302 78849 132393 78967
rect 132511 78849 132602 78967
rect 132302 61127 132602 78849
rect 132302 61009 132393 61127
rect 132511 61009 132602 61127
rect 132302 60967 132602 61009
rect 132302 60849 132393 60967
rect 132511 60849 132602 60967
rect 132302 43127 132602 60849
rect 132302 43009 132393 43127
rect 132511 43009 132602 43127
rect 132302 42967 132602 43009
rect 132302 42849 132393 42967
rect 132511 42849 132602 42967
rect 132302 25127 132602 42849
rect 132302 25009 132393 25127
rect 132511 25009 132602 25127
rect 132302 24967 132602 25009
rect 132302 24849 132393 24967
rect 132511 24849 132602 24967
rect 132302 7127 132602 24849
rect 132302 7009 132393 7127
rect 132511 7009 132602 7127
rect 132302 6967 132602 7009
rect 132302 6849 132393 6967
rect 132511 6849 132602 6967
rect 123302 -3581 123393 -3463
rect 123511 -3581 123602 -3463
rect 123302 -3623 123602 -3581
rect 123302 -3741 123393 -3623
rect 123511 -3741 123602 -3623
rect 123302 -3752 123602 -3741
rect 132302 -2993 132602 6849
rect 135902 352889 136202 352900
rect 135902 352771 135993 352889
rect 136111 352771 136202 352889
rect 135902 352729 136202 352771
rect 135902 352611 135993 352729
rect 136111 352611 136202 352729
rect 135902 334727 136202 352611
rect 135902 334609 135993 334727
rect 136111 334609 136202 334727
rect 135902 334567 136202 334609
rect 135902 334449 135993 334567
rect 136111 334449 136202 334567
rect 135902 316727 136202 334449
rect 135902 316609 135993 316727
rect 136111 316609 136202 316727
rect 135902 316567 136202 316609
rect 135902 316449 135993 316567
rect 136111 316449 136202 316567
rect 135902 298727 136202 316449
rect 135902 298609 135993 298727
rect 136111 298609 136202 298727
rect 135902 298567 136202 298609
rect 135902 298449 135993 298567
rect 136111 298449 136202 298567
rect 135902 280727 136202 298449
rect 135902 280609 135993 280727
rect 136111 280609 136202 280727
rect 135902 280567 136202 280609
rect 135902 280449 135993 280567
rect 136111 280449 136202 280567
rect 135902 262727 136202 280449
rect 135902 262609 135993 262727
rect 136111 262609 136202 262727
rect 135902 262567 136202 262609
rect 135902 262449 135993 262567
rect 136111 262449 136202 262567
rect 135902 244727 136202 262449
rect 135902 244609 135993 244727
rect 136111 244609 136202 244727
rect 135902 244567 136202 244609
rect 135902 244449 135993 244567
rect 136111 244449 136202 244567
rect 135902 226727 136202 244449
rect 135902 226609 135993 226727
rect 136111 226609 136202 226727
rect 135902 226567 136202 226609
rect 135902 226449 135993 226567
rect 136111 226449 136202 226567
rect 135902 208727 136202 226449
rect 135902 208609 135993 208727
rect 136111 208609 136202 208727
rect 135902 208567 136202 208609
rect 135902 208449 135993 208567
rect 136111 208449 136202 208567
rect 135902 190727 136202 208449
rect 135902 190609 135993 190727
rect 136111 190609 136202 190727
rect 135902 190567 136202 190609
rect 135902 190449 135993 190567
rect 136111 190449 136202 190567
rect 135902 172727 136202 190449
rect 135902 172609 135993 172727
rect 136111 172609 136202 172727
rect 135902 172567 136202 172609
rect 135902 172449 135993 172567
rect 136111 172449 136202 172567
rect 135902 154727 136202 172449
rect 135902 154609 135993 154727
rect 136111 154609 136202 154727
rect 135902 154567 136202 154609
rect 135902 154449 135993 154567
rect 136111 154449 136202 154567
rect 135902 136727 136202 154449
rect 135902 136609 135993 136727
rect 136111 136609 136202 136727
rect 135902 136567 136202 136609
rect 135902 136449 135993 136567
rect 136111 136449 136202 136567
rect 135902 118727 136202 136449
rect 135902 118609 135993 118727
rect 136111 118609 136202 118727
rect 135902 118567 136202 118609
rect 135902 118449 135993 118567
rect 136111 118449 136202 118567
rect 135902 100727 136202 118449
rect 135902 100609 135993 100727
rect 136111 100609 136202 100727
rect 135902 100567 136202 100609
rect 135902 100449 135993 100567
rect 136111 100449 136202 100567
rect 135902 82727 136202 100449
rect 135902 82609 135993 82727
rect 136111 82609 136202 82727
rect 135902 82567 136202 82609
rect 135902 82449 135993 82567
rect 136111 82449 136202 82567
rect 135902 64727 136202 82449
rect 135902 64609 135993 64727
rect 136111 64609 136202 64727
rect 135902 64567 136202 64609
rect 135902 64449 135993 64567
rect 136111 64449 136202 64567
rect 135902 46727 136202 64449
rect 135902 46609 135993 46727
rect 136111 46609 136202 46727
rect 135902 46567 136202 46609
rect 135902 46449 135993 46567
rect 136111 46449 136202 46567
rect 135902 28727 136202 46449
rect 135902 28609 135993 28727
rect 136111 28609 136202 28727
rect 135902 28567 136202 28609
rect 135902 28449 135993 28567
rect 136111 28449 136202 28567
rect 135902 10727 136202 28449
rect 135902 10609 135993 10727
rect 136111 10609 136202 10727
rect 135902 10567 136202 10609
rect 135902 10449 135993 10567
rect 136111 10449 136202 10567
rect 135902 -643 136202 10449
rect 135902 -761 135993 -643
rect 136111 -761 136202 -643
rect 135902 -803 136202 -761
rect 135902 -921 135993 -803
rect 136111 -921 136202 -803
rect 135902 -932 136202 -921
rect 137702 336527 138002 353551
rect 137702 336409 137793 336527
rect 137911 336409 138002 336527
rect 137702 336367 138002 336409
rect 137702 336249 137793 336367
rect 137911 336249 138002 336367
rect 137702 318527 138002 336249
rect 137702 318409 137793 318527
rect 137911 318409 138002 318527
rect 137702 318367 138002 318409
rect 137702 318249 137793 318367
rect 137911 318249 138002 318367
rect 137702 300527 138002 318249
rect 137702 300409 137793 300527
rect 137911 300409 138002 300527
rect 137702 300367 138002 300409
rect 137702 300249 137793 300367
rect 137911 300249 138002 300367
rect 137702 282527 138002 300249
rect 137702 282409 137793 282527
rect 137911 282409 138002 282527
rect 137702 282367 138002 282409
rect 137702 282249 137793 282367
rect 137911 282249 138002 282367
rect 137702 264527 138002 282249
rect 137702 264409 137793 264527
rect 137911 264409 138002 264527
rect 137702 264367 138002 264409
rect 137702 264249 137793 264367
rect 137911 264249 138002 264367
rect 137702 246527 138002 264249
rect 137702 246409 137793 246527
rect 137911 246409 138002 246527
rect 137702 246367 138002 246409
rect 137702 246249 137793 246367
rect 137911 246249 138002 246367
rect 137702 228527 138002 246249
rect 137702 228409 137793 228527
rect 137911 228409 138002 228527
rect 137702 228367 138002 228409
rect 137702 228249 137793 228367
rect 137911 228249 138002 228367
rect 137702 210527 138002 228249
rect 137702 210409 137793 210527
rect 137911 210409 138002 210527
rect 137702 210367 138002 210409
rect 137702 210249 137793 210367
rect 137911 210249 138002 210367
rect 137702 192527 138002 210249
rect 137702 192409 137793 192527
rect 137911 192409 138002 192527
rect 137702 192367 138002 192409
rect 137702 192249 137793 192367
rect 137911 192249 138002 192367
rect 137702 174527 138002 192249
rect 137702 174409 137793 174527
rect 137911 174409 138002 174527
rect 137702 174367 138002 174409
rect 137702 174249 137793 174367
rect 137911 174249 138002 174367
rect 137702 156527 138002 174249
rect 137702 156409 137793 156527
rect 137911 156409 138002 156527
rect 137702 156367 138002 156409
rect 137702 156249 137793 156367
rect 137911 156249 138002 156367
rect 137702 138527 138002 156249
rect 137702 138409 137793 138527
rect 137911 138409 138002 138527
rect 137702 138367 138002 138409
rect 137702 138249 137793 138367
rect 137911 138249 138002 138367
rect 137702 120527 138002 138249
rect 137702 120409 137793 120527
rect 137911 120409 138002 120527
rect 137702 120367 138002 120409
rect 137702 120249 137793 120367
rect 137911 120249 138002 120367
rect 137702 102527 138002 120249
rect 137702 102409 137793 102527
rect 137911 102409 138002 102527
rect 137702 102367 138002 102409
rect 137702 102249 137793 102367
rect 137911 102249 138002 102367
rect 137702 84527 138002 102249
rect 137702 84409 137793 84527
rect 137911 84409 138002 84527
rect 137702 84367 138002 84409
rect 137702 84249 137793 84367
rect 137911 84249 138002 84367
rect 137702 66527 138002 84249
rect 137702 66409 137793 66527
rect 137911 66409 138002 66527
rect 137702 66367 138002 66409
rect 137702 66249 137793 66367
rect 137911 66249 138002 66367
rect 137702 48527 138002 66249
rect 137702 48409 137793 48527
rect 137911 48409 138002 48527
rect 137702 48367 138002 48409
rect 137702 48249 137793 48367
rect 137911 48249 138002 48367
rect 137702 30527 138002 48249
rect 137702 30409 137793 30527
rect 137911 30409 138002 30527
rect 137702 30367 138002 30409
rect 137702 30249 137793 30367
rect 137911 30249 138002 30367
rect 137702 12527 138002 30249
rect 137702 12409 137793 12527
rect 137911 12409 138002 12527
rect 137702 12367 138002 12409
rect 137702 12249 137793 12367
rect 137911 12249 138002 12367
rect 137702 -1583 138002 12249
rect 137702 -1701 137793 -1583
rect 137911 -1701 138002 -1583
rect 137702 -1743 138002 -1701
rect 137702 -1861 137793 -1743
rect 137911 -1861 138002 -1743
rect 137702 -1872 138002 -1861
rect 139502 338327 139802 354491
rect 139502 338209 139593 338327
rect 139711 338209 139802 338327
rect 139502 338167 139802 338209
rect 139502 338049 139593 338167
rect 139711 338049 139802 338167
rect 139502 320327 139802 338049
rect 139502 320209 139593 320327
rect 139711 320209 139802 320327
rect 139502 320167 139802 320209
rect 139502 320049 139593 320167
rect 139711 320049 139802 320167
rect 139502 302327 139802 320049
rect 139502 302209 139593 302327
rect 139711 302209 139802 302327
rect 139502 302167 139802 302209
rect 139502 302049 139593 302167
rect 139711 302049 139802 302167
rect 139502 284327 139802 302049
rect 139502 284209 139593 284327
rect 139711 284209 139802 284327
rect 139502 284167 139802 284209
rect 139502 284049 139593 284167
rect 139711 284049 139802 284167
rect 139502 266327 139802 284049
rect 139502 266209 139593 266327
rect 139711 266209 139802 266327
rect 139502 266167 139802 266209
rect 139502 266049 139593 266167
rect 139711 266049 139802 266167
rect 139502 248327 139802 266049
rect 139502 248209 139593 248327
rect 139711 248209 139802 248327
rect 139502 248167 139802 248209
rect 139502 248049 139593 248167
rect 139711 248049 139802 248167
rect 139502 230327 139802 248049
rect 139502 230209 139593 230327
rect 139711 230209 139802 230327
rect 139502 230167 139802 230209
rect 139502 230049 139593 230167
rect 139711 230049 139802 230167
rect 139502 212327 139802 230049
rect 139502 212209 139593 212327
rect 139711 212209 139802 212327
rect 139502 212167 139802 212209
rect 139502 212049 139593 212167
rect 139711 212049 139802 212167
rect 139502 194327 139802 212049
rect 139502 194209 139593 194327
rect 139711 194209 139802 194327
rect 139502 194167 139802 194209
rect 139502 194049 139593 194167
rect 139711 194049 139802 194167
rect 139502 176327 139802 194049
rect 139502 176209 139593 176327
rect 139711 176209 139802 176327
rect 139502 176167 139802 176209
rect 139502 176049 139593 176167
rect 139711 176049 139802 176167
rect 139502 158327 139802 176049
rect 139502 158209 139593 158327
rect 139711 158209 139802 158327
rect 139502 158167 139802 158209
rect 139502 158049 139593 158167
rect 139711 158049 139802 158167
rect 139502 140327 139802 158049
rect 139502 140209 139593 140327
rect 139711 140209 139802 140327
rect 139502 140167 139802 140209
rect 139502 140049 139593 140167
rect 139711 140049 139802 140167
rect 139502 122327 139802 140049
rect 139502 122209 139593 122327
rect 139711 122209 139802 122327
rect 139502 122167 139802 122209
rect 139502 122049 139593 122167
rect 139711 122049 139802 122167
rect 139502 104327 139802 122049
rect 139502 104209 139593 104327
rect 139711 104209 139802 104327
rect 139502 104167 139802 104209
rect 139502 104049 139593 104167
rect 139711 104049 139802 104167
rect 139502 86327 139802 104049
rect 139502 86209 139593 86327
rect 139711 86209 139802 86327
rect 139502 86167 139802 86209
rect 139502 86049 139593 86167
rect 139711 86049 139802 86167
rect 139502 68327 139802 86049
rect 139502 68209 139593 68327
rect 139711 68209 139802 68327
rect 139502 68167 139802 68209
rect 139502 68049 139593 68167
rect 139711 68049 139802 68167
rect 139502 50327 139802 68049
rect 139502 50209 139593 50327
rect 139711 50209 139802 50327
rect 139502 50167 139802 50209
rect 139502 50049 139593 50167
rect 139711 50049 139802 50167
rect 139502 32327 139802 50049
rect 139502 32209 139593 32327
rect 139711 32209 139802 32327
rect 139502 32167 139802 32209
rect 139502 32049 139593 32167
rect 139711 32049 139802 32167
rect 139502 14327 139802 32049
rect 139502 14209 139593 14327
rect 139711 14209 139802 14327
rect 139502 14167 139802 14209
rect 139502 14049 139593 14167
rect 139711 14049 139802 14167
rect 139502 -2523 139802 14049
rect 139502 -2641 139593 -2523
rect 139711 -2641 139802 -2523
rect 139502 -2683 139802 -2641
rect 139502 -2801 139593 -2683
rect 139711 -2801 139802 -2683
rect 139502 -2812 139802 -2801
rect 141302 340127 141602 355431
rect 150302 355239 150602 355720
rect 150302 355121 150393 355239
rect 150511 355121 150602 355239
rect 150302 355079 150602 355121
rect 150302 354961 150393 355079
rect 150511 354961 150602 355079
rect 148502 354299 148802 354780
rect 148502 354181 148593 354299
rect 148711 354181 148802 354299
rect 148502 354139 148802 354181
rect 148502 354021 148593 354139
rect 148711 354021 148802 354139
rect 146702 353359 147002 353840
rect 146702 353241 146793 353359
rect 146911 353241 147002 353359
rect 146702 353199 147002 353241
rect 146702 353081 146793 353199
rect 146911 353081 147002 353199
rect 141302 340009 141393 340127
rect 141511 340009 141602 340127
rect 141302 339967 141602 340009
rect 141302 339849 141393 339967
rect 141511 339849 141602 339967
rect 141302 322127 141602 339849
rect 141302 322009 141393 322127
rect 141511 322009 141602 322127
rect 141302 321967 141602 322009
rect 141302 321849 141393 321967
rect 141511 321849 141602 321967
rect 141302 304127 141602 321849
rect 141302 304009 141393 304127
rect 141511 304009 141602 304127
rect 141302 303967 141602 304009
rect 141302 303849 141393 303967
rect 141511 303849 141602 303967
rect 141302 286127 141602 303849
rect 141302 286009 141393 286127
rect 141511 286009 141602 286127
rect 141302 285967 141602 286009
rect 141302 285849 141393 285967
rect 141511 285849 141602 285967
rect 141302 268127 141602 285849
rect 141302 268009 141393 268127
rect 141511 268009 141602 268127
rect 141302 267967 141602 268009
rect 141302 267849 141393 267967
rect 141511 267849 141602 267967
rect 141302 250127 141602 267849
rect 141302 250009 141393 250127
rect 141511 250009 141602 250127
rect 141302 249967 141602 250009
rect 141302 249849 141393 249967
rect 141511 249849 141602 249967
rect 141302 232127 141602 249849
rect 141302 232009 141393 232127
rect 141511 232009 141602 232127
rect 141302 231967 141602 232009
rect 141302 231849 141393 231967
rect 141511 231849 141602 231967
rect 141302 214127 141602 231849
rect 141302 214009 141393 214127
rect 141511 214009 141602 214127
rect 141302 213967 141602 214009
rect 141302 213849 141393 213967
rect 141511 213849 141602 213967
rect 141302 196127 141602 213849
rect 141302 196009 141393 196127
rect 141511 196009 141602 196127
rect 141302 195967 141602 196009
rect 141302 195849 141393 195967
rect 141511 195849 141602 195967
rect 141302 178127 141602 195849
rect 141302 178009 141393 178127
rect 141511 178009 141602 178127
rect 141302 177967 141602 178009
rect 141302 177849 141393 177967
rect 141511 177849 141602 177967
rect 141302 160127 141602 177849
rect 141302 160009 141393 160127
rect 141511 160009 141602 160127
rect 141302 159967 141602 160009
rect 141302 159849 141393 159967
rect 141511 159849 141602 159967
rect 141302 142127 141602 159849
rect 141302 142009 141393 142127
rect 141511 142009 141602 142127
rect 141302 141967 141602 142009
rect 141302 141849 141393 141967
rect 141511 141849 141602 141967
rect 141302 124127 141602 141849
rect 141302 124009 141393 124127
rect 141511 124009 141602 124127
rect 141302 123967 141602 124009
rect 141302 123849 141393 123967
rect 141511 123849 141602 123967
rect 141302 106127 141602 123849
rect 141302 106009 141393 106127
rect 141511 106009 141602 106127
rect 141302 105967 141602 106009
rect 141302 105849 141393 105967
rect 141511 105849 141602 105967
rect 141302 88127 141602 105849
rect 141302 88009 141393 88127
rect 141511 88009 141602 88127
rect 141302 87967 141602 88009
rect 141302 87849 141393 87967
rect 141511 87849 141602 87967
rect 141302 70127 141602 87849
rect 141302 70009 141393 70127
rect 141511 70009 141602 70127
rect 141302 69967 141602 70009
rect 141302 69849 141393 69967
rect 141511 69849 141602 69967
rect 141302 52127 141602 69849
rect 141302 52009 141393 52127
rect 141511 52009 141602 52127
rect 141302 51967 141602 52009
rect 141302 51849 141393 51967
rect 141511 51849 141602 51967
rect 141302 34127 141602 51849
rect 141302 34009 141393 34127
rect 141511 34009 141602 34127
rect 141302 33967 141602 34009
rect 141302 33849 141393 33967
rect 141511 33849 141602 33967
rect 141302 16127 141602 33849
rect 141302 16009 141393 16127
rect 141511 16009 141602 16127
rect 141302 15967 141602 16009
rect 141302 15849 141393 15967
rect 141511 15849 141602 15967
rect 132302 -3111 132393 -2993
rect 132511 -3111 132602 -2993
rect 132302 -3153 132602 -3111
rect 132302 -3271 132393 -3153
rect 132511 -3271 132602 -3153
rect 132302 -3752 132602 -3271
rect 141302 -3463 141602 15849
rect 144902 352419 145202 352900
rect 144902 352301 144993 352419
rect 145111 352301 145202 352419
rect 144902 352259 145202 352301
rect 144902 352141 144993 352259
rect 145111 352141 145202 352259
rect 144902 343727 145202 352141
rect 144902 343609 144993 343727
rect 145111 343609 145202 343727
rect 144902 343567 145202 343609
rect 144902 343449 144993 343567
rect 145111 343449 145202 343567
rect 144902 325727 145202 343449
rect 144902 325609 144993 325727
rect 145111 325609 145202 325727
rect 144902 325567 145202 325609
rect 144902 325449 144993 325567
rect 145111 325449 145202 325567
rect 144902 307727 145202 325449
rect 144902 307609 144993 307727
rect 145111 307609 145202 307727
rect 144902 307567 145202 307609
rect 144902 307449 144993 307567
rect 145111 307449 145202 307567
rect 144902 289727 145202 307449
rect 144902 289609 144993 289727
rect 145111 289609 145202 289727
rect 144902 289567 145202 289609
rect 144902 289449 144993 289567
rect 145111 289449 145202 289567
rect 144902 271727 145202 289449
rect 144902 271609 144993 271727
rect 145111 271609 145202 271727
rect 144902 271567 145202 271609
rect 144902 271449 144993 271567
rect 145111 271449 145202 271567
rect 144902 253727 145202 271449
rect 144902 253609 144993 253727
rect 145111 253609 145202 253727
rect 144902 253567 145202 253609
rect 144902 253449 144993 253567
rect 145111 253449 145202 253567
rect 144902 235727 145202 253449
rect 144902 235609 144993 235727
rect 145111 235609 145202 235727
rect 144902 235567 145202 235609
rect 144902 235449 144993 235567
rect 145111 235449 145202 235567
rect 144902 217727 145202 235449
rect 144902 217609 144993 217727
rect 145111 217609 145202 217727
rect 144902 217567 145202 217609
rect 144902 217449 144993 217567
rect 145111 217449 145202 217567
rect 144902 199727 145202 217449
rect 144902 199609 144993 199727
rect 145111 199609 145202 199727
rect 144902 199567 145202 199609
rect 144902 199449 144993 199567
rect 145111 199449 145202 199567
rect 144902 181727 145202 199449
rect 144902 181609 144993 181727
rect 145111 181609 145202 181727
rect 144902 181567 145202 181609
rect 144902 181449 144993 181567
rect 145111 181449 145202 181567
rect 144902 163727 145202 181449
rect 144902 163609 144993 163727
rect 145111 163609 145202 163727
rect 144902 163567 145202 163609
rect 144902 163449 144993 163567
rect 145111 163449 145202 163567
rect 144902 145727 145202 163449
rect 144902 145609 144993 145727
rect 145111 145609 145202 145727
rect 144902 145567 145202 145609
rect 144902 145449 144993 145567
rect 145111 145449 145202 145567
rect 144902 127727 145202 145449
rect 144902 127609 144993 127727
rect 145111 127609 145202 127727
rect 144902 127567 145202 127609
rect 144902 127449 144993 127567
rect 145111 127449 145202 127567
rect 144902 109727 145202 127449
rect 144902 109609 144993 109727
rect 145111 109609 145202 109727
rect 144902 109567 145202 109609
rect 144902 109449 144993 109567
rect 145111 109449 145202 109567
rect 144902 91727 145202 109449
rect 144902 91609 144993 91727
rect 145111 91609 145202 91727
rect 144902 91567 145202 91609
rect 144902 91449 144993 91567
rect 145111 91449 145202 91567
rect 144902 73727 145202 91449
rect 144902 73609 144993 73727
rect 145111 73609 145202 73727
rect 144902 73567 145202 73609
rect 144902 73449 144993 73567
rect 145111 73449 145202 73567
rect 144902 55727 145202 73449
rect 144902 55609 144993 55727
rect 145111 55609 145202 55727
rect 144902 55567 145202 55609
rect 144902 55449 144993 55567
rect 145111 55449 145202 55567
rect 144902 37727 145202 55449
rect 144902 37609 144993 37727
rect 145111 37609 145202 37727
rect 144902 37567 145202 37609
rect 144902 37449 144993 37567
rect 145111 37449 145202 37567
rect 144902 19727 145202 37449
rect 144902 19609 144993 19727
rect 145111 19609 145202 19727
rect 144902 19567 145202 19609
rect 144902 19449 144993 19567
rect 145111 19449 145202 19567
rect 144902 1727 145202 19449
rect 144902 1609 144993 1727
rect 145111 1609 145202 1727
rect 144902 1567 145202 1609
rect 144902 1449 144993 1567
rect 145111 1449 145202 1567
rect 144902 -173 145202 1449
rect 144902 -291 144993 -173
rect 145111 -291 145202 -173
rect 144902 -333 145202 -291
rect 144902 -451 144993 -333
rect 145111 -451 145202 -333
rect 144902 -932 145202 -451
rect 146702 345527 147002 353081
rect 146702 345409 146793 345527
rect 146911 345409 147002 345527
rect 146702 345367 147002 345409
rect 146702 345249 146793 345367
rect 146911 345249 147002 345367
rect 146702 327527 147002 345249
rect 146702 327409 146793 327527
rect 146911 327409 147002 327527
rect 146702 327367 147002 327409
rect 146702 327249 146793 327367
rect 146911 327249 147002 327367
rect 146702 309527 147002 327249
rect 146702 309409 146793 309527
rect 146911 309409 147002 309527
rect 146702 309367 147002 309409
rect 146702 309249 146793 309367
rect 146911 309249 147002 309367
rect 146702 291527 147002 309249
rect 146702 291409 146793 291527
rect 146911 291409 147002 291527
rect 146702 291367 147002 291409
rect 146702 291249 146793 291367
rect 146911 291249 147002 291367
rect 146702 273527 147002 291249
rect 146702 273409 146793 273527
rect 146911 273409 147002 273527
rect 146702 273367 147002 273409
rect 146702 273249 146793 273367
rect 146911 273249 147002 273367
rect 146702 255527 147002 273249
rect 146702 255409 146793 255527
rect 146911 255409 147002 255527
rect 146702 255367 147002 255409
rect 146702 255249 146793 255367
rect 146911 255249 147002 255367
rect 146702 237527 147002 255249
rect 146702 237409 146793 237527
rect 146911 237409 147002 237527
rect 146702 237367 147002 237409
rect 146702 237249 146793 237367
rect 146911 237249 147002 237367
rect 146702 219527 147002 237249
rect 146702 219409 146793 219527
rect 146911 219409 147002 219527
rect 146702 219367 147002 219409
rect 146702 219249 146793 219367
rect 146911 219249 147002 219367
rect 146702 201527 147002 219249
rect 146702 201409 146793 201527
rect 146911 201409 147002 201527
rect 146702 201367 147002 201409
rect 146702 201249 146793 201367
rect 146911 201249 147002 201367
rect 146702 183527 147002 201249
rect 146702 183409 146793 183527
rect 146911 183409 147002 183527
rect 146702 183367 147002 183409
rect 146702 183249 146793 183367
rect 146911 183249 147002 183367
rect 146702 165527 147002 183249
rect 146702 165409 146793 165527
rect 146911 165409 147002 165527
rect 146702 165367 147002 165409
rect 146702 165249 146793 165367
rect 146911 165249 147002 165367
rect 146702 147527 147002 165249
rect 146702 147409 146793 147527
rect 146911 147409 147002 147527
rect 146702 147367 147002 147409
rect 146702 147249 146793 147367
rect 146911 147249 147002 147367
rect 146702 129527 147002 147249
rect 146702 129409 146793 129527
rect 146911 129409 147002 129527
rect 146702 129367 147002 129409
rect 146702 129249 146793 129367
rect 146911 129249 147002 129367
rect 146702 111527 147002 129249
rect 146702 111409 146793 111527
rect 146911 111409 147002 111527
rect 146702 111367 147002 111409
rect 146702 111249 146793 111367
rect 146911 111249 147002 111367
rect 146702 93527 147002 111249
rect 146702 93409 146793 93527
rect 146911 93409 147002 93527
rect 146702 93367 147002 93409
rect 146702 93249 146793 93367
rect 146911 93249 147002 93367
rect 146702 75527 147002 93249
rect 146702 75409 146793 75527
rect 146911 75409 147002 75527
rect 146702 75367 147002 75409
rect 146702 75249 146793 75367
rect 146911 75249 147002 75367
rect 146702 57527 147002 75249
rect 146702 57409 146793 57527
rect 146911 57409 147002 57527
rect 146702 57367 147002 57409
rect 146702 57249 146793 57367
rect 146911 57249 147002 57367
rect 146702 39527 147002 57249
rect 146702 39409 146793 39527
rect 146911 39409 147002 39527
rect 146702 39367 147002 39409
rect 146702 39249 146793 39367
rect 146911 39249 147002 39367
rect 146702 21527 147002 39249
rect 146702 21409 146793 21527
rect 146911 21409 147002 21527
rect 146702 21367 147002 21409
rect 146702 21249 146793 21367
rect 146911 21249 147002 21367
rect 146702 3527 147002 21249
rect 146702 3409 146793 3527
rect 146911 3409 147002 3527
rect 146702 3367 147002 3409
rect 146702 3249 146793 3367
rect 146911 3249 147002 3367
rect 146702 -1113 147002 3249
rect 146702 -1231 146793 -1113
rect 146911 -1231 147002 -1113
rect 146702 -1273 147002 -1231
rect 146702 -1391 146793 -1273
rect 146911 -1391 147002 -1273
rect 146702 -1872 147002 -1391
rect 148502 347327 148802 354021
rect 148502 347209 148593 347327
rect 148711 347209 148802 347327
rect 148502 347167 148802 347209
rect 148502 347049 148593 347167
rect 148711 347049 148802 347167
rect 148502 329327 148802 347049
rect 148502 329209 148593 329327
rect 148711 329209 148802 329327
rect 148502 329167 148802 329209
rect 148502 329049 148593 329167
rect 148711 329049 148802 329167
rect 148502 311327 148802 329049
rect 148502 311209 148593 311327
rect 148711 311209 148802 311327
rect 148502 311167 148802 311209
rect 148502 311049 148593 311167
rect 148711 311049 148802 311167
rect 148502 293327 148802 311049
rect 148502 293209 148593 293327
rect 148711 293209 148802 293327
rect 148502 293167 148802 293209
rect 148502 293049 148593 293167
rect 148711 293049 148802 293167
rect 148502 275327 148802 293049
rect 148502 275209 148593 275327
rect 148711 275209 148802 275327
rect 148502 275167 148802 275209
rect 148502 275049 148593 275167
rect 148711 275049 148802 275167
rect 148502 257327 148802 275049
rect 148502 257209 148593 257327
rect 148711 257209 148802 257327
rect 148502 257167 148802 257209
rect 148502 257049 148593 257167
rect 148711 257049 148802 257167
rect 148502 239327 148802 257049
rect 148502 239209 148593 239327
rect 148711 239209 148802 239327
rect 148502 239167 148802 239209
rect 148502 239049 148593 239167
rect 148711 239049 148802 239167
rect 148502 221327 148802 239049
rect 148502 221209 148593 221327
rect 148711 221209 148802 221327
rect 148502 221167 148802 221209
rect 148502 221049 148593 221167
rect 148711 221049 148802 221167
rect 148502 203327 148802 221049
rect 148502 203209 148593 203327
rect 148711 203209 148802 203327
rect 148502 203167 148802 203209
rect 148502 203049 148593 203167
rect 148711 203049 148802 203167
rect 148502 185327 148802 203049
rect 148502 185209 148593 185327
rect 148711 185209 148802 185327
rect 148502 185167 148802 185209
rect 148502 185049 148593 185167
rect 148711 185049 148802 185167
rect 148502 167327 148802 185049
rect 148502 167209 148593 167327
rect 148711 167209 148802 167327
rect 148502 167167 148802 167209
rect 148502 167049 148593 167167
rect 148711 167049 148802 167167
rect 148502 149327 148802 167049
rect 148502 149209 148593 149327
rect 148711 149209 148802 149327
rect 148502 149167 148802 149209
rect 148502 149049 148593 149167
rect 148711 149049 148802 149167
rect 148502 131327 148802 149049
rect 148502 131209 148593 131327
rect 148711 131209 148802 131327
rect 148502 131167 148802 131209
rect 148502 131049 148593 131167
rect 148711 131049 148802 131167
rect 148502 113327 148802 131049
rect 148502 113209 148593 113327
rect 148711 113209 148802 113327
rect 148502 113167 148802 113209
rect 148502 113049 148593 113167
rect 148711 113049 148802 113167
rect 148502 95327 148802 113049
rect 148502 95209 148593 95327
rect 148711 95209 148802 95327
rect 148502 95167 148802 95209
rect 148502 95049 148593 95167
rect 148711 95049 148802 95167
rect 148502 77327 148802 95049
rect 148502 77209 148593 77327
rect 148711 77209 148802 77327
rect 148502 77167 148802 77209
rect 148502 77049 148593 77167
rect 148711 77049 148802 77167
rect 148502 59327 148802 77049
rect 148502 59209 148593 59327
rect 148711 59209 148802 59327
rect 148502 59167 148802 59209
rect 148502 59049 148593 59167
rect 148711 59049 148802 59167
rect 148502 41327 148802 59049
rect 148502 41209 148593 41327
rect 148711 41209 148802 41327
rect 148502 41167 148802 41209
rect 148502 41049 148593 41167
rect 148711 41049 148802 41167
rect 148502 23327 148802 41049
rect 148502 23209 148593 23327
rect 148711 23209 148802 23327
rect 148502 23167 148802 23209
rect 148502 23049 148593 23167
rect 148711 23049 148802 23167
rect 148502 5327 148802 23049
rect 148502 5209 148593 5327
rect 148711 5209 148802 5327
rect 148502 5167 148802 5209
rect 148502 5049 148593 5167
rect 148711 5049 148802 5167
rect 148502 -2053 148802 5049
rect 148502 -2171 148593 -2053
rect 148711 -2171 148802 -2053
rect 148502 -2213 148802 -2171
rect 148502 -2331 148593 -2213
rect 148711 -2331 148802 -2213
rect 148502 -2812 148802 -2331
rect 150302 349127 150602 354961
rect 159302 355709 159602 355720
rect 159302 355591 159393 355709
rect 159511 355591 159602 355709
rect 159302 355549 159602 355591
rect 159302 355431 159393 355549
rect 159511 355431 159602 355549
rect 157502 354769 157802 354780
rect 157502 354651 157593 354769
rect 157711 354651 157802 354769
rect 157502 354609 157802 354651
rect 157502 354491 157593 354609
rect 157711 354491 157802 354609
rect 155702 353829 156002 353840
rect 155702 353711 155793 353829
rect 155911 353711 156002 353829
rect 155702 353669 156002 353711
rect 155702 353551 155793 353669
rect 155911 353551 156002 353669
rect 150302 349009 150393 349127
rect 150511 349009 150602 349127
rect 150302 348967 150602 349009
rect 150302 348849 150393 348967
rect 150511 348849 150602 348967
rect 150302 331127 150602 348849
rect 150302 331009 150393 331127
rect 150511 331009 150602 331127
rect 150302 330967 150602 331009
rect 150302 330849 150393 330967
rect 150511 330849 150602 330967
rect 150302 313127 150602 330849
rect 150302 313009 150393 313127
rect 150511 313009 150602 313127
rect 150302 312967 150602 313009
rect 150302 312849 150393 312967
rect 150511 312849 150602 312967
rect 150302 295127 150602 312849
rect 150302 295009 150393 295127
rect 150511 295009 150602 295127
rect 150302 294967 150602 295009
rect 150302 294849 150393 294967
rect 150511 294849 150602 294967
rect 150302 277127 150602 294849
rect 150302 277009 150393 277127
rect 150511 277009 150602 277127
rect 150302 276967 150602 277009
rect 150302 276849 150393 276967
rect 150511 276849 150602 276967
rect 150302 259127 150602 276849
rect 150302 259009 150393 259127
rect 150511 259009 150602 259127
rect 150302 258967 150602 259009
rect 150302 258849 150393 258967
rect 150511 258849 150602 258967
rect 150302 241127 150602 258849
rect 150302 241009 150393 241127
rect 150511 241009 150602 241127
rect 150302 240967 150602 241009
rect 150302 240849 150393 240967
rect 150511 240849 150602 240967
rect 150302 223127 150602 240849
rect 150302 223009 150393 223127
rect 150511 223009 150602 223127
rect 150302 222967 150602 223009
rect 150302 222849 150393 222967
rect 150511 222849 150602 222967
rect 150302 205127 150602 222849
rect 150302 205009 150393 205127
rect 150511 205009 150602 205127
rect 150302 204967 150602 205009
rect 150302 204849 150393 204967
rect 150511 204849 150602 204967
rect 150302 187127 150602 204849
rect 150302 187009 150393 187127
rect 150511 187009 150602 187127
rect 150302 186967 150602 187009
rect 150302 186849 150393 186967
rect 150511 186849 150602 186967
rect 150302 169127 150602 186849
rect 150302 169009 150393 169127
rect 150511 169009 150602 169127
rect 150302 168967 150602 169009
rect 150302 168849 150393 168967
rect 150511 168849 150602 168967
rect 150302 151127 150602 168849
rect 150302 151009 150393 151127
rect 150511 151009 150602 151127
rect 150302 150967 150602 151009
rect 150302 150849 150393 150967
rect 150511 150849 150602 150967
rect 150302 133127 150602 150849
rect 150302 133009 150393 133127
rect 150511 133009 150602 133127
rect 150302 132967 150602 133009
rect 150302 132849 150393 132967
rect 150511 132849 150602 132967
rect 150302 115127 150602 132849
rect 150302 115009 150393 115127
rect 150511 115009 150602 115127
rect 150302 114967 150602 115009
rect 150302 114849 150393 114967
rect 150511 114849 150602 114967
rect 150302 97127 150602 114849
rect 150302 97009 150393 97127
rect 150511 97009 150602 97127
rect 150302 96967 150602 97009
rect 150302 96849 150393 96967
rect 150511 96849 150602 96967
rect 150302 79127 150602 96849
rect 150302 79009 150393 79127
rect 150511 79009 150602 79127
rect 150302 78967 150602 79009
rect 150302 78849 150393 78967
rect 150511 78849 150602 78967
rect 150302 61127 150602 78849
rect 150302 61009 150393 61127
rect 150511 61009 150602 61127
rect 150302 60967 150602 61009
rect 150302 60849 150393 60967
rect 150511 60849 150602 60967
rect 150302 43127 150602 60849
rect 150302 43009 150393 43127
rect 150511 43009 150602 43127
rect 150302 42967 150602 43009
rect 150302 42849 150393 42967
rect 150511 42849 150602 42967
rect 150302 25127 150602 42849
rect 150302 25009 150393 25127
rect 150511 25009 150602 25127
rect 150302 24967 150602 25009
rect 150302 24849 150393 24967
rect 150511 24849 150602 24967
rect 150302 7127 150602 24849
rect 150302 7009 150393 7127
rect 150511 7009 150602 7127
rect 150302 6967 150602 7009
rect 150302 6849 150393 6967
rect 150511 6849 150602 6967
rect 141302 -3581 141393 -3463
rect 141511 -3581 141602 -3463
rect 141302 -3623 141602 -3581
rect 141302 -3741 141393 -3623
rect 141511 -3741 141602 -3623
rect 141302 -3752 141602 -3741
rect 150302 -2993 150602 6849
rect 153902 352889 154202 352900
rect 153902 352771 153993 352889
rect 154111 352771 154202 352889
rect 153902 352729 154202 352771
rect 153902 352611 153993 352729
rect 154111 352611 154202 352729
rect 153902 334727 154202 352611
rect 153902 334609 153993 334727
rect 154111 334609 154202 334727
rect 153902 334567 154202 334609
rect 153902 334449 153993 334567
rect 154111 334449 154202 334567
rect 153902 316727 154202 334449
rect 153902 316609 153993 316727
rect 154111 316609 154202 316727
rect 153902 316567 154202 316609
rect 153902 316449 153993 316567
rect 154111 316449 154202 316567
rect 153902 298727 154202 316449
rect 153902 298609 153993 298727
rect 154111 298609 154202 298727
rect 153902 298567 154202 298609
rect 153902 298449 153993 298567
rect 154111 298449 154202 298567
rect 153902 280727 154202 298449
rect 153902 280609 153993 280727
rect 154111 280609 154202 280727
rect 153902 280567 154202 280609
rect 153902 280449 153993 280567
rect 154111 280449 154202 280567
rect 153902 262727 154202 280449
rect 153902 262609 153993 262727
rect 154111 262609 154202 262727
rect 153902 262567 154202 262609
rect 153902 262449 153993 262567
rect 154111 262449 154202 262567
rect 153902 244727 154202 262449
rect 153902 244609 153993 244727
rect 154111 244609 154202 244727
rect 153902 244567 154202 244609
rect 153902 244449 153993 244567
rect 154111 244449 154202 244567
rect 153902 226727 154202 244449
rect 153902 226609 153993 226727
rect 154111 226609 154202 226727
rect 153902 226567 154202 226609
rect 153902 226449 153993 226567
rect 154111 226449 154202 226567
rect 153902 208727 154202 226449
rect 153902 208609 153993 208727
rect 154111 208609 154202 208727
rect 153902 208567 154202 208609
rect 153902 208449 153993 208567
rect 154111 208449 154202 208567
rect 153902 190727 154202 208449
rect 153902 190609 153993 190727
rect 154111 190609 154202 190727
rect 153902 190567 154202 190609
rect 153902 190449 153993 190567
rect 154111 190449 154202 190567
rect 153902 172727 154202 190449
rect 153902 172609 153993 172727
rect 154111 172609 154202 172727
rect 153902 172567 154202 172609
rect 153902 172449 153993 172567
rect 154111 172449 154202 172567
rect 153902 154727 154202 172449
rect 153902 154609 153993 154727
rect 154111 154609 154202 154727
rect 153902 154567 154202 154609
rect 153902 154449 153993 154567
rect 154111 154449 154202 154567
rect 153902 136727 154202 154449
rect 153902 136609 153993 136727
rect 154111 136609 154202 136727
rect 153902 136567 154202 136609
rect 153902 136449 153993 136567
rect 154111 136449 154202 136567
rect 153902 118727 154202 136449
rect 153902 118609 153993 118727
rect 154111 118609 154202 118727
rect 153902 118567 154202 118609
rect 153902 118449 153993 118567
rect 154111 118449 154202 118567
rect 153902 100727 154202 118449
rect 153902 100609 153993 100727
rect 154111 100609 154202 100727
rect 153902 100567 154202 100609
rect 153902 100449 153993 100567
rect 154111 100449 154202 100567
rect 153902 82727 154202 100449
rect 153902 82609 153993 82727
rect 154111 82609 154202 82727
rect 153902 82567 154202 82609
rect 153902 82449 153993 82567
rect 154111 82449 154202 82567
rect 153902 64727 154202 82449
rect 153902 64609 153993 64727
rect 154111 64609 154202 64727
rect 153902 64567 154202 64609
rect 153902 64449 153993 64567
rect 154111 64449 154202 64567
rect 153902 46727 154202 64449
rect 153902 46609 153993 46727
rect 154111 46609 154202 46727
rect 153902 46567 154202 46609
rect 153902 46449 153993 46567
rect 154111 46449 154202 46567
rect 153902 28727 154202 46449
rect 153902 28609 153993 28727
rect 154111 28609 154202 28727
rect 153902 28567 154202 28609
rect 153902 28449 153993 28567
rect 154111 28449 154202 28567
rect 153902 10727 154202 28449
rect 153902 10609 153993 10727
rect 154111 10609 154202 10727
rect 153902 10567 154202 10609
rect 153902 10449 153993 10567
rect 154111 10449 154202 10567
rect 153902 -643 154202 10449
rect 153902 -761 153993 -643
rect 154111 -761 154202 -643
rect 153902 -803 154202 -761
rect 153902 -921 153993 -803
rect 154111 -921 154202 -803
rect 153902 -932 154202 -921
rect 155702 336527 156002 353551
rect 155702 336409 155793 336527
rect 155911 336409 156002 336527
rect 155702 336367 156002 336409
rect 155702 336249 155793 336367
rect 155911 336249 156002 336367
rect 155702 318527 156002 336249
rect 155702 318409 155793 318527
rect 155911 318409 156002 318527
rect 155702 318367 156002 318409
rect 155702 318249 155793 318367
rect 155911 318249 156002 318367
rect 155702 300527 156002 318249
rect 155702 300409 155793 300527
rect 155911 300409 156002 300527
rect 155702 300367 156002 300409
rect 155702 300249 155793 300367
rect 155911 300249 156002 300367
rect 155702 282527 156002 300249
rect 155702 282409 155793 282527
rect 155911 282409 156002 282527
rect 155702 282367 156002 282409
rect 155702 282249 155793 282367
rect 155911 282249 156002 282367
rect 155702 264527 156002 282249
rect 155702 264409 155793 264527
rect 155911 264409 156002 264527
rect 155702 264367 156002 264409
rect 155702 264249 155793 264367
rect 155911 264249 156002 264367
rect 155702 246527 156002 264249
rect 155702 246409 155793 246527
rect 155911 246409 156002 246527
rect 155702 246367 156002 246409
rect 155702 246249 155793 246367
rect 155911 246249 156002 246367
rect 155702 228527 156002 246249
rect 155702 228409 155793 228527
rect 155911 228409 156002 228527
rect 155702 228367 156002 228409
rect 155702 228249 155793 228367
rect 155911 228249 156002 228367
rect 155702 210527 156002 228249
rect 155702 210409 155793 210527
rect 155911 210409 156002 210527
rect 155702 210367 156002 210409
rect 155702 210249 155793 210367
rect 155911 210249 156002 210367
rect 155702 192527 156002 210249
rect 155702 192409 155793 192527
rect 155911 192409 156002 192527
rect 155702 192367 156002 192409
rect 155702 192249 155793 192367
rect 155911 192249 156002 192367
rect 155702 174527 156002 192249
rect 155702 174409 155793 174527
rect 155911 174409 156002 174527
rect 155702 174367 156002 174409
rect 155702 174249 155793 174367
rect 155911 174249 156002 174367
rect 155702 156527 156002 174249
rect 155702 156409 155793 156527
rect 155911 156409 156002 156527
rect 155702 156367 156002 156409
rect 155702 156249 155793 156367
rect 155911 156249 156002 156367
rect 155702 138527 156002 156249
rect 155702 138409 155793 138527
rect 155911 138409 156002 138527
rect 155702 138367 156002 138409
rect 155702 138249 155793 138367
rect 155911 138249 156002 138367
rect 155702 120527 156002 138249
rect 155702 120409 155793 120527
rect 155911 120409 156002 120527
rect 155702 120367 156002 120409
rect 155702 120249 155793 120367
rect 155911 120249 156002 120367
rect 155702 102527 156002 120249
rect 155702 102409 155793 102527
rect 155911 102409 156002 102527
rect 155702 102367 156002 102409
rect 155702 102249 155793 102367
rect 155911 102249 156002 102367
rect 155702 84527 156002 102249
rect 155702 84409 155793 84527
rect 155911 84409 156002 84527
rect 155702 84367 156002 84409
rect 155702 84249 155793 84367
rect 155911 84249 156002 84367
rect 155702 66527 156002 84249
rect 155702 66409 155793 66527
rect 155911 66409 156002 66527
rect 155702 66367 156002 66409
rect 155702 66249 155793 66367
rect 155911 66249 156002 66367
rect 155702 48527 156002 66249
rect 155702 48409 155793 48527
rect 155911 48409 156002 48527
rect 155702 48367 156002 48409
rect 155702 48249 155793 48367
rect 155911 48249 156002 48367
rect 155702 30527 156002 48249
rect 155702 30409 155793 30527
rect 155911 30409 156002 30527
rect 155702 30367 156002 30409
rect 155702 30249 155793 30367
rect 155911 30249 156002 30367
rect 155702 12527 156002 30249
rect 155702 12409 155793 12527
rect 155911 12409 156002 12527
rect 155702 12367 156002 12409
rect 155702 12249 155793 12367
rect 155911 12249 156002 12367
rect 155702 -1583 156002 12249
rect 155702 -1701 155793 -1583
rect 155911 -1701 156002 -1583
rect 155702 -1743 156002 -1701
rect 155702 -1861 155793 -1743
rect 155911 -1861 156002 -1743
rect 155702 -1872 156002 -1861
rect 157502 338327 157802 354491
rect 157502 338209 157593 338327
rect 157711 338209 157802 338327
rect 157502 338167 157802 338209
rect 157502 338049 157593 338167
rect 157711 338049 157802 338167
rect 157502 320327 157802 338049
rect 157502 320209 157593 320327
rect 157711 320209 157802 320327
rect 157502 320167 157802 320209
rect 157502 320049 157593 320167
rect 157711 320049 157802 320167
rect 157502 302327 157802 320049
rect 157502 302209 157593 302327
rect 157711 302209 157802 302327
rect 157502 302167 157802 302209
rect 157502 302049 157593 302167
rect 157711 302049 157802 302167
rect 157502 284327 157802 302049
rect 157502 284209 157593 284327
rect 157711 284209 157802 284327
rect 157502 284167 157802 284209
rect 157502 284049 157593 284167
rect 157711 284049 157802 284167
rect 157502 266327 157802 284049
rect 157502 266209 157593 266327
rect 157711 266209 157802 266327
rect 157502 266167 157802 266209
rect 157502 266049 157593 266167
rect 157711 266049 157802 266167
rect 157502 248327 157802 266049
rect 157502 248209 157593 248327
rect 157711 248209 157802 248327
rect 157502 248167 157802 248209
rect 157502 248049 157593 248167
rect 157711 248049 157802 248167
rect 157502 230327 157802 248049
rect 157502 230209 157593 230327
rect 157711 230209 157802 230327
rect 157502 230167 157802 230209
rect 157502 230049 157593 230167
rect 157711 230049 157802 230167
rect 157502 212327 157802 230049
rect 157502 212209 157593 212327
rect 157711 212209 157802 212327
rect 157502 212167 157802 212209
rect 157502 212049 157593 212167
rect 157711 212049 157802 212167
rect 157502 194327 157802 212049
rect 157502 194209 157593 194327
rect 157711 194209 157802 194327
rect 157502 194167 157802 194209
rect 157502 194049 157593 194167
rect 157711 194049 157802 194167
rect 157502 176327 157802 194049
rect 157502 176209 157593 176327
rect 157711 176209 157802 176327
rect 157502 176167 157802 176209
rect 157502 176049 157593 176167
rect 157711 176049 157802 176167
rect 157502 158327 157802 176049
rect 157502 158209 157593 158327
rect 157711 158209 157802 158327
rect 157502 158167 157802 158209
rect 157502 158049 157593 158167
rect 157711 158049 157802 158167
rect 157502 140327 157802 158049
rect 157502 140209 157593 140327
rect 157711 140209 157802 140327
rect 157502 140167 157802 140209
rect 157502 140049 157593 140167
rect 157711 140049 157802 140167
rect 157502 122327 157802 140049
rect 157502 122209 157593 122327
rect 157711 122209 157802 122327
rect 157502 122167 157802 122209
rect 157502 122049 157593 122167
rect 157711 122049 157802 122167
rect 157502 104327 157802 122049
rect 157502 104209 157593 104327
rect 157711 104209 157802 104327
rect 157502 104167 157802 104209
rect 157502 104049 157593 104167
rect 157711 104049 157802 104167
rect 157502 86327 157802 104049
rect 157502 86209 157593 86327
rect 157711 86209 157802 86327
rect 157502 86167 157802 86209
rect 157502 86049 157593 86167
rect 157711 86049 157802 86167
rect 157502 68327 157802 86049
rect 157502 68209 157593 68327
rect 157711 68209 157802 68327
rect 157502 68167 157802 68209
rect 157502 68049 157593 68167
rect 157711 68049 157802 68167
rect 157502 50327 157802 68049
rect 157502 50209 157593 50327
rect 157711 50209 157802 50327
rect 157502 50167 157802 50209
rect 157502 50049 157593 50167
rect 157711 50049 157802 50167
rect 157502 32327 157802 50049
rect 157502 32209 157593 32327
rect 157711 32209 157802 32327
rect 157502 32167 157802 32209
rect 157502 32049 157593 32167
rect 157711 32049 157802 32167
rect 157502 14327 157802 32049
rect 157502 14209 157593 14327
rect 157711 14209 157802 14327
rect 157502 14167 157802 14209
rect 157502 14049 157593 14167
rect 157711 14049 157802 14167
rect 157502 -2523 157802 14049
rect 157502 -2641 157593 -2523
rect 157711 -2641 157802 -2523
rect 157502 -2683 157802 -2641
rect 157502 -2801 157593 -2683
rect 157711 -2801 157802 -2683
rect 157502 -2812 157802 -2801
rect 159302 340127 159602 355431
rect 168302 355239 168602 355720
rect 168302 355121 168393 355239
rect 168511 355121 168602 355239
rect 168302 355079 168602 355121
rect 168302 354961 168393 355079
rect 168511 354961 168602 355079
rect 166502 354299 166802 354780
rect 166502 354181 166593 354299
rect 166711 354181 166802 354299
rect 166502 354139 166802 354181
rect 166502 354021 166593 354139
rect 166711 354021 166802 354139
rect 164702 353359 165002 353840
rect 164702 353241 164793 353359
rect 164911 353241 165002 353359
rect 164702 353199 165002 353241
rect 164702 353081 164793 353199
rect 164911 353081 165002 353199
rect 159302 340009 159393 340127
rect 159511 340009 159602 340127
rect 159302 339967 159602 340009
rect 159302 339849 159393 339967
rect 159511 339849 159602 339967
rect 159302 322127 159602 339849
rect 159302 322009 159393 322127
rect 159511 322009 159602 322127
rect 159302 321967 159602 322009
rect 159302 321849 159393 321967
rect 159511 321849 159602 321967
rect 159302 304127 159602 321849
rect 159302 304009 159393 304127
rect 159511 304009 159602 304127
rect 159302 303967 159602 304009
rect 159302 303849 159393 303967
rect 159511 303849 159602 303967
rect 159302 286127 159602 303849
rect 159302 286009 159393 286127
rect 159511 286009 159602 286127
rect 159302 285967 159602 286009
rect 159302 285849 159393 285967
rect 159511 285849 159602 285967
rect 159302 268127 159602 285849
rect 159302 268009 159393 268127
rect 159511 268009 159602 268127
rect 159302 267967 159602 268009
rect 159302 267849 159393 267967
rect 159511 267849 159602 267967
rect 159302 250127 159602 267849
rect 159302 250009 159393 250127
rect 159511 250009 159602 250127
rect 159302 249967 159602 250009
rect 159302 249849 159393 249967
rect 159511 249849 159602 249967
rect 159302 232127 159602 249849
rect 159302 232009 159393 232127
rect 159511 232009 159602 232127
rect 159302 231967 159602 232009
rect 159302 231849 159393 231967
rect 159511 231849 159602 231967
rect 159302 214127 159602 231849
rect 159302 214009 159393 214127
rect 159511 214009 159602 214127
rect 159302 213967 159602 214009
rect 159302 213849 159393 213967
rect 159511 213849 159602 213967
rect 159302 196127 159602 213849
rect 159302 196009 159393 196127
rect 159511 196009 159602 196127
rect 159302 195967 159602 196009
rect 159302 195849 159393 195967
rect 159511 195849 159602 195967
rect 159302 178127 159602 195849
rect 159302 178009 159393 178127
rect 159511 178009 159602 178127
rect 159302 177967 159602 178009
rect 159302 177849 159393 177967
rect 159511 177849 159602 177967
rect 159302 160127 159602 177849
rect 159302 160009 159393 160127
rect 159511 160009 159602 160127
rect 159302 159967 159602 160009
rect 159302 159849 159393 159967
rect 159511 159849 159602 159967
rect 159302 142127 159602 159849
rect 159302 142009 159393 142127
rect 159511 142009 159602 142127
rect 159302 141967 159602 142009
rect 159302 141849 159393 141967
rect 159511 141849 159602 141967
rect 159302 124127 159602 141849
rect 159302 124009 159393 124127
rect 159511 124009 159602 124127
rect 159302 123967 159602 124009
rect 159302 123849 159393 123967
rect 159511 123849 159602 123967
rect 159302 106127 159602 123849
rect 159302 106009 159393 106127
rect 159511 106009 159602 106127
rect 159302 105967 159602 106009
rect 159302 105849 159393 105967
rect 159511 105849 159602 105967
rect 159302 88127 159602 105849
rect 159302 88009 159393 88127
rect 159511 88009 159602 88127
rect 159302 87967 159602 88009
rect 159302 87849 159393 87967
rect 159511 87849 159602 87967
rect 159302 70127 159602 87849
rect 159302 70009 159393 70127
rect 159511 70009 159602 70127
rect 159302 69967 159602 70009
rect 159302 69849 159393 69967
rect 159511 69849 159602 69967
rect 159302 52127 159602 69849
rect 159302 52009 159393 52127
rect 159511 52009 159602 52127
rect 159302 51967 159602 52009
rect 159302 51849 159393 51967
rect 159511 51849 159602 51967
rect 159302 34127 159602 51849
rect 159302 34009 159393 34127
rect 159511 34009 159602 34127
rect 159302 33967 159602 34009
rect 159302 33849 159393 33967
rect 159511 33849 159602 33967
rect 159302 16127 159602 33849
rect 159302 16009 159393 16127
rect 159511 16009 159602 16127
rect 159302 15967 159602 16009
rect 159302 15849 159393 15967
rect 159511 15849 159602 15967
rect 150302 -3111 150393 -2993
rect 150511 -3111 150602 -2993
rect 150302 -3153 150602 -3111
rect 150302 -3271 150393 -3153
rect 150511 -3271 150602 -3153
rect 150302 -3752 150602 -3271
rect 159302 -3463 159602 15849
rect 162902 352419 163202 352900
rect 162902 352301 162993 352419
rect 163111 352301 163202 352419
rect 162902 352259 163202 352301
rect 162902 352141 162993 352259
rect 163111 352141 163202 352259
rect 162902 343727 163202 352141
rect 162902 343609 162993 343727
rect 163111 343609 163202 343727
rect 162902 343567 163202 343609
rect 162902 343449 162993 343567
rect 163111 343449 163202 343567
rect 162902 325727 163202 343449
rect 162902 325609 162993 325727
rect 163111 325609 163202 325727
rect 162902 325567 163202 325609
rect 162902 325449 162993 325567
rect 163111 325449 163202 325567
rect 162902 307727 163202 325449
rect 162902 307609 162993 307727
rect 163111 307609 163202 307727
rect 162902 307567 163202 307609
rect 162902 307449 162993 307567
rect 163111 307449 163202 307567
rect 162902 289727 163202 307449
rect 162902 289609 162993 289727
rect 163111 289609 163202 289727
rect 162902 289567 163202 289609
rect 162902 289449 162993 289567
rect 163111 289449 163202 289567
rect 162902 271727 163202 289449
rect 162902 271609 162993 271727
rect 163111 271609 163202 271727
rect 162902 271567 163202 271609
rect 162902 271449 162993 271567
rect 163111 271449 163202 271567
rect 162902 253727 163202 271449
rect 162902 253609 162993 253727
rect 163111 253609 163202 253727
rect 162902 253567 163202 253609
rect 162902 253449 162993 253567
rect 163111 253449 163202 253567
rect 162902 235727 163202 253449
rect 162902 235609 162993 235727
rect 163111 235609 163202 235727
rect 162902 235567 163202 235609
rect 162902 235449 162993 235567
rect 163111 235449 163202 235567
rect 162902 217727 163202 235449
rect 162902 217609 162993 217727
rect 163111 217609 163202 217727
rect 162902 217567 163202 217609
rect 162902 217449 162993 217567
rect 163111 217449 163202 217567
rect 162902 199727 163202 217449
rect 162902 199609 162993 199727
rect 163111 199609 163202 199727
rect 162902 199567 163202 199609
rect 162902 199449 162993 199567
rect 163111 199449 163202 199567
rect 162902 181727 163202 199449
rect 162902 181609 162993 181727
rect 163111 181609 163202 181727
rect 162902 181567 163202 181609
rect 162902 181449 162993 181567
rect 163111 181449 163202 181567
rect 162902 163727 163202 181449
rect 162902 163609 162993 163727
rect 163111 163609 163202 163727
rect 162902 163567 163202 163609
rect 162902 163449 162993 163567
rect 163111 163449 163202 163567
rect 162902 145727 163202 163449
rect 162902 145609 162993 145727
rect 163111 145609 163202 145727
rect 162902 145567 163202 145609
rect 162902 145449 162993 145567
rect 163111 145449 163202 145567
rect 162902 127727 163202 145449
rect 162902 127609 162993 127727
rect 163111 127609 163202 127727
rect 162902 127567 163202 127609
rect 162902 127449 162993 127567
rect 163111 127449 163202 127567
rect 162902 109727 163202 127449
rect 162902 109609 162993 109727
rect 163111 109609 163202 109727
rect 162902 109567 163202 109609
rect 162902 109449 162993 109567
rect 163111 109449 163202 109567
rect 162902 91727 163202 109449
rect 162902 91609 162993 91727
rect 163111 91609 163202 91727
rect 162902 91567 163202 91609
rect 162902 91449 162993 91567
rect 163111 91449 163202 91567
rect 162902 73727 163202 91449
rect 162902 73609 162993 73727
rect 163111 73609 163202 73727
rect 162902 73567 163202 73609
rect 162902 73449 162993 73567
rect 163111 73449 163202 73567
rect 162902 55727 163202 73449
rect 162902 55609 162993 55727
rect 163111 55609 163202 55727
rect 162902 55567 163202 55609
rect 162902 55449 162993 55567
rect 163111 55449 163202 55567
rect 162902 37727 163202 55449
rect 162902 37609 162993 37727
rect 163111 37609 163202 37727
rect 162902 37567 163202 37609
rect 162902 37449 162993 37567
rect 163111 37449 163202 37567
rect 162902 19727 163202 37449
rect 162902 19609 162993 19727
rect 163111 19609 163202 19727
rect 162902 19567 163202 19609
rect 162902 19449 162993 19567
rect 163111 19449 163202 19567
rect 162902 1727 163202 19449
rect 162902 1609 162993 1727
rect 163111 1609 163202 1727
rect 162902 1567 163202 1609
rect 162902 1449 162993 1567
rect 163111 1449 163202 1567
rect 162902 -173 163202 1449
rect 162902 -291 162993 -173
rect 163111 -291 163202 -173
rect 162902 -333 163202 -291
rect 162902 -451 162993 -333
rect 163111 -451 163202 -333
rect 162902 -932 163202 -451
rect 164702 345527 165002 353081
rect 164702 345409 164793 345527
rect 164911 345409 165002 345527
rect 164702 345367 165002 345409
rect 164702 345249 164793 345367
rect 164911 345249 165002 345367
rect 164702 327527 165002 345249
rect 164702 327409 164793 327527
rect 164911 327409 165002 327527
rect 164702 327367 165002 327409
rect 164702 327249 164793 327367
rect 164911 327249 165002 327367
rect 164702 309527 165002 327249
rect 164702 309409 164793 309527
rect 164911 309409 165002 309527
rect 164702 309367 165002 309409
rect 164702 309249 164793 309367
rect 164911 309249 165002 309367
rect 164702 291527 165002 309249
rect 164702 291409 164793 291527
rect 164911 291409 165002 291527
rect 164702 291367 165002 291409
rect 164702 291249 164793 291367
rect 164911 291249 165002 291367
rect 164702 273527 165002 291249
rect 164702 273409 164793 273527
rect 164911 273409 165002 273527
rect 164702 273367 165002 273409
rect 164702 273249 164793 273367
rect 164911 273249 165002 273367
rect 164702 255527 165002 273249
rect 164702 255409 164793 255527
rect 164911 255409 165002 255527
rect 164702 255367 165002 255409
rect 164702 255249 164793 255367
rect 164911 255249 165002 255367
rect 164702 237527 165002 255249
rect 164702 237409 164793 237527
rect 164911 237409 165002 237527
rect 164702 237367 165002 237409
rect 164702 237249 164793 237367
rect 164911 237249 165002 237367
rect 164702 219527 165002 237249
rect 164702 219409 164793 219527
rect 164911 219409 165002 219527
rect 164702 219367 165002 219409
rect 164702 219249 164793 219367
rect 164911 219249 165002 219367
rect 164702 201527 165002 219249
rect 164702 201409 164793 201527
rect 164911 201409 165002 201527
rect 164702 201367 165002 201409
rect 164702 201249 164793 201367
rect 164911 201249 165002 201367
rect 164702 183527 165002 201249
rect 164702 183409 164793 183527
rect 164911 183409 165002 183527
rect 164702 183367 165002 183409
rect 164702 183249 164793 183367
rect 164911 183249 165002 183367
rect 164702 165527 165002 183249
rect 164702 165409 164793 165527
rect 164911 165409 165002 165527
rect 164702 165367 165002 165409
rect 164702 165249 164793 165367
rect 164911 165249 165002 165367
rect 164702 147527 165002 165249
rect 164702 147409 164793 147527
rect 164911 147409 165002 147527
rect 164702 147367 165002 147409
rect 164702 147249 164793 147367
rect 164911 147249 165002 147367
rect 164702 129527 165002 147249
rect 164702 129409 164793 129527
rect 164911 129409 165002 129527
rect 164702 129367 165002 129409
rect 164702 129249 164793 129367
rect 164911 129249 165002 129367
rect 164702 111527 165002 129249
rect 164702 111409 164793 111527
rect 164911 111409 165002 111527
rect 164702 111367 165002 111409
rect 164702 111249 164793 111367
rect 164911 111249 165002 111367
rect 164702 93527 165002 111249
rect 164702 93409 164793 93527
rect 164911 93409 165002 93527
rect 164702 93367 165002 93409
rect 164702 93249 164793 93367
rect 164911 93249 165002 93367
rect 164702 75527 165002 93249
rect 164702 75409 164793 75527
rect 164911 75409 165002 75527
rect 164702 75367 165002 75409
rect 164702 75249 164793 75367
rect 164911 75249 165002 75367
rect 164702 57527 165002 75249
rect 164702 57409 164793 57527
rect 164911 57409 165002 57527
rect 164702 57367 165002 57409
rect 164702 57249 164793 57367
rect 164911 57249 165002 57367
rect 164702 39527 165002 57249
rect 164702 39409 164793 39527
rect 164911 39409 165002 39527
rect 164702 39367 165002 39409
rect 164702 39249 164793 39367
rect 164911 39249 165002 39367
rect 164702 21527 165002 39249
rect 164702 21409 164793 21527
rect 164911 21409 165002 21527
rect 164702 21367 165002 21409
rect 164702 21249 164793 21367
rect 164911 21249 165002 21367
rect 164702 3527 165002 21249
rect 164702 3409 164793 3527
rect 164911 3409 165002 3527
rect 164702 3367 165002 3409
rect 164702 3249 164793 3367
rect 164911 3249 165002 3367
rect 164702 -1113 165002 3249
rect 164702 -1231 164793 -1113
rect 164911 -1231 165002 -1113
rect 164702 -1273 165002 -1231
rect 164702 -1391 164793 -1273
rect 164911 -1391 165002 -1273
rect 164702 -1872 165002 -1391
rect 166502 347327 166802 354021
rect 166502 347209 166593 347327
rect 166711 347209 166802 347327
rect 166502 347167 166802 347209
rect 166502 347049 166593 347167
rect 166711 347049 166802 347167
rect 166502 329327 166802 347049
rect 166502 329209 166593 329327
rect 166711 329209 166802 329327
rect 166502 329167 166802 329209
rect 166502 329049 166593 329167
rect 166711 329049 166802 329167
rect 166502 311327 166802 329049
rect 166502 311209 166593 311327
rect 166711 311209 166802 311327
rect 166502 311167 166802 311209
rect 166502 311049 166593 311167
rect 166711 311049 166802 311167
rect 166502 293327 166802 311049
rect 166502 293209 166593 293327
rect 166711 293209 166802 293327
rect 166502 293167 166802 293209
rect 166502 293049 166593 293167
rect 166711 293049 166802 293167
rect 166502 275327 166802 293049
rect 166502 275209 166593 275327
rect 166711 275209 166802 275327
rect 166502 275167 166802 275209
rect 166502 275049 166593 275167
rect 166711 275049 166802 275167
rect 166502 257327 166802 275049
rect 166502 257209 166593 257327
rect 166711 257209 166802 257327
rect 166502 257167 166802 257209
rect 166502 257049 166593 257167
rect 166711 257049 166802 257167
rect 166502 239327 166802 257049
rect 166502 239209 166593 239327
rect 166711 239209 166802 239327
rect 166502 239167 166802 239209
rect 166502 239049 166593 239167
rect 166711 239049 166802 239167
rect 166502 221327 166802 239049
rect 166502 221209 166593 221327
rect 166711 221209 166802 221327
rect 166502 221167 166802 221209
rect 166502 221049 166593 221167
rect 166711 221049 166802 221167
rect 166502 203327 166802 221049
rect 166502 203209 166593 203327
rect 166711 203209 166802 203327
rect 166502 203167 166802 203209
rect 166502 203049 166593 203167
rect 166711 203049 166802 203167
rect 166502 185327 166802 203049
rect 166502 185209 166593 185327
rect 166711 185209 166802 185327
rect 166502 185167 166802 185209
rect 166502 185049 166593 185167
rect 166711 185049 166802 185167
rect 166502 167327 166802 185049
rect 166502 167209 166593 167327
rect 166711 167209 166802 167327
rect 166502 167167 166802 167209
rect 166502 167049 166593 167167
rect 166711 167049 166802 167167
rect 166502 149327 166802 167049
rect 166502 149209 166593 149327
rect 166711 149209 166802 149327
rect 166502 149167 166802 149209
rect 166502 149049 166593 149167
rect 166711 149049 166802 149167
rect 166502 131327 166802 149049
rect 166502 131209 166593 131327
rect 166711 131209 166802 131327
rect 166502 131167 166802 131209
rect 166502 131049 166593 131167
rect 166711 131049 166802 131167
rect 166502 113327 166802 131049
rect 166502 113209 166593 113327
rect 166711 113209 166802 113327
rect 166502 113167 166802 113209
rect 166502 113049 166593 113167
rect 166711 113049 166802 113167
rect 166502 95327 166802 113049
rect 166502 95209 166593 95327
rect 166711 95209 166802 95327
rect 166502 95167 166802 95209
rect 166502 95049 166593 95167
rect 166711 95049 166802 95167
rect 166502 77327 166802 95049
rect 166502 77209 166593 77327
rect 166711 77209 166802 77327
rect 166502 77167 166802 77209
rect 166502 77049 166593 77167
rect 166711 77049 166802 77167
rect 166502 59327 166802 77049
rect 166502 59209 166593 59327
rect 166711 59209 166802 59327
rect 166502 59167 166802 59209
rect 166502 59049 166593 59167
rect 166711 59049 166802 59167
rect 166502 41327 166802 59049
rect 166502 41209 166593 41327
rect 166711 41209 166802 41327
rect 166502 41167 166802 41209
rect 166502 41049 166593 41167
rect 166711 41049 166802 41167
rect 166502 23327 166802 41049
rect 166502 23209 166593 23327
rect 166711 23209 166802 23327
rect 166502 23167 166802 23209
rect 166502 23049 166593 23167
rect 166711 23049 166802 23167
rect 166502 5327 166802 23049
rect 166502 5209 166593 5327
rect 166711 5209 166802 5327
rect 166502 5167 166802 5209
rect 166502 5049 166593 5167
rect 166711 5049 166802 5167
rect 166502 -2053 166802 5049
rect 166502 -2171 166593 -2053
rect 166711 -2171 166802 -2053
rect 166502 -2213 166802 -2171
rect 166502 -2331 166593 -2213
rect 166711 -2331 166802 -2213
rect 166502 -2812 166802 -2331
rect 168302 349127 168602 354961
rect 177302 355709 177602 355720
rect 177302 355591 177393 355709
rect 177511 355591 177602 355709
rect 177302 355549 177602 355591
rect 177302 355431 177393 355549
rect 177511 355431 177602 355549
rect 175502 354769 175802 354780
rect 175502 354651 175593 354769
rect 175711 354651 175802 354769
rect 175502 354609 175802 354651
rect 175502 354491 175593 354609
rect 175711 354491 175802 354609
rect 173702 353829 174002 353840
rect 173702 353711 173793 353829
rect 173911 353711 174002 353829
rect 173702 353669 174002 353711
rect 173702 353551 173793 353669
rect 173911 353551 174002 353669
rect 168302 349009 168393 349127
rect 168511 349009 168602 349127
rect 168302 348967 168602 349009
rect 168302 348849 168393 348967
rect 168511 348849 168602 348967
rect 168302 331127 168602 348849
rect 168302 331009 168393 331127
rect 168511 331009 168602 331127
rect 168302 330967 168602 331009
rect 168302 330849 168393 330967
rect 168511 330849 168602 330967
rect 168302 313127 168602 330849
rect 168302 313009 168393 313127
rect 168511 313009 168602 313127
rect 168302 312967 168602 313009
rect 168302 312849 168393 312967
rect 168511 312849 168602 312967
rect 168302 295127 168602 312849
rect 168302 295009 168393 295127
rect 168511 295009 168602 295127
rect 168302 294967 168602 295009
rect 168302 294849 168393 294967
rect 168511 294849 168602 294967
rect 168302 277127 168602 294849
rect 168302 277009 168393 277127
rect 168511 277009 168602 277127
rect 168302 276967 168602 277009
rect 168302 276849 168393 276967
rect 168511 276849 168602 276967
rect 168302 259127 168602 276849
rect 168302 259009 168393 259127
rect 168511 259009 168602 259127
rect 168302 258967 168602 259009
rect 168302 258849 168393 258967
rect 168511 258849 168602 258967
rect 168302 241127 168602 258849
rect 168302 241009 168393 241127
rect 168511 241009 168602 241127
rect 168302 240967 168602 241009
rect 168302 240849 168393 240967
rect 168511 240849 168602 240967
rect 168302 223127 168602 240849
rect 168302 223009 168393 223127
rect 168511 223009 168602 223127
rect 168302 222967 168602 223009
rect 168302 222849 168393 222967
rect 168511 222849 168602 222967
rect 168302 205127 168602 222849
rect 168302 205009 168393 205127
rect 168511 205009 168602 205127
rect 168302 204967 168602 205009
rect 168302 204849 168393 204967
rect 168511 204849 168602 204967
rect 168302 187127 168602 204849
rect 168302 187009 168393 187127
rect 168511 187009 168602 187127
rect 168302 186967 168602 187009
rect 168302 186849 168393 186967
rect 168511 186849 168602 186967
rect 168302 169127 168602 186849
rect 168302 169009 168393 169127
rect 168511 169009 168602 169127
rect 168302 168967 168602 169009
rect 168302 168849 168393 168967
rect 168511 168849 168602 168967
rect 168302 151127 168602 168849
rect 168302 151009 168393 151127
rect 168511 151009 168602 151127
rect 168302 150967 168602 151009
rect 168302 150849 168393 150967
rect 168511 150849 168602 150967
rect 168302 133127 168602 150849
rect 168302 133009 168393 133127
rect 168511 133009 168602 133127
rect 168302 132967 168602 133009
rect 168302 132849 168393 132967
rect 168511 132849 168602 132967
rect 168302 115127 168602 132849
rect 168302 115009 168393 115127
rect 168511 115009 168602 115127
rect 168302 114967 168602 115009
rect 168302 114849 168393 114967
rect 168511 114849 168602 114967
rect 168302 97127 168602 114849
rect 168302 97009 168393 97127
rect 168511 97009 168602 97127
rect 168302 96967 168602 97009
rect 168302 96849 168393 96967
rect 168511 96849 168602 96967
rect 168302 79127 168602 96849
rect 168302 79009 168393 79127
rect 168511 79009 168602 79127
rect 168302 78967 168602 79009
rect 168302 78849 168393 78967
rect 168511 78849 168602 78967
rect 168302 61127 168602 78849
rect 168302 61009 168393 61127
rect 168511 61009 168602 61127
rect 168302 60967 168602 61009
rect 168302 60849 168393 60967
rect 168511 60849 168602 60967
rect 168302 43127 168602 60849
rect 168302 43009 168393 43127
rect 168511 43009 168602 43127
rect 168302 42967 168602 43009
rect 168302 42849 168393 42967
rect 168511 42849 168602 42967
rect 168302 25127 168602 42849
rect 168302 25009 168393 25127
rect 168511 25009 168602 25127
rect 168302 24967 168602 25009
rect 168302 24849 168393 24967
rect 168511 24849 168602 24967
rect 168302 7127 168602 24849
rect 168302 7009 168393 7127
rect 168511 7009 168602 7127
rect 168302 6967 168602 7009
rect 168302 6849 168393 6967
rect 168511 6849 168602 6967
rect 159302 -3581 159393 -3463
rect 159511 -3581 159602 -3463
rect 159302 -3623 159602 -3581
rect 159302 -3741 159393 -3623
rect 159511 -3741 159602 -3623
rect 159302 -3752 159602 -3741
rect 168302 -2993 168602 6849
rect 171902 352889 172202 352900
rect 171902 352771 171993 352889
rect 172111 352771 172202 352889
rect 171902 352729 172202 352771
rect 171902 352611 171993 352729
rect 172111 352611 172202 352729
rect 171902 334727 172202 352611
rect 171902 334609 171993 334727
rect 172111 334609 172202 334727
rect 171902 334567 172202 334609
rect 171902 334449 171993 334567
rect 172111 334449 172202 334567
rect 171902 316727 172202 334449
rect 171902 316609 171993 316727
rect 172111 316609 172202 316727
rect 171902 316567 172202 316609
rect 171902 316449 171993 316567
rect 172111 316449 172202 316567
rect 171902 298727 172202 316449
rect 171902 298609 171993 298727
rect 172111 298609 172202 298727
rect 171902 298567 172202 298609
rect 171902 298449 171993 298567
rect 172111 298449 172202 298567
rect 171902 280727 172202 298449
rect 171902 280609 171993 280727
rect 172111 280609 172202 280727
rect 171902 280567 172202 280609
rect 171902 280449 171993 280567
rect 172111 280449 172202 280567
rect 171902 262727 172202 280449
rect 171902 262609 171993 262727
rect 172111 262609 172202 262727
rect 171902 262567 172202 262609
rect 171902 262449 171993 262567
rect 172111 262449 172202 262567
rect 171902 244727 172202 262449
rect 171902 244609 171993 244727
rect 172111 244609 172202 244727
rect 171902 244567 172202 244609
rect 171902 244449 171993 244567
rect 172111 244449 172202 244567
rect 171902 226727 172202 244449
rect 171902 226609 171993 226727
rect 172111 226609 172202 226727
rect 171902 226567 172202 226609
rect 171902 226449 171993 226567
rect 172111 226449 172202 226567
rect 171902 208727 172202 226449
rect 171902 208609 171993 208727
rect 172111 208609 172202 208727
rect 171902 208567 172202 208609
rect 171902 208449 171993 208567
rect 172111 208449 172202 208567
rect 171902 190727 172202 208449
rect 171902 190609 171993 190727
rect 172111 190609 172202 190727
rect 171902 190567 172202 190609
rect 171902 190449 171993 190567
rect 172111 190449 172202 190567
rect 171902 172727 172202 190449
rect 171902 172609 171993 172727
rect 172111 172609 172202 172727
rect 171902 172567 172202 172609
rect 171902 172449 171993 172567
rect 172111 172449 172202 172567
rect 171902 154727 172202 172449
rect 171902 154609 171993 154727
rect 172111 154609 172202 154727
rect 171902 154567 172202 154609
rect 171902 154449 171993 154567
rect 172111 154449 172202 154567
rect 171902 136727 172202 154449
rect 171902 136609 171993 136727
rect 172111 136609 172202 136727
rect 171902 136567 172202 136609
rect 171902 136449 171993 136567
rect 172111 136449 172202 136567
rect 171902 118727 172202 136449
rect 171902 118609 171993 118727
rect 172111 118609 172202 118727
rect 171902 118567 172202 118609
rect 171902 118449 171993 118567
rect 172111 118449 172202 118567
rect 171902 100727 172202 118449
rect 171902 100609 171993 100727
rect 172111 100609 172202 100727
rect 171902 100567 172202 100609
rect 171902 100449 171993 100567
rect 172111 100449 172202 100567
rect 171902 82727 172202 100449
rect 171902 82609 171993 82727
rect 172111 82609 172202 82727
rect 171902 82567 172202 82609
rect 171902 82449 171993 82567
rect 172111 82449 172202 82567
rect 171902 64727 172202 82449
rect 171902 64609 171993 64727
rect 172111 64609 172202 64727
rect 171902 64567 172202 64609
rect 171902 64449 171993 64567
rect 172111 64449 172202 64567
rect 171902 46727 172202 64449
rect 171902 46609 171993 46727
rect 172111 46609 172202 46727
rect 171902 46567 172202 46609
rect 171902 46449 171993 46567
rect 172111 46449 172202 46567
rect 171902 28727 172202 46449
rect 171902 28609 171993 28727
rect 172111 28609 172202 28727
rect 171902 28567 172202 28609
rect 171902 28449 171993 28567
rect 172111 28449 172202 28567
rect 171902 10727 172202 28449
rect 171902 10609 171993 10727
rect 172111 10609 172202 10727
rect 171902 10567 172202 10609
rect 171902 10449 171993 10567
rect 172111 10449 172202 10567
rect 171902 -643 172202 10449
rect 171902 -761 171993 -643
rect 172111 -761 172202 -643
rect 171902 -803 172202 -761
rect 171902 -921 171993 -803
rect 172111 -921 172202 -803
rect 171902 -932 172202 -921
rect 173702 336527 174002 353551
rect 173702 336409 173793 336527
rect 173911 336409 174002 336527
rect 173702 336367 174002 336409
rect 173702 336249 173793 336367
rect 173911 336249 174002 336367
rect 173702 318527 174002 336249
rect 173702 318409 173793 318527
rect 173911 318409 174002 318527
rect 173702 318367 174002 318409
rect 173702 318249 173793 318367
rect 173911 318249 174002 318367
rect 173702 300527 174002 318249
rect 173702 300409 173793 300527
rect 173911 300409 174002 300527
rect 173702 300367 174002 300409
rect 173702 300249 173793 300367
rect 173911 300249 174002 300367
rect 173702 282527 174002 300249
rect 173702 282409 173793 282527
rect 173911 282409 174002 282527
rect 173702 282367 174002 282409
rect 173702 282249 173793 282367
rect 173911 282249 174002 282367
rect 173702 264527 174002 282249
rect 173702 264409 173793 264527
rect 173911 264409 174002 264527
rect 173702 264367 174002 264409
rect 173702 264249 173793 264367
rect 173911 264249 174002 264367
rect 173702 246527 174002 264249
rect 173702 246409 173793 246527
rect 173911 246409 174002 246527
rect 173702 246367 174002 246409
rect 173702 246249 173793 246367
rect 173911 246249 174002 246367
rect 173702 228527 174002 246249
rect 173702 228409 173793 228527
rect 173911 228409 174002 228527
rect 173702 228367 174002 228409
rect 173702 228249 173793 228367
rect 173911 228249 174002 228367
rect 173702 210527 174002 228249
rect 173702 210409 173793 210527
rect 173911 210409 174002 210527
rect 173702 210367 174002 210409
rect 173702 210249 173793 210367
rect 173911 210249 174002 210367
rect 173702 192527 174002 210249
rect 173702 192409 173793 192527
rect 173911 192409 174002 192527
rect 173702 192367 174002 192409
rect 173702 192249 173793 192367
rect 173911 192249 174002 192367
rect 173702 174527 174002 192249
rect 173702 174409 173793 174527
rect 173911 174409 174002 174527
rect 173702 174367 174002 174409
rect 173702 174249 173793 174367
rect 173911 174249 174002 174367
rect 173702 156527 174002 174249
rect 173702 156409 173793 156527
rect 173911 156409 174002 156527
rect 173702 156367 174002 156409
rect 173702 156249 173793 156367
rect 173911 156249 174002 156367
rect 173702 138527 174002 156249
rect 173702 138409 173793 138527
rect 173911 138409 174002 138527
rect 173702 138367 174002 138409
rect 173702 138249 173793 138367
rect 173911 138249 174002 138367
rect 173702 120527 174002 138249
rect 173702 120409 173793 120527
rect 173911 120409 174002 120527
rect 173702 120367 174002 120409
rect 173702 120249 173793 120367
rect 173911 120249 174002 120367
rect 173702 102527 174002 120249
rect 173702 102409 173793 102527
rect 173911 102409 174002 102527
rect 173702 102367 174002 102409
rect 173702 102249 173793 102367
rect 173911 102249 174002 102367
rect 173702 84527 174002 102249
rect 173702 84409 173793 84527
rect 173911 84409 174002 84527
rect 173702 84367 174002 84409
rect 173702 84249 173793 84367
rect 173911 84249 174002 84367
rect 173702 66527 174002 84249
rect 173702 66409 173793 66527
rect 173911 66409 174002 66527
rect 173702 66367 174002 66409
rect 173702 66249 173793 66367
rect 173911 66249 174002 66367
rect 173702 48527 174002 66249
rect 173702 48409 173793 48527
rect 173911 48409 174002 48527
rect 173702 48367 174002 48409
rect 173702 48249 173793 48367
rect 173911 48249 174002 48367
rect 173702 30527 174002 48249
rect 173702 30409 173793 30527
rect 173911 30409 174002 30527
rect 173702 30367 174002 30409
rect 173702 30249 173793 30367
rect 173911 30249 174002 30367
rect 173702 12527 174002 30249
rect 173702 12409 173793 12527
rect 173911 12409 174002 12527
rect 173702 12367 174002 12409
rect 173702 12249 173793 12367
rect 173911 12249 174002 12367
rect 173702 -1583 174002 12249
rect 173702 -1701 173793 -1583
rect 173911 -1701 174002 -1583
rect 173702 -1743 174002 -1701
rect 173702 -1861 173793 -1743
rect 173911 -1861 174002 -1743
rect 173702 -1872 174002 -1861
rect 175502 338327 175802 354491
rect 175502 338209 175593 338327
rect 175711 338209 175802 338327
rect 175502 338167 175802 338209
rect 175502 338049 175593 338167
rect 175711 338049 175802 338167
rect 175502 320327 175802 338049
rect 175502 320209 175593 320327
rect 175711 320209 175802 320327
rect 175502 320167 175802 320209
rect 175502 320049 175593 320167
rect 175711 320049 175802 320167
rect 175502 302327 175802 320049
rect 175502 302209 175593 302327
rect 175711 302209 175802 302327
rect 175502 302167 175802 302209
rect 175502 302049 175593 302167
rect 175711 302049 175802 302167
rect 175502 284327 175802 302049
rect 175502 284209 175593 284327
rect 175711 284209 175802 284327
rect 175502 284167 175802 284209
rect 175502 284049 175593 284167
rect 175711 284049 175802 284167
rect 175502 266327 175802 284049
rect 175502 266209 175593 266327
rect 175711 266209 175802 266327
rect 175502 266167 175802 266209
rect 175502 266049 175593 266167
rect 175711 266049 175802 266167
rect 175502 248327 175802 266049
rect 175502 248209 175593 248327
rect 175711 248209 175802 248327
rect 175502 248167 175802 248209
rect 175502 248049 175593 248167
rect 175711 248049 175802 248167
rect 175502 230327 175802 248049
rect 175502 230209 175593 230327
rect 175711 230209 175802 230327
rect 175502 230167 175802 230209
rect 175502 230049 175593 230167
rect 175711 230049 175802 230167
rect 175502 212327 175802 230049
rect 175502 212209 175593 212327
rect 175711 212209 175802 212327
rect 175502 212167 175802 212209
rect 175502 212049 175593 212167
rect 175711 212049 175802 212167
rect 175502 194327 175802 212049
rect 175502 194209 175593 194327
rect 175711 194209 175802 194327
rect 175502 194167 175802 194209
rect 175502 194049 175593 194167
rect 175711 194049 175802 194167
rect 175502 176327 175802 194049
rect 175502 176209 175593 176327
rect 175711 176209 175802 176327
rect 175502 176167 175802 176209
rect 175502 176049 175593 176167
rect 175711 176049 175802 176167
rect 175502 158327 175802 176049
rect 175502 158209 175593 158327
rect 175711 158209 175802 158327
rect 175502 158167 175802 158209
rect 175502 158049 175593 158167
rect 175711 158049 175802 158167
rect 175502 140327 175802 158049
rect 175502 140209 175593 140327
rect 175711 140209 175802 140327
rect 175502 140167 175802 140209
rect 175502 140049 175593 140167
rect 175711 140049 175802 140167
rect 175502 122327 175802 140049
rect 175502 122209 175593 122327
rect 175711 122209 175802 122327
rect 175502 122167 175802 122209
rect 175502 122049 175593 122167
rect 175711 122049 175802 122167
rect 175502 104327 175802 122049
rect 175502 104209 175593 104327
rect 175711 104209 175802 104327
rect 175502 104167 175802 104209
rect 175502 104049 175593 104167
rect 175711 104049 175802 104167
rect 175502 86327 175802 104049
rect 175502 86209 175593 86327
rect 175711 86209 175802 86327
rect 175502 86167 175802 86209
rect 175502 86049 175593 86167
rect 175711 86049 175802 86167
rect 175502 68327 175802 86049
rect 175502 68209 175593 68327
rect 175711 68209 175802 68327
rect 175502 68167 175802 68209
rect 175502 68049 175593 68167
rect 175711 68049 175802 68167
rect 175502 50327 175802 68049
rect 175502 50209 175593 50327
rect 175711 50209 175802 50327
rect 175502 50167 175802 50209
rect 175502 50049 175593 50167
rect 175711 50049 175802 50167
rect 175502 32327 175802 50049
rect 175502 32209 175593 32327
rect 175711 32209 175802 32327
rect 175502 32167 175802 32209
rect 175502 32049 175593 32167
rect 175711 32049 175802 32167
rect 175502 14327 175802 32049
rect 175502 14209 175593 14327
rect 175711 14209 175802 14327
rect 175502 14167 175802 14209
rect 175502 14049 175593 14167
rect 175711 14049 175802 14167
rect 175502 -2523 175802 14049
rect 175502 -2641 175593 -2523
rect 175711 -2641 175802 -2523
rect 175502 -2683 175802 -2641
rect 175502 -2801 175593 -2683
rect 175711 -2801 175802 -2683
rect 175502 -2812 175802 -2801
rect 177302 340127 177602 355431
rect 186302 355239 186602 355720
rect 186302 355121 186393 355239
rect 186511 355121 186602 355239
rect 186302 355079 186602 355121
rect 186302 354961 186393 355079
rect 186511 354961 186602 355079
rect 184502 354299 184802 354780
rect 184502 354181 184593 354299
rect 184711 354181 184802 354299
rect 184502 354139 184802 354181
rect 184502 354021 184593 354139
rect 184711 354021 184802 354139
rect 182702 353359 183002 353840
rect 182702 353241 182793 353359
rect 182911 353241 183002 353359
rect 182702 353199 183002 353241
rect 182702 353081 182793 353199
rect 182911 353081 183002 353199
rect 177302 340009 177393 340127
rect 177511 340009 177602 340127
rect 177302 339967 177602 340009
rect 177302 339849 177393 339967
rect 177511 339849 177602 339967
rect 177302 322127 177602 339849
rect 177302 322009 177393 322127
rect 177511 322009 177602 322127
rect 177302 321967 177602 322009
rect 177302 321849 177393 321967
rect 177511 321849 177602 321967
rect 177302 304127 177602 321849
rect 177302 304009 177393 304127
rect 177511 304009 177602 304127
rect 177302 303967 177602 304009
rect 177302 303849 177393 303967
rect 177511 303849 177602 303967
rect 177302 286127 177602 303849
rect 177302 286009 177393 286127
rect 177511 286009 177602 286127
rect 177302 285967 177602 286009
rect 177302 285849 177393 285967
rect 177511 285849 177602 285967
rect 177302 268127 177602 285849
rect 177302 268009 177393 268127
rect 177511 268009 177602 268127
rect 177302 267967 177602 268009
rect 177302 267849 177393 267967
rect 177511 267849 177602 267967
rect 177302 250127 177602 267849
rect 177302 250009 177393 250127
rect 177511 250009 177602 250127
rect 177302 249967 177602 250009
rect 177302 249849 177393 249967
rect 177511 249849 177602 249967
rect 177302 232127 177602 249849
rect 177302 232009 177393 232127
rect 177511 232009 177602 232127
rect 177302 231967 177602 232009
rect 177302 231849 177393 231967
rect 177511 231849 177602 231967
rect 177302 214127 177602 231849
rect 177302 214009 177393 214127
rect 177511 214009 177602 214127
rect 177302 213967 177602 214009
rect 177302 213849 177393 213967
rect 177511 213849 177602 213967
rect 177302 196127 177602 213849
rect 177302 196009 177393 196127
rect 177511 196009 177602 196127
rect 177302 195967 177602 196009
rect 177302 195849 177393 195967
rect 177511 195849 177602 195967
rect 177302 178127 177602 195849
rect 177302 178009 177393 178127
rect 177511 178009 177602 178127
rect 177302 177967 177602 178009
rect 177302 177849 177393 177967
rect 177511 177849 177602 177967
rect 177302 160127 177602 177849
rect 177302 160009 177393 160127
rect 177511 160009 177602 160127
rect 177302 159967 177602 160009
rect 177302 159849 177393 159967
rect 177511 159849 177602 159967
rect 177302 142127 177602 159849
rect 177302 142009 177393 142127
rect 177511 142009 177602 142127
rect 177302 141967 177602 142009
rect 177302 141849 177393 141967
rect 177511 141849 177602 141967
rect 177302 124127 177602 141849
rect 177302 124009 177393 124127
rect 177511 124009 177602 124127
rect 177302 123967 177602 124009
rect 177302 123849 177393 123967
rect 177511 123849 177602 123967
rect 177302 106127 177602 123849
rect 177302 106009 177393 106127
rect 177511 106009 177602 106127
rect 177302 105967 177602 106009
rect 177302 105849 177393 105967
rect 177511 105849 177602 105967
rect 177302 88127 177602 105849
rect 177302 88009 177393 88127
rect 177511 88009 177602 88127
rect 177302 87967 177602 88009
rect 177302 87849 177393 87967
rect 177511 87849 177602 87967
rect 177302 70127 177602 87849
rect 177302 70009 177393 70127
rect 177511 70009 177602 70127
rect 177302 69967 177602 70009
rect 177302 69849 177393 69967
rect 177511 69849 177602 69967
rect 177302 52127 177602 69849
rect 177302 52009 177393 52127
rect 177511 52009 177602 52127
rect 177302 51967 177602 52009
rect 177302 51849 177393 51967
rect 177511 51849 177602 51967
rect 177302 34127 177602 51849
rect 177302 34009 177393 34127
rect 177511 34009 177602 34127
rect 177302 33967 177602 34009
rect 177302 33849 177393 33967
rect 177511 33849 177602 33967
rect 177302 16127 177602 33849
rect 177302 16009 177393 16127
rect 177511 16009 177602 16127
rect 177302 15967 177602 16009
rect 177302 15849 177393 15967
rect 177511 15849 177602 15967
rect 168302 -3111 168393 -2993
rect 168511 -3111 168602 -2993
rect 168302 -3153 168602 -3111
rect 168302 -3271 168393 -3153
rect 168511 -3271 168602 -3153
rect 168302 -3752 168602 -3271
rect 177302 -3463 177602 15849
rect 180902 352419 181202 352900
rect 180902 352301 180993 352419
rect 181111 352301 181202 352419
rect 180902 352259 181202 352301
rect 180902 352141 180993 352259
rect 181111 352141 181202 352259
rect 180902 343727 181202 352141
rect 180902 343609 180993 343727
rect 181111 343609 181202 343727
rect 180902 343567 181202 343609
rect 180902 343449 180993 343567
rect 181111 343449 181202 343567
rect 180902 325727 181202 343449
rect 180902 325609 180993 325727
rect 181111 325609 181202 325727
rect 180902 325567 181202 325609
rect 180902 325449 180993 325567
rect 181111 325449 181202 325567
rect 180902 307727 181202 325449
rect 180902 307609 180993 307727
rect 181111 307609 181202 307727
rect 180902 307567 181202 307609
rect 180902 307449 180993 307567
rect 181111 307449 181202 307567
rect 180902 289727 181202 307449
rect 180902 289609 180993 289727
rect 181111 289609 181202 289727
rect 180902 289567 181202 289609
rect 180902 289449 180993 289567
rect 181111 289449 181202 289567
rect 180902 271727 181202 289449
rect 180902 271609 180993 271727
rect 181111 271609 181202 271727
rect 180902 271567 181202 271609
rect 180902 271449 180993 271567
rect 181111 271449 181202 271567
rect 180902 253727 181202 271449
rect 180902 253609 180993 253727
rect 181111 253609 181202 253727
rect 180902 253567 181202 253609
rect 180902 253449 180993 253567
rect 181111 253449 181202 253567
rect 180902 235727 181202 253449
rect 180902 235609 180993 235727
rect 181111 235609 181202 235727
rect 180902 235567 181202 235609
rect 180902 235449 180993 235567
rect 181111 235449 181202 235567
rect 180902 217727 181202 235449
rect 180902 217609 180993 217727
rect 181111 217609 181202 217727
rect 180902 217567 181202 217609
rect 180902 217449 180993 217567
rect 181111 217449 181202 217567
rect 180902 199727 181202 217449
rect 180902 199609 180993 199727
rect 181111 199609 181202 199727
rect 180902 199567 181202 199609
rect 180902 199449 180993 199567
rect 181111 199449 181202 199567
rect 180902 181727 181202 199449
rect 180902 181609 180993 181727
rect 181111 181609 181202 181727
rect 180902 181567 181202 181609
rect 180902 181449 180993 181567
rect 181111 181449 181202 181567
rect 180902 163727 181202 181449
rect 180902 163609 180993 163727
rect 181111 163609 181202 163727
rect 180902 163567 181202 163609
rect 180902 163449 180993 163567
rect 181111 163449 181202 163567
rect 180902 145727 181202 163449
rect 180902 145609 180993 145727
rect 181111 145609 181202 145727
rect 180902 145567 181202 145609
rect 180902 145449 180993 145567
rect 181111 145449 181202 145567
rect 180902 127727 181202 145449
rect 180902 127609 180993 127727
rect 181111 127609 181202 127727
rect 180902 127567 181202 127609
rect 180902 127449 180993 127567
rect 181111 127449 181202 127567
rect 180902 109727 181202 127449
rect 180902 109609 180993 109727
rect 181111 109609 181202 109727
rect 180902 109567 181202 109609
rect 180902 109449 180993 109567
rect 181111 109449 181202 109567
rect 180902 91727 181202 109449
rect 180902 91609 180993 91727
rect 181111 91609 181202 91727
rect 180902 91567 181202 91609
rect 180902 91449 180993 91567
rect 181111 91449 181202 91567
rect 180902 73727 181202 91449
rect 180902 73609 180993 73727
rect 181111 73609 181202 73727
rect 180902 73567 181202 73609
rect 180902 73449 180993 73567
rect 181111 73449 181202 73567
rect 180902 55727 181202 73449
rect 180902 55609 180993 55727
rect 181111 55609 181202 55727
rect 180902 55567 181202 55609
rect 180902 55449 180993 55567
rect 181111 55449 181202 55567
rect 180902 37727 181202 55449
rect 180902 37609 180993 37727
rect 181111 37609 181202 37727
rect 180902 37567 181202 37609
rect 180902 37449 180993 37567
rect 181111 37449 181202 37567
rect 180902 19727 181202 37449
rect 180902 19609 180993 19727
rect 181111 19609 181202 19727
rect 180902 19567 181202 19609
rect 180902 19449 180993 19567
rect 181111 19449 181202 19567
rect 180902 1727 181202 19449
rect 180902 1609 180993 1727
rect 181111 1609 181202 1727
rect 180902 1567 181202 1609
rect 180902 1449 180993 1567
rect 181111 1449 181202 1567
rect 180902 -173 181202 1449
rect 180902 -291 180993 -173
rect 181111 -291 181202 -173
rect 180902 -333 181202 -291
rect 180902 -451 180993 -333
rect 181111 -451 181202 -333
rect 180902 -932 181202 -451
rect 182702 345527 183002 353081
rect 182702 345409 182793 345527
rect 182911 345409 183002 345527
rect 182702 345367 183002 345409
rect 182702 345249 182793 345367
rect 182911 345249 183002 345367
rect 182702 327527 183002 345249
rect 182702 327409 182793 327527
rect 182911 327409 183002 327527
rect 182702 327367 183002 327409
rect 182702 327249 182793 327367
rect 182911 327249 183002 327367
rect 182702 309527 183002 327249
rect 182702 309409 182793 309527
rect 182911 309409 183002 309527
rect 182702 309367 183002 309409
rect 182702 309249 182793 309367
rect 182911 309249 183002 309367
rect 182702 291527 183002 309249
rect 182702 291409 182793 291527
rect 182911 291409 183002 291527
rect 182702 291367 183002 291409
rect 182702 291249 182793 291367
rect 182911 291249 183002 291367
rect 182702 273527 183002 291249
rect 182702 273409 182793 273527
rect 182911 273409 183002 273527
rect 182702 273367 183002 273409
rect 182702 273249 182793 273367
rect 182911 273249 183002 273367
rect 182702 255527 183002 273249
rect 182702 255409 182793 255527
rect 182911 255409 183002 255527
rect 182702 255367 183002 255409
rect 182702 255249 182793 255367
rect 182911 255249 183002 255367
rect 182702 237527 183002 255249
rect 182702 237409 182793 237527
rect 182911 237409 183002 237527
rect 182702 237367 183002 237409
rect 182702 237249 182793 237367
rect 182911 237249 183002 237367
rect 182702 219527 183002 237249
rect 182702 219409 182793 219527
rect 182911 219409 183002 219527
rect 182702 219367 183002 219409
rect 182702 219249 182793 219367
rect 182911 219249 183002 219367
rect 182702 201527 183002 219249
rect 182702 201409 182793 201527
rect 182911 201409 183002 201527
rect 182702 201367 183002 201409
rect 182702 201249 182793 201367
rect 182911 201249 183002 201367
rect 182702 183527 183002 201249
rect 182702 183409 182793 183527
rect 182911 183409 183002 183527
rect 182702 183367 183002 183409
rect 182702 183249 182793 183367
rect 182911 183249 183002 183367
rect 182702 165527 183002 183249
rect 182702 165409 182793 165527
rect 182911 165409 183002 165527
rect 182702 165367 183002 165409
rect 182702 165249 182793 165367
rect 182911 165249 183002 165367
rect 182702 147527 183002 165249
rect 182702 147409 182793 147527
rect 182911 147409 183002 147527
rect 182702 147367 183002 147409
rect 182702 147249 182793 147367
rect 182911 147249 183002 147367
rect 182702 129527 183002 147249
rect 182702 129409 182793 129527
rect 182911 129409 183002 129527
rect 182702 129367 183002 129409
rect 182702 129249 182793 129367
rect 182911 129249 183002 129367
rect 182702 111527 183002 129249
rect 182702 111409 182793 111527
rect 182911 111409 183002 111527
rect 182702 111367 183002 111409
rect 182702 111249 182793 111367
rect 182911 111249 183002 111367
rect 182702 93527 183002 111249
rect 182702 93409 182793 93527
rect 182911 93409 183002 93527
rect 182702 93367 183002 93409
rect 182702 93249 182793 93367
rect 182911 93249 183002 93367
rect 182702 75527 183002 93249
rect 182702 75409 182793 75527
rect 182911 75409 183002 75527
rect 182702 75367 183002 75409
rect 182702 75249 182793 75367
rect 182911 75249 183002 75367
rect 182702 57527 183002 75249
rect 182702 57409 182793 57527
rect 182911 57409 183002 57527
rect 182702 57367 183002 57409
rect 182702 57249 182793 57367
rect 182911 57249 183002 57367
rect 182702 39527 183002 57249
rect 182702 39409 182793 39527
rect 182911 39409 183002 39527
rect 182702 39367 183002 39409
rect 182702 39249 182793 39367
rect 182911 39249 183002 39367
rect 182702 21527 183002 39249
rect 182702 21409 182793 21527
rect 182911 21409 183002 21527
rect 182702 21367 183002 21409
rect 182702 21249 182793 21367
rect 182911 21249 183002 21367
rect 182702 3527 183002 21249
rect 182702 3409 182793 3527
rect 182911 3409 183002 3527
rect 182702 3367 183002 3409
rect 182702 3249 182793 3367
rect 182911 3249 183002 3367
rect 182702 -1113 183002 3249
rect 182702 -1231 182793 -1113
rect 182911 -1231 183002 -1113
rect 182702 -1273 183002 -1231
rect 182702 -1391 182793 -1273
rect 182911 -1391 183002 -1273
rect 182702 -1872 183002 -1391
rect 184502 347327 184802 354021
rect 184502 347209 184593 347327
rect 184711 347209 184802 347327
rect 184502 347167 184802 347209
rect 184502 347049 184593 347167
rect 184711 347049 184802 347167
rect 184502 329327 184802 347049
rect 184502 329209 184593 329327
rect 184711 329209 184802 329327
rect 184502 329167 184802 329209
rect 184502 329049 184593 329167
rect 184711 329049 184802 329167
rect 184502 311327 184802 329049
rect 184502 311209 184593 311327
rect 184711 311209 184802 311327
rect 184502 311167 184802 311209
rect 184502 311049 184593 311167
rect 184711 311049 184802 311167
rect 184502 293327 184802 311049
rect 184502 293209 184593 293327
rect 184711 293209 184802 293327
rect 184502 293167 184802 293209
rect 184502 293049 184593 293167
rect 184711 293049 184802 293167
rect 184502 275327 184802 293049
rect 184502 275209 184593 275327
rect 184711 275209 184802 275327
rect 184502 275167 184802 275209
rect 184502 275049 184593 275167
rect 184711 275049 184802 275167
rect 184502 257327 184802 275049
rect 184502 257209 184593 257327
rect 184711 257209 184802 257327
rect 184502 257167 184802 257209
rect 184502 257049 184593 257167
rect 184711 257049 184802 257167
rect 184502 239327 184802 257049
rect 184502 239209 184593 239327
rect 184711 239209 184802 239327
rect 184502 239167 184802 239209
rect 184502 239049 184593 239167
rect 184711 239049 184802 239167
rect 184502 221327 184802 239049
rect 184502 221209 184593 221327
rect 184711 221209 184802 221327
rect 184502 221167 184802 221209
rect 184502 221049 184593 221167
rect 184711 221049 184802 221167
rect 184502 203327 184802 221049
rect 184502 203209 184593 203327
rect 184711 203209 184802 203327
rect 184502 203167 184802 203209
rect 184502 203049 184593 203167
rect 184711 203049 184802 203167
rect 184502 185327 184802 203049
rect 184502 185209 184593 185327
rect 184711 185209 184802 185327
rect 184502 185167 184802 185209
rect 184502 185049 184593 185167
rect 184711 185049 184802 185167
rect 184502 167327 184802 185049
rect 184502 167209 184593 167327
rect 184711 167209 184802 167327
rect 184502 167167 184802 167209
rect 184502 167049 184593 167167
rect 184711 167049 184802 167167
rect 184502 149327 184802 167049
rect 184502 149209 184593 149327
rect 184711 149209 184802 149327
rect 184502 149167 184802 149209
rect 184502 149049 184593 149167
rect 184711 149049 184802 149167
rect 184502 131327 184802 149049
rect 184502 131209 184593 131327
rect 184711 131209 184802 131327
rect 184502 131167 184802 131209
rect 184502 131049 184593 131167
rect 184711 131049 184802 131167
rect 184502 113327 184802 131049
rect 184502 113209 184593 113327
rect 184711 113209 184802 113327
rect 184502 113167 184802 113209
rect 184502 113049 184593 113167
rect 184711 113049 184802 113167
rect 184502 95327 184802 113049
rect 184502 95209 184593 95327
rect 184711 95209 184802 95327
rect 184502 95167 184802 95209
rect 184502 95049 184593 95167
rect 184711 95049 184802 95167
rect 184502 77327 184802 95049
rect 184502 77209 184593 77327
rect 184711 77209 184802 77327
rect 184502 77167 184802 77209
rect 184502 77049 184593 77167
rect 184711 77049 184802 77167
rect 184502 59327 184802 77049
rect 184502 59209 184593 59327
rect 184711 59209 184802 59327
rect 184502 59167 184802 59209
rect 184502 59049 184593 59167
rect 184711 59049 184802 59167
rect 184502 41327 184802 59049
rect 184502 41209 184593 41327
rect 184711 41209 184802 41327
rect 184502 41167 184802 41209
rect 184502 41049 184593 41167
rect 184711 41049 184802 41167
rect 184502 23327 184802 41049
rect 184502 23209 184593 23327
rect 184711 23209 184802 23327
rect 184502 23167 184802 23209
rect 184502 23049 184593 23167
rect 184711 23049 184802 23167
rect 184502 5327 184802 23049
rect 184502 5209 184593 5327
rect 184711 5209 184802 5327
rect 184502 5167 184802 5209
rect 184502 5049 184593 5167
rect 184711 5049 184802 5167
rect 184502 -2053 184802 5049
rect 184502 -2171 184593 -2053
rect 184711 -2171 184802 -2053
rect 184502 -2213 184802 -2171
rect 184502 -2331 184593 -2213
rect 184711 -2331 184802 -2213
rect 184502 -2812 184802 -2331
rect 186302 349127 186602 354961
rect 195302 355709 195602 355720
rect 195302 355591 195393 355709
rect 195511 355591 195602 355709
rect 195302 355549 195602 355591
rect 195302 355431 195393 355549
rect 195511 355431 195602 355549
rect 193502 354769 193802 354780
rect 193502 354651 193593 354769
rect 193711 354651 193802 354769
rect 193502 354609 193802 354651
rect 193502 354491 193593 354609
rect 193711 354491 193802 354609
rect 191702 353829 192002 353840
rect 191702 353711 191793 353829
rect 191911 353711 192002 353829
rect 191702 353669 192002 353711
rect 191702 353551 191793 353669
rect 191911 353551 192002 353669
rect 186302 349009 186393 349127
rect 186511 349009 186602 349127
rect 186302 348967 186602 349009
rect 186302 348849 186393 348967
rect 186511 348849 186602 348967
rect 186302 331127 186602 348849
rect 186302 331009 186393 331127
rect 186511 331009 186602 331127
rect 186302 330967 186602 331009
rect 186302 330849 186393 330967
rect 186511 330849 186602 330967
rect 186302 313127 186602 330849
rect 186302 313009 186393 313127
rect 186511 313009 186602 313127
rect 186302 312967 186602 313009
rect 186302 312849 186393 312967
rect 186511 312849 186602 312967
rect 186302 295127 186602 312849
rect 186302 295009 186393 295127
rect 186511 295009 186602 295127
rect 186302 294967 186602 295009
rect 186302 294849 186393 294967
rect 186511 294849 186602 294967
rect 186302 277127 186602 294849
rect 186302 277009 186393 277127
rect 186511 277009 186602 277127
rect 186302 276967 186602 277009
rect 186302 276849 186393 276967
rect 186511 276849 186602 276967
rect 186302 259127 186602 276849
rect 186302 259009 186393 259127
rect 186511 259009 186602 259127
rect 186302 258967 186602 259009
rect 186302 258849 186393 258967
rect 186511 258849 186602 258967
rect 186302 241127 186602 258849
rect 186302 241009 186393 241127
rect 186511 241009 186602 241127
rect 186302 240967 186602 241009
rect 186302 240849 186393 240967
rect 186511 240849 186602 240967
rect 186302 223127 186602 240849
rect 186302 223009 186393 223127
rect 186511 223009 186602 223127
rect 186302 222967 186602 223009
rect 186302 222849 186393 222967
rect 186511 222849 186602 222967
rect 186302 205127 186602 222849
rect 186302 205009 186393 205127
rect 186511 205009 186602 205127
rect 186302 204967 186602 205009
rect 186302 204849 186393 204967
rect 186511 204849 186602 204967
rect 186302 187127 186602 204849
rect 186302 187009 186393 187127
rect 186511 187009 186602 187127
rect 186302 186967 186602 187009
rect 186302 186849 186393 186967
rect 186511 186849 186602 186967
rect 186302 169127 186602 186849
rect 186302 169009 186393 169127
rect 186511 169009 186602 169127
rect 186302 168967 186602 169009
rect 186302 168849 186393 168967
rect 186511 168849 186602 168967
rect 186302 151127 186602 168849
rect 186302 151009 186393 151127
rect 186511 151009 186602 151127
rect 186302 150967 186602 151009
rect 186302 150849 186393 150967
rect 186511 150849 186602 150967
rect 186302 133127 186602 150849
rect 186302 133009 186393 133127
rect 186511 133009 186602 133127
rect 186302 132967 186602 133009
rect 186302 132849 186393 132967
rect 186511 132849 186602 132967
rect 186302 115127 186602 132849
rect 186302 115009 186393 115127
rect 186511 115009 186602 115127
rect 186302 114967 186602 115009
rect 186302 114849 186393 114967
rect 186511 114849 186602 114967
rect 186302 97127 186602 114849
rect 186302 97009 186393 97127
rect 186511 97009 186602 97127
rect 186302 96967 186602 97009
rect 186302 96849 186393 96967
rect 186511 96849 186602 96967
rect 186302 79127 186602 96849
rect 186302 79009 186393 79127
rect 186511 79009 186602 79127
rect 186302 78967 186602 79009
rect 186302 78849 186393 78967
rect 186511 78849 186602 78967
rect 186302 61127 186602 78849
rect 186302 61009 186393 61127
rect 186511 61009 186602 61127
rect 186302 60967 186602 61009
rect 186302 60849 186393 60967
rect 186511 60849 186602 60967
rect 186302 43127 186602 60849
rect 186302 43009 186393 43127
rect 186511 43009 186602 43127
rect 186302 42967 186602 43009
rect 186302 42849 186393 42967
rect 186511 42849 186602 42967
rect 186302 25127 186602 42849
rect 186302 25009 186393 25127
rect 186511 25009 186602 25127
rect 186302 24967 186602 25009
rect 186302 24849 186393 24967
rect 186511 24849 186602 24967
rect 186302 7127 186602 24849
rect 186302 7009 186393 7127
rect 186511 7009 186602 7127
rect 186302 6967 186602 7009
rect 186302 6849 186393 6967
rect 186511 6849 186602 6967
rect 177302 -3581 177393 -3463
rect 177511 -3581 177602 -3463
rect 177302 -3623 177602 -3581
rect 177302 -3741 177393 -3623
rect 177511 -3741 177602 -3623
rect 177302 -3752 177602 -3741
rect 186302 -2993 186602 6849
rect 189902 352889 190202 352900
rect 189902 352771 189993 352889
rect 190111 352771 190202 352889
rect 189902 352729 190202 352771
rect 189902 352611 189993 352729
rect 190111 352611 190202 352729
rect 189902 334727 190202 352611
rect 189902 334609 189993 334727
rect 190111 334609 190202 334727
rect 189902 334567 190202 334609
rect 189902 334449 189993 334567
rect 190111 334449 190202 334567
rect 189902 316727 190202 334449
rect 189902 316609 189993 316727
rect 190111 316609 190202 316727
rect 189902 316567 190202 316609
rect 189902 316449 189993 316567
rect 190111 316449 190202 316567
rect 189902 298727 190202 316449
rect 189902 298609 189993 298727
rect 190111 298609 190202 298727
rect 189902 298567 190202 298609
rect 189902 298449 189993 298567
rect 190111 298449 190202 298567
rect 189902 280727 190202 298449
rect 189902 280609 189993 280727
rect 190111 280609 190202 280727
rect 189902 280567 190202 280609
rect 189902 280449 189993 280567
rect 190111 280449 190202 280567
rect 189902 262727 190202 280449
rect 189902 262609 189993 262727
rect 190111 262609 190202 262727
rect 189902 262567 190202 262609
rect 189902 262449 189993 262567
rect 190111 262449 190202 262567
rect 189902 244727 190202 262449
rect 189902 244609 189993 244727
rect 190111 244609 190202 244727
rect 189902 244567 190202 244609
rect 189902 244449 189993 244567
rect 190111 244449 190202 244567
rect 189902 226727 190202 244449
rect 189902 226609 189993 226727
rect 190111 226609 190202 226727
rect 189902 226567 190202 226609
rect 189902 226449 189993 226567
rect 190111 226449 190202 226567
rect 189902 208727 190202 226449
rect 189902 208609 189993 208727
rect 190111 208609 190202 208727
rect 189902 208567 190202 208609
rect 189902 208449 189993 208567
rect 190111 208449 190202 208567
rect 189902 190727 190202 208449
rect 189902 190609 189993 190727
rect 190111 190609 190202 190727
rect 189902 190567 190202 190609
rect 189902 190449 189993 190567
rect 190111 190449 190202 190567
rect 189902 172727 190202 190449
rect 189902 172609 189993 172727
rect 190111 172609 190202 172727
rect 189902 172567 190202 172609
rect 189902 172449 189993 172567
rect 190111 172449 190202 172567
rect 189902 154727 190202 172449
rect 189902 154609 189993 154727
rect 190111 154609 190202 154727
rect 189902 154567 190202 154609
rect 189902 154449 189993 154567
rect 190111 154449 190202 154567
rect 189902 136727 190202 154449
rect 189902 136609 189993 136727
rect 190111 136609 190202 136727
rect 189902 136567 190202 136609
rect 189902 136449 189993 136567
rect 190111 136449 190202 136567
rect 189902 118727 190202 136449
rect 189902 118609 189993 118727
rect 190111 118609 190202 118727
rect 189902 118567 190202 118609
rect 189902 118449 189993 118567
rect 190111 118449 190202 118567
rect 189902 100727 190202 118449
rect 189902 100609 189993 100727
rect 190111 100609 190202 100727
rect 189902 100567 190202 100609
rect 189902 100449 189993 100567
rect 190111 100449 190202 100567
rect 189902 82727 190202 100449
rect 189902 82609 189993 82727
rect 190111 82609 190202 82727
rect 189902 82567 190202 82609
rect 189902 82449 189993 82567
rect 190111 82449 190202 82567
rect 189902 64727 190202 82449
rect 189902 64609 189993 64727
rect 190111 64609 190202 64727
rect 189902 64567 190202 64609
rect 189902 64449 189993 64567
rect 190111 64449 190202 64567
rect 189902 46727 190202 64449
rect 189902 46609 189993 46727
rect 190111 46609 190202 46727
rect 189902 46567 190202 46609
rect 189902 46449 189993 46567
rect 190111 46449 190202 46567
rect 189902 28727 190202 46449
rect 189902 28609 189993 28727
rect 190111 28609 190202 28727
rect 189902 28567 190202 28609
rect 189902 28449 189993 28567
rect 190111 28449 190202 28567
rect 189902 10727 190202 28449
rect 189902 10609 189993 10727
rect 190111 10609 190202 10727
rect 189902 10567 190202 10609
rect 189902 10449 189993 10567
rect 190111 10449 190202 10567
rect 189902 -643 190202 10449
rect 189902 -761 189993 -643
rect 190111 -761 190202 -643
rect 189902 -803 190202 -761
rect 189902 -921 189993 -803
rect 190111 -921 190202 -803
rect 189902 -932 190202 -921
rect 191702 336527 192002 353551
rect 191702 336409 191793 336527
rect 191911 336409 192002 336527
rect 191702 336367 192002 336409
rect 191702 336249 191793 336367
rect 191911 336249 192002 336367
rect 191702 318527 192002 336249
rect 191702 318409 191793 318527
rect 191911 318409 192002 318527
rect 191702 318367 192002 318409
rect 191702 318249 191793 318367
rect 191911 318249 192002 318367
rect 191702 300527 192002 318249
rect 191702 300409 191793 300527
rect 191911 300409 192002 300527
rect 191702 300367 192002 300409
rect 191702 300249 191793 300367
rect 191911 300249 192002 300367
rect 191702 282527 192002 300249
rect 191702 282409 191793 282527
rect 191911 282409 192002 282527
rect 191702 282367 192002 282409
rect 191702 282249 191793 282367
rect 191911 282249 192002 282367
rect 191702 264527 192002 282249
rect 191702 264409 191793 264527
rect 191911 264409 192002 264527
rect 191702 264367 192002 264409
rect 191702 264249 191793 264367
rect 191911 264249 192002 264367
rect 191702 246527 192002 264249
rect 191702 246409 191793 246527
rect 191911 246409 192002 246527
rect 191702 246367 192002 246409
rect 191702 246249 191793 246367
rect 191911 246249 192002 246367
rect 191702 228527 192002 246249
rect 191702 228409 191793 228527
rect 191911 228409 192002 228527
rect 191702 228367 192002 228409
rect 191702 228249 191793 228367
rect 191911 228249 192002 228367
rect 191702 210527 192002 228249
rect 191702 210409 191793 210527
rect 191911 210409 192002 210527
rect 191702 210367 192002 210409
rect 191702 210249 191793 210367
rect 191911 210249 192002 210367
rect 191702 192527 192002 210249
rect 191702 192409 191793 192527
rect 191911 192409 192002 192527
rect 191702 192367 192002 192409
rect 191702 192249 191793 192367
rect 191911 192249 192002 192367
rect 191702 174527 192002 192249
rect 191702 174409 191793 174527
rect 191911 174409 192002 174527
rect 191702 174367 192002 174409
rect 191702 174249 191793 174367
rect 191911 174249 192002 174367
rect 191702 156527 192002 174249
rect 191702 156409 191793 156527
rect 191911 156409 192002 156527
rect 191702 156367 192002 156409
rect 191702 156249 191793 156367
rect 191911 156249 192002 156367
rect 191702 138527 192002 156249
rect 191702 138409 191793 138527
rect 191911 138409 192002 138527
rect 191702 138367 192002 138409
rect 191702 138249 191793 138367
rect 191911 138249 192002 138367
rect 191702 120527 192002 138249
rect 191702 120409 191793 120527
rect 191911 120409 192002 120527
rect 191702 120367 192002 120409
rect 191702 120249 191793 120367
rect 191911 120249 192002 120367
rect 191702 102527 192002 120249
rect 191702 102409 191793 102527
rect 191911 102409 192002 102527
rect 191702 102367 192002 102409
rect 191702 102249 191793 102367
rect 191911 102249 192002 102367
rect 191702 84527 192002 102249
rect 191702 84409 191793 84527
rect 191911 84409 192002 84527
rect 191702 84367 192002 84409
rect 191702 84249 191793 84367
rect 191911 84249 192002 84367
rect 191702 66527 192002 84249
rect 191702 66409 191793 66527
rect 191911 66409 192002 66527
rect 191702 66367 192002 66409
rect 191702 66249 191793 66367
rect 191911 66249 192002 66367
rect 191702 48527 192002 66249
rect 191702 48409 191793 48527
rect 191911 48409 192002 48527
rect 191702 48367 192002 48409
rect 191702 48249 191793 48367
rect 191911 48249 192002 48367
rect 191702 30527 192002 48249
rect 191702 30409 191793 30527
rect 191911 30409 192002 30527
rect 191702 30367 192002 30409
rect 191702 30249 191793 30367
rect 191911 30249 192002 30367
rect 191702 12527 192002 30249
rect 191702 12409 191793 12527
rect 191911 12409 192002 12527
rect 191702 12367 192002 12409
rect 191702 12249 191793 12367
rect 191911 12249 192002 12367
rect 191702 -1583 192002 12249
rect 191702 -1701 191793 -1583
rect 191911 -1701 192002 -1583
rect 191702 -1743 192002 -1701
rect 191702 -1861 191793 -1743
rect 191911 -1861 192002 -1743
rect 191702 -1872 192002 -1861
rect 193502 338327 193802 354491
rect 193502 338209 193593 338327
rect 193711 338209 193802 338327
rect 193502 338167 193802 338209
rect 193502 338049 193593 338167
rect 193711 338049 193802 338167
rect 193502 320327 193802 338049
rect 193502 320209 193593 320327
rect 193711 320209 193802 320327
rect 193502 320167 193802 320209
rect 193502 320049 193593 320167
rect 193711 320049 193802 320167
rect 193502 302327 193802 320049
rect 193502 302209 193593 302327
rect 193711 302209 193802 302327
rect 193502 302167 193802 302209
rect 193502 302049 193593 302167
rect 193711 302049 193802 302167
rect 193502 284327 193802 302049
rect 193502 284209 193593 284327
rect 193711 284209 193802 284327
rect 193502 284167 193802 284209
rect 193502 284049 193593 284167
rect 193711 284049 193802 284167
rect 193502 266327 193802 284049
rect 193502 266209 193593 266327
rect 193711 266209 193802 266327
rect 193502 266167 193802 266209
rect 193502 266049 193593 266167
rect 193711 266049 193802 266167
rect 193502 248327 193802 266049
rect 193502 248209 193593 248327
rect 193711 248209 193802 248327
rect 193502 248167 193802 248209
rect 193502 248049 193593 248167
rect 193711 248049 193802 248167
rect 193502 230327 193802 248049
rect 193502 230209 193593 230327
rect 193711 230209 193802 230327
rect 193502 230167 193802 230209
rect 193502 230049 193593 230167
rect 193711 230049 193802 230167
rect 193502 212327 193802 230049
rect 193502 212209 193593 212327
rect 193711 212209 193802 212327
rect 193502 212167 193802 212209
rect 193502 212049 193593 212167
rect 193711 212049 193802 212167
rect 193502 194327 193802 212049
rect 193502 194209 193593 194327
rect 193711 194209 193802 194327
rect 193502 194167 193802 194209
rect 193502 194049 193593 194167
rect 193711 194049 193802 194167
rect 193502 176327 193802 194049
rect 193502 176209 193593 176327
rect 193711 176209 193802 176327
rect 193502 176167 193802 176209
rect 193502 176049 193593 176167
rect 193711 176049 193802 176167
rect 193502 158327 193802 176049
rect 193502 158209 193593 158327
rect 193711 158209 193802 158327
rect 193502 158167 193802 158209
rect 193502 158049 193593 158167
rect 193711 158049 193802 158167
rect 193502 140327 193802 158049
rect 193502 140209 193593 140327
rect 193711 140209 193802 140327
rect 193502 140167 193802 140209
rect 193502 140049 193593 140167
rect 193711 140049 193802 140167
rect 193502 122327 193802 140049
rect 193502 122209 193593 122327
rect 193711 122209 193802 122327
rect 193502 122167 193802 122209
rect 193502 122049 193593 122167
rect 193711 122049 193802 122167
rect 193502 104327 193802 122049
rect 193502 104209 193593 104327
rect 193711 104209 193802 104327
rect 193502 104167 193802 104209
rect 193502 104049 193593 104167
rect 193711 104049 193802 104167
rect 193502 86327 193802 104049
rect 193502 86209 193593 86327
rect 193711 86209 193802 86327
rect 193502 86167 193802 86209
rect 193502 86049 193593 86167
rect 193711 86049 193802 86167
rect 193502 68327 193802 86049
rect 193502 68209 193593 68327
rect 193711 68209 193802 68327
rect 193502 68167 193802 68209
rect 193502 68049 193593 68167
rect 193711 68049 193802 68167
rect 193502 50327 193802 68049
rect 193502 50209 193593 50327
rect 193711 50209 193802 50327
rect 193502 50167 193802 50209
rect 193502 50049 193593 50167
rect 193711 50049 193802 50167
rect 193502 32327 193802 50049
rect 193502 32209 193593 32327
rect 193711 32209 193802 32327
rect 193502 32167 193802 32209
rect 193502 32049 193593 32167
rect 193711 32049 193802 32167
rect 193502 14327 193802 32049
rect 193502 14209 193593 14327
rect 193711 14209 193802 14327
rect 193502 14167 193802 14209
rect 193502 14049 193593 14167
rect 193711 14049 193802 14167
rect 193502 -2523 193802 14049
rect 193502 -2641 193593 -2523
rect 193711 -2641 193802 -2523
rect 193502 -2683 193802 -2641
rect 193502 -2801 193593 -2683
rect 193711 -2801 193802 -2683
rect 193502 -2812 193802 -2801
rect 195302 340127 195602 355431
rect 204302 355239 204602 355720
rect 204302 355121 204393 355239
rect 204511 355121 204602 355239
rect 204302 355079 204602 355121
rect 204302 354961 204393 355079
rect 204511 354961 204602 355079
rect 202502 354299 202802 354780
rect 202502 354181 202593 354299
rect 202711 354181 202802 354299
rect 202502 354139 202802 354181
rect 202502 354021 202593 354139
rect 202711 354021 202802 354139
rect 200702 353359 201002 353840
rect 200702 353241 200793 353359
rect 200911 353241 201002 353359
rect 200702 353199 201002 353241
rect 200702 353081 200793 353199
rect 200911 353081 201002 353199
rect 195302 340009 195393 340127
rect 195511 340009 195602 340127
rect 195302 339967 195602 340009
rect 195302 339849 195393 339967
rect 195511 339849 195602 339967
rect 195302 322127 195602 339849
rect 195302 322009 195393 322127
rect 195511 322009 195602 322127
rect 195302 321967 195602 322009
rect 195302 321849 195393 321967
rect 195511 321849 195602 321967
rect 195302 304127 195602 321849
rect 195302 304009 195393 304127
rect 195511 304009 195602 304127
rect 195302 303967 195602 304009
rect 195302 303849 195393 303967
rect 195511 303849 195602 303967
rect 195302 286127 195602 303849
rect 195302 286009 195393 286127
rect 195511 286009 195602 286127
rect 195302 285967 195602 286009
rect 195302 285849 195393 285967
rect 195511 285849 195602 285967
rect 195302 268127 195602 285849
rect 195302 268009 195393 268127
rect 195511 268009 195602 268127
rect 195302 267967 195602 268009
rect 195302 267849 195393 267967
rect 195511 267849 195602 267967
rect 195302 250127 195602 267849
rect 195302 250009 195393 250127
rect 195511 250009 195602 250127
rect 195302 249967 195602 250009
rect 195302 249849 195393 249967
rect 195511 249849 195602 249967
rect 195302 232127 195602 249849
rect 195302 232009 195393 232127
rect 195511 232009 195602 232127
rect 195302 231967 195602 232009
rect 195302 231849 195393 231967
rect 195511 231849 195602 231967
rect 195302 214127 195602 231849
rect 195302 214009 195393 214127
rect 195511 214009 195602 214127
rect 195302 213967 195602 214009
rect 195302 213849 195393 213967
rect 195511 213849 195602 213967
rect 195302 196127 195602 213849
rect 195302 196009 195393 196127
rect 195511 196009 195602 196127
rect 195302 195967 195602 196009
rect 195302 195849 195393 195967
rect 195511 195849 195602 195967
rect 195302 178127 195602 195849
rect 195302 178009 195393 178127
rect 195511 178009 195602 178127
rect 195302 177967 195602 178009
rect 195302 177849 195393 177967
rect 195511 177849 195602 177967
rect 195302 160127 195602 177849
rect 195302 160009 195393 160127
rect 195511 160009 195602 160127
rect 195302 159967 195602 160009
rect 195302 159849 195393 159967
rect 195511 159849 195602 159967
rect 195302 142127 195602 159849
rect 195302 142009 195393 142127
rect 195511 142009 195602 142127
rect 195302 141967 195602 142009
rect 195302 141849 195393 141967
rect 195511 141849 195602 141967
rect 195302 124127 195602 141849
rect 195302 124009 195393 124127
rect 195511 124009 195602 124127
rect 195302 123967 195602 124009
rect 195302 123849 195393 123967
rect 195511 123849 195602 123967
rect 195302 106127 195602 123849
rect 195302 106009 195393 106127
rect 195511 106009 195602 106127
rect 195302 105967 195602 106009
rect 195302 105849 195393 105967
rect 195511 105849 195602 105967
rect 195302 88127 195602 105849
rect 195302 88009 195393 88127
rect 195511 88009 195602 88127
rect 195302 87967 195602 88009
rect 195302 87849 195393 87967
rect 195511 87849 195602 87967
rect 195302 70127 195602 87849
rect 195302 70009 195393 70127
rect 195511 70009 195602 70127
rect 195302 69967 195602 70009
rect 195302 69849 195393 69967
rect 195511 69849 195602 69967
rect 195302 52127 195602 69849
rect 195302 52009 195393 52127
rect 195511 52009 195602 52127
rect 195302 51967 195602 52009
rect 195302 51849 195393 51967
rect 195511 51849 195602 51967
rect 195302 34127 195602 51849
rect 195302 34009 195393 34127
rect 195511 34009 195602 34127
rect 195302 33967 195602 34009
rect 195302 33849 195393 33967
rect 195511 33849 195602 33967
rect 195302 16127 195602 33849
rect 195302 16009 195393 16127
rect 195511 16009 195602 16127
rect 195302 15967 195602 16009
rect 195302 15849 195393 15967
rect 195511 15849 195602 15967
rect 186302 -3111 186393 -2993
rect 186511 -3111 186602 -2993
rect 186302 -3153 186602 -3111
rect 186302 -3271 186393 -3153
rect 186511 -3271 186602 -3153
rect 186302 -3752 186602 -3271
rect 195302 -3463 195602 15849
rect 198902 352419 199202 352900
rect 198902 352301 198993 352419
rect 199111 352301 199202 352419
rect 198902 352259 199202 352301
rect 198902 352141 198993 352259
rect 199111 352141 199202 352259
rect 198902 343727 199202 352141
rect 198902 343609 198993 343727
rect 199111 343609 199202 343727
rect 198902 343567 199202 343609
rect 198902 343449 198993 343567
rect 199111 343449 199202 343567
rect 198902 325727 199202 343449
rect 198902 325609 198993 325727
rect 199111 325609 199202 325727
rect 198902 325567 199202 325609
rect 198902 325449 198993 325567
rect 199111 325449 199202 325567
rect 198902 307727 199202 325449
rect 198902 307609 198993 307727
rect 199111 307609 199202 307727
rect 198902 307567 199202 307609
rect 198902 307449 198993 307567
rect 199111 307449 199202 307567
rect 198902 289727 199202 307449
rect 198902 289609 198993 289727
rect 199111 289609 199202 289727
rect 198902 289567 199202 289609
rect 198902 289449 198993 289567
rect 199111 289449 199202 289567
rect 198902 271727 199202 289449
rect 198902 271609 198993 271727
rect 199111 271609 199202 271727
rect 198902 271567 199202 271609
rect 198902 271449 198993 271567
rect 199111 271449 199202 271567
rect 198902 253727 199202 271449
rect 198902 253609 198993 253727
rect 199111 253609 199202 253727
rect 198902 253567 199202 253609
rect 198902 253449 198993 253567
rect 199111 253449 199202 253567
rect 198902 235727 199202 253449
rect 198902 235609 198993 235727
rect 199111 235609 199202 235727
rect 198902 235567 199202 235609
rect 198902 235449 198993 235567
rect 199111 235449 199202 235567
rect 198902 217727 199202 235449
rect 198902 217609 198993 217727
rect 199111 217609 199202 217727
rect 198902 217567 199202 217609
rect 198902 217449 198993 217567
rect 199111 217449 199202 217567
rect 198902 199727 199202 217449
rect 198902 199609 198993 199727
rect 199111 199609 199202 199727
rect 198902 199567 199202 199609
rect 198902 199449 198993 199567
rect 199111 199449 199202 199567
rect 198902 181727 199202 199449
rect 198902 181609 198993 181727
rect 199111 181609 199202 181727
rect 198902 181567 199202 181609
rect 198902 181449 198993 181567
rect 199111 181449 199202 181567
rect 198902 163727 199202 181449
rect 198902 163609 198993 163727
rect 199111 163609 199202 163727
rect 198902 163567 199202 163609
rect 198902 163449 198993 163567
rect 199111 163449 199202 163567
rect 198902 145727 199202 163449
rect 198902 145609 198993 145727
rect 199111 145609 199202 145727
rect 198902 145567 199202 145609
rect 198902 145449 198993 145567
rect 199111 145449 199202 145567
rect 198902 127727 199202 145449
rect 198902 127609 198993 127727
rect 199111 127609 199202 127727
rect 198902 127567 199202 127609
rect 198902 127449 198993 127567
rect 199111 127449 199202 127567
rect 198902 109727 199202 127449
rect 198902 109609 198993 109727
rect 199111 109609 199202 109727
rect 198902 109567 199202 109609
rect 198902 109449 198993 109567
rect 199111 109449 199202 109567
rect 198902 91727 199202 109449
rect 198902 91609 198993 91727
rect 199111 91609 199202 91727
rect 198902 91567 199202 91609
rect 198902 91449 198993 91567
rect 199111 91449 199202 91567
rect 198902 73727 199202 91449
rect 198902 73609 198993 73727
rect 199111 73609 199202 73727
rect 198902 73567 199202 73609
rect 198902 73449 198993 73567
rect 199111 73449 199202 73567
rect 198902 55727 199202 73449
rect 198902 55609 198993 55727
rect 199111 55609 199202 55727
rect 198902 55567 199202 55609
rect 198902 55449 198993 55567
rect 199111 55449 199202 55567
rect 198902 37727 199202 55449
rect 198902 37609 198993 37727
rect 199111 37609 199202 37727
rect 198902 37567 199202 37609
rect 198902 37449 198993 37567
rect 199111 37449 199202 37567
rect 198902 19727 199202 37449
rect 198902 19609 198993 19727
rect 199111 19609 199202 19727
rect 198902 19567 199202 19609
rect 198902 19449 198993 19567
rect 199111 19449 199202 19567
rect 198902 1727 199202 19449
rect 198902 1609 198993 1727
rect 199111 1609 199202 1727
rect 198902 1567 199202 1609
rect 198902 1449 198993 1567
rect 199111 1449 199202 1567
rect 198902 -173 199202 1449
rect 198902 -291 198993 -173
rect 199111 -291 199202 -173
rect 198902 -333 199202 -291
rect 198902 -451 198993 -333
rect 199111 -451 199202 -333
rect 198902 -932 199202 -451
rect 200702 345527 201002 353081
rect 200702 345409 200793 345527
rect 200911 345409 201002 345527
rect 200702 345367 201002 345409
rect 200702 345249 200793 345367
rect 200911 345249 201002 345367
rect 200702 327527 201002 345249
rect 200702 327409 200793 327527
rect 200911 327409 201002 327527
rect 200702 327367 201002 327409
rect 200702 327249 200793 327367
rect 200911 327249 201002 327367
rect 200702 309527 201002 327249
rect 200702 309409 200793 309527
rect 200911 309409 201002 309527
rect 200702 309367 201002 309409
rect 200702 309249 200793 309367
rect 200911 309249 201002 309367
rect 200702 291527 201002 309249
rect 200702 291409 200793 291527
rect 200911 291409 201002 291527
rect 200702 291367 201002 291409
rect 200702 291249 200793 291367
rect 200911 291249 201002 291367
rect 200702 273527 201002 291249
rect 200702 273409 200793 273527
rect 200911 273409 201002 273527
rect 200702 273367 201002 273409
rect 200702 273249 200793 273367
rect 200911 273249 201002 273367
rect 200702 255527 201002 273249
rect 200702 255409 200793 255527
rect 200911 255409 201002 255527
rect 200702 255367 201002 255409
rect 200702 255249 200793 255367
rect 200911 255249 201002 255367
rect 200702 237527 201002 255249
rect 200702 237409 200793 237527
rect 200911 237409 201002 237527
rect 200702 237367 201002 237409
rect 200702 237249 200793 237367
rect 200911 237249 201002 237367
rect 200702 219527 201002 237249
rect 200702 219409 200793 219527
rect 200911 219409 201002 219527
rect 200702 219367 201002 219409
rect 200702 219249 200793 219367
rect 200911 219249 201002 219367
rect 200702 201527 201002 219249
rect 200702 201409 200793 201527
rect 200911 201409 201002 201527
rect 200702 201367 201002 201409
rect 200702 201249 200793 201367
rect 200911 201249 201002 201367
rect 200702 183527 201002 201249
rect 200702 183409 200793 183527
rect 200911 183409 201002 183527
rect 200702 183367 201002 183409
rect 200702 183249 200793 183367
rect 200911 183249 201002 183367
rect 200702 165527 201002 183249
rect 200702 165409 200793 165527
rect 200911 165409 201002 165527
rect 200702 165367 201002 165409
rect 200702 165249 200793 165367
rect 200911 165249 201002 165367
rect 200702 147527 201002 165249
rect 200702 147409 200793 147527
rect 200911 147409 201002 147527
rect 200702 147367 201002 147409
rect 200702 147249 200793 147367
rect 200911 147249 201002 147367
rect 200702 129527 201002 147249
rect 200702 129409 200793 129527
rect 200911 129409 201002 129527
rect 200702 129367 201002 129409
rect 200702 129249 200793 129367
rect 200911 129249 201002 129367
rect 200702 111527 201002 129249
rect 200702 111409 200793 111527
rect 200911 111409 201002 111527
rect 200702 111367 201002 111409
rect 200702 111249 200793 111367
rect 200911 111249 201002 111367
rect 200702 93527 201002 111249
rect 200702 93409 200793 93527
rect 200911 93409 201002 93527
rect 200702 93367 201002 93409
rect 200702 93249 200793 93367
rect 200911 93249 201002 93367
rect 200702 75527 201002 93249
rect 200702 75409 200793 75527
rect 200911 75409 201002 75527
rect 200702 75367 201002 75409
rect 200702 75249 200793 75367
rect 200911 75249 201002 75367
rect 200702 57527 201002 75249
rect 200702 57409 200793 57527
rect 200911 57409 201002 57527
rect 200702 57367 201002 57409
rect 200702 57249 200793 57367
rect 200911 57249 201002 57367
rect 200702 39527 201002 57249
rect 200702 39409 200793 39527
rect 200911 39409 201002 39527
rect 200702 39367 201002 39409
rect 200702 39249 200793 39367
rect 200911 39249 201002 39367
rect 200702 21527 201002 39249
rect 200702 21409 200793 21527
rect 200911 21409 201002 21527
rect 200702 21367 201002 21409
rect 200702 21249 200793 21367
rect 200911 21249 201002 21367
rect 200702 3527 201002 21249
rect 200702 3409 200793 3527
rect 200911 3409 201002 3527
rect 200702 3367 201002 3409
rect 200702 3249 200793 3367
rect 200911 3249 201002 3367
rect 200702 -1113 201002 3249
rect 200702 -1231 200793 -1113
rect 200911 -1231 201002 -1113
rect 200702 -1273 201002 -1231
rect 200702 -1391 200793 -1273
rect 200911 -1391 201002 -1273
rect 200702 -1872 201002 -1391
rect 202502 347327 202802 354021
rect 202502 347209 202593 347327
rect 202711 347209 202802 347327
rect 202502 347167 202802 347209
rect 202502 347049 202593 347167
rect 202711 347049 202802 347167
rect 202502 329327 202802 347049
rect 202502 329209 202593 329327
rect 202711 329209 202802 329327
rect 202502 329167 202802 329209
rect 202502 329049 202593 329167
rect 202711 329049 202802 329167
rect 202502 311327 202802 329049
rect 202502 311209 202593 311327
rect 202711 311209 202802 311327
rect 202502 311167 202802 311209
rect 202502 311049 202593 311167
rect 202711 311049 202802 311167
rect 202502 293327 202802 311049
rect 202502 293209 202593 293327
rect 202711 293209 202802 293327
rect 202502 293167 202802 293209
rect 202502 293049 202593 293167
rect 202711 293049 202802 293167
rect 202502 275327 202802 293049
rect 202502 275209 202593 275327
rect 202711 275209 202802 275327
rect 202502 275167 202802 275209
rect 202502 275049 202593 275167
rect 202711 275049 202802 275167
rect 202502 257327 202802 275049
rect 202502 257209 202593 257327
rect 202711 257209 202802 257327
rect 202502 257167 202802 257209
rect 202502 257049 202593 257167
rect 202711 257049 202802 257167
rect 202502 239327 202802 257049
rect 202502 239209 202593 239327
rect 202711 239209 202802 239327
rect 202502 239167 202802 239209
rect 202502 239049 202593 239167
rect 202711 239049 202802 239167
rect 202502 221327 202802 239049
rect 202502 221209 202593 221327
rect 202711 221209 202802 221327
rect 202502 221167 202802 221209
rect 202502 221049 202593 221167
rect 202711 221049 202802 221167
rect 202502 203327 202802 221049
rect 202502 203209 202593 203327
rect 202711 203209 202802 203327
rect 202502 203167 202802 203209
rect 202502 203049 202593 203167
rect 202711 203049 202802 203167
rect 202502 185327 202802 203049
rect 202502 185209 202593 185327
rect 202711 185209 202802 185327
rect 202502 185167 202802 185209
rect 202502 185049 202593 185167
rect 202711 185049 202802 185167
rect 202502 167327 202802 185049
rect 202502 167209 202593 167327
rect 202711 167209 202802 167327
rect 202502 167167 202802 167209
rect 202502 167049 202593 167167
rect 202711 167049 202802 167167
rect 202502 149327 202802 167049
rect 202502 149209 202593 149327
rect 202711 149209 202802 149327
rect 202502 149167 202802 149209
rect 202502 149049 202593 149167
rect 202711 149049 202802 149167
rect 202502 131327 202802 149049
rect 202502 131209 202593 131327
rect 202711 131209 202802 131327
rect 202502 131167 202802 131209
rect 202502 131049 202593 131167
rect 202711 131049 202802 131167
rect 202502 113327 202802 131049
rect 202502 113209 202593 113327
rect 202711 113209 202802 113327
rect 202502 113167 202802 113209
rect 202502 113049 202593 113167
rect 202711 113049 202802 113167
rect 202502 95327 202802 113049
rect 202502 95209 202593 95327
rect 202711 95209 202802 95327
rect 202502 95167 202802 95209
rect 202502 95049 202593 95167
rect 202711 95049 202802 95167
rect 202502 77327 202802 95049
rect 202502 77209 202593 77327
rect 202711 77209 202802 77327
rect 202502 77167 202802 77209
rect 202502 77049 202593 77167
rect 202711 77049 202802 77167
rect 202502 59327 202802 77049
rect 202502 59209 202593 59327
rect 202711 59209 202802 59327
rect 202502 59167 202802 59209
rect 202502 59049 202593 59167
rect 202711 59049 202802 59167
rect 202502 41327 202802 59049
rect 202502 41209 202593 41327
rect 202711 41209 202802 41327
rect 202502 41167 202802 41209
rect 202502 41049 202593 41167
rect 202711 41049 202802 41167
rect 202502 23327 202802 41049
rect 202502 23209 202593 23327
rect 202711 23209 202802 23327
rect 202502 23167 202802 23209
rect 202502 23049 202593 23167
rect 202711 23049 202802 23167
rect 202502 5327 202802 23049
rect 202502 5209 202593 5327
rect 202711 5209 202802 5327
rect 202502 5167 202802 5209
rect 202502 5049 202593 5167
rect 202711 5049 202802 5167
rect 202502 -2053 202802 5049
rect 202502 -2171 202593 -2053
rect 202711 -2171 202802 -2053
rect 202502 -2213 202802 -2171
rect 202502 -2331 202593 -2213
rect 202711 -2331 202802 -2213
rect 202502 -2812 202802 -2331
rect 204302 349127 204602 354961
rect 213302 355709 213602 355720
rect 213302 355591 213393 355709
rect 213511 355591 213602 355709
rect 213302 355549 213602 355591
rect 213302 355431 213393 355549
rect 213511 355431 213602 355549
rect 211502 354769 211802 354780
rect 211502 354651 211593 354769
rect 211711 354651 211802 354769
rect 211502 354609 211802 354651
rect 211502 354491 211593 354609
rect 211711 354491 211802 354609
rect 209702 353829 210002 353840
rect 209702 353711 209793 353829
rect 209911 353711 210002 353829
rect 209702 353669 210002 353711
rect 209702 353551 209793 353669
rect 209911 353551 210002 353669
rect 204302 349009 204393 349127
rect 204511 349009 204602 349127
rect 204302 348967 204602 349009
rect 204302 348849 204393 348967
rect 204511 348849 204602 348967
rect 204302 331127 204602 348849
rect 204302 331009 204393 331127
rect 204511 331009 204602 331127
rect 204302 330967 204602 331009
rect 204302 330849 204393 330967
rect 204511 330849 204602 330967
rect 204302 313127 204602 330849
rect 204302 313009 204393 313127
rect 204511 313009 204602 313127
rect 204302 312967 204602 313009
rect 204302 312849 204393 312967
rect 204511 312849 204602 312967
rect 204302 295127 204602 312849
rect 204302 295009 204393 295127
rect 204511 295009 204602 295127
rect 204302 294967 204602 295009
rect 204302 294849 204393 294967
rect 204511 294849 204602 294967
rect 204302 277127 204602 294849
rect 204302 277009 204393 277127
rect 204511 277009 204602 277127
rect 204302 276967 204602 277009
rect 204302 276849 204393 276967
rect 204511 276849 204602 276967
rect 204302 259127 204602 276849
rect 204302 259009 204393 259127
rect 204511 259009 204602 259127
rect 204302 258967 204602 259009
rect 204302 258849 204393 258967
rect 204511 258849 204602 258967
rect 204302 241127 204602 258849
rect 204302 241009 204393 241127
rect 204511 241009 204602 241127
rect 204302 240967 204602 241009
rect 204302 240849 204393 240967
rect 204511 240849 204602 240967
rect 204302 223127 204602 240849
rect 204302 223009 204393 223127
rect 204511 223009 204602 223127
rect 204302 222967 204602 223009
rect 204302 222849 204393 222967
rect 204511 222849 204602 222967
rect 204302 205127 204602 222849
rect 204302 205009 204393 205127
rect 204511 205009 204602 205127
rect 204302 204967 204602 205009
rect 204302 204849 204393 204967
rect 204511 204849 204602 204967
rect 204302 187127 204602 204849
rect 204302 187009 204393 187127
rect 204511 187009 204602 187127
rect 204302 186967 204602 187009
rect 204302 186849 204393 186967
rect 204511 186849 204602 186967
rect 204302 169127 204602 186849
rect 204302 169009 204393 169127
rect 204511 169009 204602 169127
rect 204302 168967 204602 169009
rect 204302 168849 204393 168967
rect 204511 168849 204602 168967
rect 204302 151127 204602 168849
rect 204302 151009 204393 151127
rect 204511 151009 204602 151127
rect 204302 150967 204602 151009
rect 204302 150849 204393 150967
rect 204511 150849 204602 150967
rect 204302 133127 204602 150849
rect 204302 133009 204393 133127
rect 204511 133009 204602 133127
rect 204302 132967 204602 133009
rect 204302 132849 204393 132967
rect 204511 132849 204602 132967
rect 204302 115127 204602 132849
rect 204302 115009 204393 115127
rect 204511 115009 204602 115127
rect 204302 114967 204602 115009
rect 204302 114849 204393 114967
rect 204511 114849 204602 114967
rect 204302 97127 204602 114849
rect 204302 97009 204393 97127
rect 204511 97009 204602 97127
rect 204302 96967 204602 97009
rect 204302 96849 204393 96967
rect 204511 96849 204602 96967
rect 204302 79127 204602 96849
rect 204302 79009 204393 79127
rect 204511 79009 204602 79127
rect 204302 78967 204602 79009
rect 204302 78849 204393 78967
rect 204511 78849 204602 78967
rect 204302 61127 204602 78849
rect 204302 61009 204393 61127
rect 204511 61009 204602 61127
rect 204302 60967 204602 61009
rect 204302 60849 204393 60967
rect 204511 60849 204602 60967
rect 204302 43127 204602 60849
rect 204302 43009 204393 43127
rect 204511 43009 204602 43127
rect 204302 42967 204602 43009
rect 204302 42849 204393 42967
rect 204511 42849 204602 42967
rect 204302 25127 204602 42849
rect 204302 25009 204393 25127
rect 204511 25009 204602 25127
rect 204302 24967 204602 25009
rect 204302 24849 204393 24967
rect 204511 24849 204602 24967
rect 204302 7127 204602 24849
rect 204302 7009 204393 7127
rect 204511 7009 204602 7127
rect 204302 6967 204602 7009
rect 204302 6849 204393 6967
rect 204511 6849 204602 6967
rect 195302 -3581 195393 -3463
rect 195511 -3581 195602 -3463
rect 195302 -3623 195602 -3581
rect 195302 -3741 195393 -3623
rect 195511 -3741 195602 -3623
rect 195302 -3752 195602 -3741
rect 204302 -2993 204602 6849
rect 207902 352889 208202 352900
rect 207902 352771 207993 352889
rect 208111 352771 208202 352889
rect 207902 352729 208202 352771
rect 207902 352611 207993 352729
rect 208111 352611 208202 352729
rect 207902 334727 208202 352611
rect 207902 334609 207993 334727
rect 208111 334609 208202 334727
rect 207902 334567 208202 334609
rect 207902 334449 207993 334567
rect 208111 334449 208202 334567
rect 207902 316727 208202 334449
rect 207902 316609 207993 316727
rect 208111 316609 208202 316727
rect 207902 316567 208202 316609
rect 207902 316449 207993 316567
rect 208111 316449 208202 316567
rect 207902 298727 208202 316449
rect 207902 298609 207993 298727
rect 208111 298609 208202 298727
rect 207902 298567 208202 298609
rect 207902 298449 207993 298567
rect 208111 298449 208202 298567
rect 207902 280727 208202 298449
rect 207902 280609 207993 280727
rect 208111 280609 208202 280727
rect 207902 280567 208202 280609
rect 207902 280449 207993 280567
rect 208111 280449 208202 280567
rect 207902 262727 208202 280449
rect 207902 262609 207993 262727
rect 208111 262609 208202 262727
rect 207902 262567 208202 262609
rect 207902 262449 207993 262567
rect 208111 262449 208202 262567
rect 207902 244727 208202 262449
rect 207902 244609 207993 244727
rect 208111 244609 208202 244727
rect 207902 244567 208202 244609
rect 207902 244449 207993 244567
rect 208111 244449 208202 244567
rect 207902 226727 208202 244449
rect 207902 226609 207993 226727
rect 208111 226609 208202 226727
rect 207902 226567 208202 226609
rect 207902 226449 207993 226567
rect 208111 226449 208202 226567
rect 207902 208727 208202 226449
rect 207902 208609 207993 208727
rect 208111 208609 208202 208727
rect 207902 208567 208202 208609
rect 207902 208449 207993 208567
rect 208111 208449 208202 208567
rect 207902 190727 208202 208449
rect 207902 190609 207993 190727
rect 208111 190609 208202 190727
rect 207902 190567 208202 190609
rect 207902 190449 207993 190567
rect 208111 190449 208202 190567
rect 207902 172727 208202 190449
rect 207902 172609 207993 172727
rect 208111 172609 208202 172727
rect 207902 172567 208202 172609
rect 207902 172449 207993 172567
rect 208111 172449 208202 172567
rect 207902 154727 208202 172449
rect 207902 154609 207993 154727
rect 208111 154609 208202 154727
rect 207902 154567 208202 154609
rect 207902 154449 207993 154567
rect 208111 154449 208202 154567
rect 207902 136727 208202 154449
rect 207902 136609 207993 136727
rect 208111 136609 208202 136727
rect 207902 136567 208202 136609
rect 207902 136449 207993 136567
rect 208111 136449 208202 136567
rect 207902 118727 208202 136449
rect 207902 118609 207993 118727
rect 208111 118609 208202 118727
rect 207902 118567 208202 118609
rect 207902 118449 207993 118567
rect 208111 118449 208202 118567
rect 207902 100727 208202 118449
rect 207902 100609 207993 100727
rect 208111 100609 208202 100727
rect 207902 100567 208202 100609
rect 207902 100449 207993 100567
rect 208111 100449 208202 100567
rect 207902 82727 208202 100449
rect 207902 82609 207993 82727
rect 208111 82609 208202 82727
rect 207902 82567 208202 82609
rect 207902 82449 207993 82567
rect 208111 82449 208202 82567
rect 207902 64727 208202 82449
rect 207902 64609 207993 64727
rect 208111 64609 208202 64727
rect 207902 64567 208202 64609
rect 207902 64449 207993 64567
rect 208111 64449 208202 64567
rect 207902 46727 208202 64449
rect 207902 46609 207993 46727
rect 208111 46609 208202 46727
rect 207902 46567 208202 46609
rect 207902 46449 207993 46567
rect 208111 46449 208202 46567
rect 207902 28727 208202 46449
rect 207902 28609 207993 28727
rect 208111 28609 208202 28727
rect 207902 28567 208202 28609
rect 207902 28449 207993 28567
rect 208111 28449 208202 28567
rect 207902 10727 208202 28449
rect 207902 10609 207993 10727
rect 208111 10609 208202 10727
rect 207902 10567 208202 10609
rect 207902 10449 207993 10567
rect 208111 10449 208202 10567
rect 207902 -643 208202 10449
rect 207902 -761 207993 -643
rect 208111 -761 208202 -643
rect 207902 -803 208202 -761
rect 207902 -921 207993 -803
rect 208111 -921 208202 -803
rect 207902 -932 208202 -921
rect 209702 336527 210002 353551
rect 209702 336409 209793 336527
rect 209911 336409 210002 336527
rect 209702 336367 210002 336409
rect 209702 336249 209793 336367
rect 209911 336249 210002 336367
rect 209702 318527 210002 336249
rect 209702 318409 209793 318527
rect 209911 318409 210002 318527
rect 209702 318367 210002 318409
rect 209702 318249 209793 318367
rect 209911 318249 210002 318367
rect 209702 300527 210002 318249
rect 209702 300409 209793 300527
rect 209911 300409 210002 300527
rect 209702 300367 210002 300409
rect 209702 300249 209793 300367
rect 209911 300249 210002 300367
rect 209702 282527 210002 300249
rect 209702 282409 209793 282527
rect 209911 282409 210002 282527
rect 209702 282367 210002 282409
rect 209702 282249 209793 282367
rect 209911 282249 210002 282367
rect 209702 264527 210002 282249
rect 209702 264409 209793 264527
rect 209911 264409 210002 264527
rect 209702 264367 210002 264409
rect 209702 264249 209793 264367
rect 209911 264249 210002 264367
rect 209702 246527 210002 264249
rect 209702 246409 209793 246527
rect 209911 246409 210002 246527
rect 209702 246367 210002 246409
rect 209702 246249 209793 246367
rect 209911 246249 210002 246367
rect 209702 228527 210002 246249
rect 209702 228409 209793 228527
rect 209911 228409 210002 228527
rect 209702 228367 210002 228409
rect 209702 228249 209793 228367
rect 209911 228249 210002 228367
rect 209702 210527 210002 228249
rect 209702 210409 209793 210527
rect 209911 210409 210002 210527
rect 209702 210367 210002 210409
rect 209702 210249 209793 210367
rect 209911 210249 210002 210367
rect 209702 192527 210002 210249
rect 209702 192409 209793 192527
rect 209911 192409 210002 192527
rect 209702 192367 210002 192409
rect 209702 192249 209793 192367
rect 209911 192249 210002 192367
rect 209702 174527 210002 192249
rect 209702 174409 209793 174527
rect 209911 174409 210002 174527
rect 209702 174367 210002 174409
rect 209702 174249 209793 174367
rect 209911 174249 210002 174367
rect 209702 156527 210002 174249
rect 209702 156409 209793 156527
rect 209911 156409 210002 156527
rect 209702 156367 210002 156409
rect 209702 156249 209793 156367
rect 209911 156249 210002 156367
rect 209702 138527 210002 156249
rect 209702 138409 209793 138527
rect 209911 138409 210002 138527
rect 209702 138367 210002 138409
rect 209702 138249 209793 138367
rect 209911 138249 210002 138367
rect 209702 120527 210002 138249
rect 209702 120409 209793 120527
rect 209911 120409 210002 120527
rect 209702 120367 210002 120409
rect 209702 120249 209793 120367
rect 209911 120249 210002 120367
rect 209702 102527 210002 120249
rect 209702 102409 209793 102527
rect 209911 102409 210002 102527
rect 209702 102367 210002 102409
rect 209702 102249 209793 102367
rect 209911 102249 210002 102367
rect 209702 84527 210002 102249
rect 209702 84409 209793 84527
rect 209911 84409 210002 84527
rect 209702 84367 210002 84409
rect 209702 84249 209793 84367
rect 209911 84249 210002 84367
rect 209702 66527 210002 84249
rect 209702 66409 209793 66527
rect 209911 66409 210002 66527
rect 209702 66367 210002 66409
rect 209702 66249 209793 66367
rect 209911 66249 210002 66367
rect 209702 48527 210002 66249
rect 209702 48409 209793 48527
rect 209911 48409 210002 48527
rect 209702 48367 210002 48409
rect 209702 48249 209793 48367
rect 209911 48249 210002 48367
rect 209702 30527 210002 48249
rect 209702 30409 209793 30527
rect 209911 30409 210002 30527
rect 209702 30367 210002 30409
rect 209702 30249 209793 30367
rect 209911 30249 210002 30367
rect 209702 12527 210002 30249
rect 209702 12409 209793 12527
rect 209911 12409 210002 12527
rect 209702 12367 210002 12409
rect 209702 12249 209793 12367
rect 209911 12249 210002 12367
rect 209702 -1583 210002 12249
rect 209702 -1701 209793 -1583
rect 209911 -1701 210002 -1583
rect 209702 -1743 210002 -1701
rect 209702 -1861 209793 -1743
rect 209911 -1861 210002 -1743
rect 209702 -1872 210002 -1861
rect 211502 338327 211802 354491
rect 211502 338209 211593 338327
rect 211711 338209 211802 338327
rect 211502 338167 211802 338209
rect 211502 338049 211593 338167
rect 211711 338049 211802 338167
rect 211502 320327 211802 338049
rect 211502 320209 211593 320327
rect 211711 320209 211802 320327
rect 211502 320167 211802 320209
rect 211502 320049 211593 320167
rect 211711 320049 211802 320167
rect 211502 302327 211802 320049
rect 211502 302209 211593 302327
rect 211711 302209 211802 302327
rect 211502 302167 211802 302209
rect 211502 302049 211593 302167
rect 211711 302049 211802 302167
rect 211502 284327 211802 302049
rect 211502 284209 211593 284327
rect 211711 284209 211802 284327
rect 211502 284167 211802 284209
rect 211502 284049 211593 284167
rect 211711 284049 211802 284167
rect 211502 266327 211802 284049
rect 211502 266209 211593 266327
rect 211711 266209 211802 266327
rect 211502 266167 211802 266209
rect 211502 266049 211593 266167
rect 211711 266049 211802 266167
rect 211502 248327 211802 266049
rect 211502 248209 211593 248327
rect 211711 248209 211802 248327
rect 211502 248167 211802 248209
rect 211502 248049 211593 248167
rect 211711 248049 211802 248167
rect 211502 230327 211802 248049
rect 211502 230209 211593 230327
rect 211711 230209 211802 230327
rect 211502 230167 211802 230209
rect 211502 230049 211593 230167
rect 211711 230049 211802 230167
rect 211502 212327 211802 230049
rect 211502 212209 211593 212327
rect 211711 212209 211802 212327
rect 211502 212167 211802 212209
rect 211502 212049 211593 212167
rect 211711 212049 211802 212167
rect 211502 194327 211802 212049
rect 211502 194209 211593 194327
rect 211711 194209 211802 194327
rect 211502 194167 211802 194209
rect 211502 194049 211593 194167
rect 211711 194049 211802 194167
rect 211502 176327 211802 194049
rect 211502 176209 211593 176327
rect 211711 176209 211802 176327
rect 211502 176167 211802 176209
rect 211502 176049 211593 176167
rect 211711 176049 211802 176167
rect 211502 158327 211802 176049
rect 211502 158209 211593 158327
rect 211711 158209 211802 158327
rect 211502 158167 211802 158209
rect 211502 158049 211593 158167
rect 211711 158049 211802 158167
rect 211502 140327 211802 158049
rect 211502 140209 211593 140327
rect 211711 140209 211802 140327
rect 211502 140167 211802 140209
rect 211502 140049 211593 140167
rect 211711 140049 211802 140167
rect 211502 122327 211802 140049
rect 211502 122209 211593 122327
rect 211711 122209 211802 122327
rect 211502 122167 211802 122209
rect 211502 122049 211593 122167
rect 211711 122049 211802 122167
rect 211502 104327 211802 122049
rect 211502 104209 211593 104327
rect 211711 104209 211802 104327
rect 211502 104167 211802 104209
rect 211502 104049 211593 104167
rect 211711 104049 211802 104167
rect 211502 86327 211802 104049
rect 211502 86209 211593 86327
rect 211711 86209 211802 86327
rect 211502 86167 211802 86209
rect 211502 86049 211593 86167
rect 211711 86049 211802 86167
rect 211502 68327 211802 86049
rect 211502 68209 211593 68327
rect 211711 68209 211802 68327
rect 211502 68167 211802 68209
rect 211502 68049 211593 68167
rect 211711 68049 211802 68167
rect 211502 50327 211802 68049
rect 211502 50209 211593 50327
rect 211711 50209 211802 50327
rect 211502 50167 211802 50209
rect 211502 50049 211593 50167
rect 211711 50049 211802 50167
rect 211502 32327 211802 50049
rect 211502 32209 211593 32327
rect 211711 32209 211802 32327
rect 211502 32167 211802 32209
rect 211502 32049 211593 32167
rect 211711 32049 211802 32167
rect 211502 14327 211802 32049
rect 211502 14209 211593 14327
rect 211711 14209 211802 14327
rect 211502 14167 211802 14209
rect 211502 14049 211593 14167
rect 211711 14049 211802 14167
rect 211502 -2523 211802 14049
rect 211502 -2641 211593 -2523
rect 211711 -2641 211802 -2523
rect 211502 -2683 211802 -2641
rect 211502 -2801 211593 -2683
rect 211711 -2801 211802 -2683
rect 211502 -2812 211802 -2801
rect 213302 340127 213602 355431
rect 222302 355239 222602 355720
rect 222302 355121 222393 355239
rect 222511 355121 222602 355239
rect 222302 355079 222602 355121
rect 222302 354961 222393 355079
rect 222511 354961 222602 355079
rect 220502 354299 220802 354780
rect 220502 354181 220593 354299
rect 220711 354181 220802 354299
rect 220502 354139 220802 354181
rect 220502 354021 220593 354139
rect 220711 354021 220802 354139
rect 218702 353359 219002 353840
rect 218702 353241 218793 353359
rect 218911 353241 219002 353359
rect 218702 353199 219002 353241
rect 218702 353081 218793 353199
rect 218911 353081 219002 353199
rect 213302 340009 213393 340127
rect 213511 340009 213602 340127
rect 213302 339967 213602 340009
rect 213302 339849 213393 339967
rect 213511 339849 213602 339967
rect 213302 322127 213602 339849
rect 213302 322009 213393 322127
rect 213511 322009 213602 322127
rect 213302 321967 213602 322009
rect 213302 321849 213393 321967
rect 213511 321849 213602 321967
rect 213302 304127 213602 321849
rect 213302 304009 213393 304127
rect 213511 304009 213602 304127
rect 213302 303967 213602 304009
rect 213302 303849 213393 303967
rect 213511 303849 213602 303967
rect 213302 286127 213602 303849
rect 213302 286009 213393 286127
rect 213511 286009 213602 286127
rect 213302 285967 213602 286009
rect 213302 285849 213393 285967
rect 213511 285849 213602 285967
rect 213302 268127 213602 285849
rect 213302 268009 213393 268127
rect 213511 268009 213602 268127
rect 213302 267967 213602 268009
rect 213302 267849 213393 267967
rect 213511 267849 213602 267967
rect 213302 250127 213602 267849
rect 213302 250009 213393 250127
rect 213511 250009 213602 250127
rect 213302 249967 213602 250009
rect 213302 249849 213393 249967
rect 213511 249849 213602 249967
rect 213302 232127 213602 249849
rect 213302 232009 213393 232127
rect 213511 232009 213602 232127
rect 213302 231967 213602 232009
rect 213302 231849 213393 231967
rect 213511 231849 213602 231967
rect 213302 214127 213602 231849
rect 213302 214009 213393 214127
rect 213511 214009 213602 214127
rect 213302 213967 213602 214009
rect 213302 213849 213393 213967
rect 213511 213849 213602 213967
rect 213302 196127 213602 213849
rect 213302 196009 213393 196127
rect 213511 196009 213602 196127
rect 213302 195967 213602 196009
rect 213302 195849 213393 195967
rect 213511 195849 213602 195967
rect 213302 178127 213602 195849
rect 213302 178009 213393 178127
rect 213511 178009 213602 178127
rect 213302 177967 213602 178009
rect 213302 177849 213393 177967
rect 213511 177849 213602 177967
rect 213302 160127 213602 177849
rect 213302 160009 213393 160127
rect 213511 160009 213602 160127
rect 213302 159967 213602 160009
rect 213302 159849 213393 159967
rect 213511 159849 213602 159967
rect 213302 142127 213602 159849
rect 213302 142009 213393 142127
rect 213511 142009 213602 142127
rect 213302 141967 213602 142009
rect 213302 141849 213393 141967
rect 213511 141849 213602 141967
rect 213302 124127 213602 141849
rect 213302 124009 213393 124127
rect 213511 124009 213602 124127
rect 213302 123967 213602 124009
rect 213302 123849 213393 123967
rect 213511 123849 213602 123967
rect 213302 106127 213602 123849
rect 213302 106009 213393 106127
rect 213511 106009 213602 106127
rect 213302 105967 213602 106009
rect 213302 105849 213393 105967
rect 213511 105849 213602 105967
rect 213302 88127 213602 105849
rect 213302 88009 213393 88127
rect 213511 88009 213602 88127
rect 213302 87967 213602 88009
rect 213302 87849 213393 87967
rect 213511 87849 213602 87967
rect 213302 70127 213602 87849
rect 213302 70009 213393 70127
rect 213511 70009 213602 70127
rect 213302 69967 213602 70009
rect 213302 69849 213393 69967
rect 213511 69849 213602 69967
rect 213302 52127 213602 69849
rect 213302 52009 213393 52127
rect 213511 52009 213602 52127
rect 213302 51967 213602 52009
rect 213302 51849 213393 51967
rect 213511 51849 213602 51967
rect 213302 34127 213602 51849
rect 213302 34009 213393 34127
rect 213511 34009 213602 34127
rect 213302 33967 213602 34009
rect 213302 33849 213393 33967
rect 213511 33849 213602 33967
rect 213302 16127 213602 33849
rect 213302 16009 213393 16127
rect 213511 16009 213602 16127
rect 213302 15967 213602 16009
rect 213302 15849 213393 15967
rect 213511 15849 213602 15967
rect 204302 -3111 204393 -2993
rect 204511 -3111 204602 -2993
rect 204302 -3153 204602 -3111
rect 204302 -3271 204393 -3153
rect 204511 -3271 204602 -3153
rect 204302 -3752 204602 -3271
rect 213302 -3463 213602 15849
rect 216902 352419 217202 352900
rect 216902 352301 216993 352419
rect 217111 352301 217202 352419
rect 216902 352259 217202 352301
rect 216902 352141 216993 352259
rect 217111 352141 217202 352259
rect 216902 343727 217202 352141
rect 216902 343609 216993 343727
rect 217111 343609 217202 343727
rect 216902 343567 217202 343609
rect 216902 343449 216993 343567
rect 217111 343449 217202 343567
rect 216902 325727 217202 343449
rect 216902 325609 216993 325727
rect 217111 325609 217202 325727
rect 216902 325567 217202 325609
rect 216902 325449 216993 325567
rect 217111 325449 217202 325567
rect 216902 307727 217202 325449
rect 216902 307609 216993 307727
rect 217111 307609 217202 307727
rect 216902 307567 217202 307609
rect 216902 307449 216993 307567
rect 217111 307449 217202 307567
rect 216902 289727 217202 307449
rect 216902 289609 216993 289727
rect 217111 289609 217202 289727
rect 216902 289567 217202 289609
rect 216902 289449 216993 289567
rect 217111 289449 217202 289567
rect 216902 271727 217202 289449
rect 216902 271609 216993 271727
rect 217111 271609 217202 271727
rect 216902 271567 217202 271609
rect 216902 271449 216993 271567
rect 217111 271449 217202 271567
rect 216902 253727 217202 271449
rect 216902 253609 216993 253727
rect 217111 253609 217202 253727
rect 216902 253567 217202 253609
rect 216902 253449 216993 253567
rect 217111 253449 217202 253567
rect 216902 235727 217202 253449
rect 216902 235609 216993 235727
rect 217111 235609 217202 235727
rect 216902 235567 217202 235609
rect 216902 235449 216993 235567
rect 217111 235449 217202 235567
rect 216902 217727 217202 235449
rect 216902 217609 216993 217727
rect 217111 217609 217202 217727
rect 216902 217567 217202 217609
rect 216902 217449 216993 217567
rect 217111 217449 217202 217567
rect 216902 199727 217202 217449
rect 216902 199609 216993 199727
rect 217111 199609 217202 199727
rect 216902 199567 217202 199609
rect 216902 199449 216993 199567
rect 217111 199449 217202 199567
rect 216902 181727 217202 199449
rect 216902 181609 216993 181727
rect 217111 181609 217202 181727
rect 216902 181567 217202 181609
rect 216902 181449 216993 181567
rect 217111 181449 217202 181567
rect 216902 163727 217202 181449
rect 216902 163609 216993 163727
rect 217111 163609 217202 163727
rect 216902 163567 217202 163609
rect 216902 163449 216993 163567
rect 217111 163449 217202 163567
rect 216902 145727 217202 163449
rect 216902 145609 216993 145727
rect 217111 145609 217202 145727
rect 216902 145567 217202 145609
rect 216902 145449 216993 145567
rect 217111 145449 217202 145567
rect 216902 127727 217202 145449
rect 216902 127609 216993 127727
rect 217111 127609 217202 127727
rect 216902 127567 217202 127609
rect 216902 127449 216993 127567
rect 217111 127449 217202 127567
rect 216902 109727 217202 127449
rect 216902 109609 216993 109727
rect 217111 109609 217202 109727
rect 216902 109567 217202 109609
rect 216902 109449 216993 109567
rect 217111 109449 217202 109567
rect 216902 91727 217202 109449
rect 216902 91609 216993 91727
rect 217111 91609 217202 91727
rect 216902 91567 217202 91609
rect 216902 91449 216993 91567
rect 217111 91449 217202 91567
rect 216902 73727 217202 91449
rect 216902 73609 216993 73727
rect 217111 73609 217202 73727
rect 216902 73567 217202 73609
rect 216902 73449 216993 73567
rect 217111 73449 217202 73567
rect 216902 55727 217202 73449
rect 216902 55609 216993 55727
rect 217111 55609 217202 55727
rect 216902 55567 217202 55609
rect 216902 55449 216993 55567
rect 217111 55449 217202 55567
rect 216902 37727 217202 55449
rect 216902 37609 216993 37727
rect 217111 37609 217202 37727
rect 216902 37567 217202 37609
rect 216902 37449 216993 37567
rect 217111 37449 217202 37567
rect 216902 19727 217202 37449
rect 216902 19609 216993 19727
rect 217111 19609 217202 19727
rect 216902 19567 217202 19609
rect 216902 19449 216993 19567
rect 217111 19449 217202 19567
rect 216902 1727 217202 19449
rect 216902 1609 216993 1727
rect 217111 1609 217202 1727
rect 216902 1567 217202 1609
rect 216902 1449 216993 1567
rect 217111 1449 217202 1567
rect 216902 -173 217202 1449
rect 216902 -291 216993 -173
rect 217111 -291 217202 -173
rect 216902 -333 217202 -291
rect 216902 -451 216993 -333
rect 217111 -451 217202 -333
rect 216902 -932 217202 -451
rect 218702 345527 219002 353081
rect 218702 345409 218793 345527
rect 218911 345409 219002 345527
rect 218702 345367 219002 345409
rect 218702 345249 218793 345367
rect 218911 345249 219002 345367
rect 218702 327527 219002 345249
rect 218702 327409 218793 327527
rect 218911 327409 219002 327527
rect 218702 327367 219002 327409
rect 218702 327249 218793 327367
rect 218911 327249 219002 327367
rect 218702 309527 219002 327249
rect 218702 309409 218793 309527
rect 218911 309409 219002 309527
rect 218702 309367 219002 309409
rect 218702 309249 218793 309367
rect 218911 309249 219002 309367
rect 218702 291527 219002 309249
rect 218702 291409 218793 291527
rect 218911 291409 219002 291527
rect 218702 291367 219002 291409
rect 218702 291249 218793 291367
rect 218911 291249 219002 291367
rect 218702 273527 219002 291249
rect 218702 273409 218793 273527
rect 218911 273409 219002 273527
rect 218702 273367 219002 273409
rect 218702 273249 218793 273367
rect 218911 273249 219002 273367
rect 218702 255527 219002 273249
rect 218702 255409 218793 255527
rect 218911 255409 219002 255527
rect 218702 255367 219002 255409
rect 218702 255249 218793 255367
rect 218911 255249 219002 255367
rect 218702 237527 219002 255249
rect 218702 237409 218793 237527
rect 218911 237409 219002 237527
rect 218702 237367 219002 237409
rect 218702 237249 218793 237367
rect 218911 237249 219002 237367
rect 218702 219527 219002 237249
rect 218702 219409 218793 219527
rect 218911 219409 219002 219527
rect 218702 219367 219002 219409
rect 218702 219249 218793 219367
rect 218911 219249 219002 219367
rect 218702 201527 219002 219249
rect 218702 201409 218793 201527
rect 218911 201409 219002 201527
rect 218702 201367 219002 201409
rect 218702 201249 218793 201367
rect 218911 201249 219002 201367
rect 218702 183527 219002 201249
rect 218702 183409 218793 183527
rect 218911 183409 219002 183527
rect 218702 183367 219002 183409
rect 218702 183249 218793 183367
rect 218911 183249 219002 183367
rect 218702 165527 219002 183249
rect 218702 165409 218793 165527
rect 218911 165409 219002 165527
rect 218702 165367 219002 165409
rect 218702 165249 218793 165367
rect 218911 165249 219002 165367
rect 218702 147527 219002 165249
rect 218702 147409 218793 147527
rect 218911 147409 219002 147527
rect 218702 147367 219002 147409
rect 218702 147249 218793 147367
rect 218911 147249 219002 147367
rect 218702 129527 219002 147249
rect 218702 129409 218793 129527
rect 218911 129409 219002 129527
rect 218702 129367 219002 129409
rect 218702 129249 218793 129367
rect 218911 129249 219002 129367
rect 218702 111527 219002 129249
rect 218702 111409 218793 111527
rect 218911 111409 219002 111527
rect 218702 111367 219002 111409
rect 218702 111249 218793 111367
rect 218911 111249 219002 111367
rect 218702 93527 219002 111249
rect 218702 93409 218793 93527
rect 218911 93409 219002 93527
rect 218702 93367 219002 93409
rect 218702 93249 218793 93367
rect 218911 93249 219002 93367
rect 218702 75527 219002 93249
rect 218702 75409 218793 75527
rect 218911 75409 219002 75527
rect 218702 75367 219002 75409
rect 218702 75249 218793 75367
rect 218911 75249 219002 75367
rect 218702 57527 219002 75249
rect 218702 57409 218793 57527
rect 218911 57409 219002 57527
rect 218702 57367 219002 57409
rect 218702 57249 218793 57367
rect 218911 57249 219002 57367
rect 218702 39527 219002 57249
rect 218702 39409 218793 39527
rect 218911 39409 219002 39527
rect 218702 39367 219002 39409
rect 218702 39249 218793 39367
rect 218911 39249 219002 39367
rect 218702 21527 219002 39249
rect 218702 21409 218793 21527
rect 218911 21409 219002 21527
rect 218702 21367 219002 21409
rect 218702 21249 218793 21367
rect 218911 21249 219002 21367
rect 218702 3527 219002 21249
rect 218702 3409 218793 3527
rect 218911 3409 219002 3527
rect 218702 3367 219002 3409
rect 218702 3249 218793 3367
rect 218911 3249 219002 3367
rect 218702 -1113 219002 3249
rect 218702 -1231 218793 -1113
rect 218911 -1231 219002 -1113
rect 218702 -1273 219002 -1231
rect 218702 -1391 218793 -1273
rect 218911 -1391 219002 -1273
rect 218702 -1872 219002 -1391
rect 220502 347327 220802 354021
rect 220502 347209 220593 347327
rect 220711 347209 220802 347327
rect 220502 347167 220802 347209
rect 220502 347049 220593 347167
rect 220711 347049 220802 347167
rect 220502 329327 220802 347049
rect 220502 329209 220593 329327
rect 220711 329209 220802 329327
rect 220502 329167 220802 329209
rect 220502 329049 220593 329167
rect 220711 329049 220802 329167
rect 220502 311327 220802 329049
rect 220502 311209 220593 311327
rect 220711 311209 220802 311327
rect 220502 311167 220802 311209
rect 220502 311049 220593 311167
rect 220711 311049 220802 311167
rect 220502 293327 220802 311049
rect 220502 293209 220593 293327
rect 220711 293209 220802 293327
rect 220502 293167 220802 293209
rect 220502 293049 220593 293167
rect 220711 293049 220802 293167
rect 220502 275327 220802 293049
rect 220502 275209 220593 275327
rect 220711 275209 220802 275327
rect 220502 275167 220802 275209
rect 220502 275049 220593 275167
rect 220711 275049 220802 275167
rect 220502 257327 220802 275049
rect 220502 257209 220593 257327
rect 220711 257209 220802 257327
rect 220502 257167 220802 257209
rect 220502 257049 220593 257167
rect 220711 257049 220802 257167
rect 220502 239327 220802 257049
rect 220502 239209 220593 239327
rect 220711 239209 220802 239327
rect 220502 239167 220802 239209
rect 220502 239049 220593 239167
rect 220711 239049 220802 239167
rect 220502 221327 220802 239049
rect 220502 221209 220593 221327
rect 220711 221209 220802 221327
rect 220502 221167 220802 221209
rect 220502 221049 220593 221167
rect 220711 221049 220802 221167
rect 220502 203327 220802 221049
rect 220502 203209 220593 203327
rect 220711 203209 220802 203327
rect 220502 203167 220802 203209
rect 220502 203049 220593 203167
rect 220711 203049 220802 203167
rect 220502 185327 220802 203049
rect 220502 185209 220593 185327
rect 220711 185209 220802 185327
rect 220502 185167 220802 185209
rect 220502 185049 220593 185167
rect 220711 185049 220802 185167
rect 220502 167327 220802 185049
rect 220502 167209 220593 167327
rect 220711 167209 220802 167327
rect 220502 167167 220802 167209
rect 220502 167049 220593 167167
rect 220711 167049 220802 167167
rect 220502 149327 220802 167049
rect 220502 149209 220593 149327
rect 220711 149209 220802 149327
rect 220502 149167 220802 149209
rect 220502 149049 220593 149167
rect 220711 149049 220802 149167
rect 220502 131327 220802 149049
rect 220502 131209 220593 131327
rect 220711 131209 220802 131327
rect 220502 131167 220802 131209
rect 220502 131049 220593 131167
rect 220711 131049 220802 131167
rect 220502 113327 220802 131049
rect 220502 113209 220593 113327
rect 220711 113209 220802 113327
rect 220502 113167 220802 113209
rect 220502 113049 220593 113167
rect 220711 113049 220802 113167
rect 220502 95327 220802 113049
rect 220502 95209 220593 95327
rect 220711 95209 220802 95327
rect 220502 95167 220802 95209
rect 220502 95049 220593 95167
rect 220711 95049 220802 95167
rect 220502 77327 220802 95049
rect 220502 77209 220593 77327
rect 220711 77209 220802 77327
rect 220502 77167 220802 77209
rect 220502 77049 220593 77167
rect 220711 77049 220802 77167
rect 220502 59327 220802 77049
rect 220502 59209 220593 59327
rect 220711 59209 220802 59327
rect 220502 59167 220802 59209
rect 220502 59049 220593 59167
rect 220711 59049 220802 59167
rect 220502 41327 220802 59049
rect 220502 41209 220593 41327
rect 220711 41209 220802 41327
rect 220502 41167 220802 41209
rect 220502 41049 220593 41167
rect 220711 41049 220802 41167
rect 220502 23327 220802 41049
rect 220502 23209 220593 23327
rect 220711 23209 220802 23327
rect 220502 23167 220802 23209
rect 220502 23049 220593 23167
rect 220711 23049 220802 23167
rect 220502 5327 220802 23049
rect 220502 5209 220593 5327
rect 220711 5209 220802 5327
rect 220502 5167 220802 5209
rect 220502 5049 220593 5167
rect 220711 5049 220802 5167
rect 220502 -2053 220802 5049
rect 220502 -2171 220593 -2053
rect 220711 -2171 220802 -2053
rect 220502 -2213 220802 -2171
rect 220502 -2331 220593 -2213
rect 220711 -2331 220802 -2213
rect 220502 -2812 220802 -2331
rect 222302 349127 222602 354961
rect 231302 355709 231602 355720
rect 231302 355591 231393 355709
rect 231511 355591 231602 355709
rect 231302 355549 231602 355591
rect 231302 355431 231393 355549
rect 231511 355431 231602 355549
rect 229502 354769 229802 354780
rect 229502 354651 229593 354769
rect 229711 354651 229802 354769
rect 229502 354609 229802 354651
rect 229502 354491 229593 354609
rect 229711 354491 229802 354609
rect 227702 353829 228002 353840
rect 227702 353711 227793 353829
rect 227911 353711 228002 353829
rect 227702 353669 228002 353711
rect 227702 353551 227793 353669
rect 227911 353551 228002 353669
rect 222302 349009 222393 349127
rect 222511 349009 222602 349127
rect 222302 348967 222602 349009
rect 222302 348849 222393 348967
rect 222511 348849 222602 348967
rect 222302 331127 222602 348849
rect 222302 331009 222393 331127
rect 222511 331009 222602 331127
rect 222302 330967 222602 331009
rect 222302 330849 222393 330967
rect 222511 330849 222602 330967
rect 222302 313127 222602 330849
rect 222302 313009 222393 313127
rect 222511 313009 222602 313127
rect 222302 312967 222602 313009
rect 222302 312849 222393 312967
rect 222511 312849 222602 312967
rect 222302 295127 222602 312849
rect 222302 295009 222393 295127
rect 222511 295009 222602 295127
rect 222302 294967 222602 295009
rect 222302 294849 222393 294967
rect 222511 294849 222602 294967
rect 222302 277127 222602 294849
rect 222302 277009 222393 277127
rect 222511 277009 222602 277127
rect 222302 276967 222602 277009
rect 222302 276849 222393 276967
rect 222511 276849 222602 276967
rect 222302 259127 222602 276849
rect 222302 259009 222393 259127
rect 222511 259009 222602 259127
rect 222302 258967 222602 259009
rect 222302 258849 222393 258967
rect 222511 258849 222602 258967
rect 222302 241127 222602 258849
rect 222302 241009 222393 241127
rect 222511 241009 222602 241127
rect 222302 240967 222602 241009
rect 222302 240849 222393 240967
rect 222511 240849 222602 240967
rect 222302 223127 222602 240849
rect 222302 223009 222393 223127
rect 222511 223009 222602 223127
rect 222302 222967 222602 223009
rect 222302 222849 222393 222967
rect 222511 222849 222602 222967
rect 222302 205127 222602 222849
rect 222302 205009 222393 205127
rect 222511 205009 222602 205127
rect 222302 204967 222602 205009
rect 222302 204849 222393 204967
rect 222511 204849 222602 204967
rect 222302 187127 222602 204849
rect 222302 187009 222393 187127
rect 222511 187009 222602 187127
rect 222302 186967 222602 187009
rect 222302 186849 222393 186967
rect 222511 186849 222602 186967
rect 222302 169127 222602 186849
rect 222302 169009 222393 169127
rect 222511 169009 222602 169127
rect 222302 168967 222602 169009
rect 222302 168849 222393 168967
rect 222511 168849 222602 168967
rect 222302 151127 222602 168849
rect 222302 151009 222393 151127
rect 222511 151009 222602 151127
rect 222302 150967 222602 151009
rect 222302 150849 222393 150967
rect 222511 150849 222602 150967
rect 222302 133127 222602 150849
rect 222302 133009 222393 133127
rect 222511 133009 222602 133127
rect 222302 132967 222602 133009
rect 222302 132849 222393 132967
rect 222511 132849 222602 132967
rect 222302 115127 222602 132849
rect 222302 115009 222393 115127
rect 222511 115009 222602 115127
rect 222302 114967 222602 115009
rect 222302 114849 222393 114967
rect 222511 114849 222602 114967
rect 222302 97127 222602 114849
rect 222302 97009 222393 97127
rect 222511 97009 222602 97127
rect 222302 96967 222602 97009
rect 222302 96849 222393 96967
rect 222511 96849 222602 96967
rect 222302 79127 222602 96849
rect 222302 79009 222393 79127
rect 222511 79009 222602 79127
rect 222302 78967 222602 79009
rect 222302 78849 222393 78967
rect 222511 78849 222602 78967
rect 222302 61127 222602 78849
rect 222302 61009 222393 61127
rect 222511 61009 222602 61127
rect 222302 60967 222602 61009
rect 222302 60849 222393 60967
rect 222511 60849 222602 60967
rect 222302 43127 222602 60849
rect 222302 43009 222393 43127
rect 222511 43009 222602 43127
rect 222302 42967 222602 43009
rect 222302 42849 222393 42967
rect 222511 42849 222602 42967
rect 222302 25127 222602 42849
rect 222302 25009 222393 25127
rect 222511 25009 222602 25127
rect 222302 24967 222602 25009
rect 222302 24849 222393 24967
rect 222511 24849 222602 24967
rect 222302 7127 222602 24849
rect 222302 7009 222393 7127
rect 222511 7009 222602 7127
rect 222302 6967 222602 7009
rect 222302 6849 222393 6967
rect 222511 6849 222602 6967
rect 213302 -3581 213393 -3463
rect 213511 -3581 213602 -3463
rect 213302 -3623 213602 -3581
rect 213302 -3741 213393 -3623
rect 213511 -3741 213602 -3623
rect 213302 -3752 213602 -3741
rect 222302 -2993 222602 6849
rect 225902 352889 226202 352900
rect 225902 352771 225993 352889
rect 226111 352771 226202 352889
rect 225902 352729 226202 352771
rect 225902 352611 225993 352729
rect 226111 352611 226202 352729
rect 225902 334727 226202 352611
rect 225902 334609 225993 334727
rect 226111 334609 226202 334727
rect 225902 334567 226202 334609
rect 225902 334449 225993 334567
rect 226111 334449 226202 334567
rect 225902 316727 226202 334449
rect 225902 316609 225993 316727
rect 226111 316609 226202 316727
rect 225902 316567 226202 316609
rect 225902 316449 225993 316567
rect 226111 316449 226202 316567
rect 225902 298727 226202 316449
rect 225902 298609 225993 298727
rect 226111 298609 226202 298727
rect 225902 298567 226202 298609
rect 225902 298449 225993 298567
rect 226111 298449 226202 298567
rect 225902 280727 226202 298449
rect 225902 280609 225993 280727
rect 226111 280609 226202 280727
rect 225902 280567 226202 280609
rect 225902 280449 225993 280567
rect 226111 280449 226202 280567
rect 225902 262727 226202 280449
rect 225902 262609 225993 262727
rect 226111 262609 226202 262727
rect 225902 262567 226202 262609
rect 225902 262449 225993 262567
rect 226111 262449 226202 262567
rect 225902 244727 226202 262449
rect 225902 244609 225993 244727
rect 226111 244609 226202 244727
rect 225902 244567 226202 244609
rect 225902 244449 225993 244567
rect 226111 244449 226202 244567
rect 225902 226727 226202 244449
rect 225902 226609 225993 226727
rect 226111 226609 226202 226727
rect 225902 226567 226202 226609
rect 225902 226449 225993 226567
rect 226111 226449 226202 226567
rect 225902 208727 226202 226449
rect 225902 208609 225993 208727
rect 226111 208609 226202 208727
rect 225902 208567 226202 208609
rect 225902 208449 225993 208567
rect 226111 208449 226202 208567
rect 225902 190727 226202 208449
rect 225902 190609 225993 190727
rect 226111 190609 226202 190727
rect 225902 190567 226202 190609
rect 225902 190449 225993 190567
rect 226111 190449 226202 190567
rect 225902 172727 226202 190449
rect 225902 172609 225993 172727
rect 226111 172609 226202 172727
rect 225902 172567 226202 172609
rect 225902 172449 225993 172567
rect 226111 172449 226202 172567
rect 225902 154727 226202 172449
rect 225902 154609 225993 154727
rect 226111 154609 226202 154727
rect 225902 154567 226202 154609
rect 225902 154449 225993 154567
rect 226111 154449 226202 154567
rect 225902 136727 226202 154449
rect 225902 136609 225993 136727
rect 226111 136609 226202 136727
rect 225902 136567 226202 136609
rect 225902 136449 225993 136567
rect 226111 136449 226202 136567
rect 225902 118727 226202 136449
rect 225902 118609 225993 118727
rect 226111 118609 226202 118727
rect 225902 118567 226202 118609
rect 225902 118449 225993 118567
rect 226111 118449 226202 118567
rect 225902 100727 226202 118449
rect 225902 100609 225993 100727
rect 226111 100609 226202 100727
rect 225902 100567 226202 100609
rect 225902 100449 225993 100567
rect 226111 100449 226202 100567
rect 225902 82727 226202 100449
rect 225902 82609 225993 82727
rect 226111 82609 226202 82727
rect 225902 82567 226202 82609
rect 225902 82449 225993 82567
rect 226111 82449 226202 82567
rect 225902 64727 226202 82449
rect 225902 64609 225993 64727
rect 226111 64609 226202 64727
rect 225902 64567 226202 64609
rect 225902 64449 225993 64567
rect 226111 64449 226202 64567
rect 225902 46727 226202 64449
rect 225902 46609 225993 46727
rect 226111 46609 226202 46727
rect 225902 46567 226202 46609
rect 225902 46449 225993 46567
rect 226111 46449 226202 46567
rect 225902 28727 226202 46449
rect 225902 28609 225993 28727
rect 226111 28609 226202 28727
rect 225902 28567 226202 28609
rect 225902 28449 225993 28567
rect 226111 28449 226202 28567
rect 225902 10727 226202 28449
rect 225902 10609 225993 10727
rect 226111 10609 226202 10727
rect 225902 10567 226202 10609
rect 225902 10449 225993 10567
rect 226111 10449 226202 10567
rect 225902 -643 226202 10449
rect 225902 -761 225993 -643
rect 226111 -761 226202 -643
rect 225902 -803 226202 -761
rect 225902 -921 225993 -803
rect 226111 -921 226202 -803
rect 225902 -932 226202 -921
rect 227702 336527 228002 353551
rect 227702 336409 227793 336527
rect 227911 336409 228002 336527
rect 227702 336367 228002 336409
rect 227702 336249 227793 336367
rect 227911 336249 228002 336367
rect 227702 318527 228002 336249
rect 227702 318409 227793 318527
rect 227911 318409 228002 318527
rect 227702 318367 228002 318409
rect 227702 318249 227793 318367
rect 227911 318249 228002 318367
rect 227702 300527 228002 318249
rect 227702 300409 227793 300527
rect 227911 300409 228002 300527
rect 227702 300367 228002 300409
rect 227702 300249 227793 300367
rect 227911 300249 228002 300367
rect 227702 282527 228002 300249
rect 227702 282409 227793 282527
rect 227911 282409 228002 282527
rect 227702 282367 228002 282409
rect 227702 282249 227793 282367
rect 227911 282249 228002 282367
rect 227702 264527 228002 282249
rect 227702 264409 227793 264527
rect 227911 264409 228002 264527
rect 227702 264367 228002 264409
rect 227702 264249 227793 264367
rect 227911 264249 228002 264367
rect 227702 246527 228002 264249
rect 227702 246409 227793 246527
rect 227911 246409 228002 246527
rect 227702 246367 228002 246409
rect 227702 246249 227793 246367
rect 227911 246249 228002 246367
rect 227702 228527 228002 246249
rect 227702 228409 227793 228527
rect 227911 228409 228002 228527
rect 227702 228367 228002 228409
rect 227702 228249 227793 228367
rect 227911 228249 228002 228367
rect 227702 210527 228002 228249
rect 227702 210409 227793 210527
rect 227911 210409 228002 210527
rect 227702 210367 228002 210409
rect 227702 210249 227793 210367
rect 227911 210249 228002 210367
rect 227702 192527 228002 210249
rect 227702 192409 227793 192527
rect 227911 192409 228002 192527
rect 227702 192367 228002 192409
rect 227702 192249 227793 192367
rect 227911 192249 228002 192367
rect 227702 174527 228002 192249
rect 227702 174409 227793 174527
rect 227911 174409 228002 174527
rect 227702 174367 228002 174409
rect 227702 174249 227793 174367
rect 227911 174249 228002 174367
rect 227702 156527 228002 174249
rect 227702 156409 227793 156527
rect 227911 156409 228002 156527
rect 227702 156367 228002 156409
rect 227702 156249 227793 156367
rect 227911 156249 228002 156367
rect 227702 138527 228002 156249
rect 227702 138409 227793 138527
rect 227911 138409 228002 138527
rect 227702 138367 228002 138409
rect 227702 138249 227793 138367
rect 227911 138249 228002 138367
rect 227702 120527 228002 138249
rect 227702 120409 227793 120527
rect 227911 120409 228002 120527
rect 227702 120367 228002 120409
rect 227702 120249 227793 120367
rect 227911 120249 228002 120367
rect 227702 102527 228002 120249
rect 227702 102409 227793 102527
rect 227911 102409 228002 102527
rect 227702 102367 228002 102409
rect 227702 102249 227793 102367
rect 227911 102249 228002 102367
rect 227702 84527 228002 102249
rect 227702 84409 227793 84527
rect 227911 84409 228002 84527
rect 227702 84367 228002 84409
rect 227702 84249 227793 84367
rect 227911 84249 228002 84367
rect 227702 66527 228002 84249
rect 227702 66409 227793 66527
rect 227911 66409 228002 66527
rect 227702 66367 228002 66409
rect 227702 66249 227793 66367
rect 227911 66249 228002 66367
rect 227702 48527 228002 66249
rect 227702 48409 227793 48527
rect 227911 48409 228002 48527
rect 227702 48367 228002 48409
rect 227702 48249 227793 48367
rect 227911 48249 228002 48367
rect 227702 30527 228002 48249
rect 227702 30409 227793 30527
rect 227911 30409 228002 30527
rect 227702 30367 228002 30409
rect 227702 30249 227793 30367
rect 227911 30249 228002 30367
rect 227702 12527 228002 30249
rect 227702 12409 227793 12527
rect 227911 12409 228002 12527
rect 227702 12367 228002 12409
rect 227702 12249 227793 12367
rect 227911 12249 228002 12367
rect 227702 -1583 228002 12249
rect 227702 -1701 227793 -1583
rect 227911 -1701 228002 -1583
rect 227702 -1743 228002 -1701
rect 227702 -1861 227793 -1743
rect 227911 -1861 228002 -1743
rect 227702 -1872 228002 -1861
rect 229502 338327 229802 354491
rect 229502 338209 229593 338327
rect 229711 338209 229802 338327
rect 229502 338167 229802 338209
rect 229502 338049 229593 338167
rect 229711 338049 229802 338167
rect 229502 320327 229802 338049
rect 229502 320209 229593 320327
rect 229711 320209 229802 320327
rect 229502 320167 229802 320209
rect 229502 320049 229593 320167
rect 229711 320049 229802 320167
rect 229502 302327 229802 320049
rect 229502 302209 229593 302327
rect 229711 302209 229802 302327
rect 229502 302167 229802 302209
rect 229502 302049 229593 302167
rect 229711 302049 229802 302167
rect 229502 284327 229802 302049
rect 229502 284209 229593 284327
rect 229711 284209 229802 284327
rect 229502 284167 229802 284209
rect 229502 284049 229593 284167
rect 229711 284049 229802 284167
rect 229502 266327 229802 284049
rect 229502 266209 229593 266327
rect 229711 266209 229802 266327
rect 229502 266167 229802 266209
rect 229502 266049 229593 266167
rect 229711 266049 229802 266167
rect 229502 248327 229802 266049
rect 229502 248209 229593 248327
rect 229711 248209 229802 248327
rect 229502 248167 229802 248209
rect 229502 248049 229593 248167
rect 229711 248049 229802 248167
rect 229502 230327 229802 248049
rect 229502 230209 229593 230327
rect 229711 230209 229802 230327
rect 229502 230167 229802 230209
rect 229502 230049 229593 230167
rect 229711 230049 229802 230167
rect 229502 212327 229802 230049
rect 229502 212209 229593 212327
rect 229711 212209 229802 212327
rect 229502 212167 229802 212209
rect 229502 212049 229593 212167
rect 229711 212049 229802 212167
rect 229502 194327 229802 212049
rect 229502 194209 229593 194327
rect 229711 194209 229802 194327
rect 229502 194167 229802 194209
rect 229502 194049 229593 194167
rect 229711 194049 229802 194167
rect 229502 176327 229802 194049
rect 229502 176209 229593 176327
rect 229711 176209 229802 176327
rect 229502 176167 229802 176209
rect 229502 176049 229593 176167
rect 229711 176049 229802 176167
rect 229502 158327 229802 176049
rect 229502 158209 229593 158327
rect 229711 158209 229802 158327
rect 229502 158167 229802 158209
rect 229502 158049 229593 158167
rect 229711 158049 229802 158167
rect 229502 140327 229802 158049
rect 229502 140209 229593 140327
rect 229711 140209 229802 140327
rect 229502 140167 229802 140209
rect 229502 140049 229593 140167
rect 229711 140049 229802 140167
rect 229502 122327 229802 140049
rect 229502 122209 229593 122327
rect 229711 122209 229802 122327
rect 229502 122167 229802 122209
rect 229502 122049 229593 122167
rect 229711 122049 229802 122167
rect 229502 104327 229802 122049
rect 229502 104209 229593 104327
rect 229711 104209 229802 104327
rect 229502 104167 229802 104209
rect 229502 104049 229593 104167
rect 229711 104049 229802 104167
rect 229502 86327 229802 104049
rect 229502 86209 229593 86327
rect 229711 86209 229802 86327
rect 229502 86167 229802 86209
rect 229502 86049 229593 86167
rect 229711 86049 229802 86167
rect 229502 68327 229802 86049
rect 229502 68209 229593 68327
rect 229711 68209 229802 68327
rect 229502 68167 229802 68209
rect 229502 68049 229593 68167
rect 229711 68049 229802 68167
rect 229502 50327 229802 68049
rect 229502 50209 229593 50327
rect 229711 50209 229802 50327
rect 229502 50167 229802 50209
rect 229502 50049 229593 50167
rect 229711 50049 229802 50167
rect 229502 32327 229802 50049
rect 229502 32209 229593 32327
rect 229711 32209 229802 32327
rect 229502 32167 229802 32209
rect 229502 32049 229593 32167
rect 229711 32049 229802 32167
rect 229502 14327 229802 32049
rect 229502 14209 229593 14327
rect 229711 14209 229802 14327
rect 229502 14167 229802 14209
rect 229502 14049 229593 14167
rect 229711 14049 229802 14167
rect 229502 -2523 229802 14049
rect 229502 -2641 229593 -2523
rect 229711 -2641 229802 -2523
rect 229502 -2683 229802 -2641
rect 229502 -2801 229593 -2683
rect 229711 -2801 229802 -2683
rect 229502 -2812 229802 -2801
rect 231302 340127 231602 355431
rect 240302 355239 240602 355720
rect 240302 355121 240393 355239
rect 240511 355121 240602 355239
rect 240302 355079 240602 355121
rect 240302 354961 240393 355079
rect 240511 354961 240602 355079
rect 238502 354299 238802 354780
rect 238502 354181 238593 354299
rect 238711 354181 238802 354299
rect 238502 354139 238802 354181
rect 238502 354021 238593 354139
rect 238711 354021 238802 354139
rect 236702 353359 237002 353840
rect 236702 353241 236793 353359
rect 236911 353241 237002 353359
rect 236702 353199 237002 353241
rect 236702 353081 236793 353199
rect 236911 353081 237002 353199
rect 231302 340009 231393 340127
rect 231511 340009 231602 340127
rect 231302 339967 231602 340009
rect 231302 339849 231393 339967
rect 231511 339849 231602 339967
rect 231302 322127 231602 339849
rect 231302 322009 231393 322127
rect 231511 322009 231602 322127
rect 231302 321967 231602 322009
rect 231302 321849 231393 321967
rect 231511 321849 231602 321967
rect 231302 304127 231602 321849
rect 231302 304009 231393 304127
rect 231511 304009 231602 304127
rect 231302 303967 231602 304009
rect 231302 303849 231393 303967
rect 231511 303849 231602 303967
rect 231302 286127 231602 303849
rect 231302 286009 231393 286127
rect 231511 286009 231602 286127
rect 231302 285967 231602 286009
rect 231302 285849 231393 285967
rect 231511 285849 231602 285967
rect 231302 268127 231602 285849
rect 231302 268009 231393 268127
rect 231511 268009 231602 268127
rect 231302 267967 231602 268009
rect 231302 267849 231393 267967
rect 231511 267849 231602 267967
rect 231302 250127 231602 267849
rect 231302 250009 231393 250127
rect 231511 250009 231602 250127
rect 231302 249967 231602 250009
rect 231302 249849 231393 249967
rect 231511 249849 231602 249967
rect 231302 232127 231602 249849
rect 231302 232009 231393 232127
rect 231511 232009 231602 232127
rect 231302 231967 231602 232009
rect 231302 231849 231393 231967
rect 231511 231849 231602 231967
rect 231302 214127 231602 231849
rect 231302 214009 231393 214127
rect 231511 214009 231602 214127
rect 231302 213967 231602 214009
rect 231302 213849 231393 213967
rect 231511 213849 231602 213967
rect 231302 196127 231602 213849
rect 231302 196009 231393 196127
rect 231511 196009 231602 196127
rect 231302 195967 231602 196009
rect 231302 195849 231393 195967
rect 231511 195849 231602 195967
rect 231302 178127 231602 195849
rect 231302 178009 231393 178127
rect 231511 178009 231602 178127
rect 231302 177967 231602 178009
rect 231302 177849 231393 177967
rect 231511 177849 231602 177967
rect 231302 160127 231602 177849
rect 231302 160009 231393 160127
rect 231511 160009 231602 160127
rect 231302 159967 231602 160009
rect 231302 159849 231393 159967
rect 231511 159849 231602 159967
rect 231302 142127 231602 159849
rect 231302 142009 231393 142127
rect 231511 142009 231602 142127
rect 231302 141967 231602 142009
rect 231302 141849 231393 141967
rect 231511 141849 231602 141967
rect 231302 124127 231602 141849
rect 231302 124009 231393 124127
rect 231511 124009 231602 124127
rect 231302 123967 231602 124009
rect 231302 123849 231393 123967
rect 231511 123849 231602 123967
rect 231302 106127 231602 123849
rect 231302 106009 231393 106127
rect 231511 106009 231602 106127
rect 231302 105967 231602 106009
rect 231302 105849 231393 105967
rect 231511 105849 231602 105967
rect 231302 88127 231602 105849
rect 231302 88009 231393 88127
rect 231511 88009 231602 88127
rect 231302 87967 231602 88009
rect 231302 87849 231393 87967
rect 231511 87849 231602 87967
rect 231302 70127 231602 87849
rect 231302 70009 231393 70127
rect 231511 70009 231602 70127
rect 231302 69967 231602 70009
rect 231302 69849 231393 69967
rect 231511 69849 231602 69967
rect 231302 52127 231602 69849
rect 231302 52009 231393 52127
rect 231511 52009 231602 52127
rect 231302 51967 231602 52009
rect 231302 51849 231393 51967
rect 231511 51849 231602 51967
rect 231302 34127 231602 51849
rect 231302 34009 231393 34127
rect 231511 34009 231602 34127
rect 231302 33967 231602 34009
rect 231302 33849 231393 33967
rect 231511 33849 231602 33967
rect 231302 16127 231602 33849
rect 231302 16009 231393 16127
rect 231511 16009 231602 16127
rect 231302 15967 231602 16009
rect 231302 15849 231393 15967
rect 231511 15849 231602 15967
rect 222302 -3111 222393 -2993
rect 222511 -3111 222602 -2993
rect 222302 -3153 222602 -3111
rect 222302 -3271 222393 -3153
rect 222511 -3271 222602 -3153
rect 222302 -3752 222602 -3271
rect 231302 -3463 231602 15849
rect 234902 352419 235202 352900
rect 234902 352301 234993 352419
rect 235111 352301 235202 352419
rect 234902 352259 235202 352301
rect 234902 352141 234993 352259
rect 235111 352141 235202 352259
rect 234902 343727 235202 352141
rect 234902 343609 234993 343727
rect 235111 343609 235202 343727
rect 234902 343567 235202 343609
rect 234902 343449 234993 343567
rect 235111 343449 235202 343567
rect 234902 325727 235202 343449
rect 234902 325609 234993 325727
rect 235111 325609 235202 325727
rect 234902 325567 235202 325609
rect 234902 325449 234993 325567
rect 235111 325449 235202 325567
rect 234902 307727 235202 325449
rect 234902 307609 234993 307727
rect 235111 307609 235202 307727
rect 234902 307567 235202 307609
rect 234902 307449 234993 307567
rect 235111 307449 235202 307567
rect 234902 289727 235202 307449
rect 234902 289609 234993 289727
rect 235111 289609 235202 289727
rect 234902 289567 235202 289609
rect 234902 289449 234993 289567
rect 235111 289449 235202 289567
rect 234902 271727 235202 289449
rect 234902 271609 234993 271727
rect 235111 271609 235202 271727
rect 234902 271567 235202 271609
rect 234902 271449 234993 271567
rect 235111 271449 235202 271567
rect 234902 253727 235202 271449
rect 234902 253609 234993 253727
rect 235111 253609 235202 253727
rect 234902 253567 235202 253609
rect 234902 253449 234993 253567
rect 235111 253449 235202 253567
rect 234902 235727 235202 253449
rect 234902 235609 234993 235727
rect 235111 235609 235202 235727
rect 234902 235567 235202 235609
rect 234902 235449 234993 235567
rect 235111 235449 235202 235567
rect 234902 217727 235202 235449
rect 234902 217609 234993 217727
rect 235111 217609 235202 217727
rect 234902 217567 235202 217609
rect 234902 217449 234993 217567
rect 235111 217449 235202 217567
rect 234902 199727 235202 217449
rect 234902 199609 234993 199727
rect 235111 199609 235202 199727
rect 234902 199567 235202 199609
rect 234902 199449 234993 199567
rect 235111 199449 235202 199567
rect 234902 181727 235202 199449
rect 234902 181609 234993 181727
rect 235111 181609 235202 181727
rect 234902 181567 235202 181609
rect 234902 181449 234993 181567
rect 235111 181449 235202 181567
rect 234902 163727 235202 181449
rect 234902 163609 234993 163727
rect 235111 163609 235202 163727
rect 234902 163567 235202 163609
rect 234902 163449 234993 163567
rect 235111 163449 235202 163567
rect 234902 145727 235202 163449
rect 234902 145609 234993 145727
rect 235111 145609 235202 145727
rect 234902 145567 235202 145609
rect 234902 145449 234993 145567
rect 235111 145449 235202 145567
rect 234902 127727 235202 145449
rect 234902 127609 234993 127727
rect 235111 127609 235202 127727
rect 234902 127567 235202 127609
rect 234902 127449 234993 127567
rect 235111 127449 235202 127567
rect 234902 109727 235202 127449
rect 234902 109609 234993 109727
rect 235111 109609 235202 109727
rect 234902 109567 235202 109609
rect 234902 109449 234993 109567
rect 235111 109449 235202 109567
rect 234902 91727 235202 109449
rect 234902 91609 234993 91727
rect 235111 91609 235202 91727
rect 234902 91567 235202 91609
rect 234902 91449 234993 91567
rect 235111 91449 235202 91567
rect 234902 73727 235202 91449
rect 234902 73609 234993 73727
rect 235111 73609 235202 73727
rect 234902 73567 235202 73609
rect 234902 73449 234993 73567
rect 235111 73449 235202 73567
rect 234902 55727 235202 73449
rect 234902 55609 234993 55727
rect 235111 55609 235202 55727
rect 234902 55567 235202 55609
rect 234902 55449 234993 55567
rect 235111 55449 235202 55567
rect 234902 37727 235202 55449
rect 234902 37609 234993 37727
rect 235111 37609 235202 37727
rect 234902 37567 235202 37609
rect 234902 37449 234993 37567
rect 235111 37449 235202 37567
rect 234902 19727 235202 37449
rect 234902 19609 234993 19727
rect 235111 19609 235202 19727
rect 234902 19567 235202 19609
rect 234902 19449 234993 19567
rect 235111 19449 235202 19567
rect 234902 1727 235202 19449
rect 234902 1609 234993 1727
rect 235111 1609 235202 1727
rect 234902 1567 235202 1609
rect 234902 1449 234993 1567
rect 235111 1449 235202 1567
rect 234902 -173 235202 1449
rect 234902 -291 234993 -173
rect 235111 -291 235202 -173
rect 234902 -333 235202 -291
rect 234902 -451 234993 -333
rect 235111 -451 235202 -333
rect 234902 -932 235202 -451
rect 236702 345527 237002 353081
rect 236702 345409 236793 345527
rect 236911 345409 237002 345527
rect 236702 345367 237002 345409
rect 236702 345249 236793 345367
rect 236911 345249 237002 345367
rect 236702 327527 237002 345249
rect 236702 327409 236793 327527
rect 236911 327409 237002 327527
rect 236702 327367 237002 327409
rect 236702 327249 236793 327367
rect 236911 327249 237002 327367
rect 236702 309527 237002 327249
rect 236702 309409 236793 309527
rect 236911 309409 237002 309527
rect 236702 309367 237002 309409
rect 236702 309249 236793 309367
rect 236911 309249 237002 309367
rect 236702 291527 237002 309249
rect 236702 291409 236793 291527
rect 236911 291409 237002 291527
rect 236702 291367 237002 291409
rect 236702 291249 236793 291367
rect 236911 291249 237002 291367
rect 236702 273527 237002 291249
rect 236702 273409 236793 273527
rect 236911 273409 237002 273527
rect 236702 273367 237002 273409
rect 236702 273249 236793 273367
rect 236911 273249 237002 273367
rect 236702 255527 237002 273249
rect 236702 255409 236793 255527
rect 236911 255409 237002 255527
rect 236702 255367 237002 255409
rect 236702 255249 236793 255367
rect 236911 255249 237002 255367
rect 236702 237527 237002 255249
rect 236702 237409 236793 237527
rect 236911 237409 237002 237527
rect 236702 237367 237002 237409
rect 236702 237249 236793 237367
rect 236911 237249 237002 237367
rect 236702 219527 237002 237249
rect 236702 219409 236793 219527
rect 236911 219409 237002 219527
rect 236702 219367 237002 219409
rect 236702 219249 236793 219367
rect 236911 219249 237002 219367
rect 236702 201527 237002 219249
rect 236702 201409 236793 201527
rect 236911 201409 237002 201527
rect 236702 201367 237002 201409
rect 236702 201249 236793 201367
rect 236911 201249 237002 201367
rect 236702 183527 237002 201249
rect 236702 183409 236793 183527
rect 236911 183409 237002 183527
rect 236702 183367 237002 183409
rect 236702 183249 236793 183367
rect 236911 183249 237002 183367
rect 236702 165527 237002 183249
rect 236702 165409 236793 165527
rect 236911 165409 237002 165527
rect 236702 165367 237002 165409
rect 236702 165249 236793 165367
rect 236911 165249 237002 165367
rect 236702 147527 237002 165249
rect 236702 147409 236793 147527
rect 236911 147409 237002 147527
rect 236702 147367 237002 147409
rect 236702 147249 236793 147367
rect 236911 147249 237002 147367
rect 236702 129527 237002 147249
rect 236702 129409 236793 129527
rect 236911 129409 237002 129527
rect 236702 129367 237002 129409
rect 236702 129249 236793 129367
rect 236911 129249 237002 129367
rect 236702 111527 237002 129249
rect 236702 111409 236793 111527
rect 236911 111409 237002 111527
rect 236702 111367 237002 111409
rect 236702 111249 236793 111367
rect 236911 111249 237002 111367
rect 236702 93527 237002 111249
rect 236702 93409 236793 93527
rect 236911 93409 237002 93527
rect 236702 93367 237002 93409
rect 236702 93249 236793 93367
rect 236911 93249 237002 93367
rect 236702 75527 237002 93249
rect 236702 75409 236793 75527
rect 236911 75409 237002 75527
rect 236702 75367 237002 75409
rect 236702 75249 236793 75367
rect 236911 75249 237002 75367
rect 236702 57527 237002 75249
rect 236702 57409 236793 57527
rect 236911 57409 237002 57527
rect 236702 57367 237002 57409
rect 236702 57249 236793 57367
rect 236911 57249 237002 57367
rect 236702 39527 237002 57249
rect 236702 39409 236793 39527
rect 236911 39409 237002 39527
rect 236702 39367 237002 39409
rect 236702 39249 236793 39367
rect 236911 39249 237002 39367
rect 236702 21527 237002 39249
rect 236702 21409 236793 21527
rect 236911 21409 237002 21527
rect 236702 21367 237002 21409
rect 236702 21249 236793 21367
rect 236911 21249 237002 21367
rect 236702 3527 237002 21249
rect 236702 3409 236793 3527
rect 236911 3409 237002 3527
rect 236702 3367 237002 3409
rect 236702 3249 236793 3367
rect 236911 3249 237002 3367
rect 236702 -1113 237002 3249
rect 236702 -1231 236793 -1113
rect 236911 -1231 237002 -1113
rect 236702 -1273 237002 -1231
rect 236702 -1391 236793 -1273
rect 236911 -1391 237002 -1273
rect 236702 -1872 237002 -1391
rect 238502 347327 238802 354021
rect 238502 347209 238593 347327
rect 238711 347209 238802 347327
rect 238502 347167 238802 347209
rect 238502 347049 238593 347167
rect 238711 347049 238802 347167
rect 238502 329327 238802 347049
rect 238502 329209 238593 329327
rect 238711 329209 238802 329327
rect 238502 329167 238802 329209
rect 238502 329049 238593 329167
rect 238711 329049 238802 329167
rect 238502 311327 238802 329049
rect 238502 311209 238593 311327
rect 238711 311209 238802 311327
rect 238502 311167 238802 311209
rect 238502 311049 238593 311167
rect 238711 311049 238802 311167
rect 238502 293327 238802 311049
rect 238502 293209 238593 293327
rect 238711 293209 238802 293327
rect 238502 293167 238802 293209
rect 238502 293049 238593 293167
rect 238711 293049 238802 293167
rect 238502 275327 238802 293049
rect 238502 275209 238593 275327
rect 238711 275209 238802 275327
rect 238502 275167 238802 275209
rect 238502 275049 238593 275167
rect 238711 275049 238802 275167
rect 238502 257327 238802 275049
rect 238502 257209 238593 257327
rect 238711 257209 238802 257327
rect 238502 257167 238802 257209
rect 238502 257049 238593 257167
rect 238711 257049 238802 257167
rect 238502 239327 238802 257049
rect 238502 239209 238593 239327
rect 238711 239209 238802 239327
rect 238502 239167 238802 239209
rect 238502 239049 238593 239167
rect 238711 239049 238802 239167
rect 238502 221327 238802 239049
rect 238502 221209 238593 221327
rect 238711 221209 238802 221327
rect 238502 221167 238802 221209
rect 238502 221049 238593 221167
rect 238711 221049 238802 221167
rect 238502 203327 238802 221049
rect 238502 203209 238593 203327
rect 238711 203209 238802 203327
rect 238502 203167 238802 203209
rect 238502 203049 238593 203167
rect 238711 203049 238802 203167
rect 238502 185327 238802 203049
rect 238502 185209 238593 185327
rect 238711 185209 238802 185327
rect 238502 185167 238802 185209
rect 238502 185049 238593 185167
rect 238711 185049 238802 185167
rect 238502 167327 238802 185049
rect 238502 167209 238593 167327
rect 238711 167209 238802 167327
rect 238502 167167 238802 167209
rect 238502 167049 238593 167167
rect 238711 167049 238802 167167
rect 238502 149327 238802 167049
rect 238502 149209 238593 149327
rect 238711 149209 238802 149327
rect 238502 149167 238802 149209
rect 238502 149049 238593 149167
rect 238711 149049 238802 149167
rect 238502 131327 238802 149049
rect 238502 131209 238593 131327
rect 238711 131209 238802 131327
rect 238502 131167 238802 131209
rect 238502 131049 238593 131167
rect 238711 131049 238802 131167
rect 238502 113327 238802 131049
rect 238502 113209 238593 113327
rect 238711 113209 238802 113327
rect 238502 113167 238802 113209
rect 238502 113049 238593 113167
rect 238711 113049 238802 113167
rect 238502 95327 238802 113049
rect 238502 95209 238593 95327
rect 238711 95209 238802 95327
rect 238502 95167 238802 95209
rect 238502 95049 238593 95167
rect 238711 95049 238802 95167
rect 238502 77327 238802 95049
rect 238502 77209 238593 77327
rect 238711 77209 238802 77327
rect 238502 77167 238802 77209
rect 238502 77049 238593 77167
rect 238711 77049 238802 77167
rect 238502 59327 238802 77049
rect 238502 59209 238593 59327
rect 238711 59209 238802 59327
rect 238502 59167 238802 59209
rect 238502 59049 238593 59167
rect 238711 59049 238802 59167
rect 238502 41327 238802 59049
rect 238502 41209 238593 41327
rect 238711 41209 238802 41327
rect 238502 41167 238802 41209
rect 238502 41049 238593 41167
rect 238711 41049 238802 41167
rect 238502 23327 238802 41049
rect 238502 23209 238593 23327
rect 238711 23209 238802 23327
rect 238502 23167 238802 23209
rect 238502 23049 238593 23167
rect 238711 23049 238802 23167
rect 238502 5327 238802 23049
rect 238502 5209 238593 5327
rect 238711 5209 238802 5327
rect 238502 5167 238802 5209
rect 238502 5049 238593 5167
rect 238711 5049 238802 5167
rect 238502 -2053 238802 5049
rect 238502 -2171 238593 -2053
rect 238711 -2171 238802 -2053
rect 238502 -2213 238802 -2171
rect 238502 -2331 238593 -2213
rect 238711 -2331 238802 -2213
rect 238502 -2812 238802 -2331
rect 240302 349127 240602 354961
rect 249302 355709 249602 355720
rect 249302 355591 249393 355709
rect 249511 355591 249602 355709
rect 249302 355549 249602 355591
rect 249302 355431 249393 355549
rect 249511 355431 249602 355549
rect 247502 354769 247802 354780
rect 247502 354651 247593 354769
rect 247711 354651 247802 354769
rect 247502 354609 247802 354651
rect 247502 354491 247593 354609
rect 247711 354491 247802 354609
rect 245702 353829 246002 353840
rect 245702 353711 245793 353829
rect 245911 353711 246002 353829
rect 245702 353669 246002 353711
rect 245702 353551 245793 353669
rect 245911 353551 246002 353669
rect 240302 349009 240393 349127
rect 240511 349009 240602 349127
rect 240302 348967 240602 349009
rect 240302 348849 240393 348967
rect 240511 348849 240602 348967
rect 240302 331127 240602 348849
rect 240302 331009 240393 331127
rect 240511 331009 240602 331127
rect 240302 330967 240602 331009
rect 240302 330849 240393 330967
rect 240511 330849 240602 330967
rect 240302 313127 240602 330849
rect 240302 313009 240393 313127
rect 240511 313009 240602 313127
rect 240302 312967 240602 313009
rect 240302 312849 240393 312967
rect 240511 312849 240602 312967
rect 240302 295127 240602 312849
rect 240302 295009 240393 295127
rect 240511 295009 240602 295127
rect 240302 294967 240602 295009
rect 240302 294849 240393 294967
rect 240511 294849 240602 294967
rect 240302 277127 240602 294849
rect 240302 277009 240393 277127
rect 240511 277009 240602 277127
rect 240302 276967 240602 277009
rect 240302 276849 240393 276967
rect 240511 276849 240602 276967
rect 240302 259127 240602 276849
rect 240302 259009 240393 259127
rect 240511 259009 240602 259127
rect 240302 258967 240602 259009
rect 240302 258849 240393 258967
rect 240511 258849 240602 258967
rect 240302 241127 240602 258849
rect 240302 241009 240393 241127
rect 240511 241009 240602 241127
rect 240302 240967 240602 241009
rect 240302 240849 240393 240967
rect 240511 240849 240602 240967
rect 240302 223127 240602 240849
rect 240302 223009 240393 223127
rect 240511 223009 240602 223127
rect 240302 222967 240602 223009
rect 240302 222849 240393 222967
rect 240511 222849 240602 222967
rect 240302 205127 240602 222849
rect 240302 205009 240393 205127
rect 240511 205009 240602 205127
rect 240302 204967 240602 205009
rect 240302 204849 240393 204967
rect 240511 204849 240602 204967
rect 240302 187127 240602 204849
rect 240302 187009 240393 187127
rect 240511 187009 240602 187127
rect 240302 186967 240602 187009
rect 240302 186849 240393 186967
rect 240511 186849 240602 186967
rect 240302 169127 240602 186849
rect 240302 169009 240393 169127
rect 240511 169009 240602 169127
rect 240302 168967 240602 169009
rect 240302 168849 240393 168967
rect 240511 168849 240602 168967
rect 240302 151127 240602 168849
rect 240302 151009 240393 151127
rect 240511 151009 240602 151127
rect 240302 150967 240602 151009
rect 240302 150849 240393 150967
rect 240511 150849 240602 150967
rect 240302 133127 240602 150849
rect 240302 133009 240393 133127
rect 240511 133009 240602 133127
rect 240302 132967 240602 133009
rect 240302 132849 240393 132967
rect 240511 132849 240602 132967
rect 240302 115127 240602 132849
rect 240302 115009 240393 115127
rect 240511 115009 240602 115127
rect 240302 114967 240602 115009
rect 240302 114849 240393 114967
rect 240511 114849 240602 114967
rect 240302 97127 240602 114849
rect 240302 97009 240393 97127
rect 240511 97009 240602 97127
rect 240302 96967 240602 97009
rect 240302 96849 240393 96967
rect 240511 96849 240602 96967
rect 240302 79127 240602 96849
rect 240302 79009 240393 79127
rect 240511 79009 240602 79127
rect 240302 78967 240602 79009
rect 240302 78849 240393 78967
rect 240511 78849 240602 78967
rect 240302 61127 240602 78849
rect 240302 61009 240393 61127
rect 240511 61009 240602 61127
rect 240302 60967 240602 61009
rect 240302 60849 240393 60967
rect 240511 60849 240602 60967
rect 240302 43127 240602 60849
rect 240302 43009 240393 43127
rect 240511 43009 240602 43127
rect 240302 42967 240602 43009
rect 240302 42849 240393 42967
rect 240511 42849 240602 42967
rect 240302 25127 240602 42849
rect 240302 25009 240393 25127
rect 240511 25009 240602 25127
rect 240302 24967 240602 25009
rect 240302 24849 240393 24967
rect 240511 24849 240602 24967
rect 240302 7127 240602 24849
rect 240302 7009 240393 7127
rect 240511 7009 240602 7127
rect 240302 6967 240602 7009
rect 240302 6849 240393 6967
rect 240511 6849 240602 6967
rect 231302 -3581 231393 -3463
rect 231511 -3581 231602 -3463
rect 231302 -3623 231602 -3581
rect 231302 -3741 231393 -3623
rect 231511 -3741 231602 -3623
rect 231302 -3752 231602 -3741
rect 240302 -2993 240602 6849
rect 243902 352889 244202 352900
rect 243902 352771 243993 352889
rect 244111 352771 244202 352889
rect 243902 352729 244202 352771
rect 243902 352611 243993 352729
rect 244111 352611 244202 352729
rect 243902 334727 244202 352611
rect 243902 334609 243993 334727
rect 244111 334609 244202 334727
rect 243902 334567 244202 334609
rect 243902 334449 243993 334567
rect 244111 334449 244202 334567
rect 243902 316727 244202 334449
rect 243902 316609 243993 316727
rect 244111 316609 244202 316727
rect 243902 316567 244202 316609
rect 243902 316449 243993 316567
rect 244111 316449 244202 316567
rect 243902 298727 244202 316449
rect 243902 298609 243993 298727
rect 244111 298609 244202 298727
rect 243902 298567 244202 298609
rect 243902 298449 243993 298567
rect 244111 298449 244202 298567
rect 243902 280727 244202 298449
rect 243902 280609 243993 280727
rect 244111 280609 244202 280727
rect 243902 280567 244202 280609
rect 243902 280449 243993 280567
rect 244111 280449 244202 280567
rect 243902 262727 244202 280449
rect 243902 262609 243993 262727
rect 244111 262609 244202 262727
rect 243902 262567 244202 262609
rect 243902 262449 243993 262567
rect 244111 262449 244202 262567
rect 243902 244727 244202 262449
rect 243902 244609 243993 244727
rect 244111 244609 244202 244727
rect 243902 244567 244202 244609
rect 243902 244449 243993 244567
rect 244111 244449 244202 244567
rect 243902 226727 244202 244449
rect 243902 226609 243993 226727
rect 244111 226609 244202 226727
rect 243902 226567 244202 226609
rect 243902 226449 243993 226567
rect 244111 226449 244202 226567
rect 243902 208727 244202 226449
rect 243902 208609 243993 208727
rect 244111 208609 244202 208727
rect 243902 208567 244202 208609
rect 243902 208449 243993 208567
rect 244111 208449 244202 208567
rect 243902 190727 244202 208449
rect 243902 190609 243993 190727
rect 244111 190609 244202 190727
rect 243902 190567 244202 190609
rect 243902 190449 243993 190567
rect 244111 190449 244202 190567
rect 243902 172727 244202 190449
rect 243902 172609 243993 172727
rect 244111 172609 244202 172727
rect 243902 172567 244202 172609
rect 243902 172449 243993 172567
rect 244111 172449 244202 172567
rect 243902 154727 244202 172449
rect 243902 154609 243993 154727
rect 244111 154609 244202 154727
rect 243902 154567 244202 154609
rect 243902 154449 243993 154567
rect 244111 154449 244202 154567
rect 243902 136727 244202 154449
rect 243902 136609 243993 136727
rect 244111 136609 244202 136727
rect 243902 136567 244202 136609
rect 243902 136449 243993 136567
rect 244111 136449 244202 136567
rect 243902 118727 244202 136449
rect 243902 118609 243993 118727
rect 244111 118609 244202 118727
rect 243902 118567 244202 118609
rect 243902 118449 243993 118567
rect 244111 118449 244202 118567
rect 243902 100727 244202 118449
rect 243902 100609 243993 100727
rect 244111 100609 244202 100727
rect 243902 100567 244202 100609
rect 243902 100449 243993 100567
rect 244111 100449 244202 100567
rect 243902 82727 244202 100449
rect 243902 82609 243993 82727
rect 244111 82609 244202 82727
rect 243902 82567 244202 82609
rect 243902 82449 243993 82567
rect 244111 82449 244202 82567
rect 243902 64727 244202 82449
rect 243902 64609 243993 64727
rect 244111 64609 244202 64727
rect 243902 64567 244202 64609
rect 243902 64449 243993 64567
rect 244111 64449 244202 64567
rect 243902 46727 244202 64449
rect 243902 46609 243993 46727
rect 244111 46609 244202 46727
rect 243902 46567 244202 46609
rect 243902 46449 243993 46567
rect 244111 46449 244202 46567
rect 243902 28727 244202 46449
rect 243902 28609 243993 28727
rect 244111 28609 244202 28727
rect 243902 28567 244202 28609
rect 243902 28449 243993 28567
rect 244111 28449 244202 28567
rect 243902 10727 244202 28449
rect 243902 10609 243993 10727
rect 244111 10609 244202 10727
rect 243902 10567 244202 10609
rect 243902 10449 243993 10567
rect 244111 10449 244202 10567
rect 243902 -643 244202 10449
rect 243902 -761 243993 -643
rect 244111 -761 244202 -643
rect 243902 -803 244202 -761
rect 243902 -921 243993 -803
rect 244111 -921 244202 -803
rect 243902 -932 244202 -921
rect 245702 336527 246002 353551
rect 245702 336409 245793 336527
rect 245911 336409 246002 336527
rect 245702 336367 246002 336409
rect 245702 336249 245793 336367
rect 245911 336249 246002 336367
rect 245702 318527 246002 336249
rect 245702 318409 245793 318527
rect 245911 318409 246002 318527
rect 245702 318367 246002 318409
rect 245702 318249 245793 318367
rect 245911 318249 246002 318367
rect 245702 300527 246002 318249
rect 245702 300409 245793 300527
rect 245911 300409 246002 300527
rect 245702 300367 246002 300409
rect 245702 300249 245793 300367
rect 245911 300249 246002 300367
rect 245702 282527 246002 300249
rect 245702 282409 245793 282527
rect 245911 282409 246002 282527
rect 245702 282367 246002 282409
rect 245702 282249 245793 282367
rect 245911 282249 246002 282367
rect 245702 264527 246002 282249
rect 245702 264409 245793 264527
rect 245911 264409 246002 264527
rect 245702 264367 246002 264409
rect 245702 264249 245793 264367
rect 245911 264249 246002 264367
rect 245702 246527 246002 264249
rect 245702 246409 245793 246527
rect 245911 246409 246002 246527
rect 245702 246367 246002 246409
rect 245702 246249 245793 246367
rect 245911 246249 246002 246367
rect 245702 228527 246002 246249
rect 245702 228409 245793 228527
rect 245911 228409 246002 228527
rect 245702 228367 246002 228409
rect 245702 228249 245793 228367
rect 245911 228249 246002 228367
rect 245702 210527 246002 228249
rect 245702 210409 245793 210527
rect 245911 210409 246002 210527
rect 245702 210367 246002 210409
rect 245702 210249 245793 210367
rect 245911 210249 246002 210367
rect 245702 192527 246002 210249
rect 245702 192409 245793 192527
rect 245911 192409 246002 192527
rect 245702 192367 246002 192409
rect 245702 192249 245793 192367
rect 245911 192249 246002 192367
rect 245702 174527 246002 192249
rect 245702 174409 245793 174527
rect 245911 174409 246002 174527
rect 245702 174367 246002 174409
rect 245702 174249 245793 174367
rect 245911 174249 246002 174367
rect 245702 156527 246002 174249
rect 245702 156409 245793 156527
rect 245911 156409 246002 156527
rect 245702 156367 246002 156409
rect 245702 156249 245793 156367
rect 245911 156249 246002 156367
rect 245702 138527 246002 156249
rect 245702 138409 245793 138527
rect 245911 138409 246002 138527
rect 245702 138367 246002 138409
rect 245702 138249 245793 138367
rect 245911 138249 246002 138367
rect 245702 120527 246002 138249
rect 245702 120409 245793 120527
rect 245911 120409 246002 120527
rect 245702 120367 246002 120409
rect 245702 120249 245793 120367
rect 245911 120249 246002 120367
rect 245702 102527 246002 120249
rect 245702 102409 245793 102527
rect 245911 102409 246002 102527
rect 245702 102367 246002 102409
rect 245702 102249 245793 102367
rect 245911 102249 246002 102367
rect 245702 84527 246002 102249
rect 245702 84409 245793 84527
rect 245911 84409 246002 84527
rect 245702 84367 246002 84409
rect 245702 84249 245793 84367
rect 245911 84249 246002 84367
rect 245702 66527 246002 84249
rect 245702 66409 245793 66527
rect 245911 66409 246002 66527
rect 245702 66367 246002 66409
rect 245702 66249 245793 66367
rect 245911 66249 246002 66367
rect 245702 48527 246002 66249
rect 245702 48409 245793 48527
rect 245911 48409 246002 48527
rect 245702 48367 246002 48409
rect 245702 48249 245793 48367
rect 245911 48249 246002 48367
rect 245702 30527 246002 48249
rect 245702 30409 245793 30527
rect 245911 30409 246002 30527
rect 245702 30367 246002 30409
rect 245702 30249 245793 30367
rect 245911 30249 246002 30367
rect 245702 12527 246002 30249
rect 245702 12409 245793 12527
rect 245911 12409 246002 12527
rect 245702 12367 246002 12409
rect 245702 12249 245793 12367
rect 245911 12249 246002 12367
rect 245702 -1583 246002 12249
rect 245702 -1701 245793 -1583
rect 245911 -1701 246002 -1583
rect 245702 -1743 246002 -1701
rect 245702 -1861 245793 -1743
rect 245911 -1861 246002 -1743
rect 245702 -1872 246002 -1861
rect 247502 338327 247802 354491
rect 247502 338209 247593 338327
rect 247711 338209 247802 338327
rect 247502 338167 247802 338209
rect 247502 338049 247593 338167
rect 247711 338049 247802 338167
rect 247502 320327 247802 338049
rect 247502 320209 247593 320327
rect 247711 320209 247802 320327
rect 247502 320167 247802 320209
rect 247502 320049 247593 320167
rect 247711 320049 247802 320167
rect 247502 302327 247802 320049
rect 247502 302209 247593 302327
rect 247711 302209 247802 302327
rect 247502 302167 247802 302209
rect 247502 302049 247593 302167
rect 247711 302049 247802 302167
rect 247502 284327 247802 302049
rect 247502 284209 247593 284327
rect 247711 284209 247802 284327
rect 247502 284167 247802 284209
rect 247502 284049 247593 284167
rect 247711 284049 247802 284167
rect 247502 266327 247802 284049
rect 247502 266209 247593 266327
rect 247711 266209 247802 266327
rect 247502 266167 247802 266209
rect 247502 266049 247593 266167
rect 247711 266049 247802 266167
rect 247502 248327 247802 266049
rect 247502 248209 247593 248327
rect 247711 248209 247802 248327
rect 247502 248167 247802 248209
rect 247502 248049 247593 248167
rect 247711 248049 247802 248167
rect 247502 230327 247802 248049
rect 247502 230209 247593 230327
rect 247711 230209 247802 230327
rect 247502 230167 247802 230209
rect 247502 230049 247593 230167
rect 247711 230049 247802 230167
rect 247502 212327 247802 230049
rect 247502 212209 247593 212327
rect 247711 212209 247802 212327
rect 247502 212167 247802 212209
rect 247502 212049 247593 212167
rect 247711 212049 247802 212167
rect 247502 194327 247802 212049
rect 247502 194209 247593 194327
rect 247711 194209 247802 194327
rect 247502 194167 247802 194209
rect 247502 194049 247593 194167
rect 247711 194049 247802 194167
rect 247502 176327 247802 194049
rect 247502 176209 247593 176327
rect 247711 176209 247802 176327
rect 247502 176167 247802 176209
rect 247502 176049 247593 176167
rect 247711 176049 247802 176167
rect 247502 158327 247802 176049
rect 247502 158209 247593 158327
rect 247711 158209 247802 158327
rect 247502 158167 247802 158209
rect 247502 158049 247593 158167
rect 247711 158049 247802 158167
rect 247502 140327 247802 158049
rect 247502 140209 247593 140327
rect 247711 140209 247802 140327
rect 247502 140167 247802 140209
rect 247502 140049 247593 140167
rect 247711 140049 247802 140167
rect 247502 122327 247802 140049
rect 247502 122209 247593 122327
rect 247711 122209 247802 122327
rect 247502 122167 247802 122209
rect 247502 122049 247593 122167
rect 247711 122049 247802 122167
rect 247502 104327 247802 122049
rect 247502 104209 247593 104327
rect 247711 104209 247802 104327
rect 247502 104167 247802 104209
rect 247502 104049 247593 104167
rect 247711 104049 247802 104167
rect 247502 86327 247802 104049
rect 247502 86209 247593 86327
rect 247711 86209 247802 86327
rect 247502 86167 247802 86209
rect 247502 86049 247593 86167
rect 247711 86049 247802 86167
rect 247502 68327 247802 86049
rect 247502 68209 247593 68327
rect 247711 68209 247802 68327
rect 247502 68167 247802 68209
rect 247502 68049 247593 68167
rect 247711 68049 247802 68167
rect 247502 50327 247802 68049
rect 247502 50209 247593 50327
rect 247711 50209 247802 50327
rect 247502 50167 247802 50209
rect 247502 50049 247593 50167
rect 247711 50049 247802 50167
rect 247502 32327 247802 50049
rect 247502 32209 247593 32327
rect 247711 32209 247802 32327
rect 247502 32167 247802 32209
rect 247502 32049 247593 32167
rect 247711 32049 247802 32167
rect 247502 14327 247802 32049
rect 247502 14209 247593 14327
rect 247711 14209 247802 14327
rect 247502 14167 247802 14209
rect 247502 14049 247593 14167
rect 247711 14049 247802 14167
rect 247502 -2523 247802 14049
rect 247502 -2641 247593 -2523
rect 247711 -2641 247802 -2523
rect 247502 -2683 247802 -2641
rect 247502 -2801 247593 -2683
rect 247711 -2801 247802 -2683
rect 247502 -2812 247802 -2801
rect 249302 340127 249602 355431
rect 258302 355239 258602 355720
rect 258302 355121 258393 355239
rect 258511 355121 258602 355239
rect 258302 355079 258602 355121
rect 258302 354961 258393 355079
rect 258511 354961 258602 355079
rect 256502 354299 256802 354780
rect 256502 354181 256593 354299
rect 256711 354181 256802 354299
rect 256502 354139 256802 354181
rect 256502 354021 256593 354139
rect 256711 354021 256802 354139
rect 254702 353359 255002 353840
rect 254702 353241 254793 353359
rect 254911 353241 255002 353359
rect 254702 353199 255002 353241
rect 254702 353081 254793 353199
rect 254911 353081 255002 353199
rect 249302 340009 249393 340127
rect 249511 340009 249602 340127
rect 249302 339967 249602 340009
rect 249302 339849 249393 339967
rect 249511 339849 249602 339967
rect 249302 322127 249602 339849
rect 249302 322009 249393 322127
rect 249511 322009 249602 322127
rect 249302 321967 249602 322009
rect 249302 321849 249393 321967
rect 249511 321849 249602 321967
rect 249302 304127 249602 321849
rect 249302 304009 249393 304127
rect 249511 304009 249602 304127
rect 249302 303967 249602 304009
rect 249302 303849 249393 303967
rect 249511 303849 249602 303967
rect 249302 286127 249602 303849
rect 249302 286009 249393 286127
rect 249511 286009 249602 286127
rect 249302 285967 249602 286009
rect 249302 285849 249393 285967
rect 249511 285849 249602 285967
rect 249302 268127 249602 285849
rect 249302 268009 249393 268127
rect 249511 268009 249602 268127
rect 249302 267967 249602 268009
rect 249302 267849 249393 267967
rect 249511 267849 249602 267967
rect 249302 250127 249602 267849
rect 249302 250009 249393 250127
rect 249511 250009 249602 250127
rect 249302 249967 249602 250009
rect 249302 249849 249393 249967
rect 249511 249849 249602 249967
rect 249302 232127 249602 249849
rect 249302 232009 249393 232127
rect 249511 232009 249602 232127
rect 249302 231967 249602 232009
rect 249302 231849 249393 231967
rect 249511 231849 249602 231967
rect 249302 214127 249602 231849
rect 249302 214009 249393 214127
rect 249511 214009 249602 214127
rect 249302 213967 249602 214009
rect 249302 213849 249393 213967
rect 249511 213849 249602 213967
rect 249302 196127 249602 213849
rect 249302 196009 249393 196127
rect 249511 196009 249602 196127
rect 249302 195967 249602 196009
rect 249302 195849 249393 195967
rect 249511 195849 249602 195967
rect 249302 178127 249602 195849
rect 249302 178009 249393 178127
rect 249511 178009 249602 178127
rect 249302 177967 249602 178009
rect 249302 177849 249393 177967
rect 249511 177849 249602 177967
rect 249302 160127 249602 177849
rect 249302 160009 249393 160127
rect 249511 160009 249602 160127
rect 249302 159967 249602 160009
rect 249302 159849 249393 159967
rect 249511 159849 249602 159967
rect 249302 142127 249602 159849
rect 249302 142009 249393 142127
rect 249511 142009 249602 142127
rect 249302 141967 249602 142009
rect 249302 141849 249393 141967
rect 249511 141849 249602 141967
rect 249302 124127 249602 141849
rect 249302 124009 249393 124127
rect 249511 124009 249602 124127
rect 249302 123967 249602 124009
rect 249302 123849 249393 123967
rect 249511 123849 249602 123967
rect 249302 106127 249602 123849
rect 249302 106009 249393 106127
rect 249511 106009 249602 106127
rect 249302 105967 249602 106009
rect 249302 105849 249393 105967
rect 249511 105849 249602 105967
rect 249302 88127 249602 105849
rect 249302 88009 249393 88127
rect 249511 88009 249602 88127
rect 249302 87967 249602 88009
rect 249302 87849 249393 87967
rect 249511 87849 249602 87967
rect 249302 70127 249602 87849
rect 249302 70009 249393 70127
rect 249511 70009 249602 70127
rect 249302 69967 249602 70009
rect 249302 69849 249393 69967
rect 249511 69849 249602 69967
rect 249302 52127 249602 69849
rect 249302 52009 249393 52127
rect 249511 52009 249602 52127
rect 249302 51967 249602 52009
rect 249302 51849 249393 51967
rect 249511 51849 249602 51967
rect 249302 34127 249602 51849
rect 249302 34009 249393 34127
rect 249511 34009 249602 34127
rect 249302 33967 249602 34009
rect 249302 33849 249393 33967
rect 249511 33849 249602 33967
rect 249302 16127 249602 33849
rect 249302 16009 249393 16127
rect 249511 16009 249602 16127
rect 249302 15967 249602 16009
rect 249302 15849 249393 15967
rect 249511 15849 249602 15967
rect 240302 -3111 240393 -2993
rect 240511 -3111 240602 -2993
rect 240302 -3153 240602 -3111
rect 240302 -3271 240393 -3153
rect 240511 -3271 240602 -3153
rect 240302 -3752 240602 -3271
rect 249302 -3463 249602 15849
rect 252902 352419 253202 352900
rect 252902 352301 252993 352419
rect 253111 352301 253202 352419
rect 252902 352259 253202 352301
rect 252902 352141 252993 352259
rect 253111 352141 253202 352259
rect 252902 343727 253202 352141
rect 252902 343609 252993 343727
rect 253111 343609 253202 343727
rect 252902 343567 253202 343609
rect 252902 343449 252993 343567
rect 253111 343449 253202 343567
rect 252902 325727 253202 343449
rect 252902 325609 252993 325727
rect 253111 325609 253202 325727
rect 252902 325567 253202 325609
rect 252902 325449 252993 325567
rect 253111 325449 253202 325567
rect 252902 307727 253202 325449
rect 252902 307609 252993 307727
rect 253111 307609 253202 307727
rect 252902 307567 253202 307609
rect 252902 307449 252993 307567
rect 253111 307449 253202 307567
rect 252902 289727 253202 307449
rect 252902 289609 252993 289727
rect 253111 289609 253202 289727
rect 252902 289567 253202 289609
rect 252902 289449 252993 289567
rect 253111 289449 253202 289567
rect 252902 271727 253202 289449
rect 252902 271609 252993 271727
rect 253111 271609 253202 271727
rect 252902 271567 253202 271609
rect 252902 271449 252993 271567
rect 253111 271449 253202 271567
rect 252902 253727 253202 271449
rect 252902 253609 252993 253727
rect 253111 253609 253202 253727
rect 252902 253567 253202 253609
rect 252902 253449 252993 253567
rect 253111 253449 253202 253567
rect 252902 235727 253202 253449
rect 252902 235609 252993 235727
rect 253111 235609 253202 235727
rect 252902 235567 253202 235609
rect 252902 235449 252993 235567
rect 253111 235449 253202 235567
rect 252902 217727 253202 235449
rect 252902 217609 252993 217727
rect 253111 217609 253202 217727
rect 252902 217567 253202 217609
rect 252902 217449 252993 217567
rect 253111 217449 253202 217567
rect 252902 199727 253202 217449
rect 252902 199609 252993 199727
rect 253111 199609 253202 199727
rect 252902 199567 253202 199609
rect 252902 199449 252993 199567
rect 253111 199449 253202 199567
rect 252902 181727 253202 199449
rect 252902 181609 252993 181727
rect 253111 181609 253202 181727
rect 252902 181567 253202 181609
rect 252902 181449 252993 181567
rect 253111 181449 253202 181567
rect 252902 163727 253202 181449
rect 252902 163609 252993 163727
rect 253111 163609 253202 163727
rect 252902 163567 253202 163609
rect 252902 163449 252993 163567
rect 253111 163449 253202 163567
rect 252902 145727 253202 163449
rect 252902 145609 252993 145727
rect 253111 145609 253202 145727
rect 252902 145567 253202 145609
rect 252902 145449 252993 145567
rect 253111 145449 253202 145567
rect 252902 127727 253202 145449
rect 252902 127609 252993 127727
rect 253111 127609 253202 127727
rect 252902 127567 253202 127609
rect 252902 127449 252993 127567
rect 253111 127449 253202 127567
rect 252902 109727 253202 127449
rect 252902 109609 252993 109727
rect 253111 109609 253202 109727
rect 252902 109567 253202 109609
rect 252902 109449 252993 109567
rect 253111 109449 253202 109567
rect 252902 91727 253202 109449
rect 252902 91609 252993 91727
rect 253111 91609 253202 91727
rect 252902 91567 253202 91609
rect 252902 91449 252993 91567
rect 253111 91449 253202 91567
rect 252902 73727 253202 91449
rect 252902 73609 252993 73727
rect 253111 73609 253202 73727
rect 252902 73567 253202 73609
rect 252902 73449 252993 73567
rect 253111 73449 253202 73567
rect 252902 55727 253202 73449
rect 252902 55609 252993 55727
rect 253111 55609 253202 55727
rect 252902 55567 253202 55609
rect 252902 55449 252993 55567
rect 253111 55449 253202 55567
rect 252902 37727 253202 55449
rect 252902 37609 252993 37727
rect 253111 37609 253202 37727
rect 252902 37567 253202 37609
rect 252902 37449 252993 37567
rect 253111 37449 253202 37567
rect 252902 19727 253202 37449
rect 252902 19609 252993 19727
rect 253111 19609 253202 19727
rect 252902 19567 253202 19609
rect 252902 19449 252993 19567
rect 253111 19449 253202 19567
rect 252902 1727 253202 19449
rect 252902 1609 252993 1727
rect 253111 1609 253202 1727
rect 252902 1567 253202 1609
rect 252902 1449 252993 1567
rect 253111 1449 253202 1567
rect 252902 -173 253202 1449
rect 252902 -291 252993 -173
rect 253111 -291 253202 -173
rect 252902 -333 253202 -291
rect 252902 -451 252993 -333
rect 253111 -451 253202 -333
rect 252902 -932 253202 -451
rect 254702 345527 255002 353081
rect 254702 345409 254793 345527
rect 254911 345409 255002 345527
rect 254702 345367 255002 345409
rect 254702 345249 254793 345367
rect 254911 345249 255002 345367
rect 254702 327527 255002 345249
rect 254702 327409 254793 327527
rect 254911 327409 255002 327527
rect 254702 327367 255002 327409
rect 254702 327249 254793 327367
rect 254911 327249 255002 327367
rect 254702 309527 255002 327249
rect 254702 309409 254793 309527
rect 254911 309409 255002 309527
rect 254702 309367 255002 309409
rect 254702 309249 254793 309367
rect 254911 309249 255002 309367
rect 254702 291527 255002 309249
rect 254702 291409 254793 291527
rect 254911 291409 255002 291527
rect 254702 291367 255002 291409
rect 254702 291249 254793 291367
rect 254911 291249 255002 291367
rect 254702 273527 255002 291249
rect 254702 273409 254793 273527
rect 254911 273409 255002 273527
rect 254702 273367 255002 273409
rect 254702 273249 254793 273367
rect 254911 273249 255002 273367
rect 254702 255527 255002 273249
rect 254702 255409 254793 255527
rect 254911 255409 255002 255527
rect 254702 255367 255002 255409
rect 254702 255249 254793 255367
rect 254911 255249 255002 255367
rect 254702 237527 255002 255249
rect 254702 237409 254793 237527
rect 254911 237409 255002 237527
rect 254702 237367 255002 237409
rect 254702 237249 254793 237367
rect 254911 237249 255002 237367
rect 254702 219527 255002 237249
rect 254702 219409 254793 219527
rect 254911 219409 255002 219527
rect 254702 219367 255002 219409
rect 254702 219249 254793 219367
rect 254911 219249 255002 219367
rect 254702 201527 255002 219249
rect 254702 201409 254793 201527
rect 254911 201409 255002 201527
rect 254702 201367 255002 201409
rect 254702 201249 254793 201367
rect 254911 201249 255002 201367
rect 254702 183527 255002 201249
rect 254702 183409 254793 183527
rect 254911 183409 255002 183527
rect 254702 183367 255002 183409
rect 254702 183249 254793 183367
rect 254911 183249 255002 183367
rect 254702 165527 255002 183249
rect 254702 165409 254793 165527
rect 254911 165409 255002 165527
rect 254702 165367 255002 165409
rect 254702 165249 254793 165367
rect 254911 165249 255002 165367
rect 254702 147527 255002 165249
rect 254702 147409 254793 147527
rect 254911 147409 255002 147527
rect 254702 147367 255002 147409
rect 254702 147249 254793 147367
rect 254911 147249 255002 147367
rect 254702 129527 255002 147249
rect 254702 129409 254793 129527
rect 254911 129409 255002 129527
rect 254702 129367 255002 129409
rect 254702 129249 254793 129367
rect 254911 129249 255002 129367
rect 254702 111527 255002 129249
rect 254702 111409 254793 111527
rect 254911 111409 255002 111527
rect 254702 111367 255002 111409
rect 254702 111249 254793 111367
rect 254911 111249 255002 111367
rect 254702 93527 255002 111249
rect 254702 93409 254793 93527
rect 254911 93409 255002 93527
rect 254702 93367 255002 93409
rect 254702 93249 254793 93367
rect 254911 93249 255002 93367
rect 254702 75527 255002 93249
rect 254702 75409 254793 75527
rect 254911 75409 255002 75527
rect 254702 75367 255002 75409
rect 254702 75249 254793 75367
rect 254911 75249 255002 75367
rect 254702 57527 255002 75249
rect 254702 57409 254793 57527
rect 254911 57409 255002 57527
rect 254702 57367 255002 57409
rect 254702 57249 254793 57367
rect 254911 57249 255002 57367
rect 254702 39527 255002 57249
rect 254702 39409 254793 39527
rect 254911 39409 255002 39527
rect 254702 39367 255002 39409
rect 254702 39249 254793 39367
rect 254911 39249 255002 39367
rect 254702 21527 255002 39249
rect 254702 21409 254793 21527
rect 254911 21409 255002 21527
rect 254702 21367 255002 21409
rect 254702 21249 254793 21367
rect 254911 21249 255002 21367
rect 254702 3527 255002 21249
rect 254702 3409 254793 3527
rect 254911 3409 255002 3527
rect 254702 3367 255002 3409
rect 254702 3249 254793 3367
rect 254911 3249 255002 3367
rect 254702 -1113 255002 3249
rect 254702 -1231 254793 -1113
rect 254911 -1231 255002 -1113
rect 254702 -1273 255002 -1231
rect 254702 -1391 254793 -1273
rect 254911 -1391 255002 -1273
rect 254702 -1872 255002 -1391
rect 256502 347327 256802 354021
rect 256502 347209 256593 347327
rect 256711 347209 256802 347327
rect 256502 347167 256802 347209
rect 256502 347049 256593 347167
rect 256711 347049 256802 347167
rect 256502 329327 256802 347049
rect 256502 329209 256593 329327
rect 256711 329209 256802 329327
rect 256502 329167 256802 329209
rect 256502 329049 256593 329167
rect 256711 329049 256802 329167
rect 256502 311327 256802 329049
rect 256502 311209 256593 311327
rect 256711 311209 256802 311327
rect 256502 311167 256802 311209
rect 256502 311049 256593 311167
rect 256711 311049 256802 311167
rect 256502 293327 256802 311049
rect 256502 293209 256593 293327
rect 256711 293209 256802 293327
rect 256502 293167 256802 293209
rect 256502 293049 256593 293167
rect 256711 293049 256802 293167
rect 256502 275327 256802 293049
rect 256502 275209 256593 275327
rect 256711 275209 256802 275327
rect 256502 275167 256802 275209
rect 256502 275049 256593 275167
rect 256711 275049 256802 275167
rect 256502 257327 256802 275049
rect 256502 257209 256593 257327
rect 256711 257209 256802 257327
rect 256502 257167 256802 257209
rect 256502 257049 256593 257167
rect 256711 257049 256802 257167
rect 256502 239327 256802 257049
rect 256502 239209 256593 239327
rect 256711 239209 256802 239327
rect 256502 239167 256802 239209
rect 256502 239049 256593 239167
rect 256711 239049 256802 239167
rect 256502 221327 256802 239049
rect 256502 221209 256593 221327
rect 256711 221209 256802 221327
rect 256502 221167 256802 221209
rect 256502 221049 256593 221167
rect 256711 221049 256802 221167
rect 256502 203327 256802 221049
rect 256502 203209 256593 203327
rect 256711 203209 256802 203327
rect 256502 203167 256802 203209
rect 256502 203049 256593 203167
rect 256711 203049 256802 203167
rect 256502 185327 256802 203049
rect 256502 185209 256593 185327
rect 256711 185209 256802 185327
rect 256502 185167 256802 185209
rect 256502 185049 256593 185167
rect 256711 185049 256802 185167
rect 256502 167327 256802 185049
rect 256502 167209 256593 167327
rect 256711 167209 256802 167327
rect 256502 167167 256802 167209
rect 256502 167049 256593 167167
rect 256711 167049 256802 167167
rect 256502 149327 256802 167049
rect 256502 149209 256593 149327
rect 256711 149209 256802 149327
rect 256502 149167 256802 149209
rect 256502 149049 256593 149167
rect 256711 149049 256802 149167
rect 256502 131327 256802 149049
rect 256502 131209 256593 131327
rect 256711 131209 256802 131327
rect 256502 131167 256802 131209
rect 256502 131049 256593 131167
rect 256711 131049 256802 131167
rect 256502 113327 256802 131049
rect 256502 113209 256593 113327
rect 256711 113209 256802 113327
rect 256502 113167 256802 113209
rect 256502 113049 256593 113167
rect 256711 113049 256802 113167
rect 256502 95327 256802 113049
rect 256502 95209 256593 95327
rect 256711 95209 256802 95327
rect 256502 95167 256802 95209
rect 256502 95049 256593 95167
rect 256711 95049 256802 95167
rect 256502 77327 256802 95049
rect 256502 77209 256593 77327
rect 256711 77209 256802 77327
rect 256502 77167 256802 77209
rect 256502 77049 256593 77167
rect 256711 77049 256802 77167
rect 256502 59327 256802 77049
rect 256502 59209 256593 59327
rect 256711 59209 256802 59327
rect 256502 59167 256802 59209
rect 256502 59049 256593 59167
rect 256711 59049 256802 59167
rect 256502 41327 256802 59049
rect 256502 41209 256593 41327
rect 256711 41209 256802 41327
rect 256502 41167 256802 41209
rect 256502 41049 256593 41167
rect 256711 41049 256802 41167
rect 256502 23327 256802 41049
rect 256502 23209 256593 23327
rect 256711 23209 256802 23327
rect 256502 23167 256802 23209
rect 256502 23049 256593 23167
rect 256711 23049 256802 23167
rect 256502 5327 256802 23049
rect 256502 5209 256593 5327
rect 256711 5209 256802 5327
rect 256502 5167 256802 5209
rect 256502 5049 256593 5167
rect 256711 5049 256802 5167
rect 256502 -2053 256802 5049
rect 256502 -2171 256593 -2053
rect 256711 -2171 256802 -2053
rect 256502 -2213 256802 -2171
rect 256502 -2331 256593 -2213
rect 256711 -2331 256802 -2213
rect 256502 -2812 256802 -2331
rect 258302 349127 258602 354961
rect 267302 355709 267602 355720
rect 267302 355591 267393 355709
rect 267511 355591 267602 355709
rect 267302 355549 267602 355591
rect 267302 355431 267393 355549
rect 267511 355431 267602 355549
rect 265502 354769 265802 354780
rect 265502 354651 265593 354769
rect 265711 354651 265802 354769
rect 265502 354609 265802 354651
rect 265502 354491 265593 354609
rect 265711 354491 265802 354609
rect 263702 353829 264002 353840
rect 263702 353711 263793 353829
rect 263911 353711 264002 353829
rect 263702 353669 264002 353711
rect 263702 353551 263793 353669
rect 263911 353551 264002 353669
rect 258302 349009 258393 349127
rect 258511 349009 258602 349127
rect 258302 348967 258602 349009
rect 258302 348849 258393 348967
rect 258511 348849 258602 348967
rect 258302 331127 258602 348849
rect 258302 331009 258393 331127
rect 258511 331009 258602 331127
rect 258302 330967 258602 331009
rect 258302 330849 258393 330967
rect 258511 330849 258602 330967
rect 258302 313127 258602 330849
rect 258302 313009 258393 313127
rect 258511 313009 258602 313127
rect 258302 312967 258602 313009
rect 258302 312849 258393 312967
rect 258511 312849 258602 312967
rect 258302 295127 258602 312849
rect 258302 295009 258393 295127
rect 258511 295009 258602 295127
rect 258302 294967 258602 295009
rect 258302 294849 258393 294967
rect 258511 294849 258602 294967
rect 258302 277127 258602 294849
rect 258302 277009 258393 277127
rect 258511 277009 258602 277127
rect 258302 276967 258602 277009
rect 258302 276849 258393 276967
rect 258511 276849 258602 276967
rect 258302 259127 258602 276849
rect 258302 259009 258393 259127
rect 258511 259009 258602 259127
rect 258302 258967 258602 259009
rect 258302 258849 258393 258967
rect 258511 258849 258602 258967
rect 258302 241127 258602 258849
rect 258302 241009 258393 241127
rect 258511 241009 258602 241127
rect 258302 240967 258602 241009
rect 258302 240849 258393 240967
rect 258511 240849 258602 240967
rect 258302 223127 258602 240849
rect 258302 223009 258393 223127
rect 258511 223009 258602 223127
rect 258302 222967 258602 223009
rect 258302 222849 258393 222967
rect 258511 222849 258602 222967
rect 258302 205127 258602 222849
rect 258302 205009 258393 205127
rect 258511 205009 258602 205127
rect 258302 204967 258602 205009
rect 258302 204849 258393 204967
rect 258511 204849 258602 204967
rect 258302 187127 258602 204849
rect 258302 187009 258393 187127
rect 258511 187009 258602 187127
rect 258302 186967 258602 187009
rect 258302 186849 258393 186967
rect 258511 186849 258602 186967
rect 258302 169127 258602 186849
rect 258302 169009 258393 169127
rect 258511 169009 258602 169127
rect 258302 168967 258602 169009
rect 258302 168849 258393 168967
rect 258511 168849 258602 168967
rect 258302 151127 258602 168849
rect 258302 151009 258393 151127
rect 258511 151009 258602 151127
rect 258302 150967 258602 151009
rect 258302 150849 258393 150967
rect 258511 150849 258602 150967
rect 258302 133127 258602 150849
rect 258302 133009 258393 133127
rect 258511 133009 258602 133127
rect 258302 132967 258602 133009
rect 258302 132849 258393 132967
rect 258511 132849 258602 132967
rect 258302 115127 258602 132849
rect 258302 115009 258393 115127
rect 258511 115009 258602 115127
rect 258302 114967 258602 115009
rect 258302 114849 258393 114967
rect 258511 114849 258602 114967
rect 258302 97127 258602 114849
rect 258302 97009 258393 97127
rect 258511 97009 258602 97127
rect 258302 96967 258602 97009
rect 258302 96849 258393 96967
rect 258511 96849 258602 96967
rect 258302 79127 258602 96849
rect 258302 79009 258393 79127
rect 258511 79009 258602 79127
rect 258302 78967 258602 79009
rect 258302 78849 258393 78967
rect 258511 78849 258602 78967
rect 258302 61127 258602 78849
rect 258302 61009 258393 61127
rect 258511 61009 258602 61127
rect 258302 60967 258602 61009
rect 258302 60849 258393 60967
rect 258511 60849 258602 60967
rect 258302 43127 258602 60849
rect 258302 43009 258393 43127
rect 258511 43009 258602 43127
rect 258302 42967 258602 43009
rect 258302 42849 258393 42967
rect 258511 42849 258602 42967
rect 258302 25127 258602 42849
rect 258302 25009 258393 25127
rect 258511 25009 258602 25127
rect 258302 24967 258602 25009
rect 258302 24849 258393 24967
rect 258511 24849 258602 24967
rect 258302 7127 258602 24849
rect 258302 7009 258393 7127
rect 258511 7009 258602 7127
rect 258302 6967 258602 7009
rect 258302 6849 258393 6967
rect 258511 6849 258602 6967
rect 249302 -3581 249393 -3463
rect 249511 -3581 249602 -3463
rect 249302 -3623 249602 -3581
rect 249302 -3741 249393 -3623
rect 249511 -3741 249602 -3623
rect 249302 -3752 249602 -3741
rect 258302 -2993 258602 6849
rect 261902 352889 262202 352900
rect 261902 352771 261993 352889
rect 262111 352771 262202 352889
rect 261902 352729 262202 352771
rect 261902 352611 261993 352729
rect 262111 352611 262202 352729
rect 261902 334727 262202 352611
rect 261902 334609 261993 334727
rect 262111 334609 262202 334727
rect 261902 334567 262202 334609
rect 261902 334449 261993 334567
rect 262111 334449 262202 334567
rect 261902 316727 262202 334449
rect 261902 316609 261993 316727
rect 262111 316609 262202 316727
rect 261902 316567 262202 316609
rect 261902 316449 261993 316567
rect 262111 316449 262202 316567
rect 261902 298727 262202 316449
rect 261902 298609 261993 298727
rect 262111 298609 262202 298727
rect 261902 298567 262202 298609
rect 261902 298449 261993 298567
rect 262111 298449 262202 298567
rect 261902 280727 262202 298449
rect 261902 280609 261993 280727
rect 262111 280609 262202 280727
rect 261902 280567 262202 280609
rect 261902 280449 261993 280567
rect 262111 280449 262202 280567
rect 261902 262727 262202 280449
rect 261902 262609 261993 262727
rect 262111 262609 262202 262727
rect 261902 262567 262202 262609
rect 261902 262449 261993 262567
rect 262111 262449 262202 262567
rect 261902 244727 262202 262449
rect 261902 244609 261993 244727
rect 262111 244609 262202 244727
rect 261902 244567 262202 244609
rect 261902 244449 261993 244567
rect 262111 244449 262202 244567
rect 261902 226727 262202 244449
rect 261902 226609 261993 226727
rect 262111 226609 262202 226727
rect 261902 226567 262202 226609
rect 261902 226449 261993 226567
rect 262111 226449 262202 226567
rect 261902 208727 262202 226449
rect 261902 208609 261993 208727
rect 262111 208609 262202 208727
rect 261902 208567 262202 208609
rect 261902 208449 261993 208567
rect 262111 208449 262202 208567
rect 261902 190727 262202 208449
rect 261902 190609 261993 190727
rect 262111 190609 262202 190727
rect 261902 190567 262202 190609
rect 261902 190449 261993 190567
rect 262111 190449 262202 190567
rect 261902 172727 262202 190449
rect 261902 172609 261993 172727
rect 262111 172609 262202 172727
rect 261902 172567 262202 172609
rect 261902 172449 261993 172567
rect 262111 172449 262202 172567
rect 261902 154727 262202 172449
rect 261902 154609 261993 154727
rect 262111 154609 262202 154727
rect 261902 154567 262202 154609
rect 261902 154449 261993 154567
rect 262111 154449 262202 154567
rect 261902 136727 262202 154449
rect 261902 136609 261993 136727
rect 262111 136609 262202 136727
rect 261902 136567 262202 136609
rect 261902 136449 261993 136567
rect 262111 136449 262202 136567
rect 261902 118727 262202 136449
rect 261902 118609 261993 118727
rect 262111 118609 262202 118727
rect 261902 118567 262202 118609
rect 261902 118449 261993 118567
rect 262111 118449 262202 118567
rect 261902 100727 262202 118449
rect 261902 100609 261993 100727
rect 262111 100609 262202 100727
rect 261902 100567 262202 100609
rect 261902 100449 261993 100567
rect 262111 100449 262202 100567
rect 261902 82727 262202 100449
rect 261902 82609 261993 82727
rect 262111 82609 262202 82727
rect 261902 82567 262202 82609
rect 261902 82449 261993 82567
rect 262111 82449 262202 82567
rect 261902 64727 262202 82449
rect 261902 64609 261993 64727
rect 262111 64609 262202 64727
rect 261902 64567 262202 64609
rect 261902 64449 261993 64567
rect 262111 64449 262202 64567
rect 261902 46727 262202 64449
rect 261902 46609 261993 46727
rect 262111 46609 262202 46727
rect 261902 46567 262202 46609
rect 261902 46449 261993 46567
rect 262111 46449 262202 46567
rect 261902 28727 262202 46449
rect 261902 28609 261993 28727
rect 262111 28609 262202 28727
rect 261902 28567 262202 28609
rect 261902 28449 261993 28567
rect 262111 28449 262202 28567
rect 261902 10727 262202 28449
rect 261902 10609 261993 10727
rect 262111 10609 262202 10727
rect 261902 10567 262202 10609
rect 261902 10449 261993 10567
rect 262111 10449 262202 10567
rect 261902 -643 262202 10449
rect 261902 -761 261993 -643
rect 262111 -761 262202 -643
rect 261902 -803 262202 -761
rect 261902 -921 261993 -803
rect 262111 -921 262202 -803
rect 261902 -932 262202 -921
rect 263702 336527 264002 353551
rect 263702 336409 263793 336527
rect 263911 336409 264002 336527
rect 263702 336367 264002 336409
rect 263702 336249 263793 336367
rect 263911 336249 264002 336367
rect 263702 318527 264002 336249
rect 263702 318409 263793 318527
rect 263911 318409 264002 318527
rect 263702 318367 264002 318409
rect 263702 318249 263793 318367
rect 263911 318249 264002 318367
rect 263702 300527 264002 318249
rect 263702 300409 263793 300527
rect 263911 300409 264002 300527
rect 263702 300367 264002 300409
rect 263702 300249 263793 300367
rect 263911 300249 264002 300367
rect 263702 282527 264002 300249
rect 263702 282409 263793 282527
rect 263911 282409 264002 282527
rect 263702 282367 264002 282409
rect 263702 282249 263793 282367
rect 263911 282249 264002 282367
rect 263702 264527 264002 282249
rect 263702 264409 263793 264527
rect 263911 264409 264002 264527
rect 263702 264367 264002 264409
rect 263702 264249 263793 264367
rect 263911 264249 264002 264367
rect 263702 246527 264002 264249
rect 263702 246409 263793 246527
rect 263911 246409 264002 246527
rect 263702 246367 264002 246409
rect 263702 246249 263793 246367
rect 263911 246249 264002 246367
rect 263702 228527 264002 246249
rect 263702 228409 263793 228527
rect 263911 228409 264002 228527
rect 263702 228367 264002 228409
rect 263702 228249 263793 228367
rect 263911 228249 264002 228367
rect 263702 210527 264002 228249
rect 263702 210409 263793 210527
rect 263911 210409 264002 210527
rect 263702 210367 264002 210409
rect 263702 210249 263793 210367
rect 263911 210249 264002 210367
rect 263702 192527 264002 210249
rect 263702 192409 263793 192527
rect 263911 192409 264002 192527
rect 263702 192367 264002 192409
rect 263702 192249 263793 192367
rect 263911 192249 264002 192367
rect 263702 174527 264002 192249
rect 263702 174409 263793 174527
rect 263911 174409 264002 174527
rect 263702 174367 264002 174409
rect 263702 174249 263793 174367
rect 263911 174249 264002 174367
rect 263702 156527 264002 174249
rect 263702 156409 263793 156527
rect 263911 156409 264002 156527
rect 263702 156367 264002 156409
rect 263702 156249 263793 156367
rect 263911 156249 264002 156367
rect 263702 138527 264002 156249
rect 263702 138409 263793 138527
rect 263911 138409 264002 138527
rect 263702 138367 264002 138409
rect 263702 138249 263793 138367
rect 263911 138249 264002 138367
rect 263702 120527 264002 138249
rect 263702 120409 263793 120527
rect 263911 120409 264002 120527
rect 263702 120367 264002 120409
rect 263702 120249 263793 120367
rect 263911 120249 264002 120367
rect 263702 102527 264002 120249
rect 263702 102409 263793 102527
rect 263911 102409 264002 102527
rect 263702 102367 264002 102409
rect 263702 102249 263793 102367
rect 263911 102249 264002 102367
rect 263702 84527 264002 102249
rect 263702 84409 263793 84527
rect 263911 84409 264002 84527
rect 263702 84367 264002 84409
rect 263702 84249 263793 84367
rect 263911 84249 264002 84367
rect 263702 66527 264002 84249
rect 263702 66409 263793 66527
rect 263911 66409 264002 66527
rect 263702 66367 264002 66409
rect 263702 66249 263793 66367
rect 263911 66249 264002 66367
rect 263702 48527 264002 66249
rect 263702 48409 263793 48527
rect 263911 48409 264002 48527
rect 263702 48367 264002 48409
rect 263702 48249 263793 48367
rect 263911 48249 264002 48367
rect 263702 30527 264002 48249
rect 263702 30409 263793 30527
rect 263911 30409 264002 30527
rect 263702 30367 264002 30409
rect 263702 30249 263793 30367
rect 263911 30249 264002 30367
rect 263702 12527 264002 30249
rect 263702 12409 263793 12527
rect 263911 12409 264002 12527
rect 263702 12367 264002 12409
rect 263702 12249 263793 12367
rect 263911 12249 264002 12367
rect 263702 -1583 264002 12249
rect 263702 -1701 263793 -1583
rect 263911 -1701 264002 -1583
rect 263702 -1743 264002 -1701
rect 263702 -1861 263793 -1743
rect 263911 -1861 264002 -1743
rect 263702 -1872 264002 -1861
rect 265502 338327 265802 354491
rect 265502 338209 265593 338327
rect 265711 338209 265802 338327
rect 265502 338167 265802 338209
rect 265502 338049 265593 338167
rect 265711 338049 265802 338167
rect 265502 320327 265802 338049
rect 265502 320209 265593 320327
rect 265711 320209 265802 320327
rect 265502 320167 265802 320209
rect 265502 320049 265593 320167
rect 265711 320049 265802 320167
rect 265502 302327 265802 320049
rect 265502 302209 265593 302327
rect 265711 302209 265802 302327
rect 265502 302167 265802 302209
rect 265502 302049 265593 302167
rect 265711 302049 265802 302167
rect 265502 284327 265802 302049
rect 265502 284209 265593 284327
rect 265711 284209 265802 284327
rect 265502 284167 265802 284209
rect 265502 284049 265593 284167
rect 265711 284049 265802 284167
rect 265502 266327 265802 284049
rect 265502 266209 265593 266327
rect 265711 266209 265802 266327
rect 265502 266167 265802 266209
rect 265502 266049 265593 266167
rect 265711 266049 265802 266167
rect 265502 248327 265802 266049
rect 265502 248209 265593 248327
rect 265711 248209 265802 248327
rect 265502 248167 265802 248209
rect 265502 248049 265593 248167
rect 265711 248049 265802 248167
rect 265502 230327 265802 248049
rect 265502 230209 265593 230327
rect 265711 230209 265802 230327
rect 265502 230167 265802 230209
rect 265502 230049 265593 230167
rect 265711 230049 265802 230167
rect 265502 212327 265802 230049
rect 265502 212209 265593 212327
rect 265711 212209 265802 212327
rect 265502 212167 265802 212209
rect 265502 212049 265593 212167
rect 265711 212049 265802 212167
rect 265502 194327 265802 212049
rect 265502 194209 265593 194327
rect 265711 194209 265802 194327
rect 265502 194167 265802 194209
rect 265502 194049 265593 194167
rect 265711 194049 265802 194167
rect 265502 176327 265802 194049
rect 265502 176209 265593 176327
rect 265711 176209 265802 176327
rect 265502 176167 265802 176209
rect 265502 176049 265593 176167
rect 265711 176049 265802 176167
rect 265502 158327 265802 176049
rect 265502 158209 265593 158327
rect 265711 158209 265802 158327
rect 265502 158167 265802 158209
rect 265502 158049 265593 158167
rect 265711 158049 265802 158167
rect 265502 140327 265802 158049
rect 265502 140209 265593 140327
rect 265711 140209 265802 140327
rect 265502 140167 265802 140209
rect 265502 140049 265593 140167
rect 265711 140049 265802 140167
rect 265502 122327 265802 140049
rect 265502 122209 265593 122327
rect 265711 122209 265802 122327
rect 265502 122167 265802 122209
rect 265502 122049 265593 122167
rect 265711 122049 265802 122167
rect 265502 104327 265802 122049
rect 265502 104209 265593 104327
rect 265711 104209 265802 104327
rect 265502 104167 265802 104209
rect 265502 104049 265593 104167
rect 265711 104049 265802 104167
rect 265502 86327 265802 104049
rect 265502 86209 265593 86327
rect 265711 86209 265802 86327
rect 265502 86167 265802 86209
rect 265502 86049 265593 86167
rect 265711 86049 265802 86167
rect 265502 68327 265802 86049
rect 265502 68209 265593 68327
rect 265711 68209 265802 68327
rect 265502 68167 265802 68209
rect 265502 68049 265593 68167
rect 265711 68049 265802 68167
rect 265502 50327 265802 68049
rect 265502 50209 265593 50327
rect 265711 50209 265802 50327
rect 265502 50167 265802 50209
rect 265502 50049 265593 50167
rect 265711 50049 265802 50167
rect 265502 32327 265802 50049
rect 265502 32209 265593 32327
rect 265711 32209 265802 32327
rect 265502 32167 265802 32209
rect 265502 32049 265593 32167
rect 265711 32049 265802 32167
rect 265502 14327 265802 32049
rect 265502 14209 265593 14327
rect 265711 14209 265802 14327
rect 265502 14167 265802 14209
rect 265502 14049 265593 14167
rect 265711 14049 265802 14167
rect 265502 -2523 265802 14049
rect 265502 -2641 265593 -2523
rect 265711 -2641 265802 -2523
rect 265502 -2683 265802 -2641
rect 265502 -2801 265593 -2683
rect 265711 -2801 265802 -2683
rect 265502 -2812 265802 -2801
rect 267302 340127 267602 355431
rect 276302 355239 276602 355720
rect 276302 355121 276393 355239
rect 276511 355121 276602 355239
rect 276302 355079 276602 355121
rect 276302 354961 276393 355079
rect 276511 354961 276602 355079
rect 274502 354299 274802 354780
rect 274502 354181 274593 354299
rect 274711 354181 274802 354299
rect 274502 354139 274802 354181
rect 274502 354021 274593 354139
rect 274711 354021 274802 354139
rect 272702 353359 273002 353840
rect 272702 353241 272793 353359
rect 272911 353241 273002 353359
rect 272702 353199 273002 353241
rect 272702 353081 272793 353199
rect 272911 353081 273002 353199
rect 267302 340009 267393 340127
rect 267511 340009 267602 340127
rect 267302 339967 267602 340009
rect 267302 339849 267393 339967
rect 267511 339849 267602 339967
rect 267302 322127 267602 339849
rect 267302 322009 267393 322127
rect 267511 322009 267602 322127
rect 267302 321967 267602 322009
rect 267302 321849 267393 321967
rect 267511 321849 267602 321967
rect 267302 304127 267602 321849
rect 267302 304009 267393 304127
rect 267511 304009 267602 304127
rect 267302 303967 267602 304009
rect 267302 303849 267393 303967
rect 267511 303849 267602 303967
rect 267302 286127 267602 303849
rect 267302 286009 267393 286127
rect 267511 286009 267602 286127
rect 267302 285967 267602 286009
rect 267302 285849 267393 285967
rect 267511 285849 267602 285967
rect 267302 268127 267602 285849
rect 267302 268009 267393 268127
rect 267511 268009 267602 268127
rect 267302 267967 267602 268009
rect 267302 267849 267393 267967
rect 267511 267849 267602 267967
rect 267302 250127 267602 267849
rect 267302 250009 267393 250127
rect 267511 250009 267602 250127
rect 267302 249967 267602 250009
rect 267302 249849 267393 249967
rect 267511 249849 267602 249967
rect 267302 232127 267602 249849
rect 267302 232009 267393 232127
rect 267511 232009 267602 232127
rect 267302 231967 267602 232009
rect 267302 231849 267393 231967
rect 267511 231849 267602 231967
rect 267302 214127 267602 231849
rect 267302 214009 267393 214127
rect 267511 214009 267602 214127
rect 267302 213967 267602 214009
rect 267302 213849 267393 213967
rect 267511 213849 267602 213967
rect 267302 196127 267602 213849
rect 267302 196009 267393 196127
rect 267511 196009 267602 196127
rect 267302 195967 267602 196009
rect 267302 195849 267393 195967
rect 267511 195849 267602 195967
rect 267302 178127 267602 195849
rect 267302 178009 267393 178127
rect 267511 178009 267602 178127
rect 267302 177967 267602 178009
rect 267302 177849 267393 177967
rect 267511 177849 267602 177967
rect 267302 160127 267602 177849
rect 267302 160009 267393 160127
rect 267511 160009 267602 160127
rect 267302 159967 267602 160009
rect 267302 159849 267393 159967
rect 267511 159849 267602 159967
rect 267302 142127 267602 159849
rect 267302 142009 267393 142127
rect 267511 142009 267602 142127
rect 267302 141967 267602 142009
rect 267302 141849 267393 141967
rect 267511 141849 267602 141967
rect 267302 124127 267602 141849
rect 267302 124009 267393 124127
rect 267511 124009 267602 124127
rect 267302 123967 267602 124009
rect 267302 123849 267393 123967
rect 267511 123849 267602 123967
rect 267302 106127 267602 123849
rect 267302 106009 267393 106127
rect 267511 106009 267602 106127
rect 267302 105967 267602 106009
rect 267302 105849 267393 105967
rect 267511 105849 267602 105967
rect 267302 88127 267602 105849
rect 267302 88009 267393 88127
rect 267511 88009 267602 88127
rect 267302 87967 267602 88009
rect 267302 87849 267393 87967
rect 267511 87849 267602 87967
rect 267302 70127 267602 87849
rect 267302 70009 267393 70127
rect 267511 70009 267602 70127
rect 267302 69967 267602 70009
rect 267302 69849 267393 69967
rect 267511 69849 267602 69967
rect 267302 52127 267602 69849
rect 267302 52009 267393 52127
rect 267511 52009 267602 52127
rect 267302 51967 267602 52009
rect 267302 51849 267393 51967
rect 267511 51849 267602 51967
rect 267302 34127 267602 51849
rect 267302 34009 267393 34127
rect 267511 34009 267602 34127
rect 267302 33967 267602 34009
rect 267302 33849 267393 33967
rect 267511 33849 267602 33967
rect 267302 16127 267602 33849
rect 267302 16009 267393 16127
rect 267511 16009 267602 16127
rect 267302 15967 267602 16009
rect 267302 15849 267393 15967
rect 267511 15849 267602 15967
rect 258302 -3111 258393 -2993
rect 258511 -3111 258602 -2993
rect 258302 -3153 258602 -3111
rect 258302 -3271 258393 -3153
rect 258511 -3271 258602 -3153
rect 258302 -3752 258602 -3271
rect 267302 -3463 267602 15849
rect 270902 352419 271202 352900
rect 270902 352301 270993 352419
rect 271111 352301 271202 352419
rect 270902 352259 271202 352301
rect 270902 352141 270993 352259
rect 271111 352141 271202 352259
rect 270902 343727 271202 352141
rect 270902 343609 270993 343727
rect 271111 343609 271202 343727
rect 270902 343567 271202 343609
rect 270902 343449 270993 343567
rect 271111 343449 271202 343567
rect 270902 325727 271202 343449
rect 270902 325609 270993 325727
rect 271111 325609 271202 325727
rect 270902 325567 271202 325609
rect 270902 325449 270993 325567
rect 271111 325449 271202 325567
rect 270902 307727 271202 325449
rect 270902 307609 270993 307727
rect 271111 307609 271202 307727
rect 270902 307567 271202 307609
rect 270902 307449 270993 307567
rect 271111 307449 271202 307567
rect 270902 289727 271202 307449
rect 270902 289609 270993 289727
rect 271111 289609 271202 289727
rect 270902 289567 271202 289609
rect 270902 289449 270993 289567
rect 271111 289449 271202 289567
rect 270902 271727 271202 289449
rect 270902 271609 270993 271727
rect 271111 271609 271202 271727
rect 270902 271567 271202 271609
rect 270902 271449 270993 271567
rect 271111 271449 271202 271567
rect 270902 253727 271202 271449
rect 270902 253609 270993 253727
rect 271111 253609 271202 253727
rect 270902 253567 271202 253609
rect 270902 253449 270993 253567
rect 271111 253449 271202 253567
rect 270902 235727 271202 253449
rect 270902 235609 270993 235727
rect 271111 235609 271202 235727
rect 270902 235567 271202 235609
rect 270902 235449 270993 235567
rect 271111 235449 271202 235567
rect 270902 217727 271202 235449
rect 270902 217609 270993 217727
rect 271111 217609 271202 217727
rect 270902 217567 271202 217609
rect 270902 217449 270993 217567
rect 271111 217449 271202 217567
rect 270902 199727 271202 217449
rect 270902 199609 270993 199727
rect 271111 199609 271202 199727
rect 270902 199567 271202 199609
rect 270902 199449 270993 199567
rect 271111 199449 271202 199567
rect 270902 181727 271202 199449
rect 270902 181609 270993 181727
rect 271111 181609 271202 181727
rect 270902 181567 271202 181609
rect 270902 181449 270993 181567
rect 271111 181449 271202 181567
rect 270902 163727 271202 181449
rect 270902 163609 270993 163727
rect 271111 163609 271202 163727
rect 270902 163567 271202 163609
rect 270902 163449 270993 163567
rect 271111 163449 271202 163567
rect 270902 145727 271202 163449
rect 270902 145609 270993 145727
rect 271111 145609 271202 145727
rect 270902 145567 271202 145609
rect 270902 145449 270993 145567
rect 271111 145449 271202 145567
rect 270902 127727 271202 145449
rect 270902 127609 270993 127727
rect 271111 127609 271202 127727
rect 270902 127567 271202 127609
rect 270902 127449 270993 127567
rect 271111 127449 271202 127567
rect 270902 109727 271202 127449
rect 270902 109609 270993 109727
rect 271111 109609 271202 109727
rect 270902 109567 271202 109609
rect 270902 109449 270993 109567
rect 271111 109449 271202 109567
rect 270902 91727 271202 109449
rect 270902 91609 270993 91727
rect 271111 91609 271202 91727
rect 270902 91567 271202 91609
rect 270902 91449 270993 91567
rect 271111 91449 271202 91567
rect 270902 73727 271202 91449
rect 270902 73609 270993 73727
rect 271111 73609 271202 73727
rect 270902 73567 271202 73609
rect 270902 73449 270993 73567
rect 271111 73449 271202 73567
rect 270902 55727 271202 73449
rect 270902 55609 270993 55727
rect 271111 55609 271202 55727
rect 270902 55567 271202 55609
rect 270902 55449 270993 55567
rect 271111 55449 271202 55567
rect 270902 37727 271202 55449
rect 270902 37609 270993 37727
rect 271111 37609 271202 37727
rect 270902 37567 271202 37609
rect 270902 37449 270993 37567
rect 271111 37449 271202 37567
rect 270902 19727 271202 37449
rect 270902 19609 270993 19727
rect 271111 19609 271202 19727
rect 270902 19567 271202 19609
rect 270902 19449 270993 19567
rect 271111 19449 271202 19567
rect 270902 1727 271202 19449
rect 270902 1609 270993 1727
rect 271111 1609 271202 1727
rect 270902 1567 271202 1609
rect 270902 1449 270993 1567
rect 271111 1449 271202 1567
rect 270902 -173 271202 1449
rect 270902 -291 270993 -173
rect 271111 -291 271202 -173
rect 270902 -333 271202 -291
rect 270902 -451 270993 -333
rect 271111 -451 271202 -333
rect 270902 -932 271202 -451
rect 272702 345527 273002 353081
rect 272702 345409 272793 345527
rect 272911 345409 273002 345527
rect 272702 345367 273002 345409
rect 272702 345249 272793 345367
rect 272911 345249 273002 345367
rect 272702 327527 273002 345249
rect 272702 327409 272793 327527
rect 272911 327409 273002 327527
rect 272702 327367 273002 327409
rect 272702 327249 272793 327367
rect 272911 327249 273002 327367
rect 272702 309527 273002 327249
rect 272702 309409 272793 309527
rect 272911 309409 273002 309527
rect 272702 309367 273002 309409
rect 272702 309249 272793 309367
rect 272911 309249 273002 309367
rect 272702 291527 273002 309249
rect 272702 291409 272793 291527
rect 272911 291409 273002 291527
rect 272702 291367 273002 291409
rect 272702 291249 272793 291367
rect 272911 291249 273002 291367
rect 272702 273527 273002 291249
rect 272702 273409 272793 273527
rect 272911 273409 273002 273527
rect 272702 273367 273002 273409
rect 272702 273249 272793 273367
rect 272911 273249 273002 273367
rect 272702 255527 273002 273249
rect 272702 255409 272793 255527
rect 272911 255409 273002 255527
rect 272702 255367 273002 255409
rect 272702 255249 272793 255367
rect 272911 255249 273002 255367
rect 272702 237527 273002 255249
rect 272702 237409 272793 237527
rect 272911 237409 273002 237527
rect 272702 237367 273002 237409
rect 272702 237249 272793 237367
rect 272911 237249 273002 237367
rect 272702 219527 273002 237249
rect 272702 219409 272793 219527
rect 272911 219409 273002 219527
rect 272702 219367 273002 219409
rect 272702 219249 272793 219367
rect 272911 219249 273002 219367
rect 272702 201527 273002 219249
rect 272702 201409 272793 201527
rect 272911 201409 273002 201527
rect 272702 201367 273002 201409
rect 272702 201249 272793 201367
rect 272911 201249 273002 201367
rect 272702 183527 273002 201249
rect 272702 183409 272793 183527
rect 272911 183409 273002 183527
rect 272702 183367 273002 183409
rect 272702 183249 272793 183367
rect 272911 183249 273002 183367
rect 272702 165527 273002 183249
rect 272702 165409 272793 165527
rect 272911 165409 273002 165527
rect 272702 165367 273002 165409
rect 272702 165249 272793 165367
rect 272911 165249 273002 165367
rect 272702 147527 273002 165249
rect 272702 147409 272793 147527
rect 272911 147409 273002 147527
rect 272702 147367 273002 147409
rect 272702 147249 272793 147367
rect 272911 147249 273002 147367
rect 272702 129527 273002 147249
rect 272702 129409 272793 129527
rect 272911 129409 273002 129527
rect 272702 129367 273002 129409
rect 272702 129249 272793 129367
rect 272911 129249 273002 129367
rect 272702 111527 273002 129249
rect 272702 111409 272793 111527
rect 272911 111409 273002 111527
rect 272702 111367 273002 111409
rect 272702 111249 272793 111367
rect 272911 111249 273002 111367
rect 272702 93527 273002 111249
rect 272702 93409 272793 93527
rect 272911 93409 273002 93527
rect 272702 93367 273002 93409
rect 272702 93249 272793 93367
rect 272911 93249 273002 93367
rect 272702 75527 273002 93249
rect 272702 75409 272793 75527
rect 272911 75409 273002 75527
rect 272702 75367 273002 75409
rect 272702 75249 272793 75367
rect 272911 75249 273002 75367
rect 272702 57527 273002 75249
rect 272702 57409 272793 57527
rect 272911 57409 273002 57527
rect 272702 57367 273002 57409
rect 272702 57249 272793 57367
rect 272911 57249 273002 57367
rect 272702 39527 273002 57249
rect 272702 39409 272793 39527
rect 272911 39409 273002 39527
rect 272702 39367 273002 39409
rect 272702 39249 272793 39367
rect 272911 39249 273002 39367
rect 272702 21527 273002 39249
rect 272702 21409 272793 21527
rect 272911 21409 273002 21527
rect 272702 21367 273002 21409
rect 272702 21249 272793 21367
rect 272911 21249 273002 21367
rect 272702 3527 273002 21249
rect 272702 3409 272793 3527
rect 272911 3409 273002 3527
rect 272702 3367 273002 3409
rect 272702 3249 272793 3367
rect 272911 3249 273002 3367
rect 272702 -1113 273002 3249
rect 272702 -1231 272793 -1113
rect 272911 -1231 273002 -1113
rect 272702 -1273 273002 -1231
rect 272702 -1391 272793 -1273
rect 272911 -1391 273002 -1273
rect 272702 -1872 273002 -1391
rect 274502 347327 274802 354021
rect 274502 347209 274593 347327
rect 274711 347209 274802 347327
rect 274502 347167 274802 347209
rect 274502 347049 274593 347167
rect 274711 347049 274802 347167
rect 274502 329327 274802 347049
rect 274502 329209 274593 329327
rect 274711 329209 274802 329327
rect 274502 329167 274802 329209
rect 274502 329049 274593 329167
rect 274711 329049 274802 329167
rect 274502 311327 274802 329049
rect 274502 311209 274593 311327
rect 274711 311209 274802 311327
rect 274502 311167 274802 311209
rect 274502 311049 274593 311167
rect 274711 311049 274802 311167
rect 274502 293327 274802 311049
rect 274502 293209 274593 293327
rect 274711 293209 274802 293327
rect 274502 293167 274802 293209
rect 274502 293049 274593 293167
rect 274711 293049 274802 293167
rect 274502 275327 274802 293049
rect 274502 275209 274593 275327
rect 274711 275209 274802 275327
rect 274502 275167 274802 275209
rect 274502 275049 274593 275167
rect 274711 275049 274802 275167
rect 274502 257327 274802 275049
rect 274502 257209 274593 257327
rect 274711 257209 274802 257327
rect 274502 257167 274802 257209
rect 274502 257049 274593 257167
rect 274711 257049 274802 257167
rect 274502 239327 274802 257049
rect 274502 239209 274593 239327
rect 274711 239209 274802 239327
rect 274502 239167 274802 239209
rect 274502 239049 274593 239167
rect 274711 239049 274802 239167
rect 274502 221327 274802 239049
rect 274502 221209 274593 221327
rect 274711 221209 274802 221327
rect 274502 221167 274802 221209
rect 274502 221049 274593 221167
rect 274711 221049 274802 221167
rect 274502 203327 274802 221049
rect 274502 203209 274593 203327
rect 274711 203209 274802 203327
rect 274502 203167 274802 203209
rect 274502 203049 274593 203167
rect 274711 203049 274802 203167
rect 274502 185327 274802 203049
rect 274502 185209 274593 185327
rect 274711 185209 274802 185327
rect 274502 185167 274802 185209
rect 274502 185049 274593 185167
rect 274711 185049 274802 185167
rect 274502 167327 274802 185049
rect 274502 167209 274593 167327
rect 274711 167209 274802 167327
rect 274502 167167 274802 167209
rect 274502 167049 274593 167167
rect 274711 167049 274802 167167
rect 274502 149327 274802 167049
rect 274502 149209 274593 149327
rect 274711 149209 274802 149327
rect 274502 149167 274802 149209
rect 274502 149049 274593 149167
rect 274711 149049 274802 149167
rect 274502 131327 274802 149049
rect 274502 131209 274593 131327
rect 274711 131209 274802 131327
rect 274502 131167 274802 131209
rect 274502 131049 274593 131167
rect 274711 131049 274802 131167
rect 274502 113327 274802 131049
rect 274502 113209 274593 113327
rect 274711 113209 274802 113327
rect 274502 113167 274802 113209
rect 274502 113049 274593 113167
rect 274711 113049 274802 113167
rect 274502 95327 274802 113049
rect 274502 95209 274593 95327
rect 274711 95209 274802 95327
rect 274502 95167 274802 95209
rect 274502 95049 274593 95167
rect 274711 95049 274802 95167
rect 274502 77327 274802 95049
rect 274502 77209 274593 77327
rect 274711 77209 274802 77327
rect 274502 77167 274802 77209
rect 274502 77049 274593 77167
rect 274711 77049 274802 77167
rect 274502 59327 274802 77049
rect 274502 59209 274593 59327
rect 274711 59209 274802 59327
rect 274502 59167 274802 59209
rect 274502 59049 274593 59167
rect 274711 59049 274802 59167
rect 274502 41327 274802 59049
rect 274502 41209 274593 41327
rect 274711 41209 274802 41327
rect 274502 41167 274802 41209
rect 274502 41049 274593 41167
rect 274711 41049 274802 41167
rect 274502 23327 274802 41049
rect 274502 23209 274593 23327
rect 274711 23209 274802 23327
rect 274502 23167 274802 23209
rect 274502 23049 274593 23167
rect 274711 23049 274802 23167
rect 274502 5327 274802 23049
rect 274502 5209 274593 5327
rect 274711 5209 274802 5327
rect 274502 5167 274802 5209
rect 274502 5049 274593 5167
rect 274711 5049 274802 5167
rect 274502 -2053 274802 5049
rect 274502 -2171 274593 -2053
rect 274711 -2171 274802 -2053
rect 274502 -2213 274802 -2171
rect 274502 -2331 274593 -2213
rect 274711 -2331 274802 -2213
rect 274502 -2812 274802 -2331
rect 276302 349127 276602 354961
rect 285302 355709 285602 355720
rect 285302 355591 285393 355709
rect 285511 355591 285602 355709
rect 285302 355549 285602 355591
rect 285302 355431 285393 355549
rect 285511 355431 285602 355549
rect 283502 354769 283802 354780
rect 283502 354651 283593 354769
rect 283711 354651 283802 354769
rect 283502 354609 283802 354651
rect 283502 354491 283593 354609
rect 283711 354491 283802 354609
rect 281702 353829 282002 353840
rect 281702 353711 281793 353829
rect 281911 353711 282002 353829
rect 281702 353669 282002 353711
rect 281702 353551 281793 353669
rect 281911 353551 282002 353669
rect 276302 349009 276393 349127
rect 276511 349009 276602 349127
rect 276302 348967 276602 349009
rect 276302 348849 276393 348967
rect 276511 348849 276602 348967
rect 276302 331127 276602 348849
rect 276302 331009 276393 331127
rect 276511 331009 276602 331127
rect 276302 330967 276602 331009
rect 276302 330849 276393 330967
rect 276511 330849 276602 330967
rect 276302 313127 276602 330849
rect 276302 313009 276393 313127
rect 276511 313009 276602 313127
rect 276302 312967 276602 313009
rect 276302 312849 276393 312967
rect 276511 312849 276602 312967
rect 276302 295127 276602 312849
rect 276302 295009 276393 295127
rect 276511 295009 276602 295127
rect 276302 294967 276602 295009
rect 276302 294849 276393 294967
rect 276511 294849 276602 294967
rect 276302 277127 276602 294849
rect 276302 277009 276393 277127
rect 276511 277009 276602 277127
rect 276302 276967 276602 277009
rect 276302 276849 276393 276967
rect 276511 276849 276602 276967
rect 276302 259127 276602 276849
rect 276302 259009 276393 259127
rect 276511 259009 276602 259127
rect 276302 258967 276602 259009
rect 276302 258849 276393 258967
rect 276511 258849 276602 258967
rect 276302 241127 276602 258849
rect 276302 241009 276393 241127
rect 276511 241009 276602 241127
rect 276302 240967 276602 241009
rect 276302 240849 276393 240967
rect 276511 240849 276602 240967
rect 276302 223127 276602 240849
rect 276302 223009 276393 223127
rect 276511 223009 276602 223127
rect 276302 222967 276602 223009
rect 276302 222849 276393 222967
rect 276511 222849 276602 222967
rect 276302 205127 276602 222849
rect 276302 205009 276393 205127
rect 276511 205009 276602 205127
rect 276302 204967 276602 205009
rect 276302 204849 276393 204967
rect 276511 204849 276602 204967
rect 276302 187127 276602 204849
rect 276302 187009 276393 187127
rect 276511 187009 276602 187127
rect 276302 186967 276602 187009
rect 276302 186849 276393 186967
rect 276511 186849 276602 186967
rect 276302 169127 276602 186849
rect 276302 169009 276393 169127
rect 276511 169009 276602 169127
rect 276302 168967 276602 169009
rect 276302 168849 276393 168967
rect 276511 168849 276602 168967
rect 276302 151127 276602 168849
rect 276302 151009 276393 151127
rect 276511 151009 276602 151127
rect 276302 150967 276602 151009
rect 276302 150849 276393 150967
rect 276511 150849 276602 150967
rect 276302 133127 276602 150849
rect 276302 133009 276393 133127
rect 276511 133009 276602 133127
rect 276302 132967 276602 133009
rect 276302 132849 276393 132967
rect 276511 132849 276602 132967
rect 276302 115127 276602 132849
rect 276302 115009 276393 115127
rect 276511 115009 276602 115127
rect 276302 114967 276602 115009
rect 276302 114849 276393 114967
rect 276511 114849 276602 114967
rect 276302 97127 276602 114849
rect 276302 97009 276393 97127
rect 276511 97009 276602 97127
rect 276302 96967 276602 97009
rect 276302 96849 276393 96967
rect 276511 96849 276602 96967
rect 276302 79127 276602 96849
rect 276302 79009 276393 79127
rect 276511 79009 276602 79127
rect 276302 78967 276602 79009
rect 276302 78849 276393 78967
rect 276511 78849 276602 78967
rect 276302 61127 276602 78849
rect 276302 61009 276393 61127
rect 276511 61009 276602 61127
rect 276302 60967 276602 61009
rect 276302 60849 276393 60967
rect 276511 60849 276602 60967
rect 276302 43127 276602 60849
rect 276302 43009 276393 43127
rect 276511 43009 276602 43127
rect 276302 42967 276602 43009
rect 276302 42849 276393 42967
rect 276511 42849 276602 42967
rect 276302 25127 276602 42849
rect 276302 25009 276393 25127
rect 276511 25009 276602 25127
rect 276302 24967 276602 25009
rect 276302 24849 276393 24967
rect 276511 24849 276602 24967
rect 276302 7127 276602 24849
rect 276302 7009 276393 7127
rect 276511 7009 276602 7127
rect 276302 6967 276602 7009
rect 276302 6849 276393 6967
rect 276511 6849 276602 6967
rect 267302 -3581 267393 -3463
rect 267511 -3581 267602 -3463
rect 267302 -3623 267602 -3581
rect 267302 -3741 267393 -3623
rect 267511 -3741 267602 -3623
rect 267302 -3752 267602 -3741
rect 276302 -2993 276602 6849
rect 279902 352889 280202 352900
rect 279902 352771 279993 352889
rect 280111 352771 280202 352889
rect 279902 352729 280202 352771
rect 279902 352611 279993 352729
rect 280111 352611 280202 352729
rect 279902 334727 280202 352611
rect 279902 334609 279993 334727
rect 280111 334609 280202 334727
rect 279902 334567 280202 334609
rect 279902 334449 279993 334567
rect 280111 334449 280202 334567
rect 279902 316727 280202 334449
rect 279902 316609 279993 316727
rect 280111 316609 280202 316727
rect 279902 316567 280202 316609
rect 279902 316449 279993 316567
rect 280111 316449 280202 316567
rect 279902 298727 280202 316449
rect 279902 298609 279993 298727
rect 280111 298609 280202 298727
rect 279902 298567 280202 298609
rect 279902 298449 279993 298567
rect 280111 298449 280202 298567
rect 279902 280727 280202 298449
rect 279902 280609 279993 280727
rect 280111 280609 280202 280727
rect 279902 280567 280202 280609
rect 279902 280449 279993 280567
rect 280111 280449 280202 280567
rect 279902 262727 280202 280449
rect 279902 262609 279993 262727
rect 280111 262609 280202 262727
rect 279902 262567 280202 262609
rect 279902 262449 279993 262567
rect 280111 262449 280202 262567
rect 279902 244727 280202 262449
rect 279902 244609 279993 244727
rect 280111 244609 280202 244727
rect 279902 244567 280202 244609
rect 279902 244449 279993 244567
rect 280111 244449 280202 244567
rect 279902 226727 280202 244449
rect 279902 226609 279993 226727
rect 280111 226609 280202 226727
rect 279902 226567 280202 226609
rect 279902 226449 279993 226567
rect 280111 226449 280202 226567
rect 279902 208727 280202 226449
rect 279902 208609 279993 208727
rect 280111 208609 280202 208727
rect 279902 208567 280202 208609
rect 279902 208449 279993 208567
rect 280111 208449 280202 208567
rect 279902 190727 280202 208449
rect 279902 190609 279993 190727
rect 280111 190609 280202 190727
rect 279902 190567 280202 190609
rect 279902 190449 279993 190567
rect 280111 190449 280202 190567
rect 279902 172727 280202 190449
rect 279902 172609 279993 172727
rect 280111 172609 280202 172727
rect 279902 172567 280202 172609
rect 279902 172449 279993 172567
rect 280111 172449 280202 172567
rect 279902 154727 280202 172449
rect 279902 154609 279993 154727
rect 280111 154609 280202 154727
rect 279902 154567 280202 154609
rect 279902 154449 279993 154567
rect 280111 154449 280202 154567
rect 279902 136727 280202 154449
rect 279902 136609 279993 136727
rect 280111 136609 280202 136727
rect 279902 136567 280202 136609
rect 279902 136449 279993 136567
rect 280111 136449 280202 136567
rect 279902 118727 280202 136449
rect 279902 118609 279993 118727
rect 280111 118609 280202 118727
rect 279902 118567 280202 118609
rect 279902 118449 279993 118567
rect 280111 118449 280202 118567
rect 279902 100727 280202 118449
rect 279902 100609 279993 100727
rect 280111 100609 280202 100727
rect 279902 100567 280202 100609
rect 279902 100449 279993 100567
rect 280111 100449 280202 100567
rect 279902 82727 280202 100449
rect 279902 82609 279993 82727
rect 280111 82609 280202 82727
rect 279902 82567 280202 82609
rect 279902 82449 279993 82567
rect 280111 82449 280202 82567
rect 279902 64727 280202 82449
rect 279902 64609 279993 64727
rect 280111 64609 280202 64727
rect 279902 64567 280202 64609
rect 279902 64449 279993 64567
rect 280111 64449 280202 64567
rect 279902 46727 280202 64449
rect 279902 46609 279993 46727
rect 280111 46609 280202 46727
rect 279902 46567 280202 46609
rect 279902 46449 279993 46567
rect 280111 46449 280202 46567
rect 279902 28727 280202 46449
rect 279902 28609 279993 28727
rect 280111 28609 280202 28727
rect 279902 28567 280202 28609
rect 279902 28449 279993 28567
rect 280111 28449 280202 28567
rect 279902 10727 280202 28449
rect 279902 10609 279993 10727
rect 280111 10609 280202 10727
rect 279902 10567 280202 10609
rect 279902 10449 279993 10567
rect 280111 10449 280202 10567
rect 279902 -643 280202 10449
rect 279902 -761 279993 -643
rect 280111 -761 280202 -643
rect 279902 -803 280202 -761
rect 279902 -921 279993 -803
rect 280111 -921 280202 -803
rect 279902 -932 280202 -921
rect 281702 336527 282002 353551
rect 281702 336409 281793 336527
rect 281911 336409 282002 336527
rect 281702 336367 282002 336409
rect 281702 336249 281793 336367
rect 281911 336249 282002 336367
rect 281702 318527 282002 336249
rect 281702 318409 281793 318527
rect 281911 318409 282002 318527
rect 281702 318367 282002 318409
rect 281702 318249 281793 318367
rect 281911 318249 282002 318367
rect 281702 300527 282002 318249
rect 281702 300409 281793 300527
rect 281911 300409 282002 300527
rect 281702 300367 282002 300409
rect 281702 300249 281793 300367
rect 281911 300249 282002 300367
rect 281702 282527 282002 300249
rect 281702 282409 281793 282527
rect 281911 282409 282002 282527
rect 281702 282367 282002 282409
rect 281702 282249 281793 282367
rect 281911 282249 282002 282367
rect 281702 264527 282002 282249
rect 281702 264409 281793 264527
rect 281911 264409 282002 264527
rect 281702 264367 282002 264409
rect 281702 264249 281793 264367
rect 281911 264249 282002 264367
rect 281702 246527 282002 264249
rect 281702 246409 281793 246527
rect 281911 246409 282002 246527
rect 281702 246367 282002 246409
rect 281702 246249 281793 246367
rect 281911 246249 282002 246367
rect 281702 228527 282002 246249
rect 281702 228409 281793 228527
rect 281911 228409 282002 228527
rect 281702 228367 282002 228409
rect 281702 228249 281793 228367
rect 281911 228249 282002 228367
rect 281702 210527 282002 228249
rect 281702 210409 281793 210527
rect 281911 210409 282002 210527
rect 281702 210367 282002 210409
rect 281702 210249 281793 210367
rect 281911 210249 282002 210367
rect 281702 192527 282002 210249
rect 281702 192409 281793 192527
rect 281911 192409 282002 192527
rect 281702 192367 282002 192409
rect 281702 192249 281793 192367
rect 281911 192249 282002 192367
rect 281702 174527 282002 192249
rect 281702 174409 281793 174527
rect 281911 174409 282002 174527
rect 281702 174367 282002 174409
rect 281702 174249 281793 174367
rect 281911 174249 282002 174367
rect 281702 156527 282002 174249
rect 281702 156409 281793 156527
rect 281911 156409 282002 156527
rect 281702 156367 282002 156409
rect 281702 156249 281793 156367
rect 281911 156249 282002 156367
rect 281702 138527 282002 156249
rect 281702 138409 281793 138527
rect 281911 138409 282002 138527
rect 281702 138367 282002 138409
rect 281702 138249 281793 138367
rect 281911 138249 282002 138367
rect 281702 120527 282002 138249
rect 281702 120409 281793 120527
rect 281911 120409 282002 120527
rect 281702 120367 282002 120409
rect 281702 120249 281793 120367
rect 281911 120249 282002 120367
rect 281702 102527 282002 120249
rect 281702 102409 281793 102527
rect 281911 102409 282002 102527
rect 281702 102367 282002 102409
rect 281702 102249 281793 102367
rect 281911 102249 282002 102367
rect 281702 84527 282002 102249
rect 281702 84409 281793 84527
rect 281911 84409 282002 84527
rect 281702 84367 282002 84409
rect 281702 84249 281793 84367
rect 281911 84249 282002 84367
rect 281702 66527 282002 84249
rect 281702 66409 281793 66527
rect 281911 66409 282002 66527
rect 281702 66367 282002 66409
rect 281702 66249 281793 66367
rect 281911 66249 282002 66367
rect 281702 48527 282002 66249
rect 281702 48409 281793 48527
rect 281911 48409 282002 48527
rect 281702 48367 282002 48409
rect 281702 48249 281793 48367
rect 281911 48249 282002 48367
rect 281702 30527 282002 48249
rect 281702 30409 281793 30527
rect 281911 30409 282002 30527
rect 281702 30367 282002 30409
rect 281702 30249 281793 30367
rect 281911 30249 282002 30367
rect 281702 12527 282002 30249
rect 281702 12409 281793 12527
rect 281911 12409 282002 12527
rect 281702 12367 282002 12409
rect 281702 12249 281793 12367
rect 281911 12249 282002 12367
rect 281702 -1583 282002 12249
rect 281702 -1701 281793 -1583
rect 281911 -1701 282002 -1583
rect 281702 -1743 282002 -1701
rect 281702 -1861 281793 -1743
rect 281911 -1861 282002 -1743
rect 281702 -1872 282002 -1861
rect 283502 338327 283802 354491
rect 283502 338209 283593 338327
rect 283711 338209 283802 338327
rect 283502 338167 283802 338209
rect 283502 338049 283593 338167
rect 283711 338049 283802 338167
rect 283502 320327 283802 338049
rect 283502 320209 283593 320327
rect 283711 320209 283802 320327
rect 283502 320167 283802 320209
rect 283502 320049 283593 320167
rect 283711 320049 283802 320167
rect 283502 302327 283802 320049
rect 283502 302209 283593 302327
rect 283711 302209 283802 302327
rect 283502 302167 283802 302209
rect 283502 302049 283593 302167
rect 283711 302049 283802 302167
rect 283502 284327 283802 302049
rect 283502 284209 283593 284327
rect 283711 284209 283802 284327
rect 283502 284167 283802 284209
rect 283502 284049 283593 284167
rect 283711 284049 283802 284167
rect 283502 266327 283802 284049
rect 283502 266209 283593 266327
rect 283711 266209 283802 266327
rect 283502 266167 283802 266209
rect 283502 266049 283593 266167
rect 283711 266049 283802 266167
rect 283502 248327 283802 266049
rect 283502 248209 283593 248327
rect 283711 248209 283802 248327
rect 283502 248167 283802 248209
rect 283502 248049 283593 248167
rect 283711 248049 283802 248167
rect 283502 230327 283802 248049
rect 283502 230209 283593 230327
rect 283711 230209 283802 230327
rect 283502 230167 283802 230209
rect 283502 230049 283593 230167
rect 283711 230049 283802 230167
rect 283502 212327 283802 230049
rect 283502 212209 283593 212327
rect 283711 212209 283802 212327
rect 283502 212167 283802 212209
rect 283502 212049 283593 212167
rect 283711 212049 283802 212167
rect 283502 194327 283802 212049
rect 283502 194209 283593 194327
rect 283711 194209 283802 194327
rect 283502 194167 283802 194209
rect 283502 194049 283593 194167
rect 283711 194049 283802 194167
rect 283502 176327 283802 194049
rect 283502 176209 283593 176327
rect 283711 176209 283802 176327
rect 283502 176167 283802 176209
rect 283502 176049 283593 176167
rect 283711 176049 283802 176167
rect 283502 158327 283802 176049
rect 283502 158209 283593 158327
rect 283711 158209 283802 158327
rect 283502 158167 283802 158209
rect 283502 158049 283593 158167
rect 283711 158049 283802 158167
rect 283502 140327 283802 158049
rect 283502 140209 283593 140327
rect 283711 140209 283802 140327
rect 283502 140167 283802 140209
rect 283502 140049 283593 140167
rect 283711 140049 283802 140167
rect 283502 122327 283802 140049
rect 283502 122209 283593 122327
rect 283711 122209 283802 122327
rect 283502 122167 283802 122209
rect 283502 122049 283593 122167
rect 283711 122049 283802 122167
rect 283502 104327 283802 122049
rect 283502 104209 283593 104327
rect 283711 104209 283802 104327
rect 283502 104167 283802 104209
rect 283502 104049 283593 104167
rect 283711 104049 283802 104167
rect 283502 86327 283802 104049
rect 283502 86209 283593 86327
rect 283711 86209 283802 86327
rect 283502 86167 283802 86209
rect 283502 86049 283593 86167
rect 283711 86049 283802 86167
rect 283502 68327 283802 86049
rect 283502 68209 283593 68327
rect 283711 68209 283802 68327
rect 283502 68167 283802 68209
rect 283502 68049 283593 68167
rect 283711 68049 283802 68167
rect 283502 50327 283802 68049
rect 283502 50209 283593 50327
rect 283711 50209 283802 50327
rect 283502 50167 283802 50209
rect 283502 50049 283593 50167
rect 283711 50049 283802 50167
rect 283502 32327 283802 50049
rect 283502 32209 283593 32327
rect 283711 32209 283802 32327
rect 283502 32167 283802 32209
rect 283502 32049 283593 32167
rect 283711 32049 283802 32167
rect 283502 14327 283802 32049
rect 283502 14209 283593 14327
rect 283711 14209 283802 14327
rect 283502 14167 283802 14209
rect 283502 14049 283593 14167
rect 283711 14049 283802 14167
rect 283502 -2523 283802 14049
rect 283502 -2641 283593 -2523
rect 283711 -2641 283802 -2523
rect 283502 -2683 283802 -2641
rect 283502 -2801 283593 -2683
rect 283711 -2801 283802 -2683
rect 283502 -2812 283802 -2801
rect 285302 340127 285602 355431
rect 295950 355709 296250 355720
rect 295950 355591 296041 355709
rect 296159 355591 296250 355709
rect 295950 355549 296250 355591
rect 295950 355431 296041 355549
rect 296159 355431 296250 355549
rect 295480 355239 295780 355250
rect 295480 355121 295571 355239
rect 295689 355121 295780 355239
rect 295480 355079 295780 355121
rect 295480 354961 295571 355079
rect 295689 354961 295780 355079
rect 295010 354769 295310 354780
rect 295010 354651 295101 354769
rect 295219 354651 295310 354769
rect 295010 354609 295310 354651
rect 295010 354491 295101 354609
rect 295219 354491 295310 354609
rect 294540 354299 294840 354310
rect 294540 354181 294631 354299
rect 294749 354181 294840 354299
rect 294540 354139 294840 354181
rect 294540 354021 294631 354139
rect 294749 354021 294840 354139
rect 290702 353359 291002 353840
rect 294070 353829 294370 353840
rect 294070 353711 294161 353829
rect 294279 353711 294370 353829
rect 294070 353669 294370 353711
rect 294070 353551 294161 353669
rect 294279 353551 294370 353669
rect 290702 353241 290793 353359
rect 290911 353241 291002 353359
rect 290702 353199 291002 353241
rect 290702 353081 290793 353199
rect 290911 353081 291002 353199
rect 285302 340009 285393 340127
rect 285511 340009 285602 340127
rect 285302 339967 285602 340009
rect 285302 339849 285393 339967
rect 285511 339849 285602 339967
rect 285302 322127 285602 339849
rect 285302 322009 285393 322127
rect 285511 322009 285602 322127
rect 285302 321967 285602 322009
rect 285302 321849 285393 321967
rect 285511 321849 285602 321967
rect 285302 304127 285602 321849
rect 285302 304009 285393 304127
rect 285511 304009 285602 304127
rect 285302 303967 285602 304009
rect 285302 303849 285393 303967
rect 285511 303849 285602 303967
rect 285302 286127 285602 303849
rect 285302 286009 285393 286127
rect 285511 286009 285602 286127
rect 285302 285967 285602 286009
rect 285302 285849 285393 285967
rect 285511 285849 285602 285967
rect 285302 268127 285602 285849
rect 285302 268009 285393 268127
rect 285511 268009 285602 268127
rect 285302 267967 285602 268009
rect 285302 267849 285393 267967
rect 285511 267849 285602 267967
rect 285302 250127 285602 267849
rect 285302 250009 285393 250127
rect 285511 250009 285602 250127
rect 285302 249967 285602 250009
rect 285302 249849 285393 249967
rect 285511 249849 285602 249967
rect 285302 232127 285602 249849
rect 285302 232009 285393 232127
rect 285511 232009 285602 232127
rect 285302 231967 285602 232009
rect 285302 231849 285393 231967
rect 285511 231849 285602 231967
rect 285302 214127 285602 231849
rect 285302 214009 285393 214127
rect 285511 214009 285602 214127
rect 285302 213967 285602 214009
rect 285302 213849 285393 213967
rect 285511 213849 285602 213967
rect 285302 196127 285602 213849
rect 285302 196009 285393 196127
rect 285511 196009 285602 196127
rect 285302 195967 285602 196009
rect 285302 195849 285393 195967
rect 285511 195849 285602 195967
rect 285302 178127 285602 195849
rect 285302 178009 285393 178127
rect 285511 178009 285602 178127
rect 285302 177967 285602 178009
rect 285302 177849 285393 177967
rect 285511 177849 285602 177967
rect 285302 160127 285602 177849
rect 285302 160009 285393 160127
rect 285511 160009 285602 160127
rect 285302 159967 285602 160009
rect 285302 159849 285393 159967
rect 285511 159849 285602 159967
rect 285302 142127 285602 159849
rect 285302 142009 285393 142127
rect 285511 142009 285602 142127
rect 285302 141967 285602 142009
rect 285302 141849 285393 141967
rect 285511 141849 285602 141967
rect 285302 124127 285602 141849
rect 285302 124009 285393 124127
rect 285511 124009 285602 124127
rect 285302 123967 285602 124009
rect 285302 123849 285393 123967
rect 285511 123849 285602 123967
rect 285302 106127 285602 123849
rect 285302 106009 285393 106127
rect 285511 106009 285602 106127
rect 285302 105967 285602 106009
rect 285302 105849 285393 105967
rect 285511 105849 285602 105967
rect 285302 88127 285602 105849
rect 285302 88009 285393 88127
rect 285511 88009 285602 88127
rect 285302 87967 285602 88009
rect 285302 87849 285393 87967
rect 285511 87849 285602 87967
rect 285302 70127 285602 87849
rect 285302 70009 285393 70127
rect 285511 70009 285602 70127
rect 285302 69967 285602 70009
rect 285302 69849 285393 69967
rect 285511 69849 285602 69967
rect 285302 52127 285602 69849
rect 285302 52009 285393 52127
rect 285511 52009 285602 52127
rect 285302 51967 285602 52009
rect 285302 51849 285393 51967
rect 285511 51849 285602 51967
rect 285302 34127 285602 51849
rect 285302 34009 285393 34127
rect 285511 34009 285602 34127
rect 285302 33967 285602 34009
rect 285302 33849 285393 33967
rect 285511 33849 285602 33967
rect 285302 16127 285602 33849
rect 285302 16009 285393 16127
rect 285511 16009 285602 16127
rect 285302 15967 285602 16009
rect 285302 15849 285393 15967
rect 285511 15849 285602 15967
rect 276302 -3111 276393 -2993
rect 276511 -3111 276602 -2993
rect 276302 -3153 276602 -3111
rect 276302 -3271 276393 -3153
rect 276511 -3271 276602 -3153
rect 276302 -3752 276602 -3271
rect 285302 -3463 285602 15849
rect 288902 352419 289202 352900
rect 288902 352301 288993 352419
rect 289111 352301 289202 352419
rect 288902 352259 289202 352301
rect 288902 352141 288993 352259
rect 289111 352141 289202 352259
rect 288902 343727 289202 352141
rect 288902 343609 288993 343727
rect 289111 343609 289202 343727
rect 288902 343567 289202 343609
rect 288902 343449 288993 343567
rect 289111 343449 289202 343567
rect 288902 325727 289202 343449
rect 288902 325609 288993 325727
rect 289111 325609 289202 325727
rect 288902 325567 289202 325609
rect 288902 325449 288993 325567
rect 289111 325449 289202 325567
rect 288902 307727 289202 325449
rect 288902 307609 288993 307727
rect 289111 307609 289202 307727
rect 288902 307567 289202 307609
rect 288902 307449 288993 307567
rect 289111 307449 289202 307567
rect 288902 289727 289202 307449
rect 288902 289609 288993 289727
rect 289111 289609 289202 289727
rect 288902 289567 289202 289609
rect 288902 289449 288993 289567
rect 289111 289449 289202 289567
rect 288902 271727 289202 289449
rect 288902 271609 288993 271727
rect 289111 271609 289202 271727
rect 288902 271567 289202 271609
rect 288902 271449 288993 271567
rect 289111 271449 289202 271567
rect 288902 253727 289202 271449
rect 288902 253609 288993 253727
rect 289111 253609 289202 253727
rect 288902 253567 289202 253609
rect 288902 253449 288993 253567
rect 289111 253449 289202 253567
rect 288902 235727 289202 253449
rect 288902 235609 288993 235727
rect 289111 235609 289202 235727
rect 288902 235567 289202 235609
rect 288902 235449 288993 235567
rect 289111 235449 289202 235567
rect 288902 217727 289202 235449
rect 288902 217609 288993 217727
rect 289111 217609 289202 217727
rect 288902 217567 289202 217609
rect 288902 217449 288993 217567
rect 289111 217449 289202 217567
rect 288902 199727 289202 217449
rect 288902 199609 288993 199727
rect 289111 199609 289202 199727
rect 288902 199567 289202 199609
rect 288902 199449 288993 199567
rect 289111 199449 289202 199567
rect 288902 181727 289202 199449
rect 288902 181609 288993 181727
rect 289111 181609 289202 181727
rect 288902 181567 289202 181609
rect 288902 181449 288993 181567
rect 289111 181449 289202 181567
rect 288902 163727 289202 181449
rect 288902 163609 288993 163727
rect 289111 163609 289202 163727
rect 288902 163567 289202 163609
rect 288902 163449 288993 163567
rect 289111 163449 289202 163567
rect 288902 145727 289202 163449
rect 288902 145609 288993 145727
rect 289111 145609 289202 145727
rect 288902 145567 289202 145609
rect 288902 145449 288993 145567
rect 289111 145449 289202 145567
rect 288902 127727 289202 145449
rect 288902 127609 288993 127727
rect 289111 127609 289202 127727
rect 288902 127567 289202 127609
rect 288902 127449 288993 127567
rect 289111 127449 289202 127567
rect 288902 109727 289202 127449
rect 288902 109609 288993 109727
rect 289111 109609 289202 109727
rect 288902 109567 289202 109609
rect 288902 109449 288993 109567
rect 289111 109449 289202 109567
rect 288902 91727 289202 109449
rect 288902 91609 288993 91727
rect 289111 91609 289202 91727
rect 288902 91567 289202 91609
rect 288902 91449 288993 91567
rect 289111 91449 289202 91567
rect 288902 73727 289202 91449
rect 288902 73609 288993 73727
rect 289111 73609 289202 73727
rect 288902 73567 289202 73609
rect 288902 73449 288993 73567
rect 289111 73449 289202 73567
rect 288902 55727 289202 73449
rect 288902 55609 288993 55727
rect 289111 55609 289202 55727
rect 288902 55567 289202 55609
rect 288902 55449 288993 55567
rect 289111 55449 289202 55567
rect 288902 37727 289202 55449
rect 288902 37609 288993 37727
rect 289111 37609 289202 37727
rect 288902 37567 289202 37609
rect 288902 37449 288993 37567
rect 289111 37449 289202 37567
rect 288902 19727 289202 37449
rect 288902 19609 288993 19727
rect 289111 19609 289202 19727
rect 288902 19567 289202 19609
rect 288902 19449 288993 19567
rect 289111 19449 289202 19567
rect 288902 1727 289202 19449
rect 288902 1609 288993 1727
rect 289111 1609 289202 1727
rect 288902 1567 289202 1609
rect 288902 1449 288993 1567
rect 289111 1449 289202 1567
rect 288902 -173 289202 1449
rect 288902 -291 288993 -173
rect 289111 -291 289202 -173
rect 288902 -333 289202 -291
rect 288902 -451 288993 -333
rect 289111 -451 289202 -333
rect 288902 -932 289202 -451
rect 290702 345527 291002 353081
rect 293600 353359 293900 353370
rect 293600 353241 293691 353359
rect 293809 353241 293900 353359
rect 293600 353199 293900 353241
rect 293600 353081 293691 353199
rect 293809 353081 293900 353199
rect 293130 352889 293430 352900
rect 293130 352771 293221 352889
rect 293339 352771 293430 352889
rect 293130 352729 293430 352771
rect 293130 352611 293221 352729
rect 293339 352611 293430 352729
rect 290702 345409 290793 345527
rect 290911 345409 291002 345527
rect 290702 345367 291002 345409
rect 290702 345249 290793 345367
rect 290911 345249 291002 345367
rect 290702 327527 291002 345249
rect 290702 327409 290793 327527
rect 290911 327409 291002 327527
rect 290702 327367 291002 327409
rect 290702 327249 290793 327367
rect 290911 327249 291002 327367
rect 290702 309527 291002 327249
rect 290702 309409 290793 309527
rect 290911 309409 291002 309527
rect 290702 309367 291002 309409
rect 290702 309249 290793 309367
rect 290911 309249 291002 309367
rect 290702 291527 291002 309249
rect 290702 291409 290793 291527
rect 290911 291409 291002 291527
rect 290702 291367 291002 291409
rect 290702 291249 290793 291367
rect 290911 291249 291002 291367
rect 290702 273527 291002 291249
rect 290702 273409 290793 273527
rect 290911 273409 291002 273527
rect 290702 273367 291002 273409
rect 290702 273249 290793 273367
rect 290911 273249 291002 273367
rect 290702 255527 291002 273249
rect 290702 255409 290793 255527
rect 290911 255409 291002 255527
rect 290702 255367 291002 255409
rect 290702 255249 290793 255367
rect 290911 255249 291002 255367
rect 290702 237527 291002 255249
rect 290702 237409 290793 237527
rect 290911 237409 291002 237527
rect 290702 237367 291002 237409
rect 290702 237249 290793 237367
rect 290911 237249 291002 237367
rect 290702 219527 291002 237249
rect 290702 219409 290793 219527
rect 290911 219409 291002 219527
rect 290702 219367 291002 219409
rect 290702 219249 290793 219367
rect 290911 219249 291002 219367
rect 290702 201527 291002 219249
rect 290702 201409 290793 201527
rect 290911 201409 291002 201527
rect 290702 201367 291002 201409
rect 290702 201249 290793 201367
rect 290911 201249 291002 201367
rect 290702 183527 291002 201249
rect 290702 183409 290793 183527
rect 290911 183409 291002 183527
rect 290702 183367 291002 183409
rect 290702 183249 290793 183367
rect 290911 183249 291002 183367
rect 290702 165527 291002 183249
rect 290702 165409 290793 165527
rect 290911 165409 291002 165527
rect 290702 165367 291002 165409
rect 290702 165249 290793 165367
rect 290911 165249 291002 165367
rect 290702 147527 291002 165249
rect 290702 147409 290793 147527
rect 290911 147409 291002 147527
rect 290702 147367 291002 147409
rect 290702 147249 290793 147367
rect 290911 147249 291002 147367
rect 290702 129527 291002 147249
rect 290702 129409 290793 129527
rect 290911 129409 291002 129527
rect 290702 129367 291002 129409
rect 290702 129249 290793 129367
rect 290911 129249 291002 129367
rect 290702 111527 291002 129249
rect 290702 111409 290793 111527
rect 290911 111409 291002 111527
rect 290702 111367 291002 111409
rect 290702 111249 290793 111367
rect 290911 111249 291002 111367
rect 290702 93527 291002 111249
rect 290702 93409 290793 93527
rect 290911 93409 291002 93527
rect 290702 93367 291002 93409
rect 290702 93249 290793 93367
rect 290911 93249 291002 93367
rect 290702 75527 291002 93249
rect 290702 75409 290793 75527
rect 290911 75409 291002 75527
rect 290702 75367 291002 75409
rect 290702 75249 290793 75367
rect 290911 75249 291002 75367
rect 290702 57527 291002 75249
rect 290702 57409 290793 57527
rect 290911 57409 291002 57527
rect 290702 57367 291002 57409
rect 290702 57249 290793 57367
rect 290911 57249 291002 57367
rect 290702 39527 291002 57249
rect 290702 39409 290793 39527
rect 290911 39409 291002 39527
rect 290702 39367 291002 39409
rect 290702 39249 290793 39367
rect 290911 39249 291002 39367
rect 290702 21527 291002 39249
rect 290702 21409 290793 21527
rect 290911 21409 291002 21527
rect 290702 21367 291002 21409
rect 290702 21249 290793 21367
rect 290911 21249 291002 21367
rect 290702 3527 291002 21249
rect 290702 3409 290793 3527
rect 290911 3409 291002 3527
rect 290702 3367 291002 3409
rect 290702 3249 290793 3367
rect 290911 3249 291002 3367
rect 290702 -1113 291002 3249
rect 292660 352419 292960 352430
rect 292660 352301 292751 352419
rect 292869 352301 292960 352419
rect 292660 352259 292960 352301
rect 292660 352141 292751 352259
rect 292869 352141 292960 352259
rect 292660 343727 292960 352141
rect 292660 343609 292751 343727
rect 292869 343609 292960 343727
rect 292660 343567 292960 343609
rect 292660 343449 292751 343567
rect 292869 343449 292960 343567
rect 292660 325727 292960 343449
rect 292660 325609 292751 325727
rect 292869 325609 292960 325727
rect 292660 325567 292960 325609
rect 292660 325449 292751 325567
rect 292869 325449 292960 325567
rect 292660 307727 292960 325449
rect 292660 307609 292751 307727
rect 292869 307609 292960 307727
rect 292660 307567 292960 307609
rect 292660 307449 292751 307567
rect 292869 307449 292960 307567
rect 292660 289727 292960 307449
rect 292660 289609 292751 289727
rect 292869 289609 292960 289727
rect 292660 289567 292960 289609
rect 292660 289449 292751 289567
rect 292869 289449 292960 289567
rect 292660 271727 292960 289449
rect 292660 271609 292751 271727
rect 292869 271609 292960 271727
rect 292660 271567 292960 271609
rect 292660 271449 292751 271567
rect 292869 271449 292960 271567
rect 292660 253727 292960 271449
rect 292660 253609 292751 253727
rect 292869 253609 292960 253727
rect 292660 253567 292960 253609
rect 292660 253449 292751 253567
rect 292869 253449 292960 253567
rect 292660 235727 292960 253449
rect 292660 235609 292751 235727
rect 292869 235609 292960 235727
rect 292660 235567 292960 235609
rect 292660 235449 292751 235567
rect 292869 235449 292960 235567
rect 292660 217727 292960 235449
rect 292660 217609 292751 217727
rect 292869 217609 292960 217727
rect 292660 217567 292960 217609
rect 292660 217449 292751 217567
rect 292869 217449 292960 217567
rect 292660 199727 292960 217449
rect 292660 199609 292751 199727
rect 292869 199609 292960 199727
rect 292660 199567 292960 199609
rect 292660 199449 292751 199567
rect 292869 199449 292960 199567
rect 292660 181727 292960 199449
rect 292660 181609 292751 181727
rect 292869 181609 292960 181727
rect 292660 181567 292960 181609
rect 292660 181449 292751 181567
rect 292869 181449 292960 181567
rect 292660 163727 292960 181449
rect 292660 163609 292751 163727
rect 292869 163609 292960 163727
rect 292660 163567 292960 163609
rect 292660 163449 292751 163567
rect 292869 163449 292960 163567
rect 292660 145727 292960 163449
rect 292660 145609 292751 145727
rect 292869 145609 292960 145727
rect 292660 145567 292960 145609
rect 292660 145449 292751 145567
rect 292869 145449 292960 145567
rect 292660 127727 292960 145449
rect 292660 127609 292751 127727
rect 292869 127609 292960 127727
rect 292660 127567 292960 127609
rect 292660 127449 292751 127567
rect 292869 127449 292960 127567
rect 292660 109727 292960 127449
rect 292660 109609 292751 109727
rect 292869 109609 292960 109727
rect 292660 109567 292960 109609
rect 292660 109449 292751 109567
rect 292869 109449 292960 109567
rect 292660 91727 292960 109449
rect 292660 91609 292751 91727
rect 292869 91609 292960 91727
rect 292660 91567 292960 91609
rect 292660 91449 292751 91567
rect 292869 91449 292960 91567
rect 292660 73727 292960 91449
rect 292660 73609 292751 73727
rect 292869 73609 292960 73727
rect 292660 73567 292960 73609
rect 292660 73449 292751 73567
rect 292869 73449 292960 73567
rect 292660 55727 292960 73449
rect 292660 55609 292751 55727
rect 292869 55609 292960 55727
rect 292660 55567 292960 55609
rect 292660 55449 292751 55567
rect 292869 55449 292960 55567
rect 292660 37727 292960 55449
rect 292660 37609 292751 37727
rect 292869 37609 292960 37727
rect 292660 37567 292960 37609
rect 292660 37449 292751 37567
rect 292869 37449 292960 37567
rect 292660 19727 292960 37449
rect 292660 19609 292751 19727
rect 292869 19609 292960 19727
rect 292660 19567 292960 19609
rect 292660 19449 292751 19567
rect 292869 19449 292960 19567
rect 292660 1727 292960 19449
rect 292660 1609 292751 1727
rect 292869 1609 292960 1727
rect 292660 1567 292960 1609
rect 292660 1449 292751 1567
rect 292869 1449 292960 1567
rect 292660 -173 292960 1449
rect 292660 -291 292751 -173
rect 292869 -291 292960 -173
rect 292660 -333 292960 -291
rect 292660 -451 292751 -333
rect 292869 -451 292960 -333
rect 292660 -462 292960 -451
rect 293130 334727 293430 352611
rect 293130 334609 293221 334727
rect 293339 334609 293430 334727
rect 293130 334567 293430 334609
rect 293130 334449 293221 334567
rect 293339 334449 293430 334567
rect 293130 316727 293430 334449
rect 293130 316609 293221 316727
rect 293339 316609 293430 316727
rect 293130 316567 293430 316609
rect 293130 316449 293221 316567
rect 293339 316449 293430 316567
rect 293130 298727 293430 316449
rect 293130 298609 293221 298727
rect 293339 298609 293430 298727
rect 293130 298567 293430 298609
rect 293130 298449 293221 298567
rect 293339 298449 293430 298567
rect 293130 280727 293430 298449
rect 293130 280609 293221 280727
rect 293339 280609 293430 280727
rect 293130 280567 293430 280609
rect 293130 280449 293221 280567
rect 293339 280449 293430 280567
rect 293130 262727 293430 280449
rect 293130 262609 293221 262727
rect 293339 262609 293430 262727
rect 293130 262567 293430 262609
rect 293130 262449 293221 262567
rect 293339 262449 293430 262567
rect 293130 244727 293430 262449
rect 293130 244609 293221 244727
rect 293339 244609 293430 244727
rect 293130 244567 293430 244609
rect 293130 244449 293221 244567
rect 293339 244449 293430 244567
rect 293130 226727 293430 244449
rect 293130 226609 293221 226727
rect 293339 226609 293430 226727
rect 293130 226567 293430 226609
rect 293130 226449 293221 226567
rect 293339 226449 293430 226567
rect 293130 208727 293430 226449
rect 293130 208609 293221 208727
rect 293339 208609 293430 208727
rect 293130 208567 293430 208609
rect 293130 208449 293221 208567
rect 293339 208449 293430 208567
rect 293130 190727 293430 208449
rect 293130 190609 293221 190727
rect 293339 190609 293430 190727
rect 293130 190567 293430 190609
rect 293130 190449 293221 190567
rect 293339 190449 293430 190567
rect 293130 172727 293430 190449
rect 293130 172609 293221 172727
rect 293339 172609 293430 172727
rect 293130 172567 293430 172609
rect 293130 172449 293221 172567
rect 293339 172449 293430 172567
rect 293130 154727 293430 172449
rect 293130 154609 293221 154727
rect 293339 154609 293430 154727
rect 293130 154567 293430 154609
rect 293130 154449 293221 154567
rect 293339 154449 293430 154567
rect 293130 136727 293430 154449
rect 293130 136609 293221 136727
rect 293339 136609 293430 136727
rect 293130 136567 293430 136609
rect 293130 136449 293221 136567
rect 293339 136449 293430 136567
rect 293130 118727 293430 136449
rect 293130 118609 293221 118727
rect 293339 118609 293430 118727
rect 293130 118567 293430 118609
rect 293130 118449 293221 118567
rect 293339 118449 293430 118567
rect 293130 100727 293430 118449
rect 293130 100609 293221 100727
rect 293339 100609 293430 100727
rect 293130 100567 293430 100609
rect 293130 100449 293221 100567
rect 293339 100449 293430 100567
rect 293130 82727 293430 100449
rect 293130 82609 293221 82727
rect 293339 82609 293430 82727
rect 293130 82567 293430 82609
rect 293130 82449 293221 82567
rect 293339 82449 293430 82567
rect 293130 64727 293430 82449
rect 293130 64609 293221 64727
rect 293339 64609 293430 64727
rect 293130 64567 293430 64609
rect 293130 64449 293221 64567
rect 293339 64449 293430 64567
rect 293130 46727 293430 64449
rect 293130 46609 293221 46727
rect 293339 46609 293430 46727
rect 293130 46567 293430 46609
rect 293130 46449 293221 46567
rect 293339 46449 293430 46567
rect 293130 28727 293430 46449
rect 293130 28609 293221 28727
rect 293339 28609 293430 28727
rect 293130 28567 293430 28609
rect 293130 28449 293221 28567
rect 293339 28449 293430 28567
rect 293130 10727 293430 28449
rect 293130 10609 293221 10727
rect 293339 10609 293430 10727
rect 293130 10567 293430 10609
rect 293130 10449 293221 10567
rect 293339 10449 293430 10567
rect 293130 -643 293430 10449
rect 293130 -761 293221 -643
rect 293339 -761 293430 -643
rect 293130 -803 293430 -761
rect 293130 -921 293221 -803
rect 293339 -921 293430 -803
rect 293130 -932 293430 -921
rect 293600 345527 293900 353081
rect 293600 345409 293691 345527
rect 293809 345409 293900 345527
rect 293600 345367 293900 345409
rect 293600 345249 293691 345367
rect 293809 345249 293900 345367
rect 293600 327527 293900 345249
rect 293600 327409 293691 327527
rect 293809 327409 293900 327527
rect 293600 327367 293900 327409
rect 293600 327249 293691 327367
rect 293809 327249 293900 327367
rect 293600 309527 293900 327249
rect 293600 309409 293691 309527
rect 293809 309409 293900 309527
rect 293600 309367 293900 309409
rect 293600 309249 293691 309367
rect 293809 309249 293900 309367
rect 293600 291527 293900 309249
rect 293600 291409 293691 291527
rect 293809 291409 293900 291527
rect 293600 291367 293900 291409
rect 293600 291249 293691 291367
rect 293809 291249 293900 291367
rect 293600 273527 293900 291249
rect 293600 273409 293691 273527
rect 293809 273409 293900 273527
rect 293600 273367 293900 273409
rect 293600 273249 293691 273367
rect 293809 273249 293900 273367
rect 293600 255527 293900 273249
rect 293600 255409 293691 255527
rect 293809 255409 293900 255527
rect 293600 255367 293900 255409
rect 293600 255249 293691 255367
rect 293809 255249 293900 255367
rect 293600 237527 293900 255249
rect 293600 237409 293691 237527
rect 293809 237409 293900 237527
rect 293600 237367 293900 237409
rect 293600 237249 293691 237367
rect 293809 237249 293900 237367
rect 293600 219527 293900 237249
rect 293600 219409 293691 219527
rect 293809 219409 293900 219527
rect 293600 219367 293900 219409
rect 293600 219249 293691 219367
rect 293809 219249 293900 219367
rect 293600 201527 293900 219249
rect 293600 201409 293691 201527
rect 293809 201409 293900 201527
rect 293600 201367 293900 201409
rect 293600 201249 293691 201367
rect 293809 201249 293900 201367
rect 293600 183527 293900 201249
rect 293600 183409 293691 183527
rect 293809 183409 293900 183527
rect 293600 183367 293900 183409
rect 293600 183249 293691 183367
rect 293809 183249 293900 183367
rect 293600 165527 293900 183249
rect 293600 165409 293691 165527
rect 293809 165409 293900 165527
rect 293600 165367 293900 165409
rect 293600 165249 293691 165367
rect 293809 165249 293900 165367
rect 293600 147527 293900 165249
rect 293600 147409 293691 147527
rect 293809 147409 293900 147527
rect 293600 147367 293900 147409
rect 293600 147249 293691 147367
rect 293809 147249 293900 147367
rect 293600 129527 293900 147249
rect 293600 129409 293691 129527
rect 293809 129409 293900 129527
rect 293600 129367 293900 129409
rect 293600 129249 293691 129367
rect 293809 129249 293900 129367
rect 293600 111527 293900 129249
rect 293600 111409 293691 111527
rect 293809 111409 293900 111527
rect 293600 111367 293900 111409
rect 293600 111249 293691 111367
rect 293809 111249 293900 111367
rect 293600 93527 293900 111249
rect 293600 93409 293691 93527
rect 293809 93409 293900 93527
rect 293600 93367 293900 93409
rect 293600 93249 293691 93367
rect 293809 93249 293900 93367
rect 293600 75527 293900 93249
rect 293600 75409 293691 75527
rect 293809 75409 293900 75527
rect 293600 75367 293900 75409
rect 293600 75249 293691 75367
rect 293809 75249 293900 75367
rect 293600 57527 293900 75249
rect 293600 57409 293691 57527
rect 293809 57409 293900 57527
rect 293600 57367 293900 57409
rect 293600 57249 293691 57367
rect 293809 57249 293900 57367
rect 293600 39527 293900 57249
rect 293600 39409 293691 39527
rect 293809 39409 293900 39527
rect 293600 39367 293900 39409
rect 293600 39249 293691 39367
rect 293809 39249 293900 39367
rect 293600 21527 293900 39249
rect 293600 21409 293691 21527
rect 293809 21409 293900 21527
rect 293600 21367 293900 21409
rect 293600 21249 293691 21367
rect 293809 21249 293900 21367
rect 293600 3527 293900 21249
rect 293600 3409 293691 3527
rect 293809 3409 293900 3527
rect 293600 3367 293900 3409
rect 293600 3249 293691 3367
rect 293809 3249 293900 3367
rect 290702 -1231 290793 -1113
rect 290911 -1231 291002 -1113
rect 290702 -1273 291002 -1231
rect 290702 -1391 290793 -1273
rect 290911 -1391 291002 -1273
rect 290702 -1872 291002 -1391
rect 293600 -1113 293900 3249
rect 293600 -1231 293691 -1113
rect 293809 -1231 293900 -1113
rect 293600 -1273 293900 -1231
rect 293600 -1391 293691 -1273
rect 293809 -1391 293900 -1273
rect 293600 -1402 293900 -1391
rect 294070 336527 294370 353551
rect 294070 336409 294161 336527
rect 294279 336409 294370 336527
rect 294070 336367 294370 336409
rect 294070 336249 294161 336367
rect 294279 336249 294370 336367
rect 294070 318527 294370 336249
rect 294070 318409 294161 318527
rect 294279 318409 294370 318527
rect 294070 318367 294370 318409
rect 294070 318249 294161 318367
rect 294279 318249 294370 318367
rect 294070 300527 294370 318249
rect 294070 300409 294161 300527
rect 294279 300409 294370 300527
rect 294070 300367 294370 300409
rect 294070 300249 294161 300367
rect 294279 300249 294370 300367
rect 294070 282527 294370 300249
rect 294070 282409 294161 282527
rect 294279 282409 294370 282527
rect 294070 282367 294370 282409
rect 294070 282249 294161 282367
rect 294279 282249 294370 282367
rect 294070 264527 294370 282249
rect 294070 264409 294161 264527
rect 294279 264409 294370 264527
rect 294070 264367 294370 264409
rect 294070 264249 294161 264367
rect 294279 264249 294370 264367
rect 294070 246527 294370 264249
rect 294070 246409 294161 246527
rect 294279 246409 294370 246527
rect 294070 246367 294370 246409
rect 294070 246249 294161 246367
rect 294279 246249 294370 246367
rect 294070 228527 294370 246249
rect 294070 228409 294161 228527
rect 294279 228409 294370 228527
rect 294070 228367 294370 228409
rect 294070 228249 294161 228367
rect 294279 228249 294370 228367
rect 294070 210527 294370 228249
rect 294070 210409 294161 210527
rect 294279 210409 294370 210527
rect 294070 210367 294370 210409
rect 294070 210249 294161 210367
rect 294279 210249 294370 210367
rect 294070 192527 294370 210249
rect 294070 192409 294161 192527
rect 294279 192409 294370 192527
rect 294070 192367 294370 192409
rect 294070 192249 294161 192367
rect 294279 192249 294370 192367
rect 294070 174527 294370 192249
rect 294070 174409 294161 174527
rect 294279 174409 294370 174527
rect 294070 174367 294370 174409
rect 294070 174249 294161 174367
rect 294279 174249 294370 174367
rect 294070 156527 294370 174249
rect 294070 156409 294161 156527
rect 294279 156409 294370 156527
rect 294070 156367 294370 156409
rect 294070 156249 294161 156367
rect 294279 156249 294370 156367
rect 294070 138527 294370 156249
rect 294070 138409 294161 138527
rect 294279 138409 294370 138527
rect 294070 138367 294370 138409
rect 294070 138249 294161 138367
rect 294279 138249 294370 138367
rect 294070 120527 294370 138249
rect 294070 120409 294161 120527
rect 294279 120409 294370 120527
rect 294070 120367 294370 120409
rect 294070 120249 294161 120367
rect 294279 120249 294370 120367
rect 294070 102527 294370 120249
rect 294070 102409 294161 102527
rect 294279 102409 294370 102527
rect 294070 102367 294370 102409
rect 294070 102249 294161 102367
rect 294279 102249 294370 102367
rect 294070 84527 294370 102249
rect 294070 84409 294161 84527
rect 294279 84409 294370 84527
rect 294070 84367 294370 84409
rect 294070 84249 294161 84367
rect 294279 84249 294370 84367
rect 294070 66527 294370 84249
rect 294070 66409 294161 66527
rect 294279 66409 294370 66527
rect 294070 66367 294370 66409
rect 294070 66249 294161 66367
rect 294279 66249 294370 66367
rect 294070 48527 294370 66249
rect 294070 48409 294161 48527
rect 294279 48409 294370 48527
rect 294070 48367 294370 48409
rect 294070 48249 294161 48367
rect 294279 48249 294370 48367
rect 294070 30527 294370 48249
rect 294070 30409 294161 30527
rect 294279 30409 294370 30527
rect 294070 30367 294370 30409
rect 294070 30249 294161 30367
rect 294279 30249 294370 30367
rect 294070 12527 294370 30249
rect 294070 12409 294161 12527
rect 294279 12409 294370 12527
rect 294070 12367 294370 12409
rect 294070 12249 294161 12367
rect 294279 12249 294370 12367
rect 294070 -1583 294370 12249
rect 294070 -1701 294161 -1583
rect 294279 -1701 294370 -1583
rect 294070 -1743 294370 -1701
rect 294070 -1861 294161 -1743
rect 294279 -1861 294370 -1743
rect 294070 -1872 294370 -1861
rect 294540 347327 294840 354021
rect 294540 347209 294631 347327
rect 294749 347209 294840 347327
rect 294540 347167 294840 347209
rect 294540 347049 294631 347167
rect 294749 347049 294840 347167
rect 294540 329327 294840 347049
rect 294540 329209 294631 329327
rect 294749 329209 294840 329327
rect 294540 329167 294840 329209
rect 294540 329049 294631 329167
rect 294749 329049 294840 329167
rect 294540 311327 294840 329049
rect 294540 311209 294631 311327
rect 294749 311209 294840 311327
rect 294540 311167 294840 311209
rect 294540 311049 294631 311167
rect 294749 311049 294840 311167
rect 294540 293327 294840 311049
rect 294540 293209 294631 293327
rect 294749 293209 294840 293327
rect 294540 293167 294840 293209
rect 294540 293049 294631 293167
rect 294749 293049 294840 293167
rect 294540 275327 294840 293049
rect 294540 275209 294631 275327
rect 294749 275209 294840 275327
rect 294540 275167 294840 275209
rect 294540 275049 294631 275167
rect 294749 275049 294840 275167
rect 294540 257327 294840 275049
rect 294540 257209 294631 257327
rect 294749 257209 294840 257327
rect 294540 257167 294840 257209
rect 294540 257049 294631 257167
rect 294749 257049 294840 257167
rect 294540 239327 294840 257049
rect 294540 239209 294631 239327
rect 294749 239209 294840 239327
rect 294540 239167 294840 239209
rect 294540 239049 294631 239167
rect 294749 239049 294840 239167
rect 294540 221327 294840 239049
rect 294540 221209 294631 221327
rect 294749 221209 294840 221327
rect 294540 221167 294840 221209
rect 294540 221049 294631 221167
rect 294749 221049 294840 221167
rect 294540 203327 294840 221049
rect 294540 203209 294631 203327
rect 294749 203209 294840 203327
rect 294540 203167 294840 203209
rect 294540 203049 294631 203167
rect 294749 203049 294840 203167
rect 294540 185327 294840 203049
rect 294540 185209 294631 185327
rect 294749 185209 294840 185327
rect 294540 185167 294840 185209
rect 294540 185049 294631 185167
rect 294749 185049 294840 185167
rect 294540 167327 294840 185049
rect 294540 167209 294631 167327
rect 294749 167209 294840 167327
rect 294540 167167 294840 167209
rect 294540 167049 294631 167167
rect 294749 167049 294840 167167
rect 294540 149327 294840 167049
rect 294540 149209 294631 149327
rect 294749 149209 294840 149327
rect 294540 149167 294840 149209
rect 294540 149049 294631 149167
rect 294749 149049 294840 149167
rect 294540 131327 294840 149049
rect 294540 131209 294631 131327
rect 294749 131209 294840 131327
rect 294540 131167 294840 131209
rect 294540 131049 294631 131167
rect 294749 131049 294840 131167
rect 294540 113327 294840 131049
rect 294540 113209 294631 113327
rect 294749 113209 294840 113327
rect 294540 113167 294840 113209
rect 294540 113049 294631 113167
rect 294749 113049 294840 113167
rect 294540 95327 294840 113049
rect 294540 95209 294631 95327
rect 294749 95209 294840 95327
rect 294540 95167 294840 95209
rect 294540 95049 294631 95167
rect 294749 95049 294840 95167
rect 294540 77327 294840 95049
rect 294540 77209 294631 77327
rect 294749 77209 294840 77327
rect 294540 77167 294840 77209
rect 294540 77049 294631 77167
rect 294749 77049 294840 77167
rect 294540 59327 294840 77049
rect 294540 59209 294631 59327
rect 294749 59209 294840 59327
rect 294540 59167 294840 59209
rect 294540 59049 294631 59167
rect 294749 59049 294840 59167
rect 294540 41327 294840 59049
rect 294540 41209 294631 41327
rect 294749 41209 294840 41327
rect 294540 41167 294840 41209
rect 294540 41049 294631 41167
rect 294749 41049 294840 41167
rect 294540 23327 294840 41049
rect 294540 23209 294631 23327
rect 294749 23209 294840 23327
rect 294540 23167 294840 23209
rect 294540 23049 294631 23167
rect 294749 23049 294840 23167
rect 294540 5327 294840 23049
rect 294540 5209 294631 5327
rect 294749 5209 294840 5327
rect 294540 5167 294840 5209
rect 294540 5049 294631 5167
rect 294749 5049 294840 5167
rect 294540 -2053 294840 5049
rect 294540 -2171 294631 -2053
rect 294749 -2171 294840 -2053
rect 294540 -2213 294840 -2171
rect 294540 -2331 294631 -2213
rect 294749 -2331 294840 -2213
rect 294540 -2342 294840 -2331
rect 295010 338327 295310 354491
rect 295010 338209 295101 338327
rect 295219 338209 295310 338327
rect 295010 338167 295310 338209
rect 295010 338049 295101 338167
rect 295219 338049 295310 338167
rect 295010 320327 295310 338049
rect 295010 320209 295101 320327
rect 295219 320209 295310 320327
rect 295010 320167 295310 320209
rect 295010 320049 295101 320167
rect 295219 320049 295310 320167
rect 295010 302327 295310 320049
rect 295010 302209 295101 302327
rect 295219 302209 295310 302327
rect 295010 302167 295310 302209
rect 295010 302049 295101 302167
rect 295219 302049 295310 302167
rect 295010 284327 295310 302049
rect 295010 284209 295101 284327
rect 295219 284209 295310 284327
rect 295010 284167 295310 284209
rect 295010 284049 295101 284167
rect 295219 284049 295310 284167
rect 295010 266327 295310 284049
rect 295010 266209 295101 266327
rect 295219 266209 295310 266327
rect 295010 266167 295310 266209
rect 295010 266049 295101 266167
rect 295219 266049 295310 266167
rect 295010 248327 295310 266049
rect 295010 248209 295101 248327
rect 295219 248209 295310 248327
rect 295010 248167 295310 248209
rect 295010 248049 295101 248167
rect 295219 248049 295310 248167
rect 295010 230327 295310 248049
rect 295010 230209 295101 230327
rect 295219 230209 295310 230327
rect 295010 230167 295310 230209
rect 295010 230049 295101 230167
rect 295219 230049 295310 230167
rect 295010 212327 295310 230049
rect 295010 212209 295101 212327
rect 295219 212209 295310 212327
rect 295010 212167 295310 212209
rect 295010 212049 295101 212167
rect 295219 212049 295310 212167
rect 295010 194327 295310 212049
rect 295010 194209 295101 194327
rect 295219 194209 295310 194327
rect 295010 194167 295310 194209
rect 295010 194049 295101 194167
rect 295219 194049 295310 194167
rect 295010 176327 295310 194049
rect 295010 176209 295101 176327
rect 295219 176209 295310 176327
rect 295010 176167 295310 176209
rect 295010 176049 295101 176167
rect 295219 176049 295310 176167
rect 295010 158327 295310 176049
rect 295010 158209 295101 158327
rect 295219 158209 295310 158327
rect 295010 158167 295310 158209
rect 295010 158049 295101 158167
rect 295219 158049 295310 158167
rect 295010 140327 295310 158049
rect 295010 140209 295101 140327
rect 295219 140209 295310 140327
rect 295010 140167 295310 140209
rect 295010 140049 295101 140167
rect 295219 140049 295310 140167
rect 295010 122327 295310 140049
rect 295010 122209 295101 122327
rect 295219 122209 295310 122327
rect 295010 122167 295310 122209
rect 295010 122049 295101 122167
rect 295219 122049 295310 122167
rect 295010 104327 295310 122049
rect 295010 104209 295101 104327
rect 295219 104209 295310 104327
rect 295010 104167 295310 104209
rect 295010 104049 295101 104167
rect 295219 104049 295310 104167
rect 295010 86327 295310 104049
rect 295010 86209 295101 86327
rect 295219 86209 295310 86327
rect 295010 86167 295310 86209
rect 295010 86049 295101 86167
rect 295219 86049 295310 86167
rect 295010 68327 295310 86049
rect 295010 68209 295101 68327
rect 295219 68209 295310 68327
rect 295010 68167 295310 68209
rect 295010 68049 295101 68167
rect 295219 68049 295310 68167
rect 295010 50327 295310 68049
rect 295010 50209 295101 50327
rect 295219 50209 295310 50327
rect 295010 50167 295310 50209
rect 295010 50049 295101 50167
rect 295219 50049 295310 50167
rect 295010 32327 295310 50049
rect 295010 32209 295101 32327
rect 295219 32209 295310 32327
rect 295010 32167 295310 32209
rect 295010 32049 295101 32167
rect 295219 32049 295310 32167
rect 295010 14327 295310 32049
rect 295010 14209 295101 14327
rect 295219 14209 295310 14327
rect 295010 14167 295310 14209
rect 295010 14049 295101 14167
rect 295219 14049 295310 14167
rect 295010 -2523 295310 14049
rect 295010 -2641 295101 -2523
rect 295219 -2641 295310 -2523
rect 295010 -2683 295310 -2641
rect 295010 -2801 295101 -2683
rect 295219 -2801 295310 -2683
rect 295010 -2812 295310 -2801
rect 295480 349127 295780 354961
rect 295480 349009 295571 349127
rect 295689 349009 295780 349127
rect 295480 348967 295780 349009
rect 295480 348849 295571 348967
rect 295689 348849 295780 348967
rect 295480 331127 295780 348849
rect 295480 331009 295571 331127
rect 295689 331009 295780 331127
rect 295480 330967 295780 331009
rect 295480 330849 295571 330967
rect 295689 330849 295780 330967
rect 295480 313127 295780 330849
rect 295480 313009 295571 313127
rect 295689 313009 295780 313127
rect 295480 312967 295780 313009
rect 295480 312849 295571 312967
rect 295689 312849 295780 312967
rect 295480 295127 295780 312849
rect 295480 295009 295571 295127
rect 295689 295009 295780 295127
rect 295480 294967 295780 295009
rect 295480 294849 295571 294967
rect 295689 294849 295780 294967
rect 295480 277127 295780 294849
rect 295480 277009 295571 277127
rect 295689 277009 295780 277127
rect 295480 276967 295780 277009
rect 295480 276849 295571 276967
rect 295689 276849 295780 276967
rect 295480 259127 295780 276849
rect 295480 259009 295571 259127
rect 295689 259009 295780 259127
rect 295480 258967 295780 259009
rect 295480 258849 295571 258967
rect 295689 258849 295780 258967
rect 295480 241127 295780 258849
rect 295480 241009 295571 241127
rect 295689 241009 295780 241127
rect 295480 240967 295780 241009
rect 295480 240849 295571 240967
rect 295689 240849 295780 240967
rect 295480 223127 295780 240849
rect 295480 223009 295571 223127
rect 295689 223009 295780 223127
rect 295480 222967 295780 223009
rect 295480 222849 295571 222967
rect 295689 222849 295780 222967
rect 295480 205127 295780 222849
rect 295480 205009 295571 205127
rect 295689 205009 295780 205127
rect 295480 204967 295780 205009
rect 295480 204849 295571 204967
rect 295689 204849 295780 204967
rect 295480 187127 295780 204849
rect 295480 187009 295571 187127
rect 295689 187009 295780 187127
rect 295480 186967 295780 187009
rect 295480 186849 295571 186967
rect 295689 186849 295780 186967
rect 295480 169127 295780 186849
rect 295480 169009 295571 169127
rect 295689 169009 295780 169127
rect 295480 168967 295780 169009
rect 295480 168849 295571 168967
rect 295689 168849 295780 168967
rect 295480 151127 295780 168849
rect 295480 151009 295571 151127
rect 295689 151009 295780 151127
rect 295480 150967 295780 151009
rect 295480 150849 295571 150967
rect 295689 150849 295780 150967
rect 295480 133127 295780 150849
rect 295480 133009 295571 133127
rect 295689 133009 295780 133127
rect 295480 132967 295780 133009
rect 295480 132849 295571 132967
rect 295689 132849 295780 132967
rect 295480 115127 295780 132849
rect 295480 115009 295571 115127
rect 295689 115009 295780 115127
rect 295480 114967 295780 115009
rect 295480 114849 295571 114967
rect 295689 114849 295780 114967
rect 295480 97127 295780 114849
rect 295480 97009 295571 97127
rect 295689 97009 295780 97127
rect 295480 96967 295780 97009
rect 295480 96849 295571 96967
rect 295689 96849 295780 96967
rect 295480 79127 295780 96849
rect 295480 79009 295571 79127
rect 295689 79009 295780 79127
rect 295480 78967 295780 79009
rect 295480 78849 295571 78967
rect 295689 78849 295780 78967
rect 295480 61127 295780 78849
rect 295480 61009 295571 61127
rect 295689 61009 295780 61127
rect 295480 60967 295780 61009
rect 295480 60849 295571 60967
rect 295689 60849 295780 60967
rect 295480 43127 295780 60849
rect 295480 43009 295571 43127
rect 295689 43009 295780 43127
rect 295480 42967 295780 43009
rect 295480 42849 295571 42967
rect 295689 42849 295780 42967
rect 295480 25127 295780 42849
rect 295480 25009 295571 25127
rect 295689 25009 295780 25127
rect 295480 24967 295780 25009
rect 295480 24849 295571 24967
rect 295689 24849 295780 24967
rect 295480 7127 295780 24849
rect 295480 7009 295571 7127
rect 295689 7009 295780 7127
rect 295480 6967 295780 7009
rect 295480 6849 295571 6967
rect 295689 6849 295780 6967
rect 295480 -2993 295780 6849
rect 295480 -3111 295571 -2993
rect 295689 -3111 295780 -2993
rect 295480 -3153 295780 -3111
rect 295480 -3271 295571 -3153
rect 295689 -3271 295780 -3153
rect 295480 -3282 295780 -3271
rect 295950 340127 296250 355431
rect 295950 340009 296041 340127
rect 296159 340009 296250 340127
rect 295950 339967 296250 340009
rect 295950 339849 296041 339967
rect 296159 339849 296250 339967
rect 295950 322127 296250 339849
rect 295950 322009 296041 322127
rect 296159 322009 296250 322127
rect 295950 321967 296250 322009
rect 295950 321849 296041 321967
rect 296159 321849 296250 321967
rect 295950 304127 296250 321849
rect 295950 304009 296041 304127
rect 296159 304009 296250 304127
rect 295950 303967 296250 304009
rect 295950 303849 296041 303967
rect 296159 303849 296250 303967
rect 295950 286127 296250 303849
rect 295950 286009 296041 286127
rect 296159 286009 296250 286127
rect 295950 285967 296250 286009
rect 295950 285849 296041 285967
rect 296159 285849 296250 285967
rect 295950 268127 296250 285849
rect 295950 268009 296041 268127
rect 296159 268009 296250 268127
rect 295950 267967 296250 268009
rect 295950 267849 296041 267967
rect 296159 267849 296250 267967
rect 295950 250127 296250 267849
rect 295950 250009 296041 250127
rect 296159 250009 296250 250127
rect 295950 249967 296250 250009
rect 295950 249849 296041 249967
rect 296159 249849 296250 249967
rect 295950 232127 296250 249849
rect 295950 232009 296041 232127
rect 296159 232009 296250 232127
rect 295950 231967 296250 232009
rect 295950 231849 296041 231967
rect 296159 231849 296250 231967
rect 295950 214127 296250 231849
rect 295950 214009 296041 214127
rect 296159 214009 296250 214127
rect 295950 213967 296250 214009
rect 295950 213849 296041 213967
rect 296159 213849 296250 213967
rect 295950 196127 296250 213849
rect 295950 196009 296041 196127
rect 296159 196009 296250 196127
rect 295950 195967 296250 196009
rect 295950 195849 296041 195967
rect 296159 195849 296250 195967
rect 295950 178127 296250 195849
rect 295950 178009 296041 178127
rect 296159 178009 296250 178127
rect 295950 177967 296250 178009
rect 295950 177849 296041 177967
rect 296159 177849 296250 177967
rect 295950 160127 296250 177849
rect 295950 160009 296041 160127
rect 296159 160009 296250 160127
rect 295950 159967 296250 160009
rect 295950 159849 296041 159967
rect 296159 159849 296250 159967
rect 295950 142127 296250 159849
rect 295950 142009 296041 142127
rect 296159 142009 296250 142127
rect 295950 141967 296250 142009
rect 295950 141849 296041 141967
rect 296159 141849 296250 141967
rect 295950 124127 296250 141849
rect 295950 124009 296041 124127
rect 296159 124009 296250 124127
rect 295950 123967 296250 124009
rect 295950 123849 296041 123967
rect 296159 123849 296250 123967
rect 295950 106127 296250 123849
rect 295950 106009 296041 106127
rect 296159 106009 296250 106127
rect 295950 105967 296250 106009
rect 295950 105849 296041 105967
rect 296159 105849 296250 105967
rect 295950 88127 296250 105849
rect 295950 88009 296041 88127
rect 296159 88009 296250 88127
rect 295950 87967 296250 88009
rect 295950 87849 296041 87967
rect 296159 87849 296250 87967
rect 295950 70127 296250 87849
rect 295950 70009 296041 70127
rect 296159 70009 296250 70127
rect 295950 69967 296250 70009
rect 295950 69849 296041 69967
rect 296159 69849 296250 69967
rect 295950 52127 296250 69849
rect 295950 52009 296041 52127
rect 296159 52009 296250 52127
rect 295950 51967 296250 52009
rect 295950 51849 296041 51967
rect 296159 51849 296250 51967
rect 295950 34127 296250 51849
rect 295950 34009 296041 34127
rect 296159 34009 296250 34127
rect 295950 33967 296250 34009
rect 295950 33849 296041 33967
rect 296159 33849 296250 33967
rect 295950 16127 296250 33849
rect 295950 16009 296041 16127
rect 296159 16009 296250 16127
rect 295950 15967 296250 16009
rect 295950 15849 296041 15967
rect 296159 15849 296250 15967
rect 285302 -3581 285393 -3463
rect 285511 -3581 285602 -3463
rect 285302 -3623 285602 -3581
rect 285302 -3741 285393 -3623
rect 285511 -3741 285602 -3623
rect 285302 -3752 285602 -3741
rect 295950 -3463 296250 15849
rect 295950 -3581 296041 -3463
rect 296159 -3581 296250 -3463
rect 295950 -3623 296250 -3581
rect 295950 -3741 296041 -3623
rect 296159 -3741 296250 -3623
rect 295950 -3752 296250 -3741
<< via4 >>
rect -4197 355591 -4079 355709
rect -4197 355431 -4079 355549
rect -4197 340009 -4079 340127
rect -4197 339849 -4079 339967
rect -4197 322009 -4079 322127
rect -4197 321849 -4079 321967
rect -4197 304009 -4079 304127
rect -4197 303849 -4079 303967
rect -4197 286009 -4079 286127
rect -4197 285849 -4079 285967
rect -4197 268009 -4079 268127
rect -4197 267849 -4079 267967
rect -4197 250009 -4079 250127
rect -4197 249849 -4079 249967
rect -4197 232009 -4079 232127
rect -4197 231849 -4079 231967
rect -4197 214009 -4079 214127
rect -4197 213849 -4079 213967
rect -4197 196009 -4079 196127
rect -4197 195849 -4079 195967
rect -4197 178009 -4079 178127
rect -4197 177849 -4079 177967
rect -4197 160009 -4079 160127
rect -4197 159849 -4079 159967
rect -4197 142009 -4079 142127
rect -4197 141849 -4079 141967
rect -4197 124009 -4079 124127
rect -4197 123849 -4079 123967
rect -4197 106009 -4079 106127
rect -4197 105849 -4079 105967
rect -4197 88009 -4079 88127
rect -4197 87849 -4079 87967
rect -4197 70009 -4079 70127
rect -4197 69849 -4079 69967
rect -4197 52009 -4079 52127
rect -4197 51849 -4079 51967
rect -4197 34009 -4079 34127
rect -4197 33849 -4079 33967
rect -4197 16009 -4079 16127
rect -4197 15849 -4079 15967
rect -3727 355121 -3609 355239
rect -3727 354961 -3609 355079
rect 6393 355121 6511 355239
rect 6393 354961 6511 355079
rect -3727 349009 -3609 349127
rect -3727 348849 -3609 348967
rect -3727 331009 -3609 331127
rect -3727 330849 -3609 330967
rect -3727 313009 -3609 313127
rect -3727 312849 -3609 312967
rect -3727 295009 -3609 295127
rect -3727 294849 -3609 294967
rect -3727 277009 -3609 277127
rect -3727 276849 -3609 276967
rect -3727 259009 -3609 259127
rect -3727 258849 -3609 258967
rect -3727 241009 -3609 241127
rect -3727 240849 -3609 240967
rect -3727 223009 -3609 223127
rect -3727 222849 -3609 222967
rect -3727 205009 -3609 205127
rect -3727 204849 -3609 204967
rect -3727 187009 -3609 187127
rect -3727 186849 -3609 186967
rect -3727 169009 -3609 169127
rect -3727 168849 -3609 168967
rect -3727 151009 -3609 151127
rect -3727 150849 -3609 150967
rect -3727 133009 -3609 133127
rect -3727 132849 -3609 132967
rect -3727 115009 -3609 115127
rect -3727 114849 -3609 114967
rect -3727 97009 -3609 97127
rect -3727 96849 -3609 96967
rect -3727 79009 -3609 79127
rect -3727 78849 -3609 78967
rect -3727 61009 -3609 61127
rect -3727 60849 -3609 60967
rect -3727 43009 -3609 43127
rect -3727 42849 -3609 42967
rect -3727 25009 -3609 25127
rect -3727 24849 -3609 24967
rect -3727 7009 -3609 7127
rect -3727 6849 -3609 6967
rect -3257 354651 -3139 354769
rect -3257 354491 -3139 354609
rect -3257 338209 -3139 338327
rect -3257 338049 -3139 338167
rect -3257 320209 -3139 320327
rect -3257 320049 -3139 320167
rect -3257 302209 -3139 302327
rect -3257 302049 -3139 302167
rect -3257 284209 -3139 284327
rect -3257 284049 -3139 284167
rect -3257 266209 -3139 266327
rect -3257 266049 -3139 266167
rect -3257 248209 -3139 248327
rect -3257 248049 -3139 248167
rect -3257 230209 -3139 230327
rect -3257 230049 -3139 230167
rect -3257 212209 -3139 212327
rect -3257 212049 -3139 212167
rect -3257 194209 -3139 194327
rect -3257 194049 -3139 194167
rect -3257 176209 -3139 176327
rect -3257 176049 -3139 176167
rect -3257 158209 -3139 158327
rect -3257 158049 -3139 158167
rect -3257 140209 -3139 140327
rect -3257 140049 -3139 140167
rect -3257 122209 -3139 122327
rect -3257 122049 -3139 122167
rect -3257 104209 -3139 104327
rect -3257 104049 -3139 104167
rect -3257 86209 -3139 86327
rect -3257 86049 -3139 86167
rect -3257 68209 -3139 68327
rect -3257 68049 -3139 68167
rect -3257 50209 -3139 50327
rect -3257 50049 -3139 50167
rect -3257 32209 -3139 32327
rect -3257 32049 -3139 32167
rect -3257 14209 -3139 14327
rect -3257 14049 -3139 14167
rect -2787 354181 -2669 354299
rect -2787 354021 -2669 354139
rect 4593 354181 4711 354299
rect 4593 354021 4711 354139
rect -2787 347209 -2669 347327
rect -2787 347049 -2669 347167
rect -2787 329209 -2669 329327
rect -2787 329049 -2669 329167
rect -2787 311209 -2669 311327
rect -2787 311049 -2669 311167
rect -2787 293209 -2669 293327
rect -2787 293049 -2669 293167
rect -2787 275209 -2669 275327
rect -2787 275049 -2669 275167
rect -2787 257209 -2669 257327
rect -2787 257049 -2669 257167
rect -2787 239209 -2669 239327
rect -2787 239049 -2669 239167
rect -2787 221209 -2669 221327
rect -2787 221049 -2669 221167
rect -2787 203209 -2669 203327
rect -2787 203049 -2669 203167
rect -2787 185209 -2669 185327
rect -2787 185049 -2669 185167
rect -2787 167209 -2669 167327
rect -2787 167049 -2669 167167
rect -2787 149209 -2669 149327
rect -2787 149049 -2669 149167
rect -2787 131209 -2669 131327
rect -2787 131049 -2669 131167
rect -2787 113209 -2669 113327
rect -2787 113049 -2669 113167
rect -2787 95209 -2669 95327
rect -2787 95049 -2669 95167
rect -2787 77209 -2669 77327
rect -2787 77049 -2669 77167
rect -2787 59209 -2669 59327
rect -2787 59049 -2669 59167
rect -2787 41209 -2669 41327
rect -2787 41049 -2669 41167
rect -2787 23209 -2669 23327
rect -2787 23049 -2669 23167
rect -2787 5209 -2669 5327
rect -2787 5049 -2669 5167
rect -2317 353711 -2199 353829
rect -2317 353551 -2199 353669
rect -2317 336409 -2199 336527
rect -2317 336249 -2199 336367
rect -2317 318409 -2199 318527
rect -2317 318249 -2199 318367
rect -2317 300409 -2199 300527
rect -2317 300249 -2199 300367
rect -2317 282409 -2199 282527
rect -2317 282249 -2199 282367
rect -2317 264409 -2199 264527
rect -2317 264249 -2199 264367
rect -2317 246409 -2199 246527
rect -2317 246249 -2199 246367
rect -2317 228409 -2199 228527
rect -2317 228249 -2199 228367
rect -2317 210409 -2199 210527
rect -2317 210249 -2199 210367
rect -2317 192409 -2199 192527
rect -2317 192249 -2199 192367
rect -2317 174409 -2199 174527
rect -2317 174249 -2199 174367
rect -2317 156409 -2199 156527
rect -2317 156249 -2199 156367
rect -2317 138409 -2199 138527
rect -2317 138249 -2199 138367
rect -2317 120409 -2199 120527
rect -2317 120249 -2199 120367
rect -2317 102409 -2199 102527
rect -2317 102249 -2199 102367
rect -2317 84409 -2199 84527
rect -2317 84249 -2199 84367
rect -2317 66409 -2199 66527
rect -2317 66249 -2199 66367
rect -2317 48409 -2199 48527
rect -2317 48249 -2199 48367
rect -2317 30409 -2199 30527
rect -2317 30249 -2199 30367
rect -2317 12409 -2199 12527
rect -2317 12249 -2199 12367
rect -1847 353241 -1729 353359
rect -1847 353081 -1729 353199
rect 2793 353241 2911 353359
rect 2793 353081 2911 353199
rect -1847 345409 -1729 345527
rect -1847 345249 -1729 345367
rect -1847 327409 -1729 327527
rect -1847 327249 -1729 327367
rect -1847 309409 -1729 309527
rect -1847 309249 -1729 309367
rect -1847 291409 -1729 291527
rect -1847 291249 -1729 291367
rect -1847 273409 -1729 273527
rect -1847 273249 -1729 273367
rect -1847 255409 -1729 255527
rect -1847 255249 -1729 255367
rect -1847 237409 -1729 237527
rect -1847 237249 -1729 237367
rect -1847 219409 -1729 219527
rect -1847 219249 -1729 219367
rect -1847 201409 -1729 201527
rect -1847 201249 -1729 201367
rect -1847 183409 -1729 183527
rect -1847 183249 -1729 183367
rect -1847 165409 -1729 165527
rect -1847 165249 -1729 165367
rect -1847 147409 -1729 147527
rect -1847 147249 -1729 147367
rect -1847 129409 -1729 129527
rect -1847 129249 -1729 129367
rect -1847 111409 -1729 111527
rect -1847 111249 -1729 111367
rect -1847 93409 -1729 93527
rect -1847 93249 -1729 93367
rect -1847 75409 -1729 75527
rect -1847 75249 -1729 75367
rect -1847 57409 -1729 57527
rect -1847 57249 -1729 57367
rect -1847 39409 -1729 39527
rect -1847 39249 -1729 39367
rect -1847 21409 -1729 21527
rect -1847 21249 -1729 21367
rect -1847 3409 -1729 3527
rect -1847 3249 -1729 3367
rect -1377 352771 -1259 352889
rect -1377 352611 -1259 352729
rect -1377 334609 -1259 334727
rect -1377 334449 -1259 334567
rect -1377 316609 -1259 316727
rect -1377 316449 -1259 316567
rect -1377 298609 -1259 298727
rect -1377 298449 -1259 298567
rect -1377 280609 -1259 280727
rect -1377 280449 -1259 280567
rect -1377 262609 -1259 262727
rect -1377 262449 -1259 262567
rect -1377 244609 -1259 244727
rect -1377 244449 -1259 244567
rect -1377 226609 -1259 226727
rect -1377 226449 -1259 226567
rect -1377 208609 -1259 208727
rect -1377 208449 -1259 208567
rect -1377 190609 -1259 190727
rect -1377 190449 -1259 190567
rect -1377 172609 -1259 172727
rect -1377 172449 -1259 172567
rect -1377 154609 -1259 154727
rect -1377 154449 -1259 154567
rect -1377 136609 -1259 136727
rect -1377 136449 -1259 136567
rect -1377 118609 -1259 118727
rect -1377 118449 -1259 118567
rect -1377 100609 -1259 100727
rect -1377 100449 -1259 100567
rect -1377 82609 -1259 82727
rect -1377 82449 -1259 82567
rect -1377 64609 -1259 64727
rect -1377 64449 -1259 64567
rect -1377 46609 -1259 46727
rect -1377 46449 -1259 46567
rect -1377 28609 -1259 28727
rect -1377 28449 -1259 28567
rect -1377 10609 -1259 10727
rect -1377 10449 -1259 10567
rect -907 352301 -789 352419
rect -907 352141 -789 352259
rect -907 343609 -789 343727
rect -907 343449 -789 343567
rect -907 325609 -789 325727
rect -907 325449 -789 325567
rect -907 307609 -789 307727
rect -907 307449 -789 307567
rect -907 289609 -789 289727
rect -907 289449 -789 289567
rect -907 271609 -789 271727
rect -907 271449 -789 271567
rect -907 253609 -789 253727
rect -907 253449 -789 253567
rect -907 235609 -789 235727
rect -907 235449 -789 235567
rect -907 217609 -789 217727
rect -907 217449 -789 217567
rect -907 199609 -789 199727
rect -907 199449 -789 199567
rect -907 181609 -789 181727
rect -907 181449 -789 181567
rect -907 163609 -789 163727
rect -907 163449 -789 163567
rect -907 145609 -789 145727
rect -907 145449 -789 145567
rect -907 127609 -789 127727
rect -907 127449 -789 127567
rect -907 109609 -789 109727
rect -907 109449 -789 109567
rect -907 91609 -789 91727
rect -907 91449 -789 91567
rect -907 73609 -789 73727
rect -907 73449 -789 73567
rect -907 55609 -789 55727
rect -907 55449 -789 55567
rect -907 37609 -789 37727
rect -907 37449 -789 37567
rect -907 19609 -789 19727
rect -907 19449 -789 19567
rect -907 1609 -789 1727
rect -907 1449 -789 1567
rect -907 -291 -789 -173
rect -907 -451 -789 -333
rect 993 352301 1111 352419
rect 993 352141 1111 352259
rect 993 343609 1111 343727
rect 993 343449 1111 343567
rect 993 325609 1111 325727
rect 993 325449 1111 325567
rect 993 307609 1111 307727
rect 993 307449 1111 307567
rect 993 289609 1111 289727
rect 993 289449 1111 289567
rect 993 271609 1111 271727
rect 993 271449 1111 271567
rect 993 253609 1111 253727
rect 993 253449 1111 253567
rect 993 235609 1111 235727
rect 993 235449 1111 235567
rect 993 217609 1111 217727
rect 993 217449 1111 217567
rect 993 199609 1111 199727
rect 993 199449 1111 199567
rect 993 181609 1111 181727
rect 993 181449 1111 181567
rect 993 163609 1111 163727
rect 993 163449 1111 163567
rect 993 145609 1111 145727
rect 993 145449 1111 145567
rect 993 127609 1111 127727
rect 993 127449 1111 127567
rect 993 109609 1111 109727
rect 993 109449 1111 109567
rect 993 91609 1111 91727
rect 993 91449 1111 91567
rect 993 73609 1111 73727
rect 993 73449 1111 73567
rect 993 55609 1111 55727
rect 993 55449 1111 55567
rect 993 37609 1111 37727
rect 993 37449 1111 37567
rect 993 19609 1111 19727
rect 993 19449 1111 19567
rect 993 1609 1111 1727
rect 993 1449 1111 1567
rect 993 -291 1111 -173
rect 993 -451 1111 -333
rect -1377 -761 -1259 -643
rect -1377 -921 -1259 -803
rect 2793 345409 2911 345527
rect 2793 345249 2911 345367
rect 2793 327409 2911 327527
rect 2793 327249 2911 327367
rect 2793 309409 2911 309527
rect 2793 309249 2911 309367
rect 2793 291409 2911 291527
rect 2793 291249 2911 291367
rect 2793 273409 2911 273527
rect 2793 273249 2911 273367
rect 2793 255409 2911 255527
rect 2793 255249 2911 255367
rect 2793 237409 2911 237527
rect 2793 237249 2911 237367
rect 2793 219409 2911 219527
rect 2793 219249 2911 219367
rect 2793 201409 2911 201527
rect 2793 201249 2911 201367
rect 2793 183409 2911 183527
rect 2793 183249 2911 183367
rect 2793 165409 2911 165527
rect 2793 165249 2911 165367
rect 2793 147409 2911 147527
rect 2793 147249 2911 147367
rect 2793 129409 2911 129527
rect 2793 129249 2911 129367
rect 2793 111409 2911 111527
rect 2793 111249 2911 111367
rect 2793 93409 2911 93527
rect 2793 93249 2911 93367
rect 2793 75409 2911 75527
rect 2793 75249 2911 75367
rect 2793 57409 2911 57527
rect 2793 57249 2911 57367
rect 2793 39409 2911 39527
rect 2793 39249 2911 39367
rect 2793 21409 2911 21527
rect 2793 21249 2911 21367
rect 2793 3409 2911 3527
rect 2793 3249 2911 3367
rect -1847 -1231 -1729 -1113
rect -1847 -1391 -1729 -1273
rect 2793 -1231 2911 -1113
rect 2793 -1391 2911 -1273
rect -2317 -1701 -2199 -1583
rect -2317 -1861 -2199 -1743
rect 4593 347209 4711 347327
rect 4593 347049 4711 347167
rect 4593 329209 4711 329327
rect 4593 329049 4711 329167
rect 4593 311209 4711 311327
rect 4593 311049 4711 311167
rect 4593 293209 4711 293327
rect 4593 293049 4711 293167
rect 4593 275209 4711 275327
rect 4593 275049 4711 275167
rect 4593 257209 4711 257327
rect 4593 257049 4711 257167
rect 4593 239209 4711 239327
rect 4593 239049 4711 239167
rect 4593 221209 4711 221327
rect 4593 221049 4711 221167
rect 4593 203209 4711 203327
rect 4593 203049 4711 203167
rect 4593 185209 4711 185327
rect 4593 185049 4711 185167
rect 4593 167209 4711 167327
rect 4593 167049 4711 167167
rect 4593 149209 4711 149327
rect 4593 149049 4711 149167
rect 4593 131209 4711 131327
rect 4593 131049 4711 131167
rect 4593 113209 4711 113327
rect 4593 113049 4711 113167
rect 4593 95209 4711 95327
rect 4593 95049 4711 95167
rect 4593 77209 4711 77327
rect 4593 77049 4711 77167
rect 4593 59209 4711 59327
rect 4593 59049 4711 59167
rect 4593 41209 4711 41327
rect 4593 41049 4711 41167
rect 4593 23209 4711 23327
rect 4593 23049 4711 23167
rect 4593 5209 4711 5327
rect 4593 5049 4711 5167
rect -2787 -2171 -2669 -2053
rect -2787 -2331 -2669 -2213
rect 4593 -2171 4711 -2053
rect 4593 -2331 4711 -2213
rect -3257 -2641 -3139 -2523
rect -3257 -2801 -3139 -2683
rect 15393 355591 15511 355709
rect 15393 355431 15511 355549
rect 13593 354651 13711 354769
rect 13593 354491 13711 354609
rect 11793 353711 11911 353829
rect 11793 353551 11911 353669
rect 6393 349009 6511 349127
rect 6393 348849 6511 348967
rect 6393 331009 6511 331127
rect 6393 330849 6511 330967
rect 6393 313009 6511 313127
rect 6393 312849 6511 312967
rect 6393 295009 6511 295127
rect 6393 294849 6511 294967
rect 6393 277009 6511 277127
rect 6393 276849 6511 276967
rect 6393 259009 6511 259127
rect 6393 258849 6511 258967
rect 6393 241009 6511 241127
rect 6393 240849 6511 240967
rect 6393 223009 6511 223127
rect 6393 222849 6511 222967
rect 6393 205009 6511 205127
rect 6393 204849 6511 204967
rect 6393 187009 6511 187127
rect 6393 186849 6511 186967
rect 6393 169009 6511 169127
rect 6393 168849 6511 168967
rect 6393 151009 6511 151127
rect 6393 150849 6511 150967
rect 6393 133009 6511 133127
rect 6393 132849 6511 132967
rect 6393 115009 6511 115127
rect 6393 114849 6511 114967
rect 6393 97009 6511 97127
rect 6393 96849 6511 96967
rect 6393 79009 6511 79127
rect 6393 78849 6511 78967
rect 6393 61009 6511 61127
rect 6393 60849 6511 60967
rect 6393 43009 6511 43127
rect 6393 42849 6511 42967
rect 6393 25009 6511 25127
rect 6393 24849 6511 24967
rect 6393 7009 6511 7127
rect 6393 6849 6511 6967
rect -3727 -3111 -3609 -2993
rect -3727 -3271 -3609 -3153
rect 9993 352771 10111 352889
rect 9993 352611 10111 352729
rect 9993 334609 10111 334727
rect 9993 334449 10111 334567
rect 9993 316609 10111 316727
rect 9993 316449 10111 316567
rect 9993 298609 10111 298727
rect 9993 298449 10111 298567
rect 9993 280609 10111 280727
rect 9993 280449 10111 280567
rect 9993 262609 10111 262727
rect 9993 262449 10111 262567
rect 9993 244609 10111 244727
rect 9993 244449 10111 244567
rect 9993 226609 10111 226727
rect 9993 226449 10111 226567
rect 9993 208609 10111 208727
rect 9993 208449 10111 208567
rect 9993 190609 10111 190727
rect 9993 190449 10111 190567
rect 9993 172609 10111 172727
rect 9993 172449 10111 172567
rect 9993 154609 10111 154727
rect 9993 154449 10111 154567
rect 9993 136609 10111 136727
rect 9993 136449 10111 136567
rect 9993 118609 10111 118727
rect 9993 118449 10111 118567
rect 9993 100609 10111 100727
rect 9993 100449 10111 100567
rect 9993 82609 10111 82727
rect 9993 82449 10111 82567
rect 9993 64609 10111 64727
rect 9993 64449 10111 64567
rect 9993 46609 10111 46727
rect 9993 46449 10111 46567
rect 9993 28609 10111 28727
rect 9993 28449 10111 28567
rect 9993 10609 10111 10727
rect 9993 10449 10111 10567
rect 9993 -761 10111 -643
rect 9993 -921 10111 -803
rect 11793 336409 11911 336527
rect 11793 336249 11911 336367
rect 11793 318409 11911 318527
rect 11793 318249 11911 318367
rect 11793 300409 11911 300527
rect 11793 300249 11911 300367
rect 11793 282409 11911 282527
rect 11793 282249 11911 282367
rect 11793 264409 11911 264527
rect 11793 264249 11911 264367
rect 11793 246409 11911 246527
rect 11793 246249 11911 246367
rect 11793 228409 11911 228527
rect 11793 228249 11911 228367
rect 11793 210409 11911 210527
rect 11793 210249 11911 210367
rect 11793 192409 11911 192527
rect 11793 192249 11911 192367
rect 11793 174409 11911 174527
rect 11793 174249 11911 174367
rect 11793 156409 11911 156527
rect 11793 156249 11911 156367
rect 11793 138409 11911 138527
rect 11793 138249 11911 138367
rect 11793 120409 11911 120527
rect 11793 120249 11911 120367
rect 11793 102409 11911 102527
rect 11793 102249 11911 102367
rect 11793 84409 11911 84527
rect 11793 84249 11911 84367
rect 11793 66409 11911 66527
rect 11793 66249 11911 66367
rect 11793 48409 11911 48527
rect 11793 48249 11911 48367
rect 11793 30409 11911 30527
rect 11793 30249 11911 30367
rect 11793 12409 11911 12527
rect 11793 12249 11911 12367
rect 11793 -1701 11911 -1583
rect 11793 -1861 11911 -1743
rect 13593 338209 13711 338327
rect 13593 338049 13711 338167
rect 13593 320209 13711 320327
rect 13593 320049 13711 320167
rect 13593 302209 13711 302327
rect 13593 302049 13711 302167
rect 13593 284209 13711 284327
rect 13593 284049 13711 284167
rect 13593 266209 13711 266327
rect 13593 266049 13711 266167
rect 13593 248209 13711 248327
rect 13593 248049 13711 248167
rect 13593 230209 13711 230327
rect 13593 230049 13711 230167
rect 13593 212209 13711 212327
rect 13593 212049 13711 212167
rect 13593 194209 13711 194327
rect 13593 194049 13711 194167
rect 13593 176209 13711 176327
rect 13593 176049 13711 176167
rect 13593 158209 13711 158327
rect 13593 158049 13711 158167
rect 13593 140209 13711 140327
rect 13593 140049 13711 140167
rect 13593 122209 13711 122327
rect 13593 122049 13711 122167
rect 13593 104209 13711 104327
rect 13593 104049 13711 104167
rect 13593 86209 13711 86327
rect 13593 86049 13711 86167
rect 13593 68209 13711 68327
rect 13593 68049 13711 68167
rect 13593 50209 13711 50327
rect 13593 50049 13711 50167
rect 13593 32209 13711 32327
rect 13593 32049 13711 32167
rect 13593 14209 13711 14327
rect 13593 14049 13711 14167
rect 13593 -2641 13711 -2523
rect 13593 -2801 13711 -2683
rect 24393 355121 24511 355239
rect 24393 354961 24511 355079
rect 22593 354181 22711 354299
rect 22593 354021 22711 354139
rect 20793 353241 20911 353359
rect 20793 353081 20911 353199
rect 15393 340009 15511 340127
rect 15393 339849 15511 339967
rect 15393 322009 15511 322127
rect 15393 321849 15511 321967
rect 15393 304009 15511 304127
rect 15393 303849 15511 303967
rect 15393 286009 15511 286127
rect 15393 285849 15511 285967
rect 15393 268009 15511 268127
rect 15393 267849 15511 267967
rect 15393 250009 15511 250127
rect 15393 249849 15511 249967
rect 15393 232009 15511 232127
rect 15393 231849 15511 231967
rect 15393 214009 15511 214127
rect 15393 213849 15511 213967
rect 15393 196009 15511 196127
rect 15393 195849 15511 195967
rect 15393 178009 15511 178127
rect 15393 177849 15511 177967
rect 15393 160009 15511 160127
rect 15393 159849 15511 159967
rect 15393 142009 15511 142127
rect 15393 141849 15511 141967
rect 15393 124009 15511 124127
rect 15393 123849 15511 123967
rect 15393 106009 15511 106127
rect 15393 105849 15511 105967
rect 15393 88009 15511 88127
rect 15393 87849 15511 87967
rect 15393 70009 15511 70127
rect 15393 69849 15511 69967
rect 15393 52009 15511 52127
rect 15393 51849 15511 51967
rect 15393 34009 15511 34127
rect 15393 33849 15511 33967
rect 15393 16009 15511 16127
rect 15393 15849 15511 15967
rect 6393 -3111 6511 -2993
rect 6393 -3271 6511 -3153
rect -4197 -3581 -4079 -3463
rect -4197 -3741 -4079 -3623
rect 18993 352301 19111 352419
rect 18993 352141 19111 352259
rect 18993 343609 19111 343727
rect 18993 343449 19111 343567
rect 18993 325609 19111 325727
rect 18993 325449 19111 325567
rect 18993 307609 19111 307727
rect 18993 307449 19111 307567
rect 18993 289609 19111 289727
rect 18993 289449 19111 289567
rect 18993 271609 19111 271727
rect 18993 271449 19111 271567
rect 18993 253609 19111 253727
rect 18993 253449 19111 253567
rect 18993 235609 19111 235727
rect 18993 235449 19111 235567
rect 18993 217609 19111 217727
rect 18993 217449 19111 217567
rect 18993 199609 19111 199727
rect 18993 199449 19111 199567
rect 18993 181609 19111 181727
rect 18993 181449 19111 181567
rect 18993 163609 19111 163727
rect 18993 163449 19111 163567
rect 18993 145609 19111 145727
rect 18993 145449 19111 145567
rect 18993 127609 19111 127727
rect 18993 127449 19111 127567
rect 18993 109609 19111 109727
rect 18993 109449 19111 109567
rect 18993 91609 19111 91727
rect 18993 91449 19111 91567
rect 18993 73609 19111 73727
rect 18993 73449 19111 73567
rect 18993 55609 19111 55727
rect 18993 55449 19111 55567
rect 18993 37609 19111 37727
rect 18993 37449 19111 37567
rect 18993 19609 19111 19727
rect 18993 19449 19111 19567
rect 18993 1609 19111 1727
rect 18993 1449 19111 1567
rect 18993 -291 19111 -173
rect 18993 -451 19111 -333
rect 20793 345409 20911 345527
rect 20793 345249 20911 345367
rect 20793 327409 20911 327527
rect 20793 327249 20911 327367
rect 20793 309409 20911 309527
rect 20793 309249 20911 309367
rect 20793 291409 20911 291527
rect 20793 291249 20911 291367
rect 20793 273409 20911 273527
rect 20793 273249 20911 273367
rect 20793 255409 20911 255527
rect 20793 255249 20911 255367
rect 20793 237409 20911 237527
rect 20793 237249 20911 237367
rect 20793 219409 20911 219527
rect 20793 219249 20911 219367
rect 20793 201409 20911 201527
rect 20793 201249 20911 201367
rect 20793 183409 20911 183527
rect 20793 183249 20911 183367
rect 20793 165409 20911 165527
rect 20793 165249 20911 165367
rect 20793 147409 20911 147527
rect 20793 147249 20911 147367
rect 20793 129409 20911 129527
rect 20793 129249 20911 129367
rect 20793 111409 20911 111527
rect 20793 111249 20911 111367
rect 20793 93409 20911 93527
rect 20793 93249 20911 93367
rect 20793 75409 20911 75527
rect 20793 75249 20911 75367
rect 20793 57409 20911 57527
rect 20793 57249 20911 57367
rect 20793 39409 20911 39527
rect 20793 39249 20911 39367
rect 20793 21409 20911 21527
rect 20793 21249 20911 21367
rect 20793 3409 20911 3527
rect 20793 3249 20911 3367
rect 20793 -1231 20911 -1113
rect 20793 -1391 20911 -1273
rect 22593 347209 22711 347327
rect 22593 347049 22711 347167
rect 22593 329209 22711 329327
rect 22593 329049 22711 329167
rect 22593 311209 22711 311327
rect 22593 311049 22711 311167
rect 22593 293209 22711 293327
rect 22593 293049 22711 293167
rect 22593 275209 22711 275327
rect 22593 275049 22711 275167
rect 22593 257209 22711 257327
rect 22593 257049 22711 257167
rect 22593 239209 22711 239327
rect 22593 239049 22711 239167
rect 22593 221209 22711 221327
rect 22593 221049 22711 221167
rect 22593 203209 22711 203327
rect 22593 203049 22711 203167
rect 22593 185209 22711 185327
rect 22593 185049 22711 185167
rect 22593 167209 22711 167327
rect 22593 167049 22711 167167
rect 22593 149209 22711 149327
rect 22593 149049 22711 149167
rect 22593 131209 22711 131327
rect 22593 131049 22711 131167
rect 22593 113209 22711 113327
rect 22593 113049 22711 113167
rect 22593 95209 22711 95327
rect 22593 95049 22711 95167
rect 22593 77209 22711 77327
rect 22593 77049 22711 77167
rect 22593 59209 22711 59327
rect 22593 59049 22711 59167
rect 22593 41209 22711 41327
rect 22593 41049 22711 41167
rect 22593 23209 22711 23327
rect 22593 23049 22711 23167
rect 22593 5209 22711 5327
rect 22593 5049 22711 5167
rect 22593 -2171 22711 -2053
rect 22593 -2331 22711 -2213
rect 33393 355591 33511 355709
rect 33393 355431 33511 355549
rect 31593 354651 31711 354769
rect 31593 354491 31711 354609
rect 29793 353711 29911 353829
rect 29793 353551 29911 353669
rect 24393 349009 24511 349127
rect 24393 348849 24511 348967
rect 24393 331009 24511 331127
rect 24393 330849 24511 330967
rect 24393 313009 24511 313127
rect 24393 312849 24511 312967
rect 24393 295009 24511 295127
rect 24393 294849 24511 294967
rect 24393 277009 24511 277127
rect 24393 276849 24511 276967
rect 24393 259009 24511 259127
rect 24393 258849 24511 258967
rect 24393 241009 24511 241127
rect 24393 240849 24511 240967
rect 24393 223009 24511 223127
rect 24393 222849 24511 222967
rect 24393 205009 24511 205127
rect 24393 204849 24511 204967
rect 24393 187009 24511 187127
rect 24393 186849 24511 186967
rect 24393 169009 24511 169127
rect 24393 168849 24511 168967
rect 24393 151009 24511 151127
rect 24393 150849 24511 150967
rect 24393 133009 24511 133127
rect 24393 132849 24511 132967
rect 24393 115009 24511 115127
rect 24393 114849 24511 114967
rect 24393 97009 24511 97127
rect 24393 96849 24511 96967
rect 24393 79009 24511 79127
rect 24393 78849 24511 78967
rect 24393 61009 24511 61127
rect 24393 60849 24511 60967
rect 24393 43009 24511 43127
rect 24393 42849 24511 42967
rect 24393 25009 24511 25127
rect 24393 24849 24511 24967
rect 24393 7009 24511 7127
rect 24393 6849 24511 6967
rect 15393 -3581 15511 -3463
rect 15393 -3741 15511 -3623
rect 27993 352771 28111 352889
rect 27993 352611 28111 352729
rect 27993 334609 28111 334727
rect 27993 334449 28111 334567
rect 27993 316609 28111 316727
rect 27993 316449 28111 316567
rect 27993 298609 28111 298727
rect 27993 298449 28111 298567
rect 27993 280609 28111 280727
rect 27993 280449 28111 280567
rect 27993 262609 28111 262727
rect 27993 262449 28111 262567
rect 27993 244609 28111 244727
rect 27993 244449 28111 244567
rect 27993 226609 28111 226727
rect 27993 226449 28111 226567
rect 27993 208609 28111 208727
rect 27993 208449 28111 208567
rect 27993 190609 28111 190727
rect 27993 190449 28111 190567
rect 27993 172609 28111 172727
rect 27993 172449 28111 172567
rect 27993 154609 28111 154727
rect 27993 154449 28111 154567
rect 27993 136609 28111 136727
rect 27993 136449 28111 136567
rect 27993 118609 28111 118727
rect 27993 118449 28111 118567
rect 27993 100609 28111 100727
rect 27993 100449 28111 100567
rect 27993 82609 28111 82727
rect 27993 82449 28111 82567
rect 27993 64609 28111 64727
rect 27993 64449 28111 64567
rect 27993 46609 28111 46727
rect 27993 46449 28111 46567
rect 27993 28609 28111 28727
rect 27993 28449 28111 28567
rect 27993 10609 28111 10727
rect 27993 10449 28111 10567
rect 27993 -761 28111 -643
rect 27993 -921 28111 -803
rect 29793 336409 29911 336527
rect 29793 336249 29911 336367
rect 29793 318409 29911 318527
rect 29793 318249 29911 318367
rect 29793 300409 29911 300527
rect 29793 300249 29911 300367
rect 29793 282409 29911 282527
rect 29793 282249 29911 282367
rect 29793 264409 29911 264527
rect 29793 264249 29911 264367
rect 29793 246409 29911 246527
rect 29793 246249 29911 246367
rect 29793 228409 29911 228527
rect 29793 228249 29911 228367
rect 29793 210409 29911 210527
rect 29793 210249 29911 210367
rect 29793 192409 29911 192527
rect 29793 192249 29911 192367
rect 29793 174409 29911 174527
rect 29793 174249 29911 174367
rect 29793 156409 29911 156527
rect 29793 156249 29911 156367
rect 29793 138409 29911 138527
rect 29793 138249 29911 138367
rect 29793 120409 29911 120527
rect 29793 120249 29911 120367
rect 29793 102409 29911 102527
rect 29793 102249 29911 102367
rect 29793 84409 29911 84527
rect 29793 84249 29911 84367
rect 29793 66409 29911 66527
rect 29793 66249 29911 66367
rect 29793 48409 29911 48527
rect 29793 48249 29911 48367
rect 29793 30409 29911 30527
rect 29793 30249 29911 30367
rect 29793 12409 29911 12527
rect 29793 12249 29911 12367
rect 29793 -1701 29911 -1583
rect 29793 -1861 29911 -1743
rect 31593 338209 31711 338327
rect 31593 338049 31711 338167
rect 31593 320209 31711 320327
rect 31593 320049 31711 320167
rect 31593 302209 31711 302327
rect 31593 302049 31711 302167
rect 31593 284209 31711 284327
rect 31593 284049 31711 284167
rect 31593 266209 31711 266327
rect 31593 266049 31711 266167
rect 31593 248209 31711 248327
rect 31593 248049 31711 248167
rect 31593 230209 31711 230327
rect 31593 230049 31711 230167
rect 31593 212209 31711 212327
rect 31593 212049 31711 212167
rect 31593 194209 31711 194327
rect 31593 194049 31711 194167
rect 31593 176209 31711 176327
rect 31593 176049 31711 176167
rect 31593 158209 31711 158327
rect 31593 158049 31711 158167
rect 31593 140209 31711 140327
rect 31593 140049 31711 140167
rect 31593 122209 31711 122327
rect 31593 122049 31711 122167
rect 31593 104209 31711 104327
rect 31593 104049 31711 104167
rect 31593 86209 31711 86327
rect 31593 86049 31711 86167
rect 31593 68209 31711 68327
rect 31593 68049 31711 68167
rect 31593 50209 31711 50327
rect 31593 50049 31711 50167
rect 31593 32209 31711 32327
rect 31593 32049 31711 32167
rect 31593 14209 31711 14327
rect 31593 14049 31711 14167
rect 31593 -2641 31711 -2523
rect 31593 -2801 31711 -2683
rect 42393 355121 42511 355239
rect 42393 354961 42511 355079
rect 40593 354181 40711 354299
rect 40593 354021 40711 354139
rect 38793 353241 38911 353359
rect 38793 353081 38911 353199
rect 33393 340009 33511 340127
rect 33393 339849 33511 339967
rect 33393 322009 33511 322127
rect 33393 321849 33511 321967
rect 33393 304009 33511 304127
rect 33393 303849 33511 303967
rect 33393 286009 33511 286127
rect 33393 285849 33511 285967
rect 33393 268009 33511 268127
rect 33393 267849 33511 267967
rect 33393 250009 33511 250127
rect 33393 249849 33511 249967
rect 33393 232009 33511 232127
rect 33393 231849 33511 231967
rect 33393 214009 33511 214127
rect 33393 213849 33511 213967
rect 33393 196009 33511 196127
rect 33393 195849 33511 195967
rect 33393 178009 33511 178127
rect 33393 177849 33511 177967
rect 33393 160009 33511 160127
rect 33393 159849 33511 159967
rect 33393 142009 33511 142127
rect 33393 141849 33511 141967
rect 33393 124009 33511 124127
rect 33393 123849 33511 123967
rect 33393 106009 33511 106127
rect 33393 105849 33511 105967
rect 33393 88009 33511 88127
rect 33393 87849 33511 87967
rect 33393 70009 33511 70127
rect 33393 69849 33511 69967
rect 33393 52009 33511 52127
rect 33393 51849 33511 51967
rect 33393 34009 33511 34127
rect 33393 33849 33511 33967
rect 33393 16009 33511 16127
rect 33393 15849 33511 15967
rect 24393 -3111 24511 -2993
rect 24393 -3271 24511 -3153
rect 36993 352301 37111 352419
rect 36993 352141 37111 352259
rect 36993 343609 37111 343727
rect 36993 343449 37111 343567
rect 36993 325609 37111 325727
rect 36993 325449 37111 325567
rect 36993 307609 37111 307727
rect 36993 307449 37111 307567
rect 36993 289609 37111 289727
rect 36993 289449 37111 289567
rect 36993 271609 37111 271727
rect 36993 271449 37111 271567
rect 36993 253609 37111 253727
rect 36993 253449 37111 253567
rect 36993 235609 37111 235727
rect 36993 235449 37111 235567
rect 36993 217609 37111 217727
rect 36993 217449 37111 217567
rect 36993 199609 37111 199727
rect 36993 199449 37111 199567
rect 36993 181609 37111 181727
rect 36993 181449 37111 181567
rect 36993 163609 37111 163727
rect 36993 163449 37111 163567
rect 36993 145609 37111 145727
rect 36993 145449 37111 145567
rect 36993 127609 37111 127727
rect 36993 127449 37111 127567
rect 36993 109609 37111 109727
rect 36993 109449 37111 109567
rect 36993 91609 37111 91727
rect 36993 91449 37111 91567
rect 36993 73609 37111 73727
rect 36993 73449 37111 73567
rect 36993 55609 37111 55727
rect 36993 55449 37111 55567
rect 36993 37609 37111 37727
rect 36993 37449 37111 37567
rect 36993 19609 37111 19727
rect 36993 19449 37111 19567
rect 36993 1609 37111 1727
rect 36993 1449 37111 1567
rect 36993 -291 37111 -173
rect 36993 -451 37111 -333
rect 38793 345409 38911 345527
rect 38793 345249 38911 345367
rect 38793 327409 38911 327527
rect 38793 327249 38911 327367
rect 38793 309409 38911 309527
rect 38793 309249 38911 309367
rect 38793 291409 38911 291527
rect 38793 291249 38911 291367
rect 38793 273409 38911 273527
rect 38793 273249 38911 273367
rect 38793 255409 38911 255527
rect 38793 255249 38911 255367
rect 38793 237409 38911 237527
rect 38793 237249 38911 237367
rect 38793 219409 38911 219527
rect 38793 219249 38911 219367
rect 38793 201409 38911 201527
rect 38793 201249 38911 201367
rect 38793 183409 38911 183527
rect 38793 183249 38911 183367
rect 38793 165409 38911 165527
rect 38793 165249 38911 165367
rect 38793 147409 38911 147527
rect 38793 147249 38911 147367
rect 38793 129409 38911 129527
rect 38793 129249 38911 129367
rect 38793 111409 38911 111527
rect 38793 111249 38911 111367
rect 38793 93409 38911 93527
rect 38793 93249 38911 93367
rect 38793 75409 38911 75527
rect 38793 75249 38911 75367
rect 38793 57409 38911 57527
rect 38793 57249 38911 57367
rect 38793 39409 38911 39527
rect 38793 39249 38911 39367
rect 38793 21409 38911 21527
rect 38793 21249 38911 21367
rect 38793 3409 38911 3527
rect 38793 3249 38911 3367
rect 38793 -1231 38911 -1113
rect 38793 -1391 38911 -1273
rect 40593 347209 40711 347327
rect 40593 347049 40711 347167
rect 40593 329209 40711 329327
rect 40593 329049 40711 329167
rect 40593 311209 40711 311327
rect 40593 311049 40711 311167
rect 40593 293209 40711 293327
rect 40593 293049 40711 293167
rect 40593 275209 40711 275327
rect 40593 275049 40711 275167
rect 40593 257209 40711 257327
rect 40593 257049 40711 257167
rect 40593 239209 40711 239327
rect 40593 239049 40711 239167
rect 40593 221209 40711 221327
rect 40593 221049 40711 221167
rect 40593 203209 40711 203327
rect 40593 203049 40711 203167
rect 40593 185209 40711 185327
rect 40593 185049 40711 185167
rect 40593 167209 40711 167327
rect 40593 167049 40711 167167
rect 40593 149209 40711 149327
rect 40593 149049 40711 149167
rect 40593 131209 40711 131327
rect 40593 131049 40711 131167
rect 40593 113209 40711 113327
rect 40593 113049 40711 113167
rect 40593 95209 40711 95327
rect 40593 95049 40711 95167
rect 40593 77209 40711 77327
rect 40593 77049 40711 77167
rect 40593 59209 40711 59327
rect 40593 59049 40711 59167
rect 40593 41209 40711 41327
rect 40593 41049 40711 41167
rect 40593 23209 40711 23327
rect 40593 23049 40711 23167
rect 40593 5209 40711 5327
rect 40593 5049 40711 5167
rect 40593 -2171 40711 -2053
rect 40593 -2331 40711 -2213
rect 51393 355591 51511 355709
rect 51393 355431 51511 355549
rect 49593 354651 49711 354769
rect 49593 354491 49711 354609
rect 47793 353711 47911 353829
rect 47793 353551 47911 353669
rect 42393 349009 42511 349127
rect 42393 348849 42511 348967
rect 42393 331009 42511 331127
rect 42393 330849 42511 330967
rect 42393 313009 42511 313127
rect 42393 312849 42511 312967
rect 42393 295009 42511 295127
rect 42393 294849 42511 294967
rect 42393 277009 42511 277127
rect 42393 276849 42511 276967
rect 42393 259009 42511 259127
rect 42393 258849 42511 258967
rect 42393 241009 42511 241127
rect 42393 240849 42511 240967
rect 42393 223009 42511 223127
rect 42393 222849 42511 222967
rect 42393 205009 42511 205127
rect 42393 204849 42511 204967
rect 42393 187009 42511 187127
rect 42393 186849 42511 186967
rect 42393 169009 42511 169127
rect 42393 168849 42511 168967
rect 42393 151009 42511 151127
rect 42393 150849 42511 150967
rect 42393 133009 42511 133127
rect 42393 132849 42511 132967
rect 42393 115009 42511 115127
rect 42393 114849 42511 114967
rect 42393 97009 42511 97127
rect 42393 96849 42511 96967
rect 42393 79009 42511 79127
rect 42393 78849 42511 78967
rect 42393 61009 42511 61127
rect 42393 60849 42511 60967
rect 42393 43009 42511 43127
rect 42393 42849 42511 42967
rect 42393 25009 42511 25127
rect 42393 24849 42511 24967
rect 42393 7009 42511 7127
rect 42393 6849 42511 6967
rect 33393 -3581 33511 -3463
rect 33393 -3741 33511 -3623
rect 45993 352771 46111 352889
rect 45993 352611 46111 352729
rect 45993 334609 46111 334727
rect 45993 334449 46111 334567
rect 45993 316609 46111 316727
rect 45993 316449 46111 316567
rect 45993 298609 46111 298727
rect 45993 298449 46111 298567
rect 45993 280609 46111 280727
rect 45993 280449 46111 280567
rect 45993 262609 46111 262727
rect 45993 262449 46111 262567
rect 45993 244609 46111 244727
rect 45993 244449 46111 244567
rect 45993 226609 46111 226727
rect 45993 226449 46111 226567
rect 45993 208609 46111 208727
rect 45993 208449 46111 208567
rect 45993 190609 46111 190727
rect 45993 190449 46111 190567
rect 45993 172609 46111 172727
rect 45993 172449 46111 172567
rect 45993 154609 46111 154727
rect 45993 154449 46111 154567
rect 45993 136609 46111 136727
rect 45993 136449 46111 136567
rect 45993 118609 46111 118727
rect 45993 118449 46111 118567
rect 45993 100609 46111 100727
rect 45993 100449 46111 100567
rect 45993 82609 46111 82727
rect 45993 82449 46111 82567
rect 45993 64609 46111 64727
rect 45993 64449 46111 64567
rect 45993 46609 46111 46727
rect 45993 46449 46111 46567
rect 45993 28609 46111 28727
rect 45993 28449 46111 28567
rect 45993 10609 46111 10727
rect 45993 10449 46111 10567
rect 45993 -761 46111 -643
rect 45993 -921 46111 -803
rect 47793 336409 47911 336527
rect 47793 336249 47911 336367
rect 47793 318409 47911 318527
rect 47793 318249 47911 318367
rect 47793 300409 47911 300527
rect 47793 300249 47911 300367
rect 47793 282409 47911 282527
rect 47793 282249 47911 282367
rect 47793 264409 47911 264527
rect 47793 264249 47911 264367
rect 47793 246409 47911 246527
rect 47793 246249 47911 246367
rect 47793 228409 47911 228527
rect 47793 228249 47911 228367
rect 47793 210409 47911 210527
rect 47793 210249 47911 210367
rect 47793 192409 47911 192527
rect 47793 192249 47911 192367
rect 47793 174409 47911 174527
rect 47793 174249 47911 174367
rect 47793 156409 47911 156527
rect 47793 156249 47911 156367
rect 47793 138409 47911 138527
rect 47793 138249 47911 138367
rect 47793 120409 47911 120527
rect 47793 120249 47911 120367
rect 47793 102409 47911 102527
rect 47793 102249 47911 102367
rect 47793 84409 47911 84527
rect 47793 84249 47911 84367
rect 47793 66409 47911 66527
rect 47793 66249 47911 66367
rect 47793 48409 47911 48527
rect 47793 48249 47911 48367
rect 47793 30409 47911 30527
rect 47793 30249 47911 30367
rect 47793 12409 47911 12527
rect 47793 12249 47911 12367
rect 47793 -1701 47911 -1583
rect 47793 -1861 47911 -1743
rect 49593 338209 49711 338327
rect 49593 338049 49711 338167
rect 49593 320209 49711 320327
rect 49593 320049 49711 320167
rect 49593 302209 49711 302327
rect 49593 302049 49711 302167
rect 49593 284209 49711 284327
rect 49593 284049 49711 284167
rect 49593 266209 49711 266327
rect 49593 266049 49711 266167
rect 49593 248209 49711 248327
rect 49593 248049 49711 248167
rect 49593 230209 49711 230327
rect 49593 230049 49711 230167
rect 49593 212209 49711 212327
rect 49593 212049 49711 212167
rect 49593 194209 49711 194327
rect 49593 194049 49711 194167
rect 49593 176209 49711 176327
rect 49593 176049 49711 176167
rect 49593 158209 49711 158327
rect 49593 158049 49711 158167
rect 49593 140209 49711 140327
rect 49593 140049 49711 140167
rect 49593 122209 49711 122327
rect 49593 122049 49711 122167
rect 49593 104209 49711 104327
rect 49593 104049 49711 104167
rect 49593 86209 49711 86327
rect 49593 86049 49711 86167
rect 49593 68209 49711 68327
rect 49593 68049 49711 68167
rect 49593 50209 49711 50327
rect 49593 50049 49711 50167
rect 49593 32209 49711 32327
rect 49593 32049 49711 32167
rect 49593 14209 49711 14327
rect 49593 14049 49711 14167
rect 49593 -2641 49711 -2523
rect 49593 -2801 49711 -2683
rect 60393 355121 60511 355239
rect 60393 354961 60511 355079
rect 58593 354181 58711 354299
rect 58593 354021 58711 354139
rect 56793 353241 56911 353359
rect 56793 353081 56911 353199
rect 51393 340009 51511 340127
rect 51393 339849 51511 339967
rect 51393 322009 51511 322127
rect 51393 321849 51511 321967
rect 51393 304009 51511 304127
rect 51393 303849 51511 303967
rect 51393 286009 51511 286127
rect 51393 285849 51511 285967
rect 51393 268009 51511 268127
rect 51393 267849 51511 267967
rect 51393 250009 51511 250127
rect 51393 249849 51511 249967
rect 51393 232009 51511 232127
rect 51393 231849 51511 231967
rect 51393 214009 51511 214127
rect 51393 213849 51511 213967
rect 51393 196009 51511 196127
rect 51393 195849 51511 195967
rect 51393 178009 51511 178127
rect 51393 177849 51511 177967
rect 51393 160009 51511 160127
rect 51393 159849 51511 159967
rect 51393 142009 51511 142127
rect 51393 141849 51511 141967
rect 51393 124009 51511 124127
rect 51393 123849 51511 123967
rect 51393 106009 51511 106127
rect 51393 105849 51511 105967
rect 51393 88009 51511 88127
rect 51393 87849 51511 87967
rect 51393 70009 51511 70127
rect 51393 69849 51511 69967
rect 51393 52009 51511 52127
rect 51393 51849 51511 51967
rect 51393 34009 51511 34127
rect 51393 33849 51511 33967
rect 51393 16009 51511 16127
rect 51393 15849 51511 15967
rect 42393 -3111 42511 -2993
rect 42393 -3271 42511 -3153
rect 54993 352301 55111 352419
rect 54993 352141 55111 352259
rect 54993 343609 55111 343727
rect 54993 343449 55111 343567
rect 54993 325609 55111 325727
rect 54993 325449 55111 325567
rect 54993 307609 55111 307727
rect 54993 307449 55111 307567
rect 54993 289609 55111 289727
rect 54993 289449 55111 289567
rect 54993 271609 55111 271727
rect 54993 271449 55111 271567
rect 54993 253609 55111 253727
rect 54993 253449 55111 253567
rect 54993 235609 55111 235727
rect 54993 235449 55111 235567
rect 54993 217609 55111 217727
rect 54993 217449 55111 217567
rect 54993 199609 55111 199727
rect 54993 199449 55111 199567
rect 54993 181609 55111 181727
rect 54993 181449 55111 181567
rect 54993 163609 55111 163727
rect 54993 163449 55111 163567
rect 54993 145609 55111 145727
rect 54993 145449 55111 145567
rect 54993 127609 55111 127727
rect 54993 127449 55111 127567
rect 54993 109609 55111 109727
rect 54993 109449 55111 109567
rect 54993 91609 55111 91727
rect 54993 91449 55111 91567
rect 54993 73609 55111 73727
rect 54993 73449 55111 73567
rect 54993 55609 55111 55727
rect 54993 55449 55111 55567
rect 54993 37609 55111 37727
rect 54993 37449 55111 37567
rect 54993 19609 55111 19727
rect 54993 19449 55111 19567
rect 54993 1609 55111 1727
rect 54993 1449 55111 1567
rect 54993 -291 55111 -173
rect 54993 -451 55111 -333
rect 56793 345409 56911 345527
rect 56793 345249 56911 345367
rect 56793 327409 56911 327527
rect 56793 327249 56911 327367
rect 56793 309409 56911 309527
rect 56793 309249 56911 309367
rect 56793 291409 56911 291527
rect 56793 291249 56911 291367
rect 56793 273409 56911 273527
rect 56793 273249 56911 273367
rect 56793 255409 56911 255527
rect 56793 255249 56911 255367
rect 56793 237409 56911 237527
rect 56793 237249 56911 237367
rect 56793 219409 56911 219527
rect 56793 219249 56911 219367
rect 56793 201409 56911 201527
rect 56793 201249 56911 201367
rect 56793 183409 56911 183527
rect 56793 183249 56911 183367
rect 56793 165409 56911 165527
rect 56793 165249 56911 165367
rect 56793 147409 56911 147527
rect 56793 147249 56911 147367
rect 56793 129409 56911 129527
rect 56793 129249 56911 129367
rect 56793 111409 56911 111527
rect 56793 111249 56911 111367
rect 56793 93409 56911 93527
rect 56793 93249 56911 93367
rect 56793 75409 56911 75527
rect 56793 75249 56911 75367
rect 56793 57409 56911 57527
rect 56793 57249 56911 57367
rect 56793 39409 56911 39527
rect 56793 39249 56911 39367
rect 56793 21409 56911 21527
rect 56793 21249 56911 21367
rect 56793 3409 56911 3527
rect 56793 3249 56911 3367
rect 56793 -1231 56911 -1113
rect 56793 -1391 56911 -1273
rect 58593 347209 58711 347327
rect 58593 347049 58711 347167
rect 58593 329209 58711 329327
rect 58593 329049 58711 329167
rect 58593 311209 58711 311327
rect 58593 311049 58711 311167
rect 58593 293209 58711 293327
rect 58593 293049 58711 293167
rect 58593 275209 58711 275327
rect 58593 275049 58711 275167
rect 58593 257209 58711 257327
rect 58593 257049 58711 257167
rect 58593 239209 58711 239327
rect 58593 239049 58711 239167
rect 58593 221209 58711 221327
rect 58593 221049 58711 221167
rect 58593 203209 58711 203327
rect 58593 203049 58711 203167
rect 58593 185209 58711 185327
rect 58593 185049 58711 185167
rect 58593 167209 58711 167327
rect 58593 167049 58711 167167
rect 58593 149209 58711 149327
rect 58593 149049 58711 149167
rect 58593 131209 58711 131327
rect 58593 131049 58711 131167
rect 58593 113209 58711 113327
rect 58593 113049 58711 113167
rect 58593 95209 58711 95327
rect 58593 95049 58711 95167
rect 58593 77209 58711 77327
rect 58593 77049 58711 77167
rect 58593 59209 58711 59327
rect 58593 59049 58711 59167
rect 58593 41209 58711 41327
rect 58593 41049 58711 41167
rect 58593 23209 58711 23327
rect 58593 23049 58711 23167
rect 58593 5209 58711 5327
rect 58593 5049 58711 5167
rect 58593 -2171 58711 -2053
rect 58593 -2331 58711 -2213
rect 69393 355591 69511 355709
rect 69393 355431 69511 355549
rect 67593 354651 67711 354769
rect 67593 354491 67711 354609
rect 65793 353711 65911 353829
rect 65793 353551 65911 353669
rect 60393 349009 60511 349127
rect 60393 348849 60511 348967
rect 60393 331009 60511 331127
rect 60393 330849 60511 330967
rect 60393 313009 60511 313127
rect 60393 312849 60511 312967
rect 60393 295009 60511 295127
rect 60393 294849 60511 294967
rect 60393 277009 60511 277127
rect 60393 276849 60511 276967
rect 60393 259009 60511 259127
rect 60393 258849 60511 258967
rect 60393 241009 60511 241127
rect 60393 240849 60511 240967
rect 60393 223009 60511 223127
rect 60393 222849 60511 222967
rect 60393 205009 60511 205127
rect 60393 204849 60511 204967
rect 60393 187009 60511 187127
rect 60393 186849 60511 186967
rect 60393 169009 60511 169127
rect 60393 168849 60511 168967
rect 60393 151009 60511 151127
rect 60393 150849 60511 150967
rect 60393 133009 60511 133127
rect 60393 132849 60511 132967
rect 60393 115009 60511 115127
rect 60393 114849 60511 114967
rect 60393 97009 60511 97127
rect 60393 96849 60511 96967
rect 60393 79009 60511 79127
rect 60393 78849 60511 78967
rect 60393 61009 60511 61127
rect 60393 60849 60511 60967
rect 60393 43009 60511 43127
rect 60393 42849 60511 42967
rect 60393 25009 60511 25127
rect 60393 24849 60511 24967
rect 60393 7009 60511 7127
rect 60393 6849 60511 6967
rect 51393 -3581 51511 -3463
rect 51393 -3741 51511 -3623
rect 63993 352771 64111 352889
rect 63993 352611 64111 352729
rect 63993 334609 64111 334727
rect 63993 334449 64111 334567
rect 63993 316609 64111 316727
rect 63993 316449 64111 316567
rect 63993 298609 64111 298727
rect 63993 298449 64111 298567
rect 63993 280609 64111 280727
rect 63993 280449 64111 280567
rect 63993 262609 64111 262727
rect 63993 262449 64111 262567
rect 63993 244609 64111 244727
rect 63993 244449 64111 244567
rect 63993 226609 64111 226727
rect 63993 226449 64111 226567
rect 63993 208609 64111 208727
rect 63993 208449 64111 208567
rect 63993 190609 64111 190727
rect 63993 190449 64111 190567
rect 63993 172609 64111 172727
rect 63993 172449 64111 172567
rect 63993 154609 64111 154727
rect 63993 154449 64111 154567
rect 63993 136609 64111 136727
rect 63993 136449 64111 136567
rect 63993 118609 64111 118727
rect 63993 118449 64111 118567
rect 63993 100609 64111 100727
rect 63993 100449 64111 100567
rect 63993 82609 64111 82727
rect 63993 82449 64111 82567
rect 63993 64609 64111 64727
rect 63993 64449 64111 64567
rect 63993 46609 64111 46727
rect 63993 46449 64111 46567
rect 63993 28609 64111 28727
rect 63993 28449 64111 28567
rect 63993 10609 64111 10727
rect 63993 10449 64111 10567
rect 63993 -761 64111 -643
rect 63993 -921 64111 -803
rect 65793 336409 65911 336527
rect 65793 336249 65911 336367
rect 65793 318409 65911 318527
rect 65793 318249 65911 318367
rect 65793 300409 65911 300527
rect 65793 300249 65911 300367
rect 65793 282409 65911 282527
rect 65793 282249 65911 282367
rect 65793 264409 65911 264527
rect 65793 264249 65911 264367
rect 65793 246409 65911 246527
rect 65793 246249 65911 246367
rect 65793 228409 65911 228527
rect 65793 228249 65911 228367
rect 65793 210409 65911 210527
rect 65793 210249 65911 210367
rect 65793 192409 65911 192527
rect 65793 192249 65911 192367
rect 65793 174409 65911 174527
rect 65793 174249 65911 174367
rect 65793 156409 65911 156527
rect 65793 156249 65911 156367
rect 65793 138409 65911 138527
rect 65793 138249 65911 138367
rect 65793 120409 65911 120527
rect 65793 120249 65911 120367
rect 65793 102409 65911 102527
rect 65793 102249 65911 102367
rect 65793 84409 65911 84527
rect 65793 84249 65911 84367
rect 65793 66409 65911 66527
rect 65793 66249 65911 66367
rect 65793 48409 65911 48527
rect 65793 48249 65911 48367
rect 65793 30409 65911 30527
rect 65793 30249 65911 30367
rect 65793 12409 65911 12527
rect 65793 12249 65911 12367
rect 65793 -1701 65911 -1583
rect 65793 -1861 65911 -1743
rect 67593 338209 67711 338327
rect 67593 338049 67711 338167
rect 67593 320209 67711 320327
rect 67593 320049 67711 320167
rect 67593 302209 67711 302327
rect 67593 302049 67711 302167
rect 67593 284209 67711 284327
rect 67593 284049 67711 284167
rect 67593 266209 67711 266327
rect 67593 266049 67711 266167
rect 67593 248209 67711 248327
rect 67593 248049 67711 248167
rect 67593 230209 67711 230327
rect 67593 230049 67711 230167
rect 67593 212209 67711 212327
rect 67593 212049 67711 212167
rect 67593 194209 67711 194327
rect 67593 194049 67711 194167
rect 67593 176209 67711 176327
rect 67593 176049 67711 176167
rect 67593 158209 67711 158327
rect 67593 158049 67711 158167
rect 67593 140209 67711 140327
rect 67593 140049 67711 140167
rect 67593 122209 67711 122327
rect 67593 122049 67711 122167
rect 67593 104209 67711 104327
rect 67593 104049 67711 104167
rect 67593 86209 67711 86327
rect 67593 86049 67711 86167
rect 67593 68209 67711 68327
rect 67593 68049 67711 68167
rect 67593 50209 67711 50327
rect 67593 50049 67711 50167
rect 67593 32209 67711 32327
rect 67593 32049 67711 32167
rect 67593 14209 67711 14327
rect 67593 14049 67711 14167
rect 67593 -2641 67711 -2523
rect 67593 -2801 67711 -2683
rect 78393 355121 78511 355239
rect 78393 354961 78511 355079
rect 76593 354181 76711 354299
rect 76593 354021 76711 354139
rect 74793 353241 74911 353359
rect 74793 353081 74911 353199
rect 69393 340009 69511 340127
rect 69393 339849 69511 339967
rect 69393 322009 69511 322127
rect 69393 321849 69511 321967
rect 69393 304009 69511 304127
rect 69393 303849 69511 303967
rect 69393 286009 69511 286127
rect 69393 285849 69511 285967
rect 69393 268009 69511 268127
rect 69393 267849 69511 267967
rect 69393 250009 69511 250127
rect 69393 249849 69511 249967
rect 69393 232009 69511 232127
rect 69393 231849 69511 231967
rect 69393 214009 69511 214127
rect 69393 213849 69511 213967
rect 69393 196009 69511 196127
rect 69393 195849 69511 195967
rect 69393 178009 69511 178127
rect 69393 177849 69511 177967
rect 69393 160009 69511 160127
rect 69393 159849 69511 159967
rect 69393 142009 69511 142127
rect 69393 141849 69511 141967
rect 69393 124009 69511 124127
rect 69393 123849 69511 123967
rect 69393 106009 69511 106127
rect 69393 105849 69511 105967
rect 69393 88009 69511 88127
rect 69393 87849 69511 87967
rect 69393 70009 69511 70127
rect 69393 69849 69511 69967
rect 69393 52009 69511 52127
rect 69393 51849 69511 51967
rect 69393 34009 69511 34127
rect 69393 33849 69511 33967
rect 69393 16009 69511 16127
rect 69393 15849 69511 15967
rect 60393 -3111 60511 -2993
rect 60393 -3271 60511 -3153
rect 72993 352301 73111 352419
rect 72993 352141 73111 352259
rect 72993 343609 73111 343727
rect 72993 343449 73111 343567
rect 72993 325609 73111 325727
rect 72993 325449 73111 325567
rect 72993 307609 73111 307727
rect 72993 307449 73111 307567
rect 72993 289609 73111 289727
rect 72993 289449 73111 289567
rect 72993 271609 73111 271727
rect 72993 271449 73111 271567
rect 72993 253609 73111 253727
rect 72993 253449 73111 253567
rect 72993 235609 73111 235727
rect 72993 235449 73111 235567
rect 72993 217609 73111 217727
rect 72993 217449 73111 217567
rect 72993 199609 73111 199727
rect 72993 199449 73111 199567
rect 72993 181609 73111 181727
rect 72993 181449 73111 181567
rect 72993 163609 73111 163727
rect 72993 163449 73111 163567
rect 72993 145609 73111 145727
rect 72993 145449 73111 145567
rect 72993 127609 73111 127727
rect 72993 127449 73111 127567
rect 72993 109609 73111 109727
rect 72993 109449 73111 109567
rect 72993 91609 73111 91727
rect 72993 91449 73111 91567
rect 72993 73609 73111 73727
rect 72993 73449 73111 73567
rect 72993 55609 73111 55727
rect 72993 55449 73111 55567
rect 72993 37609 73111 37727
rect 72993 37449 73111 37567
rect 72993 19609 73111 19727
rect 72993 19449 73111 19567
rect 72993 1609 73111 1727
rect 72993 1449 73111 1567
rect 72993 -291 73111 -173
rect 72993 -451 73111 -333
rect 74793 345409 74911 345527
rect 74793 345249 74911 345367
rect 74793 327409 74911 327527
rect 74793 327249 74911 327367
rect 74793 309409 74911 309527
rect 74793 309249 74911 309367
rect 74793 291409 74911 291527
rect 74793 291249 74911 291367
rect 74793 273409 74911 273527
rect 74793 273249 74911 273367
rect 74793 255409 74911 255527
rect 74793 255249 74911 255367
rect 74793 237409 74911 237527
rect 74793 237249 74911 237367
rect 74793 219409 74911 219527
rect 74793 219249 74911 219367
rect 74793 201409 74911 201527
rect 74793 201249 74911 201367
rect 74793 183409 74911 183527
rect 74793 183249 74911 183367
rect 74793 165409 74911 165527
rect 74793 165249 74911 165367
rect 74793 147409 74911 147527
rect 74793 147249 74911 147367
rect 74793 129409 74911 129527
rect 74793 129249 74911 129367
rect 74793 111409 74911 111527
rect 74793 111249 74911 111367
rect 74793 93409 74911 93527
rect 74793 93249 74911 93367
rect 74793 75409 74911 75527
rect 74793 75249 74911 75367
rect 74793 57409 74911 57527
rect 74793 57249 74911 57367
rect 74793 39409 74911 39527
rect 74793 39249 74911 39367
rect 74793 21409 74911 21527
rect 74793 21249 74911 21367
rect 74793 3409 74911 3527
rect 74793 3249 74911 3367
rect 74793 -1231 74911 -1113
rect 74793 -1391 74911 -1273
rect 76593 347209 76711 347327
rect 76593 347049 76711 347167
rect 76593 329209 76711 329327
rect 76593 329049 76711 329167
rect 76593 311209 76711 311327
rect 76593 311049 76711 311167
rect 76593 293209 76711 293327
rect 76593 293049 76711 293167
rect 76593 275209 76711 275327
rect 76593 275049 76711 275167
rect 76593 257209 76711 257327
rect 76593 257049 76711 257167
rect 76593 239209 76711 239327
rect 76593 239049 76711 239167
rect 76593 221209 76711 221327
rect 76593 221049 76711 221167
rect 76593 203209 76711 203327
rect 76593 203049 76711 203167
rect 76593 185209 76711 185327
rect 76593 185049 76711 185167
rect 76593 167209 76711 167327
rect 76593 167049 76711 167167
rect 76593 149209 76711 149327
rect 76593 149049 76711 149167
rect 76593 131209 76711 131327
rect 76593 131049 76711 131167
rect 76593 113209 76711 113327
rect 76593 113049 76711 113167
rect 76593 95209 76711 95327
rect 76593 95049 76711 95167
rect 76593 77209 76711 77327
rect 76593 77049 76711 77167
rect 76593 59209 76711 59327
rect 76593 59049 76711 59167
rect 76593 41209 76711 41327
rect 76593 41049 76711 41167
rect 76593 23209 76711 23327
rect 76593 23049 76711 23167
rect 76593 5209 76711 5327
rect 76593 5049 76711 5167
rect 76593 -2171 76711 -2053
rect 76593 -2331 76711 -2213
rect 87393 355591 87511 355709
rect 87393 355431 87511 355549
rect 85593 354651 85711 354769
rect 85593 354491 85711 354609
rect 83793 353711 83911 353829
rect 83793 353551 83911 353669
rect 78393 349009 78511 349127
rect 78393 348849 78511 348967
rect 78393 331009 78511 331127
rect 78393 330849 78511 330967
rect 78393 313009 78511 313127
rect 78393 312849 78511 312967
rect 78393 295009 78511 295127
rect 78393 294849 78511 294967
rect 78393 277009 78511 277127
rect 78393 276849 78511 276967
rect 78393 259009 78511 259127
rect 78393 258849 78511 258967
rect 78393 241009 78511 241127
rect 78393 240849 78511 240967
rect 78393 223009 78511 223127
rect 78393 222849 78511 222967
rect 78393 205009 78511 205127
rect 78393 204849 78511 204967
rect 78393 187009 78511 187127
rect 78393 186849 78511 186967
rect 78393 169009 78511 169127
rect 78393 168849 78511 168967
rect 78393 151009 78511 151127
rect 78393 150849 78511 150967
rect 78393 133009 78511 133127
rect 78393 132849 78511 132967
rect 78393 115009 78511 115127
rect 78393 114849 78511 114967
rect 78393 97009 78511 97127
rect 78393 96849 78511 96967
rect 78393 79009 78511 79127
rect 78393 78849 78511 78967
rect 78393 61009 78511 61127
rect 78393 60849 78511 60967
rect 78393 43009 78511 43127
rect 78393 42849 78511 42967
rect 78393 25009 78511 25127
rect 78393 24849 78511 24967
rect 78393 7009 78511 7127
rect 78393 6849 78511 6967
rect 69393 -3581 69511 -3463
rect 69393 -3741 69511 -3623
rect 81993 352771 82111 352889
rect 81993 352611 82111 352729
rect 81993 334609 82111 334727
rect 81993 334449 82111 334567
rect 81993 316609 82111 316727
rect 81993 316449 82111 316567
rect 81993 298609 82111 298727
rect 81993 298449 82111 298567
rect 81993 280609 82111 280727
rect 81993 280449 82111 280567
rect 81993 262609 82111 262727
rect 81993 262449 82111 262567
rect 81993 244609 82111 244727
rect 81993 244449 82111 244567
rect 81993 226609 82111 226727
rect 81993 226449 82111 226567
rect 81993 208609 82111 208727
rect 81993 208449 82111 208567
rect 81993 190609 82111 190727
rect 81993 190449 82111 190567
rect 81993 172609 82111 172727
rect 81993 172449 82111 172567
rect 81993 154609 82111 154727
rect 81993 154449 82111 154567
rect 81993 136609 82111 136727
rect 81993 136449 82111 136567
rect 81993 118609 82111 118727
rect 81993 118449 82111 118567
rect 81993 100609 82111 100727
rect 81993 100449 82111 100567
rect 81993 82609 82111 82727
rect 81993 82449 82111 82567
rect 81993 64609 82111 64727
rect 81993 64449 82111 64567
rect 81993 46609 82111 46727
rect 81993 46449 82111 46567
rect 81993 28609 82111 28727
rect 81993 28449 82111 28567
rect 81993 10609 82111 10727
rect 81993 10449 82111 10567
rect 81993 -761 82111 -643
rect 81993 -921 82111 -803
rect 83793 336409 83911 336527
rect 83793 336249 83911 336367
rect 83793 318409 83911 318527
rect 83793 318249 83911 318367
rect 83793 300409 83911 300527
rect 83793 300249 83911 300367
rect 83793 282409 83911 282527
rect 83793 282249 83911 282367
rect 83793 264409 83911 264527
rect 83793 264249 83911 264367
rect 83793 246409 83911 246527
rect 83793 246249 83911 246367
rect 83793 228409 83911 228527
rect 83793 228249 83911 228367
rect 83793 210409 83911 210527
rect 83793 210249 83911 210367
rect 83793 192409 83911 192527
rect 83793 192249 83911 192367
rect 83793 174409 83911 174527
rect 83793 174249 83911 174367
rect 83793 156409 83911 156527
rect 83793 156249 83911 156367
rect 83793 138409 83911 138527
rect 83793 138249 83911 138367
rect 83793 120409 83911 120527
rect 83793 120249 83911 120367
rect 83793 102409 83911 102527
rect 83793 102249 83911 102367
rect 83793 84409 83911 84527
rect 83793 84249 83911 84367
rect 83793 66409 83911 66527
rect 83793 66249 83911 66367
rect 83793 48409 83911 48527
rect 83793 48249 83911 48367
rect 83793 30409 83911 30527
rect 83793 30249 83911 30367
rect 83793 12409 83911 12527
rect 83793 12249 83911 12367
rect 83793 -1701 83911 -1583
rect 83793 -1861 83911 -1743
rect 85593 338209 85711 338327
rect 85593 338049 85711 338167
rect 85593 320209 85711 320327
rect 85593 320049 85711 320167
rect 85593 302209 85711 302327
rect 85593 302049 85711 302167
rect 85593 284209 85711 284327
rect 85593 284049 85711 284167
rect 85593 266209 85711 266327
rect 85593 266049 85711 266167
rect 85593 248209 85711 248327
rect 85593 248049 85711 248167
rect 85593 230209 85711 230327
rect 85593 230049 85711 230167
rect 85593 212209 85711 212327
rect 85593 212049 85711 212167
rect 85593 194209 85711 194327
rect 85593 194049 85711 194167
rect 85593 176209 85711 176327
rect 85593 176049 85711 176167
rect 85593 158209 85711 158327
rect 85593 158049 85711 158167
rect 85593 140209 85711 140327
rect 85593 140049 85711 140167
rect 85593 122209 85711 122327
rect 85593 122049 85711 122167
rect 85593 104209 85711 104327
rect 85593 104049 85711 104167
rect 85593 86209 85711 86327
rect 85593 86049 85711 86167
rect 85593 68209 85711 68327
rect 85593 68049 85711 68167
rect 85593 50209 85711 50327
rect 85593 50049 85711 50167
rect 85593 32209 85711 32327
rect 85593 32049 85711 32167
rect 85593 14209 85711 14327
rect 85593 14049 85711 14167
rect 85593 -2641 85711 -2523
rect 85593 -2801 85711 -2683
rect 96393 355121 96511 355239
rect 96393 354961 96511 355079
rect 94593 354181 94711 354299
rect 94593 354021 94711 354139
rect 92793 353241 92911 353359
rect 92793 353081 92911 353199
rect 87393 340009 87511 340127
rect 87393 339849 87511 339967
rect 87393 322009 87511 322127
rect 87393 321849 87511 321967
rect 87393 304009 87511 304127
rect 87393 303849 87511 303967
rect 87393 286009 87511 286127
rect 87393 285849 87511 285967
rect 87393 268009 87511 268127
rect 87393 267849 87511 267967
rect 87393 250009 87511 250127
rect 87393 249849 87511 249967
rect 87393 232009 87511 232127
rect 87393 231849 87511 231967
rect 87393 214009 87511 214127
rect 87393 213849 87511 213967
rect 87393 196009 87511 196127
rect 87393 195849 87511 195967
rect 87393 178009 87511 178127
rect 87393 177849 87511 177967
rect 87393 160009 87511 160127
rect 87393 159849 87511 159967
rect 87393 142009 87511 142127
rect 87393 141849 87511 141967
rect 87393 124009 87511 124127
rect 87393 123849 87511 123967
rect 87393 106009 87511 106127
rect 87393 105849 87511 105967
rect 87393 88009 87511 88127
rect 87393 87849 87511 87967
rect 87393 70009 87511 70127
rect 87393 69849 87511 69967
rect 87393 52009 87511 52127
rect 87393 51849 87511 51967
rect 87393 34009 87511 34127
rect 87393 33849 87511 33967
rect 87393 16009 87511 16127
rect 87393 15849 87511 15967
rect 78393 -3111 78511 -2993
rect 78393 -3271 78511 -3153
rect 90993 352301 91111 352419
rect 90993 352141 91111 352259
rect 90993 343609 91111 343727
rect 90993 343449 91111 343567
rect 90993 325609 91111 325727
rect 90993 325449 91111 325567
rect 90993 307609 91111 307727
rect 90993 307449 91111 307567
rect 90993 289609 91111 289727
rect 90993 289449 91111 289567
rect 90993 271609 91111 271727
rect 90993 271449 91111 271567
rect 90993 253609 91111 253727
rect 90993 253449 91111 253567
rect 90993 235609 91111 235727
rect 90993 235449 91111 235567
rect 90993 217609 91111 217727
rect 90993 217449 91111 217567
rect 90993 199609 91111 199727
rect 90993 199449 91111 199567
rect 90993 181609 91111 181727
rect 90993 181449 91111 181567
rect 90993 163609 91111 163727
rect 90993 163449 91111 163567
rect 90993 145609 91111 145727
rect 90993 145449 91111 145567
rect 90993 127609 91111 127727
rect 90993 127449 91111 127567
rect 90993 109609 91111 109727
rect 90993 109449 91111 109567
rect 90993 91609 91111 91727
rect 90993 91449 91111 91567
rect 90993 73609 91111 73727
rect 90993 73449 91111 73567
rect 90993 55609 91111 55727
rect 90993 55449 91111 55567
rect 90993 37609 91111 37727
rect 90993 37449 91111 37567
rect 90993 19609 91111 19727
rect 90993 19449 91111 19567
rect 90993 1609 91111 1727
rect 90993 1449 91111 1567
rect 90993 -291 91111 -173
rect 90993 -451 91111 -333
rect 92793 345409 92911 345527
rect 92793 345249 92911 345367
rect 92793 327409 92911 327527
rect 92793 327249 92911 327367
rect 92793 309409 92911 309527
rect 92793 309249 92911 309367
rect 92793 291409 92911 291527
rect 92793 291249 92911 291367
rect 92793 273409 92911 273527
rect 92793 273249 92911 273367
rect 92793 255409 92911 255527
rect 92793 255249 92911 255367
rect 92793 237409 92911 237527
rect 92793 237249 92911 237367
rect 92793 219409 92911 219527
rect 92793 219249 92911 219367
rect 92793 201409 92911 201527
rect 92793 201249 92911 201367
rect 92793 183409 92911 183527
rect 92793 183249 92911 183367
rect 92793 165409 92911 165527
rect 92793 165249 92911 165367
rect 92793 147409 92911 147527
rect 92793 147249 92911 147367
rect 92793 129409 92911 129527
rect 92793 129249 92911 129367
rect 92793 111409 92911 111527
rect 92793 111249 92911 111367
rect 92793 93409 92911 93527
rect 92793 93249 92911 93367
rect 92793 75409 92911 75527
rect 92793 75249 92911 75367
rect 92793 57409 92911 57527
rect 92793 57249 92911 57367
rect 92793 39409 92911 39527
rect 92793 39249 92911 39367
rect 92793 21409 92911 21527
rect 92793 21249 92911 21367
rect 92793 3409 92911 3527
rect 92793 3249 92911 3367
rect 92793 -1231 92911 -1113
rect 92793 -1391 92911 -1273
rect 94593 347209 94711 347327
rect 94593 347049 94711 347167
rect 94593 329209 94711 329327
rect 94593 329049 94711 329167
rect 94593 311209 94711 311327
rect 94593 311049 94711 311167
rect 94593 293209 94711 293327
rect 94593 293049 94711 293167
rect 94593 275209 94711 275327
rect 94593 275049 94711 275167
rect 94593 257209 94711 257327
rect 94593 257049 94711 257167
rect 94593 239209 94711 239327
rect 94593 239049 94711 239167
rect 94593 221209 94711 221327
rect 94593 221049 94711 221167
rect 94593 203209 94711 203327
rect 94593 203049 94711 203167
rect 94593 185209 94711 185327
rect 94593 185049 94711 185167
rect 94593 167209 94711 167327
rect 94593 167049 94711 167167
rect 94593 149209 94711 149327
rect 94593 149049 94711 149167
rect 94593 131209 94711 131327
rect 94593 131049 94711 131167
rect 94593 113209 94711 113327
rect 94593 113049 94711 113167
rect 94593 95209 94711 95327
rect 94593 95049 94711 95167
rect 94593 77209 94711 77327
rect 94593 77049 94711 77167
rect 94593 59209 94711 59327
rect 94593 59049 94711 59167
rect 94593 41209 94711 41327
rect 94593 41049 94711 41167
rect 94593 23209 94711 23327
rect 94593 23049 94711 23167
rect 94593 5209 94711 5327
rect 94593 5049 94711 5167
rect 94593 -2171 94711 -2053
rect 94593 -2331 94711 -2213
rect 105393 355591 105511 355709
rect 105393 355431 105511 355549
rect 103593 354651 103711 354769
rect 103593 354491 103711 354609
rect 101793 353711 101911 353829
rect 101793 353551 101911 353669
rect 96393 349009 96511 349127
rect 96393 348849 96511 348967
rect 96393 331009 96511 331127
rect 96393 330849 96511 330967
rect 96393 313009 96511 313127
rect 96393 312849 96511 312967
rect 96393 295009 96511 295127
rect 96393 294849 96511 294967
rect 96393 277009 96511 277127
rect 96393 276849 96511 276967
rect 96393 259009 96511 259127
rect 96393 258849 96511 258967
rect 96393 241009 96511 241127
rect 96393 240849 96511 240967
rect 96393 223009 96511 223127
rect 96393 222849 96511 222967
rect 96393 205009 96511 205127
rect 96393 204849 96511 204967
rect 96393 187009 96511 187127
rect 96393 186849 96511 186967
rect 96393 169009 96511 169127
rect 96393 168849 96511 168967
rect 96393 151009 96511 151127
rect 96393 150849 96511 150967
rect 96393 133009 96511 133127
rect 96393 132849 96511 132967
rect 96393 115009 96511 115127
rect 96393 114849 96511 114967
rect 96393 97009 96511 97127
rect 96393 96849 96511 96967
rect 96393 79009 96511 79127
rect 96393 78849 96511 78967
rect 96393 61009 96511 61127
rect 96393 60849 96511 60967
rect 96393 43009 96511 43127
rect 96393 42849 96511 42967
rect 96393 25009 96511 25127
rect 96393 24849 96511 24967
rect 96393 7009 96511 7127
rect 96393 6849 96511 6967
rect 87393 -3581 87511 -3463
rect 87393 -3741 87511 -3623
rect 99993 352771 100111 352889
rect 99993 352611 100111 352729
rect 99993 334609 100111 334727
rect 99993 334449 100111 334567
rect 99993 316609 100111 316727
rect 99993 316449 100111 316567
rect 99993 298609 100111 298727
rect 99993 298449 100111 298567
rect 99993 280609 100111 280727
rect 99993 280449 100111 280567
rect 99993 262609 100111 262727
rect 99993 262449 100111 262567
rect 99993 244609 100111 244727
rect 99993 244449 100111 244567
rect 99993 226609 100111 226727
rect 99993 226449 100111 226567
rect 99993 208609 100111 208727
rect 99993 208449 100111 208567
rect 99993 190609 100111 190727
rect 99993 190449 100111 190567
rect 99993 172609 100111 172727
rect 99993 172449 100111 172567
rect 99993 154609 100111 154727
rect 99993 154449 100111 154567
rect 99993 136609 100111 136727
rect 99993 136449 100111 136567
rect 99993 118609 100111 118727
rect 99993 118449 100111 118567
rect 99993 100609 100111 100727
rect 99993 100449 100111 100567
rect 99993 82609 100111 82727
rect 99993 82449 100111 82567
rect 99993 64609 100111 64727
rect 99993 64449 100111 64567
rect 99993 46609 100111 46727
rect 99993 46449 100111 46567
rect 99993 28609 100111 28727
rect 99993 28449 100111 28567
rect 99993 10609 100111 10727
rect 99993 10449 100111 10567
rect 99993 -761 100111 -643
rect 99993 -921 100111 -803
rect 101793 336409 101911 336527
rect 101793 336249 101911 336367
rect 101793 318409 101911 318527
rect 101793 318249 101911 318367
rect 101793 300409 101911 300527
rect 101793 300249 101911 300367
rect 101793 282409 101911 282527
rect 101793 282249 101911 282367
rect 101793 264409 101911 264527
rect 101793 264249 101911 264367
rect 101793 246409 101911 246527
rect 101793 246249 101911 246367
rect 101793 228409 101911 228527
rect 101793 228249 101911 228367
rect 101793 210409 101911 210527
rect 101793 210249 101911 210367
rect 101793 192409 101911 192527
rect 101793 192249 101911 192367
rect 101793 174409 101911 174527
rect 101793 174249 101911 174367
rect 101793 156409 101911 156527
rect 101793 156249 101911 156367
rect 101793 138409 101911 138527
rect 101793 138249 101911 138367
rect 101793 120409 101911 120527
rect 101793 120249 101911 120367
rect 101793 102409 101911 102527
rect 101793 102249 101911 102367
rect 101793 84409 101911 84527
rect 101793 84249 101911 84367
rect 101793 66409 101911 66527
rect 101793 66249 101911 66367
rect 101793 48409 101911 48527
rect 101793 48249 101911 48367
rect 101793 30409 101911 30527
rect 101793 30249 101911 30367
rect 101793 12409 101911 12527
rect 101793 12249 101911 12367
rect 101793 -1701 101911 -1583
rect 101793 -1861 101911 -1743
rect 103593 338209 103711 338327
rect 103593 338049 103711 338167
rect 103593 320209 103711 320327
rect 103593 320049 103711 320167
rect 103593 302209 103711 302327
rect 103593 302049 103711 302167
rect 103593 284209 103711 284327
rect 103593 284049 103711 284167
rect 103593 266209 103711 266327
rect 103593 266049 103711 266167
rect 103593 248209 103711 248327
rect 103593 248049 103711 248167
rect 103593 230209 103711 230327
rect 103593 230049 103711 230167
rect 103593 212209 103711 212327
rect 103593 212049 103711 212167
rect 103593 194209 103711 194327
rect 103593 194049 103711 194167
rect 103593 176209 103711 176327
rect 103593 176049 103711 176167
rect 103593 158209 103711 158327
rect 103593 158049 103711 158167
rect 103593 140209 103711 140327
rect 103593 140049 103711 140167
rect 103593 122209 103711 122327
rect 103593 122049 103711 122167
rect 103593 104209 103711 104327
rect 103593 104049 103711 104167
rect 103593 86209 103711 86327
rect 103593 86049 103711 86167
rect 103593 68209 103711 68327
rect 103593 68049 103711 68167
rect 103593 50209 103711 50327
rect 103593 50049 103711 50167
rect 103593 32209 103711 32327
rect 103593 32049 103711 32167
rect 103593 14209 103711 14327
rect 103593 14049 103711 14167
rect 103593 -2641 103711 -2523
rect 103593 -2801 103711 -2683
rect 114393 355121 114511 355239
rect 114393 354961 114511 355079
rect 112593 354181 112711 354299
rect 112593 354021 112711 354139
rect 110793 353241 110911 353359
rect 110793 353081 110911 353199
rect 105393 340009 105511 340127
rect 105393 339849 105511 339967
rect 105393 322009 105511 322127
rect 105393 321849 105511 321967
rect 105393 304009 105511 304127
rect 105393 303849 105511 303967
rect 105393 286009 105511 286127
rect 105393 285849 105511 285967
rect 105393 268009 105511 268127
rect 105393 267849 105511 267967
rect 105393 250009 105511 250127
rect 105393 249849 105511 249967
rect 105393 232009 105511 232127
rect 105393 231849 105511 231967
rect 105393 214009 105511 214127
rect 105393 213849 105511 213967
rect 105393 196009 105511 196127
rect 105393 195849 105511 195967
rect 105393 178009 105511 178127
rect 105393 177849 105511 177967
rect 105393 160009 105511 160127
rect 105393 159849 105511 159967
rect 105393 142009 105511 142127
rect 105393 141849 105511 141967
rect 105393 124009 105511 124127
rect 105393 123849 105511 123967
rect 105393 106009 105511 106127
rect 105393 105849 105511 105967
rect 105393 88009 105511 88127
rect 105393 87849 105511 87967
rect 105393 70009 105511 70127
rect 105393 69849 105511 69967
rect 105393 52009 105511 52127
rect 105393 51849 105511 51967
rect 105393 34009 105511 34127
rect 105393 33849 105511 33967
rect 105393 16009 105511 16127
rect 105393 15849 105511 15967
rect 96393 -3111 96511 -2993
rect 96393 -3271 96511 -3153
rect 108993 352301 109111 352419
rect 108993 352141 109111 352259
rect 108993 343609 109111 343727
rect 108993 343449 109111 343567
rect 108993 325609 109111 325727
rect 108993 325449 109111 325567
rect 108993 307609 109111 307727
rect 108993 307449 109111 307567
rect 108993 289609 109111 289727
rect 108993 289449 109111 289567
rect 108993 271609 109111 271727
rect 108993 271449 109111 271567
rect 108993 253609 109111 253727
rect 108993 253449 109111 253567
rect 108993 235609 109111 235727
rect 108993 235449 109111 235567
rect 108993 217609 109111 217727
rect 108993 217449 109111 217567
rect 108993 199609 109111 199727
rect 108993 199449 109111 199567
rect 108993 181609 109111 181727
rect 108993 181449 109111 181567
rect 108993 163609 109111 163727
rect 108993 163449 109111 163567
rect 108993 145609 109111 145727
rect 108993 145449 109111 145567
rect 108993 127609 109111 127727
rect 108993 127449 109111 127567
rect 108993 109609 109111 109727
rect 108993 109449 109111 109567
rect 108993 91609 109111 91727
rect 108993 91449 109111 91567
rect 108993 73609 109111 73727
rect 108993 73449 109111 73567
rect 108993 55609 109111 55727
rect 108993 55449 109111 55567
rect 108993 37609 109111 37727
rect 108993 37449 109111 37567
rect 108993 19609 109111 19727
rect 108993 19449 109111 19567
rect 108993 1609 109111 1727
rect 108993 1449 109111 1567
rect 108993 -291 109111 -173
rect 108993 -451 109111 -333
rect 110793 345409 110911 345527
rect 110793 345249 110911 345367
rect 110793 327409 110911 327527
rect 110793 327249 110911 327367
rect 110793 309409 110911 309527
rect 110793 309249 110911 309367
rect 110793 291409 110911 291527
rect 110793 291249 110911 291367
rect 110793 273409 110911 273527
rect 110793 273249 110911 273367
rect 110793 255409 110911 255527
rect 110793 255249 110911 255367
rect 110793 237409 110911 237527
rect 110793 237249 110911 237367
rect 110793 219409 110911 219527
rect 110793 219249 110911 219367
rect 110793 201409 110911 201527
rect 110793 201249 110911 201367
rect 110793 183409 110911 183527
rect 110793 183249 110911 183367
rect 110793 165409 110911 165527
rect 110793 165249 110911 165367
rect 110793 147409 110911 147527
rect 110793 147249 110911 147367
rect 110793 129409 110911 129527
rect 110793 129249 110911 129367
rect 110793 111409 110911 111527
rect 110793 111249 110911 111367
rect 110793 93409 110911 93527
rect 110793 93249 110911 93367
rect 110793 75409 110911 75527
rect 110793 75249 110911 75367
rect 110793 57409 110911 57527
rect 110793 57249 110911 57367
rect 110793 39409 110911 39527
rect 110793 39249 110911 39367
rect 110793 21409 110911 21527
rect 110793 21249 110911 21367
rect 110793 3409 110911 3527
rect 110793 3249 110911 3367
rect 110793 -1231 110911 -1113
rect 110793 -1391 110911 -1273
rect 112593 347209 112711 347327
rect 112593 347049 112711 347167
rect 112593 329209 112711 329327
rect 112593 329049 112711 329167
rect 112593 311209 112711 311327
rect 112593 311049 112711 311167
rect 112593 293209 112711 293327
rect 112593 293049 112711 293167
rect 112593 275209 112711 275327
rect 112593 275049 112711 275167
rect 112593 257209 112711 257327
rect 112593 257049 112711 257167
rect 112593 239209 112711 239327
rect 112593 239049 112711 239167
rect 112593 221209 112711 221327
rect 112593 221049 112711 221167
rect 112593 203209 112711 203327
rect 112593 203049 112711 203167
rect 112593 185209 112711 185327
rect 112593 185049 112711 185167
rect 112593 167209 112711 167327
rect 112593 167049 112711 167167
rect 112593 149209 112711 149327
rect 112593 149049 112711 149167
rect 112593 131209 112711 131327
rect 112593 131049 112711 131167
rect 112593 113209 112711 113327
rect 112593 113049 112711 113167
rect 112593 95209 112711 95327
rect 112593 95049 112711 95167
rect 112593 77209 112711 77327
rect 112593 77049 112711 77167
rect 112593 59209 112711 59327
rect 112593 59049 112711 59167
rect 112593 41209 112711 41327
rect 112593 41049 112711 41167
rect 112593 23209 112711 23327
rect 112593 23049 112711 23167
rect 112593 5209 112711 5327
rect 112593 5049 112711 5167
rect 112593 -2171 112711 -2053
rect 112593 -2331 112711 -2213
rect 123393 355591 123511 355709
rect 123393 355431 123511 355549
rect 121593 354651 121711 354769
rect 121593 354491 121711 354609
rect 119793 353711 119911 353829
rect 119793 353551 119911 353669
rect 114393 349009 114511 349127
rect 114393 348849 114511 348967
rect 114393 331009 114511 331127
rect 114393 330849 114511 330967
rect 114393 313009 114511 313127
rect 114393 312849 114511 312967
rect 114393 295009 114511 295127
rect 114393 294849 114511 294967
rect 114393 277009 114511 277127
rect 114393 276849 114511 276967
rect 114393 259009 114511 259127
rect 114393 258849 114511 258967
rect 114393 241009 114511 241127
rect 114393 240849 114511 240967
rect 114393 223009 114511 223127
rect 114393 222849 114511 222967
rect 114393 205009 114511 205127
rect 114393 204849 114511 204967
rect 114393 187009 114511 187127
rect 114393 186849 114511 186967
rect 114393 169009 114511 169127
rect 114393 168849 114511 168967
rect 114393 151009 114511 151127
rect 114393 150849 114511 150967
rect 114393 133009 114511 133127
rect 114393 132849 114511 132967
rect 114393 115009 114511 115127
rect 114393 114849 114511 114967
rect 114393 97009 114511 97127
rect 114393 96849 114511 96967
rect 114393 79009 114511 79127
rect 114393 78849 114511 78967
rect 114393 61009 114511 61127
rect 114393 60849 114511 60967
rect 114393 43009 114511 43127
rect 114393 42849 114511 42967
rect 114393 25009 114511 25127
rect 114393 24849 114511 24967
rect 114393 7009 114511 7127
rect 114393 6849 114511 6967
rect 105393 -3581 105511 -3463
rect 105393 -3741 105511 -3623
rect 117993 352771 118111 352889
rect 117993 352611 118111 352729
rect 117993 334609 118111 334727
rect 117993 334449 118111 334567
rect 117993 316609 118111 316727
rect 117993 316449 118111 316567
rect 117993 298609 118111 298727
rect 117993 298449 118111 298567
rect 117993 280609 118111 280727
rect 117993 280449 118111 280567
rect 117993 262609 118111 262727
rect 117993 262449 118111 262567
rect 117993 244609 118111 244727
rect 117993 244449 118111 244567
rect 117993 226609 118111 226727
rect 117993 226449 118111 226567
rect 117993 208609 118111 208727
rect 117993 208449 118111 208567
rect 117993 190609 118111 190727
rect 117993 190449 118111 190567
rect 117993 172609 118111 172727
rect 117993 172449 118111 172567
rect 117993 154609 118111 154727
rect 117993 154449 118111 154567
rect 117993 136609 118111 136727
rect 117993 136449 118111 136567
rect 117993 118609 118111 118727
rect 117993 118449 118111 118567
rect 117993 100609 118111 100727
rect 117993 100449 118111 100567
rect 117993 82609 118111 82727
rect 117993 82449 118111 82567
rect 117993 64609 118111 64727
rect 117993 64449 118111 64567
rect 117993 46609 118111 46727
rect 117993 46449 118111 46567
rect 117993 28609 118111 28727
rect 117993 28449 118111 28567
rect 117993 10609 118111 10727
rect 117993 10449 118111 10567
rect 117993 -761 118111 -643
rect 117993 -921 118111 -803
rect 119793 336409 119911 336527
rect 119793 336249 119911 336367
rect 119793 318409 119911 318527
rect 119793 318249 119911 318367
rect 119793 300409 119911 300527
rect 119793 300249 119911 300367
rect 119793 282409 119911 282527
rect 119793 282249 119911 282367
rect 119793 264409 119911 264527
rect 119793 264249 119911 264367
rect 119793 246409 119911 246527
rect 119793 246249 119911 246367
rect 119793 228409 119911 228527
rect 119793 228249 119911 228367
rect 119793 210409 119911 210527
rect 119793 210249 119911 210367
rect 119793 192409 119911 192527
rect 119793 192249 119911 192367
rect 119793 174409 119911 174527
rect 119793 174249 119911 174367
rect 119793 156409 119911 156527
rect 119793 156249 119911 156367
rect 119793 138409 119911 138527
rect 119793 138249 119911 138367
rect 119793 120409 119911 120527
rect 119793 120249 119911 120367
rect 119793 102409 119911 102527
rect 119793 102249 119911 102367
rect 119793 84409 119911 84527
rect 119793 84249 119911 84367
rect 119793 66409 119911 66527
rect 119793 66249 119911 66367
rect 119793 48409 119911 48527
rect 119793 48249 119911 48367
rect 119793 30409 119911 30527
rect 119793 30249 119911 30367
rect 119793 12409 119911 12527
rect 119793 12249 119911 12367
rect 119793 -1701 119911 -1583
rect 119793 -1861 119911 -1743
rect 121593 338209 121711 338327
rect 121593 338049 121711 338167
rect 121593 320209 121711 320327
rect 121593 320049 121711 320167
rect 121593 302209 121711 302327
rect 121593 302049 121711 302167
rect 121593 284209 121711 284327
rect 121593 284049 121711 284167
rect 121593 266209 121711 266327
rect 121593 266049 121711 266167
rect 121593 248209 121711 248327
rect 121593 248049 121711 248167
rect 121593 230209 121711 230327
rect 121593 230049 121711 230167
rect 121593 212209 121711 212327
rect 121593 212049 121711 212167
rect 121593 194209 121711 194327
rect 121593 194049 121711 194167
rect 121593 176209 121711 176327
rect 121593 176049 121711 176167
rect 121593 158209 121711 158327
rect 121593 158049 121711 158167
rect 121593 140209 121711 140327
rect 121593 140049 121711 140167
rect 121593 122209 121711 122327
rect 121593 122049 121711 122167
rect 121593 104209 121711 104327
rect 121593 104049 121711 104167
rect 121593 86209 121711 86327
rect 121593 86049 121711 86167
rect 121593 68209 121711 68327
rect 121593 68049 121711 68167
rect 121593 50209 121711 50327
rect 121593 50049 121711 50167
rect 121593 32209 121711 32327
rect 121593 32049 121711 32167
rect 121593 14209 121711 14327
rect 121593 14049 121711 14167
rect 121593 -2641 121711 -2523
rect 121593 -2801 121711 -2683
rect 132393 355121 132511 355239
rect 132393 354961 132511 355079
rect 130593 354181 130711 354299
rect 130593 354021 130711 354139
rect 128793 353241 128911 353359
rect 128793 353081 128911 353199
rect 123393 340009 123511 340127
rect 123393 339849 123511 339967
rect 123393 322009 123511 322127
rect 123393 321849 123511 321967
rect 123393 304009 123511 304127
rect 123393 303849 123511 303967
rect 123393 286009 123511 286127
rect 123393 285849 123511 285967
rect 123393 268009 123511 268127
rect 123393 267849 123511 267967
rect 123393 250009 123511 250127
rect 123393 249849 123511 249967
rect 123393 232009 123511 232127
rect 123393 231849 123511 231967
rect 123393 214009 123511 214127
rect 123393 213849 123511 213967
rect 123393 196009 123511 196127
rect 123393 195849 123511 195967
rect 123393 178009 123511 178127
rect 123393 177849 123511 177967
rect 123393 160009 123511 160127
rect 123393 159849 123511 159967
rect 123393 142009 123511 142127
rect 123393 141849 123511 141967
rect 123393 124009 123511 124127
rect 123393 123849 123511 123967
rect 123393 106009 123511 106127
rect 123393 105849 123511 105967
rect 123393 88009 123511 88127
rect 123393 87849 123511 87967
rect 123393 70009 123511 70127
rect 123393 69849 123511 69967
rect 123393 52009 123511 52127
rect 123393 51849 123511 51967
rect 123393 34009 123511 34127
rect 123393 33849 123511 33967
rect 123393 16009 123511 16127
rect 123393 15849 123511 15967
rect 114393 -3111 114511 -2993
rect 114393 -3271 114511 -3153
rect 126993 352301 127111 352419
rect 126993 352141 127111 352259
rect 126993 343609 127111 343727
rect 126993 343449 127111 343567
rect 126993 325609 127111 325727
rect 126993 325449 127111 325567
rect 126993 307609 127111 307727
rect 126993 307449 127111 307567
rect 126993 289609 127111 289727
rect 126993 289449 127111 289567
rect 126993 271609 127111 271727
rect 126993 271449 127111 271567
rect 126993 253609 127111 253727
rect 126993 253449 127111 253567
rect 126993 235609 127111 235727
rect 126993 235449 127111 235567
rect 126993 217609 127111 217727
rect 126993 217449 127111 217567
rect 126993 199609 127111 199727
rect 126993 199449 127111 199567
rect 126993 181609 127111 181727
rect 126993 181449 127111 181567
rect 126993 163609 127111 163727
rect 126993 163449 127111 163567
rect 126993 145609 127111 145727
rect 126993 145449 127111 145567
rect 126993 127609 127111 127727
rect 126993 127449 127111 127567
rect 126993 109609 127111 109727
rect 126993 109449 127111 109567
rect 126993 91609 127111 91727
rect 126993 91449 127111 91567
rect 126993 73609 127111 73727
rect 126993 73449 127111 73567
rect 126993 55609 127111 55727
rect 126993 55449 127111 55567
rect 126993 37609 127111 37727
rect 126993 37449 127111 37567
rect 126993 19609 127111 19727
rect 126993 19449 127111 19567
rect 126993 1609 127111 1727
rect 126993 1449 127111 1567
rect 126993 -291 127111 -173
rect 126993 -451 127111 -333
rect 128793 345409 128911 345527
rect 128793 345249 128911 345367
rect 128793 327409 128911 327527
rect 128793 327249 128911 327367
rect 128793 309409 128911 309527
rect 128793 309249 128911 309367
rect 128793 291409 128911 291527
rect 128793 291249 128911 291367
rect 128793 273409 128911 273527
rect 128793 273249 128911 273367
rect 128793 255409 128911 255527
rect 128793 255249 128911 255367
rect 128793 237409 128911 237527
rect 128793 237249 128911 237367
rect 128793 219409 128911 219527
rect 128793 219249 128911 219367
rect 128793 201409 128911 201527
rect 128793 201249 128911 201367
rect 128793 183409 128911 183527
rect 128793 183249 128911 183367
rect 128793 165409 128911 165527
rect 128793 165249 128911 165367
rect 128793 147409 128911 147527
rect 128793 147249 128911 147367
rect 128793 129409 128911 129527
rect 128793 129249 128911 129367
rect 128793 111409 128911 111527
rect 128793 111249 128911 111367
rect 128793 93409 128911 93527
rect 128793 93249 128911 93367
rect 128793 75409 128911 75527
rect 128793 75249 128911 75367
rect 128793 57409 128911 57527
rect 128793 57249 128911 57367
rect 128793 39409 128911 39527
rect 128793 39249 128911 39367
rect 128793 21409 128911 21527
rect 128793 21249 128911 21367
rect 128793 3409 128911 3527
rect 128793 3249 128911 3367
rect 128793 -1231 128911 -1113
rect 128793 -1391 128911 -1273
rect 130593 347209 130711 347327
rect 130593 347049 130711 347167
rect 130593 329209 130711 329327
rect 130593 329049 130711 329167
rect 130593 311209 130711 311327
rect 130593 311049 130711 311167
rect 130593 293209 130711 293327
rect 130593 293049 130711 293167
rect 130593 275209 130711 275327
rect 130593 275049 130711 275167
rect 130593 257209 130711 257327
rect 130593 257049 130711 257167
rect 130593 239209 130711 239327
rect 130593 239049 130711 239167
rect 130593 221209 130711 221327
rect 130593 221049 130711 221167
rect 130593 203209 130711 203327
rect 130593 203049 130711 203167
rect 130593 185209 130711 185327
rect 130593 185049 130711 185167
rect 130593 167209 130711 167327
rect 130593 167049 130711 167167
rect 130593 149209 130711 149327
rect 130593 149049 130711 149167
rect 130593 131209 130711 131327
rect 130593 131049 130711 131167
rect 130593 113209 130711 113327
rect 130593 113049 130711 113167
rect 130593 95209 130711 95327
rect 130593 95049 130711 95167
rect 130593 77209 130711 77327
rect 130593 77049 130711 77167
rect 130593 59209 130711 59327
rect 130593 59049 130711 59167
rect 130593 41209 130711 41327
rect 130593 41049 130711 41167
rect 130593 23209 130711 23327
rect 130593 23049 130711 23167
rect 130593 5209 130711 5327
rect 130593 5049 130711 5167
rect 130593 -2171 130711 -2053
rect 130593 -2331 130711 -2213
rect 141393 355591 141511 355709
rect 141393 355431 141511 355549
rect 139593 354651 139711 354769
rect 139593 354491 139711 354609
rect 137793 353711 137911 353829
rect 137793 353551 137911 353669
rect 132393 349009 132511 349127
rect 132393 348849 132511 348967
rect 132393 331009 132511 331127
rect 132393 330849 132511 330967
rect 132393 313009 132511 313127
rect 132393 312849 132511 312967
rect 132393 295009 132511 295127
rect 132393 294849 132511 294967
rect 132393 277009 132511 277127
rect 132393 276849 132511 276967
rect 132393 259009 132511 259127
rect 132393 258849 132511 258967
rect 132393 241009 132511 241127
rect 132393 240849 132511 240967
rect 132393 223009 132511 223127
rect 132393 222849 132511 222967
rect 132393 205009 132511 205127
rect 132393 204849 132511 204967
rect 132393 187009 132511 187127
rect 132393 186849 132511 186967
rect 132393 169009 132511 169127
rect 132393 168849 132511 168967
rect 132393 151009 132511 151127
rect 132393 150849 132511 150967
rect 132393 133009 132511 133127
rect 132393 132849 132511 132967
rect 132393 115009 132511 115127
rect 132393 114849 132511 114967
rect 132393 97009 132511 97127
rect 132393 96849 132511 96967
rect 132393 79009 132511 79127
rect 132393 78849 132511 78967
rect 132393 61009 132511 61127
rect 132393 60849 132511 60967
rect 132393 43009 132511 43127
rect 132393 42849 132511 42967
rect 132393 25009 132511 25127
rect 132393 24849 132511 24967
rect 132393 7009 132511 7127
rect 132393 6849 132511 6967
rect 123393 -3581 123511 -3463
rect 123393 -3741 123511 -3623
rect 135993 352771 136111 352889
rect 135993 352611 136111 352729
rect 135993 334609 136111 334727
rect 135993 334449 136111 334567
rect 135993 316609 136111 316727
rect 135993 316449 136111 316567
rect 135993 298609 136111 298727
rect 135993 298449 136111 298567
rect 135993 280609 136111 280727
rect 135993 280449 136111 280567
rect 135993 262609 136111 262727
rect 135993 262449 136111 262567
rect 135993 244609 136111 244727
rect 135993 244449 136111 244567
rect 135993 226609 136111 226727
rect 135993 226449 136111 226567
rect 135993 208609 136111 208727
rect 135993 208449 136111 208567
rect 135993 190609 136111 190727
rect 135993 190449 136111 190567
rect 135993 172609 136111 172727
rect 135993 172449 136111 172567
rect 135993 154609 136111 154727
rect 135993 154449 136111 154567
rect 135993 136609 136111 136727
rect 135993 136449 136111 136567
rect 135993 118609 136111 118727
rect 135993 118449 136111 118567
rect 135993 100609 136111 100727
rect 135993 100449 136111 100567
rect 135993 82609 136111 82727
rect 135993 82449 136111 82567
rect 135993 64609 136111 64727
rect 135993 64449 136111 64567
rect 135993 46609 136111 46727
rect 135993 46449 136111 46567
rect 135993 28609 136111 28727
rect 135993 28449 136111 28567
rect 135993 10609 136111 10727
rect 135993 10449 136111 10567
rect 135993 -761 136111 -643
rect 135993 -921 136111 -803
rect 137793 336409 137911 336527
rect 137793 336249 137911 336367
rect 137793 318409 137911 318527
rect 137793 318249 137911 318367
rect 137793 300409 137911 300527
rect 137793 300249 137911 300367
rect 137793 282409 137911 282527
rect 137793 282249 137911 282367
rect 137793 264409 137911 264527
rect 137793 264249 137911 264367
rect 137793 246409 137911 246527
rect 137793 246249 137911 246367
rect 137793 228409 137911 228527
rect 137793 228249 137911 228367
rect 137793 210409 137911 210527
rect 137793 210249 137911 210367
rect 137793 192409 137911 192527
rect 137793 192249 137911 192367
rect 137793 174409 137911 174527
rect 137793 174249 137911 174367
rect 137793 156409 137911 156527
rect 137793 156249 137911 156367
rect 137793 138409 137911 138527
rect 137793 138249 137911 138367
rect 137793 120409 137911 120527
rect 137793 120249 137911 120367
rect 137793 102409 137911 102527
rect 137793 102249 137911 102367
rect 137793 84409 137911 84527
rect 137793 84249 137911 84367
rect 137793 66409 137911 66527
rect 137793 66249 137911 66367
rect 137793 48409 137911 48527
rect 137793 48249 137911 48367
rect 137793 30409 137911 30527
rect 137793 30249 137911 30367
rect 137793 12409 137911 12527
rect 137793 12249 137911 12367
rect 137793 -1701 137911 -1583
rect 137793 -1861 137911 -1743
rect 139593 338209 139711 338327
rect 139593 338049 139711 338167
rect 139593 320209 139711 320327
rect 139593 320049 139711 320167
rect 139593 302209 139711 302327
rect 139593 302049 139711 302167
rect 139593 284209 139711 284327
rect 139593 284049 139711 284167
rect 139593 266209 139711 266327
rect 139593 266049 139711 266167
rect 139593 248209 139711 248327
rect 139593 248049 139711 248167
rect 139593 230209 139711 230327
rect 139593 230049 139711 230167
rect 139593 212209 139711 212327
rect 139593 212049 139711 212167
rect 139593 194209 139711 194327
rect 139593 194049 139711 194167
rect 139593 176209 139711 176327
rect 139593 176049 139711 176167
rect 139593 158209 139711 158327
rect 139593 158049 139711 158167
rect 139593 140209 139711 140327
rect 139593 140049 139711 140167
rect 139593 122209 139711 122327
rect 139593 122049 139711 122167
rect 139593 104209 139711 104327
rect 139593 104049 139711 104167
rect 139593 86209 139711 86327
rect 139593 86049 139711 86167
rect 139593 68209 139711 68327
rect 139593 68049 139711 68167
rect 139593 50209 139711 50327
rect 139593 50049 139711 50167
rect 139593 32209 139711 32327
rect 139593 32049 139711 32167
rect 139593 14209 139711 14327
rect 139593 14049 139711 14167
rect 139593 -2641 139711 -2523
rect 139593 -2801 139711 -2683
rect 150393 355121 150511 355239
rect 150393 354961 150511 355079
rect 148593 354181 148711 354299
rect 148593 354021 148711 354139
rect 146793 353241 146911 353359
rect 146793 353081 146911 353199
rect 141393 340009 141511 340127
rect 141393 339849 141511 339967
rect 141393 322009 141511 322127
rect 141393 321849 141511 321967
rect 141393 304009 141511 304127
rect 141393 303849 141511 303967
rect 141393 286009 141511 286127
rect 141393 285849 141511 285967
rect 141393 268009 141511 268127
rect 141393 267849 141511 267967
rect 141393 250009 141511 250127
rect 141393 249849 141511 249967
rect 141393 232009 141511 232127
rect 141393 231849 141511 231967
rect 141393 214009 141511 214127
rect 141393 213849 141511 213967
rect 141393 196009 141511 196127
rect 141393 195849 141511 195967
rect 141393 178009 141511 178127
rect 141393 177849 141511 177967
rect 141393 160009 141511 160127
rect 141393 159849 141511 159967
rect 141393 142009 141511 142127
rect 141393 141849 141511 141967
rect 141393 124009 141511 124127
rect 141393 123849 141511 123967
rect 141393 106009 141511 106127
rect 141393 105849 141511 105967
rect 141393 88009 141511 88127
rect 141393 87849 141511 87967
rect 141393 70009 141511 70127
rect 141393 69849 141511 69967
rect 141393 52009 141511 52127
rect 141393 51849 141511 51967
rect 141393 34009 141511 34127
rect 141393 33849 141511 33967
rect 141393 16009 141511 16127
rect 141393 15849 141511 15967
rect 132393 -3111 132511 -2993
rect 132393 -3271 132511 -3153
rect 144993 352301 145111 352419
rect 144993 352141 145111 352259
rect 144993 343609 145111 343727
rect 144993 343449 145111 343567
rect 144993 325609 145111 325727
rect 144993 325449 145111 325567
rect 144993 307609 145111 307727
rect 144993 307449 145111 307567
rect 144993 289609 145111 289727
rect 144993 289449 145111 289567
rect 144993 271609 145111 271727
rect 144993 271449 145111 271567
rect 144993 253609 145111 253727
rect 144993 253449 145111 253567
rect 144993 235609 145111 235727
rect 144993 235449 145111 235567
rect 144993 217609 145111 217727
rect 144993 217449 145111 217567
rect 144993 199609 145111 199727
rect 144993 199449 145111 199567
rect 144993 181609 145111 181727
rect 144993 181449 145111 181567
rect 144993 163609 145111 163727
rect 144993 163449 145111 163567
rect 144993 145609 145111 145727
rect 144993 145449 145111 145567
rect 144993 127609 145111 127727
rect 144993 127449 145111 127567
rect 144993 109609 145111 109727
rect 144993 109449 145111 109567
rect 144993 91609 145111 91727
rect 144993 91449 145111 91567
rect 144993 73609 145111 73727
rect 144993 73449 145111 73567
rect 144993 55609 145111 55727
rect 144993 55449 145111 55567
rect 144993 37609 145111 37727
rect 144993 37449 145111 37567
rect 144993 19609 145111 19727
rect 144993 19449 145111 19567
rect 144993 1609 145111 1727
rect 144993 1449 145111 1567
rect 144993 -291 145111 -173
rect 144993 -451 145111 -333
rect 146793 345409 146911 345527
rect 146793 345249 146911 345367
rect 146793 327409 146911 327527
rect 146793 327249 146911 327367
rect 146793 309409 146911 309527
rect 146793 309249 146911 309367
rect 146793 291409 146911 291527
rect 146793 291249 146911 291367
rect 146793 273409 146911 273527
rect 146793 273249 146911 273367
rect 146793 255409 146911 255527
rect 146793 255249 146911 255367
rect 146793 237409 146911 237527
rect 146793 237249 146911 237367
rect 146793 219409 146911 219527
rect 146793 219249 146911 219367
rect 146793 201409 146911 201527
rect 146793 201249 146911 201367
rect 146793 183409 146911 183527
rect 146793 183249 146911 183367
rect 146793 165409 146911 165527
rect 146793 165249 146911 165367
rect 146793 147409 146911 147527
rect 146793 147249 146911 147367
rect 146793 129409 146911 129527
rect 146793 129249 146911 129367
rect 146793 111409 146911 111527
rect 146793 111249 146911 111367
rect 146793 93409 146911 93527
rect 146793 93249 146911 93367
rect 146793 75409 146911 75527
rect 146793 75249 146911 75367
rect 146793 57409 146911 57527
rect 146793 57249 146911 57367
rect 146793 39409 146911 39527
rect 146793 39249 146911 39367
rect 146793 21409 146911 21527
rect 146793 21249 146911 21367
rect 146793 3409 146911 3527
rect 146793 3249 146911 3367
rect 146793 -1231 146911 -1113
rect 146793 -1391 146911 -1273
rect 148593 347209 148711 347327
rect 148593 347049 148711 347167
rect 148593 329209 148711 329327
rect 148593 329049 148711 329167
rect 148593 311209 148711 311327
rect 148593 311049 148711 311167
rect 148593 293209 148711 293327
rect 148593 293049 148711 293167
rect 148593 275209 148711 275327
rect 148593 275049 148711 275167
rect 148593 257209 148711 257327
rect 148593 257049 148711 257167
rect 148593 239209 148711 239327
rect 148593 239049 148711 239167
rect 148593 221209 148711 221327
rect 148593 221049 148711 221167
rect 148593 203209 148711 203327
rect 148593 203049 148711 203167
rect 148593 185209 148711 185327
rect 148593 185049 148711 185167
rect 148593 167209 148711 167327
rect 148593 167049 148711 167167
rect 148593 149209 148711 149327
rect 148593 149049 148711 149167
rect 148593 131209 148711 131327
rect 148593 131049 148711 131167
rect 148593 113209 148711 113327
rect 148593 113049 148711 113167
rect 148593 95209 148711 95327
rect 148593 95049 148711 95167
rect 148593 77209 148711 77327
rect 148593 77049 148711 77167
rect 148593 59209 148711 59327
rect 148593 59049 148711 59167
rect 148593 41209 148711 41327
rect 148593 41049 148711 41167
rect 148593 23209 148711 23327
rect 148593 23049 148711 23167
rect 148593 5209 148711 5327
rect 148593 5049 148711 5167
rect 148593 -2171 148711 -2053
rect 148593 -2331 148711 -2213
rect 159393 355591 159511 355709
rect 159393 355431 159511 355549
rect 157593 354651 157711 354769
rect 157593 354491 157711 354609
rect 155793 353711 155911 353829
rect 155793 353551 155911 353669
rect 150393 349009 150511 349127
rect 150393 348849 150511 348967
rect 150393 331009 150511 331127
rect 150393 330849 150511 330967
rect 150393 313009 150511 313127
rect 150393 312849 150511 312967
rect 150393 295009 150511 295127
rect 150393 294849 150511 294967
rect 150393 277009 150511 277127
rect 150393 276849 150511 276967
rect 150393 259009 150511 259127
rect 150393 258849 150511 258967
rect 150393 241009 150511 241127
rect 150393 240849 150511 240967
rect 150393 223009 150511 223127
rect 150393 222849 150511 222967
rect 150393 205009 150511 205127
rect 150393 204849 150511 204967
rect 150393 187009 150511 187127
rect 150393 186849 150511 186967
rect 150393 169009 150511 169127
rect 150393 168849 150511 168967
rect 150393 151009 150511 151127
rect 150393 150849 150511 150967
rect 150393 133009 150511 133127
rect 150393 132849 150511 132967
rect 150393 115009 150511 115127
rect 150393 114849 150511 114967
rect 150393 97009 150511 97127
rect 150393 96849 150511 96967
rect 150393 79009 150511 79127
rect 150393 78849 150511 78967
rect 150393 61009 150511 61127
rect 150393 60849 150511 60967
rect 150393 43009 150511 43127
rect 150393 42849 150511 42967
rect 150393 25009 150511 25127
rect 150393 24849 150511 24967
rect 150393 7009 150511 7127
rect 150393 6849 150511 6967
rect 141393 -3581 141511 -3463
rect 141393 -3741 141511 -3623
rect 153993 352771 154111 352889
rect 153993 352611 154111 352729
rect 153993 334609 154111 334727
rect 153993 334449 154111 334567
rect 153993 316609 154111 316727
rect 153993 316449 154111 316567
rect 153993 298609 154111 298727
rect 153993 298449 154111 298567
rect 153993 280609 154111 280727
rect 153993 280449 154111 280567
rect 153993 262609 154111 262727
rect 153993 262449 154111 262567
rect 153993 244609 154111 244727
rect 153993 244449 154111 244567
rect 153993 226609 154111 226727
rect 153993 226449 154111 226567
rect 153993 208609 154111 208727
rect 153993 208449 154111 208567
rect 153993 190609 154111 190727
rect 153993 190449 154111 190567
rect 153993 172609 154111 172727
rect 153993 172449 154111 172567
rect 153993 154609 154111 154727
rect 153993 154449 154111 154567
rect 153993 136609 154111 136727
rect 153993 136449 154111 136567
rect 153993 118609 154111 118727
rect 153993 118449 154111 118567
rect 153993 100609 154111 100727
rect 153993 100449 154111 100567
rect 153993 82609 154111 82727
rect 153993 82449 154111 82567
rect 153993 64609 154111 64727
rect 153993 64449 154111 64567
rect 153993 46609 154111 46727
rect 153993 46449 154111 46567
rect 153993 28609 154111 28727
rect 153993 28449 154111 28567
rect 153993 10609 154111 10727
rect 153993 10449 154111 10567
rect 153993 -761 154111 -643
rect 153993 -921 154111 -803
rect 155793 336409 155911 336527
rect 155793 336249 155911 336367
rect 155793 318409 155911 318527
rect 155793 318249 155911 318367
rect 155793 300409 155911 300527
rect 155793 300249 155911 300367
rect 155793 282409 155911 282527
rect 155793 282249 155911 282367
rect 155793 264409 155911 264527
rect 155793 264249 155911 264367
rect 155793 246409 155911 246527
rect 155793 246249 155911 246367
rect 155793 228409 155911 228527
rect 155793 228249 155911 228367
rect 155793 210409 155911 210527
rect 155793 210249 155911 210367
rect 155793 192409 155911 192527
rect 155793 192249 155911 192367
rect 155793 174409 155911 174527
rect 155793 174249 155911 174367
rect 155793 156409 155911 156527
rect 155793 156249 155911 156367
rect 155793 138409 155911 138527
rect 155793 138249 155911 138367
rect 155793 120409 155911 120527
rect 155793 120249 155911 120367
rect 155793 102409 155911 102527
rect 155793 102249 155911 102367
rect 155793 84409 155911 84527
rect 155793 84249 155911 84367
rect 155793 66409 155911 66527
rect 155793 66249 155911 66367
rect 155793 48409 155911 48527
rect 155793 48249 155911 48367
rect 155793 30409 155911 30527
rect 155793 30249 155911 30367
rect 155793 12409 155911 12527
rect 155793 12249 155911 12367
rect 155793 -1701 155911 -1583
rect 155793 -1861 155911 -1743
rect 157593 338209 157711 338327
rect 157593 338049 157711 338167
rect 157593 320209 157711 320327
rect 157593 320049 157711 320167
rect 157593 302209 157711 302327
rect 157593 302049 157711 302167
rect 157593 284209 157711 284327
rect 157593 284049 157711 284167
rect 157593 266209 157711 266327
rect 157593 266049 157711 266167
rect 157593 248209 157711 248327
rect 157593 248049 157711 248167
rect 157593 230209 157711 230327
rect 157593 230049 157711 230167
rect 157593 212209 157711 212327
rect 157593 212049 157711 212167
rect 157593 194209 157711 194327
rect 157593 194049 157711 194167
rect 157593 176209 157711 176327
rect 157593 176049 157711 176167
rect 157593 158209 157711 158327
rect 157593 158049 157711 158167
rect 157593 140209 157711 140327
rect 157593 140049 157711 140167
rect 157593 122209 157711 122327
rect 157593 122049 157711 122167
rect 157593 104209 157711 104327
rect 157593 104049 157711 104167
rect 157593 86209 157711 86327
rect 157593 86049 157711 86167
rect 157593 68209 157711 68327
rect 157593 68049 157711 68167
rect 157593 50209 157711 50327
rect 157593 50049 157711 50167
rect 157593 32209 157711 32327
rect 157593 32049 157711 32167
rect 157593 14209 157711 14327
rect 157593 14049 157711 14167
rect 157593 -2641 157711 -2523
rect 157593 -2801 157711 -2683
rect 168393 355121 168511 355239
rect 168393 354961 168511 355079
rect 166593 354181 166711 354299
rect 166593 354021 166711 354139
rect 164793 353241 164911 353359
rect 164793 353081 164911 353199
rect 159393 340009 159511 340127
rect 159393 339849 159511 339967
rect 159393 322009 159511 322127
rect 159393 321849 159511 321967
rect 159393 304009 159511 304127
rect 159393 303849 159511 303967
rect 159393 286009 159511 286127
rect 159393 285849 159511 285967
rect 159393 268009 159511 268127
rect 159393 267849 159511 267967
rect 159393 250009 159511 250127
rect 159393 249849 159511 249967
rect 159393 232009 159511 232127
rect 159393 231849 159511 231967
rect 159393 214009 159511 214127
rect 159393 213849 159511 213967
rect 159393 196009 159511 196127
rect 159393 195849 159511 195967
rect 159393 178009 159511 178127
rect 159393 177849 159511 177967
rect 159393 160009 159511 160127
rect 159393 159849 159511 159967
rect 159393 142009 159511 142127
rect 159393 141849 159511 141967
rect 159393 124009 159511 124127
rect 159393 123849 159511 123967
rect 159393 106009 159511 106127
rect 159393 105849 159511 105967
rect 159393 88009 159511 88127
rect 159393 87849 159511 87967
rect 159393 70009 159511 70127
rect 159393 69849 159511 69967
rect 159393 52009 159511 52127
rect 159393 51849 159511 51967
rect 159393 34009 159511 34127
rect 159393 33849 159511 33967
rect 159393 16009 159511 16127
rect 159393 15849 159511 15967
rect 150393 -3111 150511 -2993
rect 150393 -3271 150511 -3153
rect 162993 352301 163111 352419
rect 162993 352141 163111 352259
rect 162993 343609 163111 343727
rect 162993 343449 163111 343567
rect 162993 325609 163111 325727
rect 162993 325449 163111 325567
rect 162993 307609 163111 307727
rect 162993 307449 163111 307567
rect 162993 289609 163111 289727
rect 162993 289449 163111 289567
rect 162993 271609 163111 271727
rect 162993 271449 163111 271567
rect 162993 253609 163111 253727
rect 162993 253449 163111 253567
rect 162993 235609 163111 235727
rect 162993 235449 163111 235567
rect 162993 217609 163111 217727
rect 162993 217449 163111 217567
rect 162993 199609 163111 199727
rect 162993 199449 163111 199567
rect 162993 181609 163111 181727
rect 162993 181449 163111 181567
rect 162993 163609 163111 163727
rect 162993 163449 163111 163567
rect 162993 145609 163111 145727
rect 162993 145449 163111 145567
rect 162993 127609 163111 127727
rect 162993 127449 163111 127567
rect 162993 109609 163111 109727
rect 162993 109449 163111 109567
rect 162993 91609 163111 91727
rect 162993 91449 163111 91567
rect 162993 73609 163111 73727
rect 162993 73449 163111 73567
rect 162993 55609 163111 55727
rect 162993 55449 163111 55567
rect 162993 37609 163111 37727
rect 162993 37449 163111 37567
rect 162993 19609 163111 19727
rect 162993 19449 163111 19567
rect 162993 1609 163111 1727
rect 162993 1449 163111 1567
rect 162993 -291 163111 -173
rect 162993 -451 163111 -333
rect 164793 345409 164911 345527
rect 164793 345249 164911 345367
rect 164793 327409 164911 327527
rect 164793 327249 164911 327367
rect 164793 309409 164911 309527
rect 164793 309249 164911 309367
rect 164793 291409 164911 291527
rect 164793 291249 164911 291367
rect 164793 273409 164911 273527
rect 164793 273249 164911 273367
rect 164793 255409 164911 255527
rect 164793 255249 164911 255367
rect 164793 237409 164911 237527
rect 164793 237249 164911 237367
rect 164793 219409 164911 219527
rect 164793 219249 164911 219367
rect 164793 201409 164911 201527
rect 164793 201249 164911 201367
rect 164793 183409 164911 183527
rect 164793 183249 164911 183367
rect 164793 165409 164911 165527
rect 164793 165249 164911 165367
rect 164793 147409 164911 147527
rect 164793 147249 164911 147367
rect 164793 129409 164911 129527
rect 164793 129249 164911 129367
rect 164793 111409 164911 111527
rect 164793 111249 164911 111367
rect 164793 93409 164911 93527
rect 164793 93249 164911 93367
rect 164793 75409 164911 75527
rect 164793 75249 164911 75367
rect 164793 57409 164911 57527
rect 164793 57249 164911 57367
rect 164793 39409 164911 39527
rect 164793 39249 164911 39367
rect 164793 21409 164911 21527
rect 164793 21249 164911 21367
rect 164793 3409 164911 3527
rect 164793 3249 164911 3367
rect 164793 -1231 164911 -1113
rect 164793 -1391 164911 -1273
rect 166593 347209 166711 347327
rect 166593 347049 166711 347167
rect 166593 329209 166711 329327
rect 166593 329049 166711 329167
rect 166593 311209 166711 311327
rect 166593 311049 166711 311167
rect 166593 293209 166711 293327
rect 166593 293049 166711 293167
rect 166593 275209 166711 275327
rect 166593 275049 166711 275167
rect 166593 257209 166711 257327
rect 166593 257049 166711 257167
rect 166593 239209 166711 239327
rect 166593 239049 166711 239167
rect 166593 221209 166711 221327
rect 166593 221049 166711 221167
rect 166593 203209 166711 203327
rect 166593 203049 166711 203167
rect 166593 185209 166711 185327
rect 166593 185049 166711 185167
rect 166593 167209 166711 167327
rect 166593 167049 166711 167167
rect 166593 149209 166711 149327
rect 166593 149049 166711 149167
rect 166593 131209 166711 131327
rect 166593 131049 166711 131167
rect 166593 113209 166711 113327
rect 166593 113049 166711 113167
rect 166593 95209 166711 95327
rect 166593 95049 166711 95167
rect 166593 77209 166711 77327
rect 166593 77049 166711 77167
rect 166593 59209 166711 59327
rect 166593 59049 166711 59167
rect 166593 41209 166711 41327
rect 166593 41049 166711 41167
rect 166593 23209 166711 23327
rect 166593 23049 166711 23167
rect 166593 5209 166711 5327
rect 166593 5049 166711 5167
rect 166593 -2171 166711 -2053
rect 166593 -2331 166711 -2213
rect 177393 355591 177511 355709
rect 177393 355431 177511 355549
rect 175593 354651 175711 354769
rect 175593 354491 175711 354609
rect 173793 353711 173911 353829
rect 173793 353551 173911 353669
rect 168393 349009 168511 349127
rect 168393 348849 168511 348967
rect 168393 331009 168511 331127
rect 168393 330849 168511 330967
rect 168393 313009 168511 313127
rect 168393 312849 168511 312967
rect 168393 295009 168511 295127
rect 168393 294849 168511 294967
rect 168393 277009 168511 277127
rect 168393 276849 168511 276967
rect 168393 259009 168511 259127
rect 168393 258849 168511 258967
rect 168393 241009 168511 241127
rect 168393 240849 168511 240967
rect 168393 223009 168511 223127
rect 168393 222849 168511 222967
rect 168393 205009 168511 205127
rect 168393 204849 168511 204967
rect 168393 187009 168511 187127
rect 168393 186849 168511 186967
rect 168393 169009 168511 169127
rect 168393 168849 168511 168967
rect 168393 151009 168511 151127
rect 168393 150849 168511 150967
rect 168393 133009 168511 133127
rect 168393 132849 168511 132967
rect 168393 115009 168511 115127
rect 168393 114849 168511 114967
rect 168393 97009 168511 97127
rect 168393 96849 168511 96967
rect 168393 79009 168511 79127
rect 168393 78849 168511 78967
rect 168393 61009 168511 61127
rect 168393 60849 168511 60967
rect 168393 43009 168511 43127
rect 168393 42849 168511 42967
rect 168393 25009 168511 25127
rect 168393 24849 168511 24967
rect 168393 7009 168511 7127
rect 168393 6849 168511 6967
rect 159393 -3581 159511 -3463
rect 159393 -3741 159511 -3623
rect 171993 352771 172111 352889
rect 171993 352611 172111 352729
rect 171993 334609 172111 334727
rect 171993 334449 172111 334567
rect 171993 316609 172111 316727
rect 171993 316449 172111 316567
rect 171993 298609 172111 298727
rect 171993 298449 172111 298567
rect 171993 280609 172111 280727
rect 171993 280449 172111 280567
rect 171993 262609 172111 262727
rect 171993 262449 172111 262567
rect 171993 244609 172111 244727
rect 171993 244449 172111 244567
rect 171993 226609 172111 226727
rect 171993 226449 172111 226567
rect 171993 208609 172111 208727
rect 171993 208449 172111 208567
rect 171993 190609 172111 190727
rect 171993 190449 172111 190567
rect 171993 172609 172111 172727
rect 171993 172449 172111 172567
rect 171993 154609 172111 154727
rect 171993 154449 172111 154567
rect 171993 136609 172111 136727
rect 171993 136449 172111 136567
rect 171993 118609 172111 118727
rect 171993 118449 172111 118567
rect 171993 100609 172111 100727
rect 171993 100449 172111 100567
rect 171993 82609 172111 82727
rect 171993 82449 172111 82567
rect 171993 64609 172111 64727
rect 171993 64449 172111 64567
rect 171993 46609 172111 46727
rect 171993 46449 172111 46567
rect 171993 28609 172111 28727
rect 171993 28449 172111 28567
rect 171993 10609 172111 10727
rect 171993 10449 172111 10567
rect 171993 -761 172111 -643
rect 171993 -921 172111 -803
rect 173793 336409 173911 336527
rect 173793 336249 173911 336367
rect 173793 318409 173911 318527
rect 173793 318249 173911 318367
rect 173793 300409 173911 300527
rect 173793 300249 173911 300367
rect 173793 282409 173911 282527
rect 173793 282249 173911 282367
rect 173793 264409 173911 264527
rect 173793 264249 173911 264367
rect 173793 246409 173911 246527
rect 173793 246249 173911 246367
rect 173793 228409 173911 228527
rect 173793 228249 173911 228367
rect 173793 210409 173911 210527
rect 173793 210249 173911 210367
rect 173793 192409 173911 192527
rect 173793 192249 173911 192367
rect 173793 174409 173911 174527
rect 173793 174249 173911 174367
rect 173793 156409 173911 156527
rect 173793 156249 173911 156367
rect 173793 138409 173911 138527
rect 173793 138249 173911 138367
rect 173793 120409 173911 120527
rect 173793 120249 173911 120367
rect 173793 102409 173911 102527
rect 173793 102249 173911 102367
rect 173793 84409 173911 84527
rect 173793 84249 173911 84367
rect 173793 66409 173911 66527
rect 173793 66249 173911 66367
rect 173793 48409 173911 48527
rect 173793 48249 173911 48367
rect 173793 30409 173911 30527
rect 173793 30249 173911 30367
rect 173793 12409 173911 12527
rect 173793 12249 173911 12367
rect 173793 -1701 173911 -1583
rect 173793 -1861 173911 -1743
rect 175593 338209 175711 338327
rect 175593 338049 175711 338167
rect 175593 320209 175711 320327
rect 175593 320049 175711 320167
rect 175593 302209 175711 302327
rect 175593 302049 175711 302167
rect 175593 284209 175711 284327
rect 175593 284049 175711 284167
rect 175593 266209 175711 266327
rect 175593 266049 175711 266167
rect 175593 248209 175711 248327
rect 175593 248049 175711 248167
rect 175593 230209 175711 230327
rect 175593 230049 175711 230167
rect 175593 212209 175711 212327
rect 175593 212049 175711 212167
rect 175593 194209 175711 194327
rect 175593 194049 175711 194167
rect 175593 176209 175711 176327
rect 175593 176049 175711 176167
rect 175593 158209 175711 158327
rect 175593 158049 175711 158167
rect 175593 140209 175711 140327
rect 175593 140049 175711 140167
rect 175593 122209 175711 122327
rect 175593 122049 175711 122167
rect 175593 104209 175711 104327
rect 175593 104049 175711 104167
rect 175593 86209 175711 86327
rect 175593 86049 175711 86167
rect 175593 68209 175711 68327
rect 175593 68049 175711 68167
rect 175593 50209 175711 50327
rect 175593 50049 175711 50167
rect 175593 32209 175711 32327
rect 175593 32049 175711 32167
rect 175593 14209 175711 14327
rect 175593 14049 175711 14167
rect 175593 -2641 175711 -2523
rect 175593 -2801 175711 -2683
rect 186393 355121 186511 355239
rect 186393 354961 186511 355079
rect 184593 354181 184711 354299
rect 184593 354021 184711 354139
rect 182793 353241 182911 353359
rect 182793 353081 182911 353199
rect 177393 340009 177511 340127
rect 177393 339849 177511 339967
rect 177393 322009 177511 322127
rect 177393 321849 177511 321967
rect 177393 304009 177511 304127
rect 177393 303849 177511 303967
rect 177393 286009 177511 286127
rect 177393 285849 177511 285967
rect 177393 268009 177511 268127
rect 177393 267849 177511 267967
rect 177393 250009 177511 250127
rect 177393 249849 177511 249967
rect 177393 232009 177511 232127
rect 177393 231849 177511 231967
rect 177393 214009 177511 214127
rect 177393 213849 177511 213967
rect 177393 196009 177511 196127
rect 177393 195849 177511 195967
rect 177393 178009 177511 178127
rect 177393 177849 177511 177967
rect 177393 160009 177511 160127
rect 177393 159849 177511 159967
rect 177393 142009 177511 142127
rect 177393 141849 177511 141967
rect 177393 124009 177511 124127
rect 177393 123849 177511 123967
rect 177393 106009 177511 106127
rect 177393 105849 177511 105967
rect 177393 88009 177511 88127
rect 177393 87849 177511 87967
rect 177393 70009 177511 70127
rect 177393 69849 177511 69967
rect 177393 52009 177511 52127
rect 177393 51849 177511 51967
rect 177393 34009 177511 34127
rect 177393 33849 177511 33967
rect 177393 16009 177511 16127
rect 177393 15849 177511 15967
rect 168393 -3111 168511 -2993
rect 168393 -3271 168511 -3153
rect 180993 352301 181111 352419
rect 180993 352141 181111 352259
rect 180993 343609 181111 343727
rect 180993 343449 181111 343567
rect 180993 325609 181111 325727
rect 180993 325449 181111 325567
rect 180993 307609 181111 307727
rect 180993 307449 181111 307567
rect 180993 289609 181111 289727
rect 180993 289449 181111 289567
rect 180993 271609 181111 271727
rect 180993 271449 181111 271567
rect 180993 253609 181111 253727
rect 180993 253449 181111 253567
rect 180993 235609 181111 235727
rect 180993 235449 181111 235567
rect 180993 217609 181111 217727
rect 180993 217449 181111 217567
rect 180993 199609 181111 199727
rect 180993 199449 181111 199567
rect 180993 181609 181111 181727
rect 180993 181449 181111 181567
rect 180993 163609 181111 163727
rect 180993 163449 181111 163567
rect 180993 145609 181111 145727
rect 180993 145449 181111 145567
rect 180993 127609 181111 127727
rect 180993 127449 181111 127567
rect 180993 109609 181111 109727
rect 180993 109449 181111 109567
rect 180993 91609 181111 91727
rect 180993 91449 181111 91567
rect 180993 73609 181111 73727
rect 180993 73449 181111 73567
rect 180993 55609 181111 55727
rect 180993 55449 181111 55567
rect 180993 37609 181111 37727
rect 180993 37449 181111 37567
rect 180993 19609 181111 19727
rect 180993 19449 181111 19567
rect 180993 1609 181111 1727
rect 180993 1449 181111 1567
rect 180993 -291 181111 -173
rect 180993 -451 181111 -333
rect 182793 345409 182911 345527
rect 182793 345249 182911 345367
rect 182793 327409 182911 327527
rect 182793 327249 182911 327367
rect 182793 309409 182911 309527
rect 182793 309249 182911 309367
rect 182793 291409 182911 291527
rect 182793 291249 182911 291367
rect 182793 273409 182911 273527
rect 182793 273249 182911 273367
rect 182793 255409 182911 255527
rect 182793 255249 182911 255367
rect 182793 237409 182911 237527
rect 182793 237249 182911 237367
rect 182793 219409 182911 219527
rect 182793 219249 182911 219367
rect 182793 201409 182911 201527
rect 182793 201249 182911 201367
rect 182793 183409 182911 183527
rect 182793 183249 182911 183367
rect 182793 165409 182911 165527
rect 182793 165249 182911 165367
rect 182793 147409 182911 147527
rect 182793 147249 182911 147367
rect 182793 129409 182911 129527
rect 182793 129249 182911 129367
rect 182793 111409 182911 111527
rect 182793 111249 182911 111367
rect 182793 93409 182911 93527
rect 182793 93249 182911 93367
rect 182793 75409 182911 75527
rect 182793 75249 182911 75367
rect 182793 57409 182911 57527
rect 182793 57249 182911 57367
rect 182793 39409 182911 39527
rect 182793 39249 182911 39367
rect 182793 21409 182911 21527
rect 182793 21249 182911 21367
rect 182793 3409 182911 3527
rect 182793 3249 182911 3367
rect 182793 -1231 182911 -1113
rect 182793 -1391 182911 -1273
rect 184593 347209 184711 347327
rect 184593 347049 184711 347167
rect 184593 329209 184711 329327
rect 184593 329049 184711 329167
rect 184593 311209 184711 311327
rect 184593 311049 184711 311167
rect 184593 293209 184711 293327
rect 184593 293049 184711 293167
rect 184593 275209 184711 275327
rect 184593 275049 184711 275167
rect 184593 257209 184711 257327
rect 184593 257049 184711 257167
rect 184593 239209 184711 239327
rect 184593 239049 184711 239167
rect 184593 221209 184711 221327
rect 184593 221049 184711 221167
rect 184593 203209 184711 203327
rect 184593 203049 184711 203167
rect 184593 185209 184711 185327
rect 184593 185049 184711 185167
rect 184593 167209 184711 167327
rect 184593 167049 184711 167167
rect 184593 149209 184711 149327
rect 184593 149049 184711 149167
rect 184593 131209 184711 131327
rect 184593 131049 184711 131167
rect 184593 113209 184711 113327
rect 184593 113049 184711 113167
rect 184593 95209 184711 95327
rect 184593 95049 184711 95167
rect 184593 77209 184711 77327
rect 184593 77049 184711 77167
rect 184593 59209 184711 59327
rect 184593 59049 184711 59167
rect 184593 41209 184711 41327
rect 184593 41049 184711 41167
rect 184593 23209 184711 23327
rect 184593 23049 184711 23167
rect 184593 5209 184711 5327
rect 184593 5049 184711 5167
rect 184593 -2171 184711 -2053
rect 184593 -2331 184711 -2213
rect 195393 355591 195511 355709
rect 195393 355431 195511 355549
rect 193593 354651 193711 354769
rect 193593 354491 193711 354609
rect 191793 353711 191911 353829
rect 191793 353551 191911 353669
rect 186393 349009 186511 349127
rect 186393 348849 186511 348967
rect 186393 331009 186511 331127
rect 186393 330849 186511 330967
rect 186393 313009 186511 313127
rect 186393 312849 186511 312967
rect 186393 295009 186511 295127
rect 186393 294849 186511 294967
rect 186393 277009 186511 277127
rect 186393 276849 186511 276967
rect 186393 259009 186511 259127
rect 186393 258849 186511 258967
rect 186393 241009 186511 241127
rect 186393 240849 186511 240967
rect 186393 223009 186511 223127
rect 186393 222849 186511 222967
rect 186393 205009 186511 205127
rect 186393 204849 186511 204967
rect 186393 187009 186511 187127
rect 186393 186849 186511 186967
rect 186393 169009 186511 169127
rect 186393 168849 186511 168967
rect 186393 151009 186511 151127
rect 186393 150849 186511 150967
rect 186393 133009 186511 133127
rect 186393 132849 186511 132967
rect 186393 115009 186511 115127
rect 186393 114849 186511 114967
rect 186393 97009 186511 97127
rect 186393 96849 186511 96967
rect 186393 79009 186511 79127
rect 186393 78849 186511 78967
rect 186393 61009 186511 61127
rect 186393 60849 186511 60967
rect 186393 43009 186511 43127
rect 186393 42849 186511 42967
rect 186393 25009 186511 25127
rect 186393 24849 186511 24967
rect 186393 7009 186511 7127
rect 186393 6849 186511 6967
rect 177393 -3581 177511 -3463
rect 177393 -3741 177511 -3623
rect 189993 352771 190111 352889
rect 189993 352611 190111 352729
rect 189993 334609 190111 334727
rect 189993 334449 190111 334567
rect 189993 316609 190111 316727
rect 189993 316449 190111 316567
rect 189993 298609 190111 298727
rect 189993 298449 190111 298567
rect 189993 280609 190111 280727
rect 189993 280449 190111 280567
rect 189993 262609 190111 262727
rect 189993 262449 190111 262567
rect 189993 244609 190111 244727
rect 189993 244449 190111 244567
rect 189993 226609 190111 226727
rect 189993 226449 190111 226567
rect 189993 208609 190111 208727
rect 189993 208449 190111 208567
rect 189993 190609 190111 190727
rect 189993 190449 190111 190567
rect 189993 172609 190111 172727
rect 189993 172449 190111 172567
rect 189993 154609 190111 154727
rect 189993 154449 190111 154567
rect 189993 136609 190111 136727
rect 189993 136449 190111 136567
rect 189993 118609 190111 118727
rect 189993 118449 190111 118567
rect 189993 100609 190111 100727
rect 189993 100449 190111 100567
rect 189993 82609 190111 82727
rect 189993 82449 190111 82567
rect 189993 64609 190111 64727
rect 189993 64449 190111 64567
rect 189993 46609 190111 46727
rect 189993 46449 190111 46567
rect 189993 28609 190111 28727
rect 189993 28449 190111 28567
rect 189993 10609 190111 10727
rect 189993 10449 190111 10567
rect 189993 -761 190111 -643
rect 189993 -921 190111 -803
rect 191793 336409 191911 336527
rect 191793 336249 191911 336367
rect 191793 318409 191911 318527
rect 191793 318249 191911 318367
rect 191793 300409 191911 300527
rect 191793 300249 191911 300367
rect 191793 282409 191911 282527
rect 191793 282249 191911 282367
rect 191793 264409 191911 264527
rect 191793 264249 191911 264367
rect 191793 246409 191911 246527
rect 191793 246249 191911 246367
rect 191793 228409 191911 228527
rect 191793 228249 191911 228367
rect 191793 210409 191911 210527
rect 191793 210249 191911 210367
rect 191793 192409 191911 192527
rect 191793 192249 191911 192367
rect 191793 174409 191911 174527
rect 191793 174249 191911 174367
rect 191793 156409 191911 156527
rect 191793 156249 191911 156367
rect 191793 138409 191911 138527
rect 191793 138249 191911 138367
rect 191793 120409 191911 120527
rect 191793 120249 191911 120367
rect 191793 102409 191911 102527
rect 191793 102249 191911 102367
rect 191793 84409 191911 84527
rect 191793 84249 191911 84367
rect 191793 66409 191911 66527
rect 191793 66249 191911 66367
rect 191793 48409 191911 48527
rect 191793 48249 191911 48367
rect 191793 30409 191911 30527
rect 191793 30249 191911 30367
rect 191793 12409 191911 12527
rect 191793 12249 191911 12367
rect 191793 -1701 191911 -1583
rect 191793 -1861 191911 -1743
rect 193593 338209 193711 338327
rect 193593 338049 193711 338167
rect 193593 320209 193711 320327
rect 193593 320049 193711 320167
rect 193593 302209 193711 302327
rect 193593 302049 193711 302167
rect 193593 284209 193711 284327
rect 193593 284049 193711 284167
rect 193593 266209 193711 266327
rect 193593 266049 193711 266167
rect 193593 248209 193711 248327
rect 193593 248049 193711 248167
rect 193593 230209 193711 230327
rect 193593 230049 193711 230167
rect 193593 212209 193711 212327
rect 193593 212049 193711 212167
rect 193593 194209 193711 194327
rect 193593 194049 193711 194167
rect 193593 176209 193711 176327
rect 193593 176049 193711 176167
rect 193593 158209 193711 158327
rect 193593 158049 193711 158167
rect 193593 140209 193711 140327
rect 193593 140049 193711 140167
rect 193593 122209 193711 122327
rect 193593 122049 193711 122167
rect 193593 104209 193711 104327
rect 193593 104049 193711 104167
rect 193593 86209 193711 86327
rect 193593 86049 193711 86167
rect 193593 68209 193711 68327
rect 193593 68049 193711 68167
rect 193593 50209 193711 50327
rect 193593 50049 193711 50167
rect 193593 32209 193711 32327
rect 193593 32049 193711 32167
rect 193593 14209 193711 14327
rect 193593 14049 193711 14167
rect 193593 -2641 193711 -2523
rect 193593 -2801 193711 -2683
rect 204393 355121 204511 355239
rect 204393 354961 204511 355079
rect 202593 354181 202711 354299
rect 202593 354021 202711 354139
rect 200793 353241 200911 353359
rect 200793 353081 200911 353199
rect 195393 340009 195511 340127
rect 195393 339849 195511 339967
rect 195393 322009 195511 322127
rect 195393 321849 195511 321967
rect 195393 304009 195511 304127
rect 195393 303849 195511 303967
rect 195393 286009 195511 286127
rect 195393 285849 195511 285967
rect 195393 268009 195511 268127
rect 195393 267849 195511 267967
rect 195393 250009 195511 250127
rect 195393 249849 195511 249967
rect 195393 232009 195511 232127
rect 195393 231849 195511 231967
rect 195393 214009 195511 214127
rect 195393 213849 195511 213967
rect 195393 196009 195511 196127
rect 195393 195849 195511 195967
rect 195393 178009 195511 178127
rect 195393 177849 195511 177967
rect 195393 160009 195511 160127
rect 195393 159849 195511 159967
rect 195393 142009 195511 142127
rect 195393 141849 195511 141967
rect 195393 124009 195511 124127
rect 195393 123849 195511 123967
rect 195393 106009 195511 106127
rect 195393 105849 195511 105967
rect 195393 88009 195511 88127
rect 195393 87849 195511 87967
rect 195393 70009 195511 70127
rect 195393 69849 195511 69967
rect 195393 52009 195511 52127
rect 195393 51849 195511 51967
rect 195393 34009 195511 34127
rect 195393 33849 195511 33967
rect 195393 16009 195511 16127
rect 195393 15849 195511 15967
rect 186393 -3111 186511 -2993
rect 186393 -3271 186511 -3153
rect 198993 352301 199111 352419
rect 198993 352141 199111 352259
rect 198993 343609 199111 343727
rect 198993 343449 199111 343567
rect 198993 325609 199111 325727
rect 198993 325449 199111 325567
rect 198993 307609 199111 307727
rect 198993 307449 199111 307567
rect 198993 289609 199111 289727
rect 198993 289449 199111 289567
rect 198993 271609 199111 271727
rect 198993 271449 199111 271567
rect 198993 253609 199111 253727
rect 198993 253449 199111 253567
rect 198993 235609 199111 235727
rect 198993 235449 199111 235567
rect 198993 217609 199111 217727
rect 198993 217449 199111 217567
rect 198993 199609 199111 199727
rect 198993 199449 199111 199567
rect 198993 181609 199111 181727
rect 198993 181449 199111 181567
rect 198993 163609 199111 163727
rect 198993 163449 199111 163567
rect 198993 145609 199111 145727
rect 198993 145449 199111 145567
rect 198993 127609 199111 127727
rect 198993 127449 199111 127567
rect 198993 109609 199111 109727
rect 198993 109449 199111 109567
rect 198993 91609 199111 91727
rect 198993 91449 199111 91567
rect 198993 73609 199111 73727
rect 198993 73449 199111 73567
rect 198993 55609 199111 55727
rect 198993 55449 199111 55567
rect 198993 37609 199111 37727
rect 198993 37449 199111 37567
rect 198993 19609 199111 19727
rect 198993 19449 199111 19567
rect 198993 1609 199111 1727
rect 198993 1449 199111 1567
rect 198993 -291 199111 -173
rect 198993 -451 199111 -333
rect 200793 345409 200911 345527
rect 200793 345249 200911 345367
rect 200793 327409 200911 327527
rect 200793 327249 200911 327367
rect 200793 309409 200911 309527
rect 200793 309249 200911 309367
rect 200793 291409 200911 291527
rect 200793 291249 200911 291367
rect 200793 273409 200911 273527
rect 200793 273249 200911 273367
rect 200793 255409 200911 255527
rect 200793 255249 200911 255367
rect 200793 237409 200911 237527
rect 200793 237249 200911 237367
rect 200793 219409 200911 219527
rect 200793 219249 200911 219367
rect 200793 201409 200911 201527
rect 200793 201249 200911 201367
rect 200793 183409 200911 183527
rect 200793 183249 200911 183367
rect 200793 165409 200911 165527
rect 200793 165249 200911 165367
rect 200793 147409 200911 147527
rect 200793 147249 200911 147367
rect 200793 129409 200911 129527
rect 200793 129249 200911 129367
rect 200793 111409 200911 111527
rect 200793 111249 200911 111367
rect 200793 93409 200911 93527
rect 200793 93249 200911 93367
rect 200793 75409 200911 75527
rect 200793 75249 200911 75367
rect 200793 57409 200911 57527
rect 200793 57249 200911 57367
rect 200793 39409 200911 39527
rect 200793 39249 200911 39367
rect 200793 21409 200911 21527
rect 200793 21249 200911 21367
rect 200793 3409 200911 3527
rect 200793 3249 200911 3367
rect 200793 -1231 200911 -1113
rect 200793 -1391 200911 -1273
rect 202593 347209 202711 347327
rect 202593 347049 202711 347167
rect 202593 329209 202711 329327
rect 202593 329049 202711 329167
rect 202593 311209 202711 311327
rect 202593 311049 202711 311167
rect 202593 293209 202711 293327
rect 202593 293049 202711 293167
rect 202593 275209 202711 275327
rect 202593 275049 202711 275167
rect 202593 257209 202711 257327
rect 202593 257049 202711 257167
rect 202593 239209 202711 239327
rect 202593 239049 202711 239167
rect 202593 221209 202711 221327
rect 202593 221049 202711 221167
rect 202593 203209 202711 203327
rect 202593 203049 202711 203167
rect 202593 185209 202711 185327
rect 202593 185049 202711 185167
rect 202593 167209 202711 167327
rect 202593 167049 202711 167167
rect 202593 149209 202711 149327
rect 202593 149049 202711 149167
rect 202593 131209 202711 131327
rect 202593 131049 202711 131167
rect 202593 113209 202711 113327
rect 202593 113049 202711 113167
rect 202593 95209 202711 95327
rect 202593 95049 202711 95167
rect 202593 77209 202711 77327
rect 202593 77049 202711 77167
rect 202593 59209 202711 59327
rect 202593 59049 202711 59167
rect 202593 41209 202711 41327
rect 202593 41049 202711 41167
rect 202593 23209 202711 23327
rect 202593 23049 202711 23167
rect 202593 5209 202711 5327
rect 202593 5049 202711 5167
rect 202593 -2171 202711 -2053
rect 202593 -2331 202711 -2213
rect 213393 355591 213511 355709
rect 213393 355431 213511 355549
rect 211593 354651 211711 354769
rect 211593 354491 211711 354609
rect 209793 353711 209911 353829
rect 209793 353551 209911 353669
rect 204393 349009 204511 349127
rect 204393 348849 204511 348967
rect 204393 331009 204511 331127
rect 204393 330849 204511 330967
rect 204393 313009 204511 313127
rect 204393 312849 204511 312967
rect 204393 295009 204511 295127
rect 204393 294849 204511 294967
rect 204393 277009 204511 277127
rect 204393 276849 204511 276967
rect 204393 259009 204511 259127
rect 204393 258849 204511 258967
rect 204393 241009 204511 241127
rect 204393 240849 204511 240967
rect 204393 223009 204511 223127
rect 204393 222849 204511 222967
rect 204393 205009 204511 205127
rect 204393 204849 204511 204967
rect 204393 187009 204511 187127
rect 204393 186849 204511 186967
rect 204393 169009 204511 169127
rect 204393 168849 204511 168967
rect 204393 151009 204511 151127
rect 204393 150849 204511 150967
rect 204393 133009 204511 133127
rect 204393 132849 204511 132967
rect 204393 115009 204511 115127
rect 204393 114849 204511 114967
rect 204393 97009 204511 97127
rect 204393 96849 204511 96967
rect 204393 79009 204511 79127
rect 204393 78849 204511 78967
rect 204393 61009 204511 61127
rect 204393 60849 204511 60967
rect 204393 43009 204511 43127
rect 204393 42849 204511 42967
rect 204393 25009 204511 25127
rect 204393 24849 204511 24967
rect 204393 7009 204511 7127
rect 204393 6849 204511 6967
rect 195393 -3581 195511 -3463
rect 195393 -3741 195511 -3623
rect 207993 352771 208111 352889
rect 207993 352611 208111 352729
rect 207993 334609 208111 334727
rect 207993 334449 208111 334567
rect 207993 316609 208111 316727
rect 207993 316449 208111 316567
rect 207993 298609 208111 298727
rect 207993 298449 208111 298567
rect 207993 280609 208111 280727
rect 207993 280449 208111 280567
rect 207993 262609 208111 262727
rect 207993 262449 208111 262567
rect 207993 244609 208111 244727
rect 207993 244449 208111 244567
rect 207993 226609 208111 226727
rect 207993 226449 208111 226567
rect 207993 208609 208111 208727
rect 207993 208449 208111 208567
rect 207993 190609 208111 190727
rect 207993 190449 208111 190567
rect 207993 172609 208111 172727
rect 207993 172449 208111 172567
rect 207993 154609 208111 154727
rect 207993 154449 208111 154567
rect 207993 136609 208111 136727
rect 207993 136449 208111 136567
rect 207993 118609 208111 118727
rect 207993 118449 208111 118567
rect 207993 100609 208111 100727
rect 207993 100449 208111 100567
rect 207993 82609 208111 82727
rect 207993 82449 208111 82567
rect 207993 64609 208111 64727
rect 207993 64449 208111 64567
rect 207993 46609 208111 46727
rect 207993 46449 208111 46567
rect 207993 28609 208111 28727
rect 207993 28449 208111 28567
rect 207993 10609 208111 10727
rect 207993 10449 208111 10567
rect 207993 -761 208111 -643
rect 207993 -921 208111 -803
rect 209793 336409 209911 336527
rect 209793 336249 209911 336367
rect 209793 318409 209911 318527
rect 209793 318249 209911 318367
rect 209793 300409 209911 300527
rect 209793 300249 209911 300367
rect 209793 282409 209911 282527
rect 209793 282249 209911 282367
rect 209793 264409 209911 264527
rect 209793 264249 209911 264367
rect 209793 246409 209911 246527
rect 209793 246249 209911 246367
rect 209793 228409 209911 228527
rect 209793 228249 209911 228367
rect 209793 210409 209911 210527
rect 209793 210249 209911 210367
rect 209793 192409 209911 192527
rect 209793 192249 209911 192367
rect 209793 174409 209911 174527
rect 209793 174249 209911 174367
rect 209793 156409 209911 156527
rect 209793 156249 209911 156367
rect 209793 138409 209911 138527
rect 209793 138249 209911 138367
rect 209793 120409 209911 120527
rect 209793 120249 209911 120367
rect 209793 102409 209911 102527
rect 209793 102249 209911 102367
rect 209793 84409 209911 84527
rect 209793 84249 209911 84367
rect 209793 66409 209911 66527
rect 209793 66249 209911 66367
rect 209793 48409 209911 48527
rect 209793 48249 209911 48367
rect 209793 30409 209911 30527
rect 209793 30249 209911 30367
rect 209793 12409 209911 12527
rect 209793 12249 209911 12367
rect 209793 -1701 209911 -1583
rect 209793 -1861 209911 -1743
rect 211593 338209 211711 338327
rect 211593 338049 211711 338167
rect 211593 320209 211711 320327
rect 211593 320049 211711 320167
rect 211593 302209 211711 302327
rect 211593 302049 211711 302167
rect 211593 284209 211711 284327
rect 211593 284049 211711 284167
rect 211593 266209 211711 266327
rect 211593 266049 211711 266167
rect 211593 248209 211711 248327
rect 211593 248049 211711 248167
rect 211593 230209 211711 230327
rect 211593 230049 211711 230167
rect 211593 212209 211711 212327
rect 211593 212049 211711 212167
rect 211593 194209 211711 194327
rect 211593 194049 211711 194167
rect 211593 176209 211711 176327
rect 211593 176049 211711 176167
rect 211593 158209 211711 158327
rect 211593 158049 211711 158167
rect 211593 140209 211711 140327
rect 211593 140049 211711 140167
rect 211593 122209 211711 122327
rect 211593 122049 211711 122167
rect 211593 104209 211711 104327
rect 211593 104049 211711 104167
rect 211593 86209 211711 86327
rect 211593 86049 211711 86167
rect 211593 68209 211711 68327
rect 211593 68049 211711 68167
rect 211593 50209 211711 50327
rect 211593 50049 211711 50167
rect 211593 32209 211711 32327
rect 211593 32049 211711 32167
rect 211593 14209 211711 14327
rect 211593 14049 211711 14167
rect 211593 -2641 211711 -2523
rect 211593 -2801 211711 -2683
rect 222393 355121 222511 355239
rect 222393 354961 222511 355079
rect 220593 354181 220711 354299
rect 220593 354021 220711 354139
rect 218793 353241 218911 353359
rect 218793 353081 218911 353199
rect 213393 340009 213511 340127
rect 213393 339849 213511 339967
rect 213393 322009 213511 322127
rect 213393 321849 213511 321967
rect 213393 304009 213511 304127
rect 213393 303849 213511 303967
rect 213393 286009 213511 286127
rect 213393 285849 213511 285967
rect 213393 268009 213511 268127
rect 213393 267849 213511 267967
rect 213393 250009 213511 250127
rect 213393 249849 213511 249967
rect 213393 232009 213511 232127
rect 213393 231849 213511 231967
rect 213393 214009 213511 214127
rect 213393 213849 213511 213967
rect 213393 196009 213511 196127
rect 213393 195849 213511 195967
rect 213393 178009 213511 178127
rect 213393 177849 213511 177967
rect 213393 160009 213511 160127
rect 213393 159849 213511 159967
rect 213393 142009 213511 142127
rect 213393 141849 213511 141967
rect 213393 124009 213511 124127
rect 213393 123849 213511 123967
rect 213393 106009 213511 106127
rect 213393 105849 213511 105967
rect 213393 88009 213511 88127
rect 213393 87849 213511 87967
rect 213393 70009 213511 70127
rect 213393 69849 213511 69967
rect 213393 52009 213511 52127
rect 213393 51849 213511 51967
rect 213393 34009 213511 34127
rect 213393 33849 213511 33967
rect 213393 16009 213511 16127
rect 213393 15849 213511 15967
rect 204393 -3111 204511 -2993
rect 204393 -3271 204511 -3153
rect 216993 352301 217111 352419
rect 216993 352141 217111 352259
rect 216993 343609 217111 343727
rect 216993 343449 217111 343567
rect 216993 325609 217111 325727
rect 216993 325449 217111 325567
rect 216993 307609 217111 307727
rect 216993 307449 217111 307567
rect 216993 289609 217111 289727
rect 216993 289449 217111 289567
rect 216993 271609 217111 271727
rect 216993 271449 217111 271567
rect 216993 253609 217111 253727
rect 216993 253449 217111 253567
rect 216993 235609 217111 235727
rect 216993 235449 217111 235567
rect 216993 217609 217111 217727
rect 216993 217449 217111 217567
rect 216993 199609 217111 199727
rect 216993 199449 217111 199567
rect 216993 181609 217111 181727
rect 216993 181449 217111 181567
rect 216993 163609 217111 163727
rect 216993 163449 217111 163567
rect 216993 145609 217111 145727
rect 216993 145449 217111 145567
rect 216993 127609 217111 127727
rect 216993 127449 217111 127567
rect 216993 109609 217111 109727
rect 216993 109449 217111 109567
rect 216993 91609 217111 91727
rect 216993 91449 217111 91567
rect 216993 73609 217111 73727
rect 216993 73449 217111 73567
rect 216993 55609 217111 55727
rect 216993 55449 217111 55567
rect 216993 37609 217111 37727
rect 216993 37449 217111 37567
rect 216993 19609 217111 19727
rect 216993 19449 217111 19567
rect 216993 1609 217111 1727
rect 216993 1449 217111 1567
rect 216993 -291 217111 -173
rect 216993 -451 217111 -333
rect 218793 345409 218911 345527
rect 218793 345249 218911 345367
rect 218793 327409 218911 327527
rect 218793 327249 218911 327367
rect 218793 309409 218911 309527
rect 218793 309249 218911 309367
rect 218793 291409 218911 291527
rect 218793 291249 218911 291367
rect 218793 273409 218911 273527
rect 218793 273249 218911 273367
rect 218793 255409 218911 255527
rect 218793 255249 218911 255367
rect 218793 237409 218911 237527
rect 218793 237249 218911 237367
rect 218793 219409 218911 219527
rect 218793 219249 218911 219367
rect 218793 201409 218911 201527
rect 218793 201249 218911 201367
rect 218793 183409 218911 183527
rect 218793 183249 218911 183367
rect 218793 165409 218911 165527
rect 218793 165249 218911 165367
rect 218793 147409 218911 147527
rect 218793 147249 218911 147367
rect 218793 129409 218911 129527
rect 218793 129249 218911 129367
rect 218793 111409 218911 111527
rect 218793 111249 218911 111367
rect 218793 93409 218911 93527
rect 218793 93249 218911 93367
rect 218793 75409 218911 75527
rect 218793 75249 218911 75367
rect 218793 57409 218911 57527
rect 218793 57249 218911 57367
rect 218793 39409 218911 39527
rect 218793 39249 218911 39367
rect 218793 21409 218911 21527
rect 218793 21249 218911 21367
rect 218793 3409 218911 3527
rect 218793 3249 218911 3367
rect 218793 -1231 218911 -1113
rect 218793 -1391 218911 -1273
rect 220593 347209 220711 347327
rect 220593 347049 220711 347167
rect 220593 329209 220711 329327
rect 220593 329049 220711 329167
rect 220593 311209 220711 311327
rect 220593 311049 220711 311167
rect 220593 293209 220711 293327
rect 220593 293049 220711 293167
rect 220593 275209 220711 275327
rect 220593 275049 220711 275167
rect 220593 257209 220711 257327
rect 220593 257049 220711 257167
rect 220593 239209 220711 239327
rect 220593 239049 220711 239167
rect 220593 221209 220711 221327
rect 220593 221049 220711 221167
rect 220593 203209 220711 203327
rect 220593 203049 220711 203167
rect 220593 185209 220711 185327
rect 220593 185049 220711 185167
rect 220593 167209 220711 167327
rect 220593 167049 220711 167167
rect 220593 149209 220711 149327
rect 220593 149049 220711 149167
rect 220593 131209 220711 131327
rect 220593 131049 220711 131167
rect 220593 113209 220711 113327
rect 220593 113049 220711 113167
rect 220593 95209 220711 95327
rect 220593 95049 220711 95167
rect 220593 77209 220711 77327
rect 220593 77049 220711 77167
rect 220593 59209 220711 59327
rect 220593 59049 220711 59167
rect 220593 41209 220711 41327
rect 220593 41049 220711 41167
rect 220593 23209 220711 23327
rect 220593 23049 220711 23167
rect 220593 5209 220711 5327
rect 220593 5049 220711 5167
rect 220593 -2171 220711 -2053
rect 220593 -2331 220711 -2213
rect 231393 355591 231511 355709
rect 231393 355431 231511 355549
rect 229593 354651 229711 354769
rect 229593 354491 229711 354609
rect 227793 353711 227911 353829
rect 227793 353551 227911 353669
rect 222393 349009 222511 349127
rect 222393 348849 222511 348967
rect 222393 331009 222511 331127
rect 222393 330849 222511 330967
rect 222393 313009 222511 313127
rect 222393 312849 222511 312967
rect 222393 295009 222511 295127
rect 222393 294849 222511 294967
rect 222393 277009 222511 277127
rect 222393 276849 222511 276967
rect 222393 259009 222511 259127
rect 222393 258849 222511 258967
rect 222393 241009 222511 241127
rect 222393 240849 222511 240967
rect 222393 223009 222511 223127
rect 222393 222849 222511 222967
rect 222393 205009 222511 205127
rect 222393 204849 222511 204967
rect 222393 187009 222511 187127
rect 222393 186849 222511 186967
rect 222393 169009 222511 169127
rect 222393 168849 222511 168967
rect 222393 151009 222511 151127
rect 222393 150849 222511 150967
rect 222393 133009 222511 133127
rect 222393 132849 222511 132967
rect 222393 115009 222511 115127
rect 222393 114849 222511 114967
rect 222393 97009 222511 97127
rect 222393 96849 222511 96967
rect 222393 79009 222511 79127
rect 222393 78849 222511 78967
rect 222393 61009 222511 61127
rect 222393 60849 222511 60967
rect 222393 43009 222511 43127
rect 222393 42849 222511 42967
rect 222393 25009 222511 25127
rect 222393 24849 222511 24967
rect 222393 7009 222511 7127
rect 222393 6849 222511 6967
rect 213393 -3581 213511 -3463
rect 213393 -3741 213511 -3623
rect 225993 352771 226111 352889
rect 225993 352611 226111 352729
rect 225993 334609 226111 334727
rect 225993 334449 226111 334567
rect 225993 316609 226111 316727
rect 225993 316449 226111 316567
rect 225993 298609 226111 298727
rect 225993 298449 226111 298567
rect 225993 280609 226111 280727
rect 225993 280449 226111 280567
rect 225993 262609 226111 262727
rect 225993 262449 226111 262567
rect 225993 244609 226111 244727
rect 225993 244449 226111 244567
rect 225993 226609 226111 226727
rect 225993 226449 226111 226567
rect 225993 208609 226111 208727
rect 225993 208449 226111 208567
rect 225993 190609 226111 190727
rect 225993 190449 226111 190567
rect 225993 172609 226111 172727
rect 225993 172449 226111 172567
rect 225993 154609 226111 154727
rect 225993 154449 226111 154567
rect 225993 136609 226111 136727
rect 225993 136449 226111 136567
rect 225993 118609 226111 118727
rect 225993 118449 226111 118567
rect 225993 100609 226111 100727
rect 225993 100449 226111 100567
rect 225993 82609 226111 82727
rect 225993 82449 226111 82567
rect 225993 64609 226111 64727
rect 225993 64449 226111 64567
rect 225993 46609 226111 46727
rect 225993 46449 226111 46567
rect 225993 28609 226111 28727
rect 225993 28449 226111 28567
rect 225993 10609 226111 10727
rect 225993 10449 226111 10567
rect 225993 -761 226111 -643
rect 225993 -921 226111 -803
rect 227793 336409 227911 336527
rect 227793 336249 227911 336367
rect 227793 318409 227911 318527
rect 227793 318249 227911 318367
rect 227793 300409 227911 300527
rect 227793 300249 227911 300367
rect 227793 282409 227911 282527
rect 227793 282249 227911 282367
rect 227793 264409 227911 264527
rect 227793 264249 227911 264367
rect 227793 246409 227911 246527
rect 227793 246249 227911 246367
rect 227793 228409 227911 228527
rect 227793 228249 227911 228367
rect 227793 210409 227911 210527
rect 227793 210249 227911 210367
rect 227793 192409 227911 192527
rect 227793 192249 227911 192367
rect 227793 174409 227911 174527
rect 227793 174249 227911 174367
rect 227793 156409 227911 156527
rect 227793 156249 227911 156367
rect 227793 138409 227911 138527
rect 227793 138249 227911 138367
rect 227793 120409 227911 120527
rect 227793 120249 227911 120367
rect 227793 102409 227911 102527
rect 227793 102249 227911 102367
rect 227793 84409 227911 84527
rect 227793 84249 227911 84367
rect 227793 66409 227911 66527
rect 227793 66249 227911 66367
rect 227793 48409 227911 48527
rect 227793 48249 227911 48367
rect 227793 30409 227911 30527
rect 227793 30249 227911 30367
rect 227793 12409 227911 12527
rect 227793 12249 227911 12367
rect 227793 -1701 227911 -1583
rect 227793 -1861 227911 -1743
rect 229593 338209 229711 338327
rect 229593 338049 229711 338167
rect 229593 320209 229711 320327
rect 229593 320049 229711 320167
rect 229593 302209 229711 302327
rect 229593 302049 229711 302167
rect 229593 284209 229711 284327
rect 229593 284049 229711 284167
rect 229593 266209 229711 266327
rect 229593 266049 229711 266167
rect 229593 248209 229711 248327
rect 229593 248049 229711 248167
rect 229593 230209 229711 230327
rect 229593 230049 229711 230167
rect 229593 212209 229711 212327
rect 229593 212049 229711 212167
rect 229593 194209 229711 194327
rect 229593 194049 229711 194167
rect 229593 176209 229711 176327
rect 229593 176049 229711 176167
rect 229593 158209 229711 158327
rect 229593 158049 229711 158167
rect 229593 140209 229711 140327
rect 229593 140049 229711 140167
rect 229593 122209 229711 122327
rect 229593 122049 229711 122167
rect 229593 104209 229711 104327
rect 229593 104049 229711 104167
rect 229593 86209 229711 86327
rect 229593 86049 229711 86167
rect 229593 68209 229711 68327
rect 229593 68049 229711 68167
rect 229593 50209 229711 50327
rect 229593 50049 229711 50167
rect 229593 32209 229711 32327
rect 229593 32049 229711 32167
rect 229593 14209 229711 14327
rect 229593 14049 229711 14167
rect 229593 -2641 229711 -2523
rect 229593 -2801 229711 -2683
rect 240393 355121 240511 355239
rect 240393 354961 240511 355079
rect 238593 354181 238711 354299
rect 238593 354021 238711 354139
rect 236793 353241 236911 353359
rect 236793 353081 236911 353199
rect 231393 340009 231511 340127
rect 231393 339849 231511 339967
rect 231393 322009 231511 322127
rect 231393 321849 231511 321967
rect 231393 304009 231511 304127
rect 231393 303849 231511 303967
rect 231393 286009 231511 286127
rect 231393 285849 231511 285967
rect 231393 268009 231511 268127
rect 231393 267849 231511 267967
rect 231393 250009 231511 250127
rect 231393 249849 231511 249967
rect 231393 232009 231511 232127
rect 231393 231849 231511 231967
rect 231393 214009 231511 214127
rect 231393 213849 231511 213967
rect 231393 196009 231511 196127
rect 231393 195849 231511 195967
rect 231393 178009 231511 178127
rect 231393 177849 231511 177967
rect 231393 160009 231511 160127
rect 231393 159849 231511 159967
rect 231393 142009 231511 142127
rect 231393 141849 231511 141967
rect 231393 124009 231511 124127
rect 231393 123849 231511 123967
rect 231393 106009 231511 106127
rect 231393 105849 231511 105967
rect 231393 88009 231511 88127
rect 231393 87849 231511 87967
rect 231393 70009 231511 70127
rect 231393 69849 231511 69967
rect 231393 52009 231511 52127
rect 231393 51849 231511 51967
rect 231393 34009 231511 34127
rect 231393 33849 231511 33967
rect 231393 16009 231511 16127
rect 231393 15849 231511 15967
rect 222393 -3111 222511 -2993
rect 222393 -3271 222511 -3153
rect 234993 352301 235111 352419
rect 234993 352141 235111 352259
rect 234993 343609 235111 343727
rect 234993 343449 235111 343567
rect 234993 325609 235111 325727
rect 234993 325449 235111 325567
rect 234993 307609 235111 307727
rect 234993 307449 235111 307567
rect 234993 289609 235111 289727
rect 234993 289449 235111 289567
rect 234993 271609 235111 271727
rect 234993 271449 235111 271567
rect 234993 253609 235111 253727
rect 234993 253449 235111 253567
rect 234993 235609 235111 235727
rect 234993 235449 235111 235567
rect 234993 217609 235111 217727
rect 234993 217449 235111 217567
rect 234993 199609 235111 199727
rect 234993 199449 235111 199567
rect 234993 181609 235111 181727
rect 234993 181449 235111 181567
rect 234993 163609 235111 163727
rect 234993 163449 235111 163567
rect 234993 145609 235111 145727
rect 234993 145449 235111 145567
rect 234993 127609 235111 127727
rect 234993 127449 235111 127567
rect 234993 109609 235111 109727
rect 234993 109449 235111 109567
rect 234993 91609 235111 91727
rect 234993 91449 235111 91567
rect 234993 73609 235111 73727
rect 234993 73449 235111 73567
rect 234993 55609 235111 55727
rect 234993 55449 235111 55567
rect 234993 37609 235111 37727
rect 234993 37449 235111 37567
rect 234993 19609 235111 19727
rect 234993 19449 235111 19567
rect 234993 1609 235111 1727
rect 234993 1449 235111 1567
rect 234993 -291 235111 -173
rect 234993 -451 235111 -333
rect 236793 345409 236911 345527
rect 236793 345249 236911 345367
rect 236793 327409 236911 327527
rect 236793 327249 236911 327367
rect 236793 309409 236911 309527
rect 236793 309249 236911 309367
rect 236793 291409 236911 291527
rect 236793 291249 236911 291367
rect 236793 273409 236911 273527
rect 236793 273249 236911 273367
rect 236793 255409 236911 255527
rect 236793 255249 236911 255367
rect 236793 237409 236911 237527
rect 236793 237249 236911 237367
rect 236793 219409 236911 219527
rect 236793 219249 236911 219367
rect 236793 201409 236911 201527
rect 236793 201249 236911 201367
rect 236793 183409 236911 183527
rect 236793 183249 236911 183367
rect 236793 165409 236911 165527
rect 236793 165249 236911 165367
rect 236793 147409 236911 147527
rect 236793 147249 236911 147367
rect 236793 129409 236911 129527
rect 236793 129249 236911 129367
rect 236793 111409 236911 111527
rect 236793 111249 236911 111367
rect 236793 93409 236911 93527
rect 236793 93249 236911 93367
rect 236793 75409 236911 75527
rect 236793 75249 236911 75367
rect 236793 57409 236911 57527
rect 236793 57249 236911 57367
rect 236793 39409 236911 39527
rect 236793 39249 236911 39367
rect 236793 21409 236911 21527
rect 236793 21249 236911 21367
rect 236793 3409 236911 3527
rect 236793 3249 236911 3367
rect 236793 -1231 236911 -1113
rect 236793 -1391 236911 -1273
rect 238593 347209 238711 347327
rect 238593 347049 238711 347167
rect 238593 329209 238711 329327
rect 238593 329049 238711 329167
rect 238593 311209 238711 311327
rect 238593 311049 238711 311167
rect 238593 293209 238711 293327
rect 238593 293049 238711 293167
rect 238593 275209 238711 275327
rect 238593 275049 238711 275167
rect 238593 257209 238711 257327
rect 238593 257049 238711 257167
rect 238593 239209 238711 239327
rect 238593 239049 238711 239167
rect 238593 221209 238711 221327
rect 238593 221049 238711 221167
rect 238593 203209 238711 203327
rect 238593 203049 238711 203167
rect 238593 185209 238711 185327
rect 238593 185049 238711 185167
rect 238593 167209 238711 167327
rect 238593 167049 238711 167167
rect 238593 149209 238711 149327
rect 238593 149049 238711 149167
rect 238593 131209 238711 131327
rect 238593 131049 238711 131167
rect 238593 113209 238711 113327
rect 238593 113049 238711 113167
rect 238593 95209 238711 95327
rect 238593 95049 238711 95167
rect 238593 77209 238711 77327
rect 238593 77049 238711 77167
rect 238593 59209 238711 59327
rect 238593 59049 238711 59167
rect 238593 41209 238711 41327
rect 238593 41049 238711 41167
rect 238593 23209 238711 23327
rect 238593 23049 238711 23167
rect 238593 5209 238711 5327
rect 238593 5049 238711 5167
rect 238593 -2171 238711 -2053
rect 238593 -2331 238711 -2213
rect 249393 355591 249511 355709
rect 249393 355431 249511 355549
rect 247593 354651 247711 354769
rect 247593 354491 247711 354609
rect 245793 353711 245911 353829
rect 245793 353551 245911 353669
rect 240393 349009 240511 349127
rect 240393 348849 240511 348967
rect 240393 331009 240511 331127
rect 240393 330849 240511 330967
rect 240393 313009 240511 313127
rect 240393 312849 240511 312967
rect 240393 295009 240511 295127
rect 240393 294849 240511 294967
rect 240393 277009 240511 277127
rect 240393 276849 240511 276967
rect 240393 259009 240511 259127
rect 240393 258849 240511 258967
rect 240393 241009 240511 241127
rect 240393 240849 240511 240967
rect 240393 223009 240511 223127
rect 240393 222849 240511 222967
rect 240393 205009 240511 205127
rect 240393 204849 240511 204967
rect 240393 187009 240511 187127
rect 240393 186849 240511 186967
rect 240393 169009 240511 169127
rect 240393 168849 240511 168967
rect 240393 151009 240511 151127
rect 240393 150849 240511 150967
rect 240393 133009 240511 133127
rect 240393 132849 240511 132967
rect 240393 115009 240511 115127
rect 240393 114849 240511 114967
rect 240393 97009 240511 97127
rect 240393 96849 240511 96967
rect 240393 79009 240511 79127
rect 240393 78849 240511 78967
rect 240393 61009 240511 61127
rect 240393 60849 240511 60967
rect 240393 43009 240511 43127
rect 240393 42849 240511 42967
rect 240393 25009 240511 25127
rect 240393 24849 240511 24967
rect 240393 7009 240511 7127
rect 240393 6849 240511 6967
rect 231393 -3581 231511 -3463
rect 231393 -3741 231511 -3623
rect 243993 352771 244111 352889
rect 243993 352611 244111 352729
rect 243993 334609 244111 334727
rect 243993 334449 244111 334567
rect 243993 316609 244111 316727
rect 243993 316449 244111 316567
rect 243993 298609 244111 298727
rect 243993 298449 244111 298567
rect 243993 280609 244111 280727
rect 243993 280449 244111 280567
rect 243993 262609 244111 262727
rect 243993 262449 244111 262567
rect 243993 244609 244111 244727
rect 243993 244449 244111 244567
rect 243993 226609 244111 226727
rect 243993 226449 244111 226567
rect 243993 208609 244111 208727
rect 243993 208449 244111 208567
rect 243993 190609 244111 190727
rect 243993 190449 244111 190567
rect 243993 172609 244111 172727
rect 243993 172449 244111 172567
rect 243993 154609 244111 154727
rect 243993 154449 244111 154567
rect 243993 136609 244111 136727
rect 243993 136449 244111 136567
rect 243993 118609 244111 118727
rect 243993 118449 244111 118567
rect 243993 100609 244111 100727
rect 243993 100449 244111 100567
rect 243993 82609 244111 82727
rect 243993 82449 244111 82567
rect 243993 64609 244111 64727
rect 243993 64449 244111 64567
rect 243993 46609 244111 46727
rect 243993 46449 244111 46567
rect 243993 28609 244111 28727
rect 243993 28449 244111 28567
rect 243993 10609 244111 10727
rect 243993 10449 244111 10567
rect 243993 -761 244111 -643
rect 243993 -921 244111 -803
rect 245793 336409 245911 336527
rect 245793 336249 245911 336367
rect 245793 318409 245911 318527
rect 245793 318249 245911 318367
rect 245793 300409 245911 300527
rect 245793 300249 245911 300367
rect 245793 282409 245911 282527
rect 245793 282249 245911 282367
rect 245793 264409 245911 264527
rect 245793 264249 245911 264367
rect 245793 246409 245911 246527
rect 245793 246249 245911 246367
rect 245793 228409 245911 228527
rect 245793 228249 245911 228367
rect 245793 210409 245911 210527
rect 245793 210249 245911 210367
rect 245793 192409 245911 192527
rect 245793 192249 245911 192367
rect 245793 174409 245911 174527
rect 245793 174249 245911 174367
rect 245793 156409 245911 156527
rect 245793 156249 245911 156367
rect 245793 138409 245911 138527
rect 245793 138249 245911 138367
rect 245793 120409 245911 120527
rect 245793 120249 245911 120367
rect 245793 102409 245911 102527
rect 245793 102249 245911 102367
rect 245793 84409 245911 84527
rect 245793 84249 245911 84367
rect 245793 66409 245911 66527
rect 245793 66249 245911 66367
rect 245793 48409 245911 48527
rect 245793 48249 245911 48367
rect 245793 30409 245911 30527
rect 245793 30249 245911 30367
rect 245793 12409 245911 12527
rect 245793 12249 245911 12367
rect 245793 -1701 245911 -1583
rect 245793 -1861 245911 -1743
rect 247593 338209 247711 338327
rect 247593 338049 247711 338167
rect 247593 320209 247711 320327
rect 247593 320049 247711 320167
rect 247593 302209 247711 302327
rect 247593 302049 247711 302167
rect 247593 284209 247711 284327
rect 247593 284049 247711 284167
rect 247593 266209 247711 266327
rect 247593 266049 247711 266167
rect 247593 248209 247711 248327
rect 247593 248049 247711 248167
rect 247593 230209 247711 230327
rect 247593 230049 247711 230167
rect 247593 212209 247711 212327
rect 247593 212049 247711 212167
rect 247593 194209 247711 194327
rect 247593 194049 247711 194167
rect 247593 176209 247711 176327
rect 247593 176049 247711 176167
rect 247593 158209 247711 158327
rect 247593 158049 247711 158167
rect 247593 140209 247711 140327
rect 247593 140049 247711 140167
rect 247593 122209 247711 122327
rect 247593 122049 247711 122167
rect 247593 104209 247711 104327
rect 247593 104049 247711 104167
rect 247593 86209 247711 86327
rect 247593 86049 247711 86167
rect 247593 68209 247711 68327
rect 247593 68049 247711 68167
rect 247593 50209 247711 50327
rect 247593 50049 247711 50167
rect 247593 32209 247711 32327
rect 247593 32049 247711 32167
rect 247593 14209 247711 14327
rect 247593 14049 247711 14167
rect 247593 -2641 247711 -2523
rect 247593 -2801 247711 -2683
rect 258393 355121 258511 355239
rect 258393 354961 258511 355079
rect 256593 354181 256711 354299
rect 256593 354021 256711 354139
rect 254793 353241 254911 353359
rect 254793 353081 254911 353199
rect 249393 340009 249511 340127
rect 249393 339849 249511 339967
rect 249393 322009 249511 322127
rect 249393 321849 249511 321967
rect 249393 304009 249511 304127
rect 249393 303849 249511 303967
rect 249393 286009 249511 286127
rect 249393 285849 249511 285967
rect 249393 268009 249511 268127
rect 249393 267849 249511 267967
rect 249393 250009 249511 250127
rect 249393 249849 249511 249967
rect 249393 232009 249511 232127
rect 249393 231849 249511 231967
rect 249393 214009 249511 214127
rect 249393 213849 249511 213967
rect 249393 196009 249511 196127
rect 249393 195849 249511 195967
rect 249393 178009 249511 178127
rect 249393 177849 249511 177967
rect 249393 160009 249511 160127
rect 249393 159849 249511 159967
rect 249393 142009 249511 142127
rect 249393 141849 249511 141967
rect 249393 124009 249511 124127
rect 249393 123849 249511 123967
rect 249393 106009 249511 106127
rect 249393 105849 249511 105967
rect 249393 88009 249511 88127
rect 249393 87849 249511 87967
rect 249393 70009 249511 70127
rect 249393 69849 249511 69967
rect 249393 52009 249511 52127
rect 249393 51849 249511 51967
rect 249393 34009 249511 34127
rect 249393 33849 249511 33967
rect 249393 16009 249511 16127
rect 249393 15849 249511 15967
rect 240393 -3111 240511 -2993
rect 240393 -3271 240511 -3153
rect 252993 352301 253111 352419
rect 252993 352141 253111 352259
rect 252993 343609 253111 343727
rect 252993 343449 253111 343567
rect 252993 325609 253111 325727
rect 252993 325449 253111 325567
rect 252993 307609 253111 307727
rect 252993 307449 253111 307567
rect 252993 289609 253111 289727
rect 252993 289449 253111 289567
rect 252993 271609 253111 271727
rect 252993 271449 253111 271567
rect 252993 253609 253111 253727
rect 252993 253449 253111 253567
rect 252993 235609 253111 235727
rect 252993 235449 253111 235567
rect 252993 217609 253111 217727
rect 252993 217449 253111 217567
rect 252993 199609 253111 199727
rect 252993 199449 253111 199567
rect 252993 181609 253111 181727
rect 252993 181449 253111 181567
rect 252993 163609 253111 163727
rect 252993 163449 253111 163567
rect 252993 145609 253111 145727
rect 252993 145449 253111 145567
rect 252993 127609 253111 127727
rect 252993 127449 253111 127567
rect 252993 109609 253111 109727
rect 252993 109449 253111 109567
rect 252993 91609 253111 91727
rect 252993 91449 253111 91567
rect 252993 73609 253111 73727
rect 252993 73449 253111 73567
rect 252993 55609 253111 55727
rect 252993 55449 253111 55567
rect 252993 37609 253111 37727
rect 252993 37449 253111 37567
rect 252993 19609 253111 19727
rect 252993 19449 253111 19567
rect 252993 1609 253111 1727
rect 252993 1449 253111 1567
rect 252993 -291 253111 -173
rect 252993 -451 253111 -333
rect 254793 345409 254911 345527
rect 254793 345249 254911 345367
rect 254793 327409 254911 327527
rect 254793 327249 254911 327367
rect 254793 309409 254911 309527
rect 254793 309249 254911 309367
rect 254793 291409 254911 291527
rect 254793 291249 254911 291367
rect 254793 273409 254911 273527
rect 254793 273249 254911 273367
rect 254793 255409 254911 255527
rect 254793 255249 254911 255367
rect 254793 237409 254911 237527
rect 254793 237249 254911 237367
rect 254793 219409 254911 219527
rect 254793 219249 254911 219367
rect 254793 201409 254911 201527
rect 254793 201249 254911 201367
rect 254793 183409 254911 183527
rect 254793 183249 254911 183367
rect 254793 165409 254911 165527
rect 254793 165249 254911 165367
rect 254793 147409 254911 147527
rect 254793 147249 254911 147367
rect 254793 129409 254911 129527
rect 254793 129249 254911 129367
rect 254793 111409 254911 111527
rect 254793 111249 254911 111367
rect 254793 93409 254911 93527
rect 254793 93249 254911 93367
rect 254793 75409 254911 75527
rect 254793 75249 254911 75367
rect 254793 57409 254911 57527
rect 254793 57249 254911 57367
rect 254793 39409 254911 39527
rect 254793 39249 254911 39367
rect 254793 21409 254911 21527
rect 254793 21249 254911 21367
rect 254793 3409 254911 3527
rect 254793 3249 254911 3367
rect 254793 -1231 254911 -1113
rect 254793 -1391 254911 -1273
rect 256593 347209 256711 347327
rect 256593 347049 256711 347167
rect 256593 329209 256711 329327
rect 256593 329049 256711 329167
rect 256593 311209 256711 311327
rect 256593 311049 256711 311167
rect 256593 293209 256711 293327
rect 256593 293049 256711 293167
rect 256593 275209 256711 275327
rect 256593 275049 256711 275167
rect 256593 257209 256711 257327
rect 256593 257049 256711 257167
rect 256593 239209 256711 239327
rect 256593 239049 256711 239167
rect 256593 221209 256711 221327
rect 256593 221049 256711 221167
rect 256593 203209 256711 203327
rect 256593 203049 256711 203167
rect 256593 185209 256711 185327
rect 256593 185049 256711 185167
rect 256593 167209 256711 167327
rect 256593 167049 256711 167167
rect 256593 149209 256711 149327
rect 256593 149049 256711 149167
rect 256593 131209 256711 131327
rect 256593 131049 256711 131167
rect 256593 113209 256711 113327
rect 256593 113049 256711 113167
rect 256593 95209 256711 95327
rect 256593 95049 256711 95167
rect 256593 77209 256711 77327
rect 256593 77049 256711 77167
rect 256593 59209 256711 59327
rect 256593 59049 256711 59167
rect 256593 41209 256711 41327
rect 256593 41049 256711 41167
rect 256593 23209 256711 23327
rect 256593 23049 256711 23167
rect 256593 5209 256711 5327
rect 256593 5049 256711 5167
rect 256593 -2171 256711 -2053
rect 256593 -2331 256711 -2213
rect 267393 355591 267511 355709
rect 267393 355431 267511 355549
rect 265593 354651 265711 354769
rect 265593 354491 265711 354609
rect 263793 353711 263911 353829
rect 263793 353551 263911 353669
rect 258393 349009 258511 349127
rect 258393 348849 258511 348967
rect 258393 331009 258511 331127
rect 258393 330849 258511 330967
rect 258393 313009 258511 313127
rect 258393 312849 258511 312967
rect 258393 295009 258511 295127
rect 258393 294849 258511 294967
rect 258393 277009 258511 277127
rect 258393 276849 258511 276967
rect 258393 259009 258511 259127
rect 258393 258849 258511 258967
rect 258393 241009 258511 241127
rect 258393 240849 258511 240967
rect 258393 223009 258511 223127
rect 258393 222849 258511 222967
rect 258393 205009 258511 205127
rect 258393 204849 258511 204967
rect 258393 187009 258511 187127
rect 258393 186849 258511 186967
rect 258393 169009 258511 169127
rect 258393 168849 258511 168967
rect 258393 151009 258511 151127
rect 258393 150849 258511 150967
rect 258393 133009 258511 133127
rect 258393 132849 258511 132967
rect 258393 115009 258511 115127
rect 258393 114849 258511 114967
rect 258393 97009 258511 97127
rect 258393 96849 258511 96967
rect 258393 79009 258511 79127
rect 258393 78849 258511 78967
rect 258393 61009 258511 61127
rect 258393 60849 258511 60967
rect 258393 43009 258511 43127
rect 258393 42849 258511 42967
rect 258393 25009 258511 25127
rect 258393 24849 258511 24967
rect 258393 7009 258511 7127
rect 258393 6849 258511 6967
rect 249393 -3581 249511 -3463
rect 249393 -3741 249511 -3623
rect 261993 352771 262111 352889
rect 261993 352611 262111 352729
rect 261993 334609 262111 334727
rect 261993 334449 262111 334567
rect 261993 316609 262111 316727
rect 261993 316449 262111 316567
rect 261993 298609 262111 298727
rect 261993 298449 262111 298567
rect 261993 280609 262111 280727
rect 261993 280449 262111 280567
rect 261993 262609 262111 262727
rect 261993 262449 262111 262567
rect 261993 244609 262111 244727
rect 261993 244449 262111 244567
rect 261993 226609 262111 226727
rect 261993 226449 262111 226567
rect 261993 208609 262111 208727
rect 261993 208449 262111 208567
rect 261993 190609 262111 190727
rect 261993 190449 262111 190567
rect 261993 172609 262111 172727
rect 261993 172449 262111 172567
rect 261993 154609 262111 154727
rect 261993 154449 262111 154567
rect 261993 136609 262111 136727
rect 261993 136449 262111 136567
rect 261993 118609 262111 118727
rect 261993 118449 262111 118567
rect 261993 100609 262111 100727
rect 261993 100449 262111 100567
rect 261993 82609 262111 82727
rect 261993 82449 262111 82567
rect 261993 64609 262111 64727
rect 261993 64449 262111 64567
rect 261993 46609 262111 46727
rect 261993 46449 262111 46567
rect 261993 28609 262111 28727
rect 261993 28449 262111 28567
rect 261993 10609 262111 10727
rect 261993 10449 262111 10567
rect 261993 -761 262111 -643
rect 261993 -921 262111 -803
rect 263793 336409 263911 336527
rect 263793 336249 263911 336367
rect 263793 318409 263911 318527
rect 263793 318249 263911 318367
rect 263793 300409 263911 300527
rect 263793 300249 263911 300367
rect 263793 282409 263911 282527
rect 263793 282249 263911 282367
rect 263793 264409 263911 264527
rect 263793 264249 263911 264367
rect 263793 246409 263911 246527
rect 263793 246249 263911 246367
rect 263793 228409 263911 228527
rect 263793 228249 263911 228367
rect 263793 210409 263911 210527
rect 263793 210249 263911 210367
rect 263793 192409 263911 192527
rect 263793 192249 263911 192367
rect 263793 174409 263911 174527
rect 263793 174249 263911 174367
rect 263793 156409 263911 156527
rect 263793 156249 263911 156367
rect 263793 138409 263911 138527
rect 263793 138249 263911 138367
rect 263793 120409 263911 120527
rect 263793 120249 263911 120367
rect 263793 102409 263911 102527
rect 263793 102249 263911 102367
rect 263793 84409 263911 84527
rect 263793 84249 263911 84367
rect 263793 66409 263911 66527
rect 263793 66249 263911 66367
rect 263793 48409 263911 48527
rect 263793 48249 263911 48367
rect 263793 30409 263911 30527
rect 263793 30249 263911 30367
rect 263793 12409 263911 12527
rect 263793 12249 263911 12367
rect 263793 -1701 263911 -1583
rect 263793 -1861 263911 -1743
rect 265593 338209 265711 338327
rect 265593 338049 265711 338167
rect 265593 320209 265711 320327
rect 265593 320049 265711 320167
rect 265593 302209 265711 302327
rect 265593 302049 265711 302167
rect 265593 284209 265711 284327
rect 265593 284049 265711 284167
rect 265593 266209 265711 266327
rect 265593 266049 265711 266167
rect 265593 248209 265711 248327
rect 265593 248049 265711 248167
rect 265593 230209 265711 230327
rect 265593 230049 265711 230167
rect 265593 212209 265711 212327
rect 265593 212049 265711 212167
rect 265593 194209 265711 194327
rect 265593 194049 265711 194167
rect 265593 176209 265711 176327
rect 265593 176049 265711 176167
rect 265593 158209 265711 158327
rect 265593 158049 265711 158167
rect 265593 140209 265711 140327
rect 265593 140049 265711 140167
rect 265593 122209 265711 122327
rect 265593 122049 265711 122167
rect 265593 104209 265711 104327
rect 265593 104049 265711 104167
rect 265593 86209 265711 86327
rect 265593 86049 265711 86167
rect 265593 68209 265711 68327
rect 265593 68049 265711 68167
rect 265593 50209 265711 50327
rect 265593 50049 265711 50167
rect 265593 32209 265711 32327
rect 265593 32049 265711 32167
rect 265593 14209 265711 14327
rect 265593 14049 265711 14167
rect 265593 -2641 265711 -2523
rect 265593 -2801 265711 -2683
rect 276393 355121 276511 355239
rect 276393 354961 276511 355079
rect 274593 354181 274711 354299
rect 274593 354021 274711 354139
rect 272793 353241 272911 353359
rect 272793 353081 272911 353199
rect 267393 340009 267511 340127
rect 267393 339849 267511 339967
rect 267393 322009 267511 322127
rect 267393 321849 267511 321967
rect 267393 304009 267511 304127
rect 267393 303849 267511 303967
rect 267393 286009 267511 286127
rect 267393 285849 267511 285967
rect 267393 268009 267511 268127
rect 267393 267849 267511 267967
rect 267393 250009 267511 250127
rect 267393 249849 267511 249967
rect 267393 232009 267511 232127
rect 267393 231849 267511 231967
rect 267393 214009 267511 214127
rect 267393 213849 267511 213967
rect 267393 196009 267511 196127
rect 267393 195849 267511 195967
rect 267393 178009 267511 178127
rect 267393 177849 267511 177967
rect 267393 160009 267511 160127
rect 267393 159849 267511 159967
rect 267393 142009 267511 142127
rect 267393 141849 267511 141967
rect 267393 124009 267511 124127
rect 267393 123849 267511 123967
rect 267393 106009 267511 106127
rect 267393 105849 267511 105967
rect 267393 88009 267511 88127
rect 267393 87849 267511 87967
rect 267393 70009 267511 70127
rect 267393 69849 267511 69967
rect 267393 52009 267511 52127
rect 267393 51849 267511 51967
rect 267393 34009 267511 34127
rect 267393 33849 267511 33967
rect 267393 16009 267511 16127
rect 267393 15849 267511 15967
rect 258393 -3111 258511 -2993
rect 258393 -3271 258511 -3153
rect 270993 352301 271111 352419
rect 270993 352141 271111 352259
rect 270993 343609 271111 343727
rect 270993 343449 271111 343567
rect 270993 325609 271111 325727
rect 270993 325449 271111 325567
rect 270993 307609 271111 307727
rect 270993 307449 271111 307567
rect 270993 289609 271111 289727
rect 270993 289449 271111 289567
rect 270993 271609 271111 271727
rect 270993 271449 271111 271567
rect 270993 253609 271111 253727
rect 270993 253449 271111 253567
rect 270993 235609 271111 235727
rect 270993 235449 271111 235567
rect 270993 217609 271111 217727
rect 270993 217449 271111 217567
rect 270993 199609 271111 199727
rect 270993 199449 271111 199567
rect 270993 181609 271111 181727
rect 270993 181449 271111 181567
rect 270993 163609 271111 163727
rect 270993 163449 271111 163567
rect 270993 145609 271111 145727
rect 270993 145449 271111 145567
rect 270993 127609 271111 127727
rect 270993 127449 271111 127567
rect 270993 109609 271111 109727
rect 270993 109449 271111 109567
rect 270993 91609 271111 91727
rect 270993 91449 271111 91567
rect 270993 73609 271111 73727
rect 270993 73449 271111 73567
rect 270993 55609 271111 55727
rect 270993 55449 271111 55567
rect 270993 37609 271111 37727
rect 270993 37449 271111 37567
rect 270993 19609 271111 19727
rect 270993 19449 271111 19567
rect 270993 1609 271111 1727
rect 270993 1449 271111 1567
rect 270993 -291 271111 -173
rect 270993 -451 271111 -333
rect 272793 345409 272911 345527
rect 272793 345249 272911 345367
rect 272793 327409 272911 327527
rect 272793 327249 272911 327367
rect 272793 309409 272911 309527
rect 272793 309249 272911 309367
rect 272793 291409 272911 291527
rect 272793 291249 272911 291367
rect 272793 273409 272911 273527
rect 272793 273249 272911 273367
rect 272793 255409 272911 255527
rect 272793 255249 272911 255367
rect 272793 237409 272911 237527
rect 272793 237249 272911 237367
rect 272793 219409 272911 219527
rect 272793 219249 272911 219367
rect 272793 201409 272911 201527
rect 272793 201249 272911 201367
rect 272793 183409 272911 183527
rect 272793 183249 272911 183367
rect 272793 165409 272911 165527
rect 272793 165249 272911 165367
rect 272793 147409 272911 147527
rect 272793 147249 272911 147367
rect 272793 129409 272911 129527
rect 272793 129249 272911 129367
rect 272793 111409 272911 111527
rect 272793 111249 272911 111367
rect 272793 93409 272911 93527
rect 272793 93249 272911 93367
rect 272793 75409 272911 75527
rect 272793 75249 272911 75367
rect 272793 57409 272911 57527
rect 272793 57249 272911 57367
rect 272793 39409 272911 39527
rect 272793 39249 272911 39367
rect 272793 21409 272911 21527
rect 272793 21249 272911 21367
rect 272793 3409 272911 3527
rect 272793 3249 272911 3367
rect 272793 -1231 272911 -1113
rect 272793 -1391 272911 -1273
rect 274593 347209 274711 347327
rect 274593 347049 274711 347167
rect 274593 329209 274711 329327
rect 274593 329049 274711 329167
rect 274593 311209 274711 311327
rect 274593 311049 274711 311167
rect 274593 293209 274711 293327
rect 274593 293049 274711 293167
rect 274593 275209 274711 275327
rect 274593 275049 274711 275167
rect 274593 257209 274711 257327
rect 274593 257049 274711 257167
rect 274593 239209 274711 239327
rect 274593 239049 274711 239167
rect 274593 221209 274711 221327
rect 274593 221049 274711 221167
rect 274593 203209 274711 203327
rect 274593 203049 274711 203167
rect 274593 185209 274711 185327
rect 274593 185049 274711 185167
rect 274593 167209 274711 167327
rect 274593 167049 274711 167167
rect 274593 149209 274711 149327
rect 274593 149049 274711 149167
rect 274593 131209 274711 131327
rect 274593 131049 274711 131167
rect 274593 113209 274711 113327
rect 274593 113049 274711 113167
rect 274593 95209 274711 95327
rect 274593 95049 274711 95167
rect 274593 77209 274711 77327
rect 274593 77049 274711 77167
rect 274593 59209 274711 59327
rect 274593 59049 274711 59167
rect 274593 41209 274711 41327
rect 274593 41049 274711 41167
rect 274593 23209 274711 23327
rect 274593 23049 274711 23167
rect 274593 5209 274711 5327
rect 274593 5049 274711 5167
rect 274593 -2171 274711 -2053
rect 274593 -2331 274711 -2213
rect 285393 355591 285511 355709
rect 285393 355431 285511 355549
rect 283593 354651 283711 354769
rect 283593 354491 283711 354609
rect 281793 353711 281911 353829
rect 281793 353551 281911 353669
rect 276393 349009 276511 349127
rect 276393 348849 276511 348967
rect 276393 331009 276511 331127
rect 276393 330849 276511 330967
rect 276393 313009 276511 313127
rect 276393 312849 276511 312967
rect 276393 295009 276511 295127
rect 276393 294849 276511 294967
rect 276393 277009 276511 277127
rect 276393 276849 276511 276967
rect 276393 259009 276511 259127
rect 276393 258849 276511 258967
rect 276393 241009 276511 241127
rect 276393 240849 276511 240967
rect 276393 223009 276511 223127
rect 276393 222849 276511 222967
rect 276393 205009 276511 205127
rect 276393 204849 276511 204967
rect 276393 187009 276511 187127
rect 276393 186849 276511 186967
rect 276393 169009 276511 169127
rect 276393 168849 276511 168967
rect 276393 151009 276511 151127
rect 276393 150849 276511 150967
rect 276393 133009 276511 133127
rect 276393 132849 276511 132967
rect 276393 115009 276511 115127
rect 276393 114849 276511 114967
rect 276393 97009 276511 97127
rect 276393 96849 276511 96967
rect 276393 79009 276511 79127
rect 276393 78849 276511 78967
rect 276393 61009 276511 61127
rect 276393 60849 276511 60967
rect 276393 43009 276511 43127
rect 276393 42849 276511 42967
rect 276393 25009 276511 25127
rect 276393 24849 276511 24967
rect 276393 7009 276511 7127
rect 276393 6849 276511 6967
rect 267393 -3581 267511 -3463
rect 267393 -3741 267511 -3623
rect 279993 352771 280111 352889
rect 279993 352611 280111 352729
rect 279993 334609 280111 334727
rect 279993 334449 280111 334567
rect 279993 316609 280111 316727
rect 279993 316449 280111 316567
rect 279993 298609 280111 298727
rect 279993 298449 280111 298567
rect 279993 280609 280111 280727
rect 279993 280449 280111 280567
rect 279993 262609 280111 262727
rect 279993 262449 280111 262567
rect 279993 244609 280111 244727
rect 279993 244449 280111 244567
rect 279993 226609 280111 226727
rect 279993 226449 280111 226567
rect 279993 208609 280111 208727
rect 279993 208449 280111 208567
rect 279993 190609 280111 190727
rect 279993 190449 280111 190567
rect 279993 172609 280111 172727
rect 279993 172449 280111 172567
rect 279993 154609 280111 154727
rect 279993 154449 280111 154567
rect 279993 136609 280111 136727
rect 279993 136449 280111 136567
rect 279993 118609 280111 118727
rect 279993 118449 280111 118567
rect 279993 100609 280111 100727
rect 279993 100449 280111 100567
rect 279993 82609 280111 82727
rect 279993 82449 280111 82567
rect 279993 64609 280111 64727
rect 279993 64449 280111 64567
rect 279993 46609 280111 46727
rect 279993 46449 280111 46567
rect 279993 28609 280111 28727
rect 279993 28449 280111 28567
rect 279993 10609 280111 10727
rect 279993 10449 280111 10567
rect 279993 -761 280111 -643
rect 279993 -921 280111 -803
rect 281793 336409 281911 336527
rect 281793 336249 281911 336367
rect 281793 318409 281911 318527
rect 281793 318249 281911 318367
rect 281793 300409 281911 300527
rect 281793 300249 281911 300367
rect 281793 282409 281911 282527
rect 281793 282249 281911 282367
rect 281793 264409 281911 264527
rect 281793 264249 281911 264367
rect 281793 246409 281911 246527
rect 281793 246249 281911 246367
rect 281793 228409 281911 228527
rect 281793 228249 281911 228367
rect 281793 210409 281911 210527
rect 281793 210249 281911 210367
rect 281793 192409 281911 192527
rect 281793 192249 281911 192367
rect 281793 174409 281911 174527
rect 281793 174249 281911 174367
rect 281793 156409 281911 156527
rect 281793 156249 281911 156367
rect 281793 138409 281911 138527
rect 281793 138249 281911 138367
rect 281793 120409 281911 120527
rect 281793 120249 281911 120367
rect 281793 102409 281911 102527
rect 281793 102249 281911 102367
rect 281793 84409 281911 84527
rect 281793 84249 281911 84367
rect 281793 66409 281911 66527
rect 281793 66249 281911 66367
rect 281793 48409 281911 48527
rect 281793 48249 281911 48367
rect 281793 30409 281911 30527
rect 281793 30249 281911 30367
rect 281793 12409 281911 12527
rect 281793 12249 281911 12367
rect 281793 -1701 281911 -1583
rect 281793 -1861 281911 -1743
rect 283593 338209 283711 338327
rect 283593 338049 283711 338167
rect 283593 320209 283711 320327
rect 283593 320049 283711 320167
rect 283593 302209 283711 302327
rect 283593 302049 283711 302167
rect 283593 284209 283711 284327
rect 283593 284049 283711 284167
rect 283593 266209 283711 266327
rect 283593 266049 283711 266167
rect 283593 248209 283711 248327
rect 283593 248049 283711 248167
rect 283593 230209 283711 230327
rect 283593 230049 283711 230167
rect 283593 212209 283711 212327
rect 283593 212049 283711 212167
rect 283593 194209 283711 194327
rect 283593 194049 283711 194167
rect 283593 176209 283711 176327
rect 283593 176049 283711 176167
rect 283593 158209 283711 158327
rect 283593 158049 283711 158167
rect 283593 140209 283711 140327
rect 283593 140049 283711 140167
rect 283593 122209 283711 122327
rect 283593 122049 283711 122167
rect 283593 104209 283711 104327
rect 283593 104049 283711 104167
rect 283593 86209 283711 86327
rect 283593 86049 283711 86167
rect 283593 68209 283711 68327
rect 283593 68049 283711 68167
rect 283593 50209 283711 50327
rect 283593 50049 283711 50167
rect 283593 32209 283711 32327
rect 283593 32049 283711 32167
rect 283593 14209 283711 14327
rect 283593 14049 283711 14167
rect 283593 -2641 283711 -2523
rect 283593 -2801 283711 -2683
rect 296041 355591 296159 355709
rect 296041 355431 296159 355549
rect 295571 355121 295689 355239
rect 295571 354961 295689 355079
rect 295101 354651 295219 354769
rect 295101 354491 295219 354609
rect 294631 354181 294749 354299
rect 294631 354021 294749 354139
rect 294161 353711 294279 353829
rect 294161 353551 294279 353669
rect 290793 353241 290911 353359
rect 290793 353081 290911 353199
rect 285393 340009 285511 340127
rect 285393 339849 285511 339967
rect 285393 322009 285511 322127
rect 285393 321849 285511 321967
rect 285393 304009 285511 304127
rect 285393 303849 285511 303967
rect 285393 286009 285511 286127
rect 285393 285849 285511 285967
rect 285393 268009 285511 268127
rect 285393 267849 285511 267967
rect 285393 250009 285511 250127
rect 285393 249849 285511 249967
rect 285393 232009 285511 232127
rect 285393 231849 285511 231967
rect 285393 214009 285511 214127
rect 285393 213849 285511 213967
rect 285393 196009 285511 196127
rect 285393 195849 285511 195967
rect 285393 178009 285511 178127
rect 285393 177849 285511 177967
rect 285393 160009 285511 160127
rect 285393 159849 285511 159967
rect 285393 142009 285511 142127
rect 285393 141849 285511 141967
rect 285393 124009 285511 124127
rect 285393 123849 285511 123967
rect 285393 106009 285511 106127
rect 285393 105849 285511 105967
rect 285393 88009 285511 88127
rect 285393 87849 285511 87967
rect 285393 70009 285511 70127
rect 285393 69849 285511 69967
rect 285393 52009 285511 52127
rect 285393 51849 285511 51967
rect 285393 34009 285511 34127
rect 285393 33849 285511 33967
rect 285393 16009 285511 16127
rect 285393 15849 285511 15967
rect 276393 -3111 276511 -2993
rect 276393 -3271 276511 -3153
rect 288993 352301 289111 352419
rect 288993 352141 289111 352259
rect 288993 343609 289111 343727
rect 288993 343449 289111 343567
rect 288993 325609 289111 325727
rect 288993 325449 289111 325567
rect 288993 307609 289111 307727
rect 288993 307449 289111 307567
rect 288993 289609 289111 289727
rect 288993 289449 289111 289567
rect 288993 271609 289111 271727
rect 288993 271449 289111 271567
rect 288993 253609 289111 253727
rect 288993 253449 289111 253567
rect 288993 235609 289111 235727
rect 288993 235449 289111 235567
rect 288993 217609 289111 217727
rect 288993 217449 289111 217567
rect 288993 199609 289111 199727
rect 288993 199449 289111 199567
rect 288993 181609 289111 181727
rect 288993 181449 289111 181567
rect 288993 163609 289111 163727
rect 288993 163449 289111 163567
rect 288993 145609 289111 145727
rect 288993 145449 289111 145567
rect 288993 127609 289111 127727
rect 288993 127449 289111 127567
rect 288993 109609 289111 109727
rect 288993 109449 289111 109567
rect 288993 91609 289111 91727
rect 288993 91449 289111 91567
rect 288993 73609 289111 73727
rect 288993 73449 289111 73567
rect 288993 55609 289111 55727
rect 288993 55449 289111 55567
rect 288993 37609 289111 37727
rect 288993 37449 289111 37567
rect 288993 19609 289111 19727
rect 288993 19449 289111 19567
rect 288993 1609 289111 1727
rect 288993 1449 289111 1567
rect 288993 -291 289111 -173
rect 288993 -451 289111 -333
rect 293691 353241 293809 353359
rect 293691 353081 293809 353199
rect 293221 352771 293339 352889
rect 293221 352611 293339 352729
rect 290793 345409 290911 345527
rect 290793 345249 290911 345367
rect 290793 327409 290911 327527
rect 290793 327249 290911 327367
rect 290793 309409 290911 309527
rect 290793 309249 290911 309367
rect 290793 291409 290911 291527
rect 290793 291249 290911 291367
rect 290793 273409 290911 273527
rect 290793 273249 290911 273367
rect 290793 255409 290911 255527
rect 290793 255249 290911 255367
rect 290793 237409 290911 237527
rect 290793 237249 290911 237367
rect 290793 219409 290911 219527
rect 290793 219249 290911 219367
rect 290793 201409 290911 201527
rect 290793 201249 290911 201367
rect 290793 183409 290911 183527
rect 290793 183249 290911 183367
rect 290793 165409 290911 165527
rect 290793 165249 290911 165367
rect 290793 147409 290911 147527
rect 290793 147249 290911 147367
rect 290793 129409 290911 129527
rect 290793 129249 290911 129367
rect 290793 111409 290911 111527
rect 290793 111249 290911 111367
rect 290793 93409 290911 93527
rect 290793 93249 290911 93367
rect 290793 75409 290911 75527
rect 290793 75249 290911 75367
rect 290793 57409 290911 57527
rect 290793 57249 290911 57367
rect 290793 39409 290911 39527
rect 290793 39249 290911 39367
rect 290793 21409 290911 21527
rect 290793 21249 290911 21367
rect 290793 3409 290911 3527
rect 290793 3249 290911 3367
rect 292751 352301 292869 352419
rect 292751 352141 292869 352259
rect 292751 343609 292869 343727
rect 292751 343449 292869 343567
rect 292751 325609 292869 325727
rect 292751 325449 292869 325567
rect 292751 307609 292869 307727
rect 292751 307449 292869 307567
rect 292751 289609 292869 289727
rect 292751 289449 292869 289567
rect 292751 271609 292869 271727
rect 292751 271449 292869 271567
rect 292751 253609 292869 253727
rect 292751 253449 292869 253567
rect 292751 235609 292869 235727
rect 292751 235449 292869 235567
rect 292751 217609 292869 217727
rect 292751 217449 292869 217567
rect 292751 199609 292869 199727
rect 292751 199449 292869 199567
rect 292751 181609 292869 181727
rect 292751 181449 292869 181567
rect 292751 163609 292869 163727
rect 292751 163449 292869 163567
rect 292751 145609 292869 145727
rect 292751 145449 292869 145567
rect 292751 127609 292869 127727
rect 292751 127449 292869 127567
rect 292751 109609 292869 109727
rect 292751 109449 292869 109567
rect 292751 91609 292869 91727
rect 292751 91449 292869 91567
rect 292751 73609 292869 73727
rect 292751 73449 292869 73567
rect 292751 55609 292869 55727
rect 292751 55449 292869 55567
rect 292751 37609 292869 37727
rect 292751 37449 292869 37567
rect 292751 19609 292869 19727
rect 292751 19449 292869 19567
rect 292751 1609 292869 1727
rect 292751 1449 292869 1567
rect 292751 -291 292869 -173
rect 292751 -451 292869 -333
rect 293221 334609 293339 334727
rect 293221 334449 293339 334567
rect 293221 316609 293339 316727
rect 293221 316449 293339 316567
rect 293221 298609 293339 298727
rect 293221 298449 293339 298567
rect 293221 280609 293339 280727
rect 293221 280449 293339 280567
rect 293221 262609 293339 262727
rect 293221 262449 293339 262567
rect 293221 244609 293339 244727
rect 293221 244449 293339 244567
rect 293221 226609 293339 226727
rect 293221 226449 293339 226567
rect 293221 208609 293339 208727
rect 293221 208449 293339 208567
rect 293221 190609 293339 190727
rect 293221 190449 293339 190567
rect 293221 172609 293339 172727
rect 293221 172449 293339 172567
rect 293221 154609 293339 154727
rect 293221 154449 293339 154567
rect 293221 136609 293339 136727
rect 293221 136449 293339 136567
rect 293221 118609 293339 118727
rect 293221 118449 293339 118567
rect 293221 100609 293339 100727
rect 293221 100449 293339 100567
rect 293221 82609 293339 82727
rect 293221 82449 293339 82567
rect 293221 64609 293339 64727
rect 293221 64449 293339 64567
rect 293221 46609 293339 46727
rect 293221 46449 293339 46567
rect 293221 28609 293339 28727
rect 293221 28449 293339 28567
rect 293221 10609 293339 10727
rect 293221 10449 293339 10567
rect 293221 -761 293339 -643
rect 293221 -921 293339 -803
rect 293691 345409 293809 345527
rect 293691 345249 293809 345367
rect 293691 327409 293809 327527
rect 293691 327249 293809 327367
rect 293691 309409 293809 309527
rect 293691 309249 293809 309367
rect 293691 291409 293809 291527
rect 293691 291249 293809 291367
rect 293691 273409 293809 273527
rect 293691 273249 293809 273367
rect 293691 255409 293809 255527
rect 293691 255249 293809 255367
rect 293691 237409 293809 237527
rect 293691 237249 293809 237367
rect 293691 219409 293809 219527
rect 293691 219249 293809 219367
rect 293691 201409 293809 201527
rect 293691 201249 293809 201367
rect 293691 183409 293809 183527
rect 293691 183249 293809 183367
rect 293691 165409 293809 165527
rect 293691 165249 293809 165367
rect 293691 147409 293809 147527
rect 293691 147249 293809 147367
rect 293691 129409 293809 129527
rect 293691 129249 293809 129367
rect 293691 111409 293809 111527
rect 293691 111249 293809 111367
rect 293691 93409 293809 93527
rect 293691 93249 293809 93367
rect 293691 75409 293809 75527
rect 293691 75249 293809 75367
rect 293691 57409 293809 57527
rect 293691 57249 293809 57367
rect 293691 39409 293809 39527
rect 293691 39249 293809 39367
rect 293691 21409 293809 21527
rect 293691 21249 293809 21367
rect 293691 3409 293809 3527
rect 293691 3249 293809 3367
rect 290793 -1231 290911 -1113
rect 290793 -1391 290911 -1273
rect 293691 -1231 293809 -1113
rect 293691 -1391 293809 -1273
rect 294161 336409 294279 336527
rect 294161 336249 294279 336367
rect 294161 318409 294279 318527
rect 294161 318249 294279 318367
rect 294161 300409 294279 300527
rect 294161 300249 294279 300367
rect 294161 282409 294279 282527
rect 294161 282249 294279 282367
rect 294161 264409 294279 264527
rect 294161 264249 294279 264367
rect 294161 246409 294279 246527
rect 294161 246249 294279 246367
rect 294161 228409 294279 228527
rect 294161 228249 294279 228367
rect 294161 210409 294279 210527
rect 294161 210249 294279 210367
rect 294161 192409 294279 192527
rect 294161 192249 294279 192367
rect 294161 174409 294279 174527
rect 294161 174249 294279 174367
rect 294161 156409 294279 156527
rect 294161 156249 294279 156367
rect 294161 138409 294279 138527
rect 294161 138249 294279 138367
rect 294161 120409 294279 120527
rect 294161 120249 294279 120367
rect 294161 102409 294279 102527
rect 294161 102249 294279 102367
rect 294161 84409 294279 84527
rect 294161 84249 294279 84367
rect 294161 66409 294279 66527
rect 294161 66249 294279 66367
rect 294161 48409 294279 48527
rect 294161 48249 294279 48367
rect 294161 30409 294279 30527
rect 294161 30249 294279 30367
rect 294161 12409 294279 12527
rect 294161 12249 294279 12367
rect 294161 -1701 294279 -1583
rect 294161 -1861 294279 -1743
rect 294631 347209 294749 347327
rect 294631 347049 294749 347167
rect 294631 329209 294749 329327
rect 294631 329049 294749 329167
rect 294631 311209 294749 311327
rect 294631 311049 294749 311167
rect 294631 293209 294749 293327
rect 294631 293049 294749 293167
rect 294631 275209 294749 275327
rect 294631 275049 294749 275167
rect 294631 257209 294749 257327
rect 294631 257049 294749 257167
rect 294631 239209 294749 239327
rect 294631 239049 294749 239167
rect 294631 221209 294749 221327
rect 294631 221049 294749 221167
rect 294631 203209 294749 203327
rect 294631 203049 294749 203167
rect 294631 185209 294749 185327
rect 294631 185049 294749 185167
rect 294631 167209 294749 167327
rect 294631 167049 294749 167167
rect 294631 149209 294749 149327
rect 294631 149049 294749 149167
rect 294631 131209 294749 131327
rect 294631 131049 294749 131167
rect 294631 113209 294749 113327
rect 294631 113049 294749 113167
rect 294631 95209 294749 95327
rect 294631 95049 294749 95167
rect 294631 77209 294749 77327
rect 294631 77049 294749 77167
rect 294631 59209 294749 59327
rect 294631 59049 294749 59167
rect 294631 41209 294749 41327
rect 294631 41049 294749 41167
rect 294631 23209 294749 23327
rect 294631 23049 294749 23167
rect 294631 5209 294749 5327
rect 294631 5049 294749 5167
rect 294631 -2171 294749 -2053
rect 294631 -2331 294749 -2213
rect 295101 338209 295219 338327
rect 295101 338049 295219 338167
rect 295101 320209 295219 320327
rect 295101 320049 295219 320167
rect 295101 302209 295219 302327
rect 295101 302049 295219 302167
rect 295101 284209 295219 284327
rect 295101 284049 295219 284167
rect 295101 266209 295219 266327
rect 295101 266049 295219 266167
rect 295101 248209 295219 248327
rect 295101 248049 295219 248167
rect 295101 230209 295219 230327
rect 295101 230049 295219 230167
rect 295101 212209 295219 212327
rect 295101 212049 295219 212167
rect 295101 194209 295219 194327
rect 295101 194049 295219 194167
rect 295101 176209 295219 176327
rect 295101 176049 295219 176167
rect 295101 158209 295219 158327
rect 295101 158049 295219 158167
rect 295101 140209 295219 140327
rect 295101 140049 295219 140167
rect 295101 122209 295219 122327
rect 295101 122049 295219 122167
rect 295101 104209 295219 104327
rect 295101 104049 295219 104167
rect 295101 86209 295219 86327
rect 295101 86049 295219 86167
rect 295101 68209 295219 68327
rect 295101 68049 295219 68167
rect 295101 50209 295219 50327
rect 295101 50049 295219 50167
rect 295101 32209 295219 32327
rect 295101 32049 295219 32167
rect 295101 14209 295219 14327
rect 295101 14049 295219 14167
rect 295101 -2641 295219 -2523
rect 295101 -2801 295219 -2683
rect 295571 349009 295689 349127
rect 295571 348849 295689 348967
rect 295571 331009 295689 331127
rect 295571 330849 295689 330967
rect 295571 313009 295689 313127
rect 295571 312849 295689 312967
rect 295571 295009 295689 295127
rect 295571 294849 295689 294967
rect 295571 277009 295689 277127
rect 295571 276849 295689 276967
rect 295571 259009 295689 259127
rect 295571 258849 295689 258967
rect 295571 241009 295689 241127
rect 295571 240849 295689 240967
rect 295571 223009 295689 223127
rect 295571 222849 295689 222967
rect 295571 205009 295689 205127
rect 295571 204849 295689 204967
rect 295571 187009 295689 187127
rect 295571 186849 295689 186967
rect 295571 169009 295689 169127
rect 295571 168849 295689 168967
rect 295571 151009 295689 151127
rect 295571 150849 295689 150967
rect 295571 133009 295689 133127
rect 295571 132849 295689 132967
rect 295571 115009 295689 115127
rect 295571 114849 295689 114967
rect 295571 97009 295689 97127
rect 295571 96849 295689 96967
rect 295571 79009 295689 79127
rect 295571 78849 295689 78967
rect 295571 61009 295689 61127
rect 295571 60849 295689 60967
rect 295571 43009 295689 43127
rect 295571 42849 295689 42967
rect 295571 25009 295689 25127
rect 295571 24849 295689 24967
rect 295571 7009 295689 7127
rect 295571 6849 295689 6967
rect 295571 -3111 295689 -2993
rect 295571 -3271 295689 -3153
rect 296041 340009 296159 340127
rect 296041 339849 296159 339967
rect 296041 322009 296159 322127
rect 296041 321849 296159 321967
rect 296041 304009 296159 304127
rect 296041 303849 296159 303967
rect 296041 286009 296159 286127
rect 296041 285849 296159 285967
rect 296041 268009 296159 268127
rect 296041 267849 296159 267967
rect 296041 250009 296159 250127
rect 296041 249849 296159 249967
rect 296041 232009 296159 232127
rect 296041 231849 296159 231967
rect 296041 214009 296159 214127
rect 296041 213849 296159 213967
rect 296041 196009 296159 196127
rect 296041 195849 296159 195967
rect 296041 178009 296159 178127
rect 296041 177849 296159 177967
rect 296041 160009 296159 160127
rect 296041 159849 296159 159967
rect 296041 142009 296159 142127
rect 296041 141849 296159 141967
rect 296041 124009 296159 124127
rect 296041 123849 296159 123967
rect 296041 106009 296159 106127
rect 296041 105849 296159 105967
rect 296041 88009 296159 88127
rect 296041 87849 296159 87967
rect 296041 70009 296159 70127
rect 296041 69849 296159 69967
rect 296041 52009 296159 52127
rect 296041 51849 296159 51967
rect 296041 34009 296159 34127
rect 296041 33849 296159 33967
rect 296041 16009 296159 16127
rect 296041 15849 296159 15967
rect 285393 -3581 285511 -3463
rect 285393 -3741 285511 -3623
rect 296041 -3581 296159 -3463
rect 296041 -3741 296159 -3623
<< metal5 >>
rect -4288 355720 -3988 355721
rect 15302 355720 15602 355721
rect 33302 355720 33602 355721
rect 51302 355720 51602 355721
rect 69302 355720 69602 355721
rect 87302 355720 87602 355721
rect 105302 355720 105602 355721
rect 123302 355720 123602 355721
rect 141302 355720 141602 355721
rect 159302 355720 159602 355721
rect 177302 355720 177602 355721
rect 195302 355720 195602 355721
rect 213302 355720 213602 355721
rect 231302 355720 231602 355721
rect 249302 355720 249602 355721
rect 267302 355720 267602 355721
rect 285302 355720 285602 355721
rect 295950 355720 296250 355721
rect -4288 355709 296250 355720
rect -4288 355591 -4197 355709
rect -4079 355591 15393 355709
rect 15511 355591 33393 355709
rect 33511 355591 51393 355709
rect 51511 355591 69393 355709
rect 69511 355591 87393 355709
rect 87511 355591 105393 355709
rect 105511 355591 123393 355709
rect 123511 355591 141393 355709
rect 141511 355591 159393 355709
rect 159511 355591 177393 355709
rect 177511 355591 195393 355709
rect 195511 355591 213393 355709
rect 213511 355591 231393 355709
rect 231511 355591 249393 355709
rect 249511 355591 267393 355709
rect 267511 355591 285393 355709
rect 285511 355591 296041 355709
rect 296159 355591 296250 355709
rect -4288 355549 296250 355591
rect -4288 355431 -4197 355549
rect -4079 355431 15393 355549
rect 15511 355431 33393 355549
rect 33511 355431 51393 355549
rect 51511 355431 69393 355549
rect 69511 355431 87393 355549
rect 87511 355431 105393 355549
rect 105511 355431 123393 355549
rect 123511 355431 141393 355549
rect 141511 355431 159393 355549
rect 159511 355431 177393 355549
rect 177511 355431 195393 355549
rect 195511 355431 213393 355549
rect 213511 355431 231393 355549
rect 231511 355431 249393 355549
rect 249511 355431 267393 355549
rect 267511 355431 285393 355549
rect 285511 355431 296041 355549
rect 296159 355431 296250 355549
rect -4288 355420 296250 355431
rect -4288 355419 -3988 355420
rect 15302 355419 15602 355420
rect 33302 355419 33602 355420
rect 51302 355419 51602 355420
rect 69302 355419 69602 355420
rect 87302 355419 87602 355420
rect 105302 355419 105602 355420
rect 123302 355419 123602 355420
rect 141302 355419 141602 355420
rect 159302 355419 159602 355420
rect 177302 355419 177602 355420
rect 195302 355419 195602 355420
rect 213302 355419 213602 355420
rect 231302 355419 231602 355420
rect 249302 355419 249602 355420
rect 267302 355419 267602 355420
rect 285302 355419 285602 355420
rect 295950 355419 296250 355420
rect -3818 355250 -3518 355251
rect 6302 355250 6602 355251
rect 24302 355250 24602 355251
rect 42302 355250 42602 355251
rect 60302 355250 60602 355251
rect 78302 355250 78602 355251
rect 96302 355250 96602 355251
rect 114302 355250 114602 355251
rect 132302 355250 132602 355251
rect 150302 355250 150602 355251
rect 168302 355250 168602 355251
rect 186302 355250 186602 355251
rect 204302 355250 204602 355251
rect 222302 355250 222602 355251
rect 240302 355250 240602 355251
rect 258302 355250 258602 355251
rect 276302 355250 276602 355251
rect 295480 355250 295780 355251
rect -3818 355239 295780 355250
rect -3818 355121 -3727 355239
rect -3609 355121 6393 355239
rect 6511 355121 24393 355239
rect 24511 355121 42393 355239
rect 42511 355121 60393 355239
rect 60511 355121 78393 355239
rect 78511 355121 96393 355239
rect 96511 355121 114393 355239
rect 114511 355121 132393 355239
rect 132511 355121 150393 355239
rect 150511 355121 168393 355239
rect 168511 355121 186393 355239
rect 186511 355121 204393 355239
rect 204511 355121 222393 355239
rect 222511 355121 240393 355239
rect 240511 355121 258393 355239
rect 258511 355121 276393 355239
rect 276511 355121 295571 355239
rect 295689 355121 295780 355239
rect -3818 355079 295780 355121
rect -3818 354961 -3727 355079
rect -3609 354961 6393 355079
rect 6511 354961 24393 355079
rect 24511 354961 42393 355079
rect 42511 354961 60393 355079
rect 60511 354961 78393 355079
rect 78511 354961 96393 355079
rect 96511 354961 114393 355079
rect 114511 354961 132393 355079
rect 132511 354961 150393 355079
rect 150511 354961 168393 355079
rect 168511 354961 186393 355079
rect 186511 354961 204393 355079
rect 204511 354961 222393 355079
rect 222511 354961 240393 355079
rect 240511 354961 258393 355079
rect 258511 354961 276393 355079
rect 276511 354961 295571 355079
rect 295689 354961 295780 355079
rect -3818 354950 295780 354961
rect -3818 354949 -3518 354950
rect 6302 354949 6602 354950
rect 24302 354949 24602 354950
rect 42302 354949 42602 354950
rect 60302 354949 60602 354950
rect 78302 354949 78602 354950
rect 96302 354949 96602 354950
rect 114302 354949 114602 354950
rect 132302 354949 132602 354950
rect 150302 354949 150602 354950
rect 168302 354949 168602 354950
rect 186302 354949 186602 354950
rect 204302 354949 204602 354950
rect 222302 354949 222602 354950
rect 240302 354949 240602 354950
rect 258302 354949 258602 354950
rect 276302 354949 276602 354950
rect 295480 354949 295780 354950
rect -3348 354780 -3048 354781
rect 13502 354780 13802 354781
rect 31502 354780 31802 354781
rect 49502 354780 49802 354781
rect 67502 354780 67802 354781
rect 85502 354780 85802 354781
rect 103502 354780 103802 354781
rect 121502 354780 121802 354781
rect 139502 354780 139802 354781
rect 157502 354780 157802 354781
rect 175502 354780 175802 354781
rect 193502 354780 193802 354781
rect 211502 354780 211802 354781
rect 229502 354780 229802 354781
rect 247502 354780 247802 354781
rect 265502 354780 265802 354781
rect 283502 354780 283802 354781
rect 295010 354780 295310 354781
rect -3348 354769 295310 354780
rect -3348 354651 -3257 354769
rect -3139 354651 13593 354769
rect 13711 354651 31593 354769
rect 31711 354651 49593 354769
rect 49711 354651 67593 354769
rect 67711 354651 85593 354769
rect 85711 354651 103593 354769
rect 103711 354651 121593 354769
rect 121711 354651 139593 354769
rect 139711 354651 157593 354769
rect 157711 354651 175593 354769
rect 175711 354651 193593 354769
rect 193711 354651 211593 354769
rect 211711 354651 229593 354769
rect 229711 354651 247593 354769
rect 247711 354651 265593 354769
rect 265711 354651 283593 354769
rect 283711 354651 295101 354769
rect 295219 354651 295310 354769
rect -3348 354609 295310 354651
rect -3348 354491 -3257 354609
rect -3139 354491 13593 354609
rect 13711 354491 31593 354609
rect 31711 354491 49593 354609
rect 49711 354491 67593 354609
rect 67711 354491 85593 354609
rect 85711 354491 103593 354609
rect 103711 354491 121593 354609
rect 121711 354491 139593 354609
rect 139711 354491 157593 354609
rect 157711 354491 175593 354609
rect 175711 354491 193593 354609
rect 193711 354491 211593 354609
rect 211711 354491 229593 354609
rect 229711 354491 247593 354609
rect 247711 354491 265593 354609
rect 265711 354491 283593 354609
rect 283711 354491 295101 354609
rect 295219 354491 295310 354609
rect -3348 354480 295310 354491
rect -3348 354479 -3048 354480
rect 13502 354479 13802 354480
rect 31502 354479 31802 354480
rect 49502 354479 49802 354480
rect 67502 354479 67802 354480
rect 85502 354479 85802 354480
rect 103502 354479 103802 354480
rect 121502 354479 121802 354480
rect 139502 354479 139802 354480
rect 157502 354479 157802 354480
rect 175502 354479 175802 354480
rect 193502 354479 193802 354480
rect 211502 354479 211802 354480
rect 229502 354479 229802 354480
rect 247502 354479 247802 354480
rect 265502 354479 265802 354480
rect 283502 354479 283802 354480
rect 295010 354479 295310 354480
rect -2878 354310 -2578 354311
rect 4502 354310 4802 354311
rect 22502 354310 22802 354311
rect 40502 354310 40802 354311
rect 58502 354310 58802 354311
rect 76502 354310 76802 354311
rect 94502 354310 94802 354311
rect 112502 354310 112802 354311
rect 130502 354310 130802 354311
rect 148502 354310 148802 354311
rect 166502 354310 166802 354311
rect 184502 354310 184802 354311
rect 202502 354310 202802 354311
rect 220502 354310 220802 354311
rect 238502 354310 238802 354311
rect 256502 354310 256802 354311
rect 274502 354310 274802 354311
rect 294540 354310 294840 354311
rect -2878 354299 294840 354310
rect -2878 354181 -2787 354299
rect -2669 354181 4593 354299
rect 4711 354181 22593 354299
rect 22711 354181 40593 354299
rect 40711 354181 58593 354299
rect 58711 354181 76593 354299
rect 76711 354181 94593 354299
rect 94711 354181 112593 354299
rect 112711 354181 130593 354299
rect 130711 354181 148593 354299
rect 148711 354181 166593 354299
rect 166711 354181 184593 354299
rect 184711 354181 202593 354299
rect 202711 354181 220593 354299
rect 220711 354181 238593 354299
rect 238711 354181 256593 354299
rect 256711 354181 274593 354299
rect 274711 354181 294631 354299
rect 294749 354181 294840 354299
rect -2878 354139 294840 354181
rect -2878 354021 -2787 354139
rect -2669 354021 4593 354139
rect 4711 354021 22593 354139
rect 22711 354021 40593 354139
rect 40711 354021 58593 354139
rect 58711 354021 76593 354139
rect 76711 354021 94593 354139
rect 94711 354021 112593 354139
rect 112711 354021 130593 354139
rect 130711 354021 148593 354139
rect 148711 354021 166593 354139
rect 166711 354021 184593 354139
rect 184711 354021 202593 354139
rect 202711 354021 220593 354139
rect 220711 354021 238593 354139
rect 238711 354021 256593 354139
rect 256711 354021 274593 354139
rect 274711 354021 294631 354139
rect 294749 354021 294840 354139
rect -2878 354010 294840 354021
rect -2878 354009 -2578 354010
rect 4502 354009 4802 354010
rect 22502 354009 22802 354010
rect 40502 354009 40802 354010
rect 58502 354009 58802 354010
rect 76502 354009 76802 354010
rect 94502 354009 94802 354010
rect 112502 354009 112802 354010
rect 130502 354009 130802 354010
rect 148502 354009 148802 354010
rect 166502 354009 166802 354010
rect 184502 354009 184802 354010
rect 202502 354009 202802 354010
rect 220502 354009 220802 354010
rect 238502 354009 238802 354010
rect 256502 354009 256802 354010
rect 274502 354009 274802 354010
rect 294540 354009 294840 354010
rect -2408 353840 -2108 353841
rect 11702 353840 12002 353841
rect 29702 353840 30002 353841
rect 47702 353840 48002 353841
rect 65702 353840 66002 353841
rect 83702 353840 84002 353841
rect 101702 353840 102002 353841
rect 119702 353840 120002 353841
rect 137702 353840 138002 353841
rect 155702 353840 156002 353841
rect 173702 353840 174002 353841
rect 191702 353840 192002 353841
rect 209702 353840 210002 353841
rect 227702 353840 228002 353841
rect 245702 353840 246002 353841
rect 263702 353840 264002 353841
rect 281702 353840 282002 353841
rect 294070 353840 294370 353841
rect -2408 353829 294370 353840
rect -2408 353711 -2317 353829
rect -2199 353711 11793 353829
rect 11911 353711 29793 353829
rect 29911 353711 47793 353829
rect 47911 353711 65793 353829
rect 65911 353711 83793 353829
rect 83911 353711 101793 353829
rect 101911 353711 119793 353829
rect 119911 353711 137793 353829
rect 137911 353711 155793 353829
rect 155911 353711 173793 353829
rect 173911 353711 191793 353829
rect 191911 353711 209793 353829
rect 209911 353711 227793 353829
rect 227911 353711 245793 353829
rect 245911 353711 263793 353829
rect 263911 353711 281793 353829
rect 281911 353711 294161 353829
rect 294279 353711 294370 353829
rect -2408 353669 294370 353711
rect -2408 353551 -2317 353669
rect -2199 353551 11793 353669
rect 11911 353551 29793 353669
rect 29911 353551 47793 353669
rect 47911 353551 65793 353669
rect 65911 353551 83793 353669
rect 83911 353551 101793 353669
rect 101911 353551 119793 353669
rect 119911 353551 137793 353669
rect 137911 353551 155793 353669
rect 155911 353551 173793 353669
rect 173911 353551 191793 353669
rect 191911 353551 209793 353669
rect 209911 353551 227793 353669
rect 227911 353551 245793 353669
rect 245911 353551 263793 353669
rect 263911 353551 281793 353669
rect 281911 353551 294161 353669
rect 294279 353551 294370 353669
rect -2408 353540 294370 353551
rect -2408 353539 -2108 353540
rect 11702 353539 12002 353540
rect 29702 353539 30002 353540
rect 47702 353539 48002 353540
rect 65702 353539 66002 353540
rect 83702 353539 84002 353540
rect 101702 353539 102002 353540
rect 119702 353539 120002 353540
rect 137702 353539 138002 353540
rect 155702 353539 156002 353540
rect 173702 353539 174002 353540
rect 191702 353539 192002 353540
rect 209702 353539 210002 353540
rect 227702 353539 228002 353540
rect 245702 353539 246002 353540
rect 263702 353539 264002 353540
rect 281702 353539 282002 353540
rect 294070 353539 294370 353540
rect -1938 353370 -1638 353371
rect 2702 353370 3002 353371
rect 20702 353370 21002 353371
rect 38702 353370 39002 353371
rect 56702 353370 57002 353371
rect 74702 353370 75002 353371
rect 92702 353370 93002 353371
rect 110702 353370 111002 353371
rect 128702 353370 129002 353371
rect 146702 353370 147002 353371
rect 164702 353370 165002 353371
rect 182702 353370 183002 353371
rect 200702 353370 201002 353371
rect 218702 353370 219002 353371
rect 236702 353370 237002 353371
rect 254702 353370 255002 353371
rect 272702 353370 273002 353371
rect 290702 353370 291002 353371
rect 293600 353370 293900 353371
rect -1938 353359 293900 353370
rect -1938 353241 -1847 353359
rect -1729 353241 2793 353359
rect 2911 353241 20793 353359
rect 20911 353241 38793 353359
rect 38911 353241 56793 353359
rect 56911 353241 74793 353359
rect 74911 353241 92793 353359
rect 92911 353241 110793 353359
rect 110911 353241 128793 353359
rect 128911 353241 146793 353359
rect 146911 353241 164793 353359
rect 164911 353241 182793 353359
rect 182911 353241 200793 353359
rect 200911 353241 218793 353359
rect 218911 353241 236793 353359
rect 236911 353241 254793 353359
rect 254911 353241 272793 353359
rect 272911 353241 290793 353359
rect 290911 353241 293691 353359
rect 293809 353241 293900 353359
rect -1938 353199 293900 353241
rect -1938 353081 -1847 353199
rect -1729 353081 2793 353199
rect 2911 353081 20793 353199
rect 20911 353081 38793 353199
rect 38911 353081 56793 353199
rect 56911 353081 74793 353199
rect 74911 353081 92793 353199
rect 92911 353081 110793 353199
rect 110911 353081 128793 353199
rect 128911 353081 146793 353199
rect 146911 353081 164793 353199
rect 164911 353081 182793 353199
rect 182911 353081 200793 353199
rect 200911 353081 218793 353199
rect 218911 353081 236793 353199
rect 236911 353081 254793 353199
rect 254911 353081 272793 353199
rect 272911 353081 290793 353199
rect 290911 353081 293691 353199
rect 293809 353081 293900 353199
rect -1938 353070 293900 353081
rect -1938 353069 -1638 353070
rect 2702 353069 3002 353070
rect 20702 353069 21002 353070
rect 38702 353069 39002 353070
rect 56702 353069 57002 353070
rect 74702 353069 75002 353070
rect 92702 353069 93002 353070
rect 110702 353069 111002 353070
rect 128702 353069 129002 353070
rect 146702 353069 147002 353070
rect 164702 353069 165002 353070
rect 182702 353069 183002 353070
rect 200702 353069 201002 353070
rect 218702 353069 219002 353070
rect 236702 353069 237002 353070
rect 254702 353069 255002 353070
rect 272702 353069 273002 353070
rect 290702 353069 291002 353070
rect 293600 353069 293900 353070
rect -1468 352900 -1168 352901
rect 9902 352900 10202 352901
rect 27902 352900 28202 352901
rect 45902 352900 46202 352901
rect 63902 352900 64202 352901
rect 81902 352900 82202 352901
rect 99902 352900 100202 352901
rect 117902 352900 118202 352901
rect 135902 352900 136202 352901
rect 153902 352900 154202 352901
rect 171902 352900 172202 352901
rect 189902 352900 190202 352901
rect 207902 352900 208202 352901
rect 225902 352900 226202 352901
rect 243902 352900 244202 352901
rect 261902 352900 262202 352901
rect 279902 352900 280202 352901
rect 293130 352900 293430 352901
rect -1468 352889 293430 352900
rect -1468 352771 -1377 352889
rect -1259 352771 9993 352889
rect 10111 352771 27993 352889
rect 28111 352771 45993 352889
rect 46111 352771 63993 352889
rect 64111 352771 81993 352889
rect 82111 352771 99993 352889
rect 100111 352771 117993 352889
rect 118111 352771 135993 352889
rect 136111 352771 153993 352889
rect 154111 352771 171993 352889
rect 172111 352771 189993 352889
rect 190111 352771 207993 352889
rect 208111 352771 225993 352889
rect 226111 352771 243993 352889
rect 244111 352771 261993 352889
rect 262111 352771 279993 352889
rect 280111 352771 293221 352889
rect 293339 352771 293430 352889
rect -1468 352729 293430 352771
rect -1468 352611 -1377 352729
rect -1259 352611 9993 352729
rect 10111 352611 27993 352729
rect 28111 352611 45993 352729
rect 46111 352611 63993 352729
rect 64111 352611 81993 352729
rect 82111 352611 99993 352729
rect 100111 352611 117993 352729
rect 118111 352611 135993 352729
rect 136111 352611 153993 352729
rect 154111 352611 171993 352729
rect 172111 352611 189993 352729
rect 190111 352611 207993 352729
rect 208111 352611 225993 352729
rect 226111 352611 243993 352729
rect 244111 352611 261993 352729
rect 262111 352611 279993 352729
rect 280111 352611 293221 352729
rect 293339 352611 293430 352729
rect -1468 352600 293430 352611
rect -1468 352599 -1168 352600
rect 9902 352599 10202 352600
rect 27902 352599 28202 352600
rect 45902 352599 46202 352600
rect 63902 352599 64202 352600
rect 81902 352599 82202 352600
rect 99902 352599 100202 352600
rect 117902 352599 118202 352600
rect 135902 352599 136202 352600
rect 153902 352599 154202 352600
rect 171902 352599 172202 352600
rect 189902 352599 190202 352600
rect 207902 352599 208202 352600
rect 225902 352599 226202 352600
rect 243902 352599 244202 352600
rect 261902 352599 262202 352600
rect 279902 352599 280202 352600
rect 293130 352599 293430 352600
rect -998 352430 -698 352431
rect 902 352430 1202 352431
rect 18902 352430 19202 352431
rect 36902 352430 37202 352431
rect 54902 352430 55202 352431
rect 72902 352430 73202 352431
rect 90902 352430 91202 352431
rect 108902 352430 109202 352431
rect 126902 352430 127202 352431
rect 144902 352430 145202 352431
rect 162902 352430 163202 352431
rect 180902 352430 181202 352431
rect 198902 352430 199202 352431
rect 216902 352430 217202 352431
rect 234902 352430 235202 352431
rect 252902 352430 253202 352431
rect 270902 352430 271202 352431
rect 288902 352430 289202 352431
rect 292660 352430 292960 352431
rect -998 352419 292960 352430
rect -998 352301 -907 352419
rect -789 352301 993 352419
rect 1111 352301 18993 352419
rect 19111 352301 36993 352419
rect 37111 352301 54993 352419
rect 55111 352301 72993 352419
rect 73111 352301 90993 352419
rect 91111 352301 108993 352419
rect 109111 352301 126993 352419
rect 127111 352301 144993 352419
rect 145111 352301 162993 352419
rect 163111 352301 180993 352419
rect 181111 352301 198993 352419
rect 199111 352301 216993 352419
rect 217111 352301 234993 352419
rect 235111 352301 252993 352419
rect 253111 352301 270993 352419
rect 271111 352301 288993 352419
rect 289111 352301 292751 352419
rect 292869 352301 292960 352419
rect -998 352259 292960 352301
rect -998 352141 -907 352259
rect -789 352141 993 352259
rect 1111 352141 18993 352259
rect 19111 352141 36993 352259
rect 37111 352141 54993 352259
rect 55111 352141 72993 352259
rect 73111 352141 90993 352259
rect 91111 352141 108993 352259
rect 109111 352141 126993 352259
rect 127111 352141 144993 352259
rect 145111 352141 162993 352259
rect 163111 352141 180993 352259
rect 181111 352141 198993 352259
rect 199111 352141 216993 352259
rect 217111 352141 234993 352259
rect 235111 352141 252993 352259
rect 253111 352141 270993 352259
rect 271111 352141 288993 352259
rect 289111 352141 292751 352259
rect 292869 352141 292960 352259
rect -998 352130 292960 352141
rect -998 352129 -698 352130
rect 902 352129 1202 352130
rect 18902 352129 19202 352130
rect 36902 352129 37202 352130
rect 54902 352129 55202 352130
rect 72902 352129 73202 352130
rect 90902 352129 91202 352130
rect 108902 352129 109202 352130
rect 126902 352129 127202 352130
rect 144902 352129 145202 352130
rect 162902 352129 163202 352130
rect 180902 352129 181202 352130
rect 198902 352129 199202 352130
rect 216902 352129 217202 352130
rect 234902 352129 235202 352130
rect 252902 352129 253202 352130
rect 270902 352129 271202 352130
rect 288902 352129 289202 352130
rect 292660 352129 292960 352130
rect -3818 349138 -3518 349139
rect 6302 349138 6602 349139
rect 24302 349138 24602 349139
rect 42302 349138 42602 349139
rect 60302 349138 60602 349139
rect 78302 349138 78602 349139
rect 96302 349138 96602 349139
rect 114302 349138 114602 349139
rect 132302 349138 132602 349139
rect 150302 349138 150602 349139
rect 168302 349138 168602 349139
rect 186302 349138 186602 349139
rect 204302 349138 204602 349139
rect 222302 349138 222602 349139
rect 240302 349138 240602 349139
rect 258302 349138 258602 349139
rect 276302 349138 276602 349139
rect 295480 349138 295780 349139
rect -4288 349127 296250 349138
rect -4288 349009 -3727 349127
rect -3609 349009 6393 349127
rect 6511 349009 24393 349127
rect 24511 349009 42393 349127
rect 42511 349009 60393 349127
rect 60511 349009 78393 349127
rect 78511 349009 96393 349127
rect 96511 349009 114393 349127
rect 114511 349009 132393 349127
rect 132511 349009 150393 349127
rect 150511 349009 168393 349127
rect 168511 349009 186393 349127
rect 186511 349009 204393 349127
rect 204511 349009 222393 349127
rect 222511 349009 240393 349127
rect 240511 349009 258393 349127
rect 258511 349009 276393 349127
rect 276511 349009 295571 349127
rect 295689 349009 296250 349127
rect -4288 348967 296250 349009
rect -4288 348849 -3727 348967
rect -3609 348849 6393 348967
rect 6511 348849 24393 348967
rect 24511 348849 42393 348967
rect 42511 348849 60393 348967
rect 60511 348849 78393 348967
rect 78511 348849 96393 348967
rect 96511 348849 114393 348967
rect 114511 348849 132393 348967
rect 132511 348849 150393 348967
rect 150511 348849 168393 348967
rect 168511 348849 186393 348967
rect 186511 348849 204393 348967
rect 204511 348849 222393 348967
rect 222511 348849 240393 348967
rect 240511 348849 258393 348967
rect 258511 348849 276393 348967
rect 276511 348849 295571 348967
rect 295689 348849 296250 348967
rect -4288 348838 296250 348849
rect -3818 348837 -3518 348838
rect 6302 348837 6602 348838
rect 24302 348837 24602 348838
rect 42302 348837 42602 348838
rect 60302 348837 60602 348838
rect 78302 348837 78602 348838
rect 96302 348837 96602 348838
rect 114302 348837 114602 348838
rect 132302 348837 132602 348838
rect 150302 348837 150602 348838
rect 168302 348837 168602 348838
rect 186302 348837 186602 348838
rect 204302 348837 204602 348838
rect 222302 348837 222602 348838
rect 240302 348837 240602 348838
rect 258302 348837 258602 348838
rect 276302 348837 276602 348838
rect 295480 348837 295780 348838
rect -2878 347338 -2578 347339
rect 4502 347338 4802 347339
rect 22502 347338 22802 347339
rect 40502 347338 40802 347339
rect 58502 347338 58802 347339
rect 76502 347338 76802 347339
rect 94502 347338 94802 347339
rect 112502 347338 112802 347339
rect 130502 347338 130802 347339
rect 148502 347338 148802 347339
rect 166502 347338 166802 347339
rect 184502 347338 184802 347339
rect 202502 347338 202802 347339
rect 220502 347338 220802 347339
rect 238502 347338 238802 347339
rect 256502 347338 256802 347339
rect 274502 347338 274802 347339
rect 294540 347338 294840 347339
rect -3348 347327 295310 347338
rect -3348 347209 -2787 347327
rect -2669 347209 4593 347327
rect 4711 347209 22593 347327
rect 22711 347209 40593 347327
rect 40711 347209 58593 347327
rect 58711 347209 76593 347327
rect 76711 347209 94593 347327
rect 94711 347209 112593 347327
rect 112711 347209 130593 347327
rect 130711 347209 148593 347327
rect 148711 347209 166593 347327
rect 166711 347209 184593 347327
rect 184711 347209 202593 347327
rect 202711 347209 220593 347327
rect 220711 347209 238593 347327
rect 238711 347209 256593 347327
rect 256711 347209 274593 347327
rect 274711 347209 294631 347327
rect 294749 347209 295310 347327
rect -3348 347167 295310 347209
rect -3348 347049 -2787 347167
rect -2669 347049 4593 347167
rect 4711 347049 22593 347167
rect 22711 347049 40593 347167
rect 40711 347049 58593 347167
rect 58711 347049 76593 347167
rect 76711 347049 94593 347167
rect 94711 347049 112593 347167
rect 112711 347049 130593 347167
rect 130711 347049 148593 347167
rect 148711 347049 166593 347167
rect 166711 347049 184593 347167
rect 184711 347049 202593 347167
rect 202711 347049 220593 347167
rect 220711 347049 238593 347167
rect 238711 347049 256593 347167
rect 256711 347049 274593 347167
rect 274711 347049 294631 347167
rect 294749 347049 295310 347167
rect -3348 347038 295310 347049
rect -2878 347037 -2578 347038
rect 4502 347037 4802 347038
rect 22502 347037 22802 347038
rect 40502 347037 40802 347038
rect 58502 347037 58802 347038
rect 76502 347037 76802 347038
rect 94502 347037 94802 347038
rect 112502 347037 112802 347038
rect 130502 347037 130802 347038
rect 148502 347037 148802 347038
rect 166502 347037 166802 347038
rect 184502 347037 184802 347038
rect 202502 347037 202802 347038
rect 220502 347037 220802 347038
rect 238502 347037 238802 347038
rect 256502 347037 256802 347038
rect 274502 347037 274802 347038
rect 294540 347037 294840 347038
rect -1938 345538 -1638 345539
rect 2702 345538 3002 345539
rect 20702 345538 21002 345539
rect 38702 345538 39002 345539
rect 56702 345538 57002 345539
rect 74702 345538 75002 345539
rect 92702 345538 93002 345539
rect 110702 345538 111002 345539
rect 128702 345538 129002 345539
rect 146702 345538 147002 345539
rect 164702 345538 165002 345539
rect 182702 345538 183002 345539
rect 200702 345538 201002 345539
rect 218702 345538 219002 345539
rect 236702 345538 237002 345539
rect 254702 345538 255002 345539
rect 272702 345538 273002 345539
rect 290702 345538 291002 345539
rect 293600 345538 293900 345539
rect -2408 345527 294370 345538
rect -2408 345409 -1847 345527
rect -1729 345409 2793 345527
rect 2911 345409 20793 345527
rect 20911 345409 38793 345527
rect 38911 345409 56793 345527
rect 56911 345409 74793 345527
rect 74911 345409 92793 345527
rect 92911 345409 110793 345527
rect 110911 345409 128793 345527
rect 128911 345409 146793 345527
rect 146911 345409 164793 345527
rect 164911 345409 182793 345527
rect 182911 345409 200793 345527
rect 200911 345409 218793 345527
rect 218911 345409 236793 345527
rect 236911 345409 254793 345527
rect 254911 345409 272793 345527
rect 272911 345409 290793 345527
rect 290911 345409 293691 345527
rect 293809 345409 294370 345527
rect -2408 345367 294370 345409
rect -2408 345249 -1847 345367
rect -1729 345249 2793 345367
rect 2911 345249 20793 345367
rect 20911 345249 38793 345367
rect 38911 345249 56793 345367
rect 56911 345249 74793 345367
rect 74911 345249 92793 345367
rect 92911 345249 110793 345367
rect 110911 345249 128793 345367
rect 128911 345249 146793 345367
rect 146911 345249 164793 345367
rect 164911 345249 182793 345367
rect 182911 345249 200793 345367
rect 200911 345249 218793 345367
rect 218911 345249 236793 345367
rect 236911 345249 254793 345367
rect 254911 345249 272793 345367
rect 272911 345249 290793 345367
rect 290911 345249 293691 345367
rect 293809 345249 294370 345367
rect -2408 345238 294370 345249
rect -1938 345237 -1638 345238
rect 2702 345237 3002 345238
rect 20702 345237 21002 345238
rect 38702 345237 39002 345238
rect 56702 345237 57002 345238
rect 74702 345237 75002 345238
rect 92702 345237 93002 345238
rect 110702 345237 111002 345238
rect 128702 345237 129002 345238
rect 146702 345237 147002 345238
rect 164702 345237 165002 345238
rect 182702 345237 183002 345238
rect 200702 345237 201002 345238
rect 218702 345237 219002 345238
rect 236702 345237 237002 345238
rect 254702 345237 255002 345238
rect 272702 345237 273002 345238
rect 290702 345237 291002 345238
rect 293600 345237 293900 345238
rect -998 343738 -698 343739
rect 902 343738 1202 343739
rect 18902 343738 19202 343739
rect 36902 343738 37202 343739
rect 54902 343738 55202 343739
rect 72902 343738 73202 343739
rect 90902 343738 91202 343739
rect 108902 343738 109202 343739
rect 126902 343738 127202 343739
rect 144902 343738 145202 343739
rect 162902 343738 163202 343739
rect 180902 343738 181202 343739
rect 198902 343738 199202 343739
rect 216902 343738 217202 343739
rect 234902 343738 235202 343739
rect 252902 343738 253202 343739
rect 270902 343738 271202 343739
rect 288902 343738 289202 343739
rect 292660 343738 292960 343739
rect -1468 343727 293430 343738
rect -1468 343609 -907 343727
rect -789 343609 993 343727
rect 1111 343609 18993 343727
rect 19111 343609 36993 343727
rect 37111 343609 54993 343727
rect 55111 343609 72993 343727
rect 73111 343609 90993 343727
rect 91111 343609 108993 343727
rect 109111 343609 126993 343727
rect 127111 343609 144993 343727
rect 145111 343609 162993 343727
rect 163111 343609 180993 343727
rect 181111 343609 198993 343727
rect 199111 343609 216993 343727
rect 217111 343609 234993 343727
rect 235111 343609 252993 343727
rect 253111 343609 270993 343727
rect 271111 343609 288993 343727
rect 289111 343609 292751 343727
rect 292869 343609 293430 343727
rect -1468 343567 293430 343609
rect -1468 343449 -907 343567
rect -789 343449 993 343567
rect 1111 343449 18993 343567
rect 19111 343449 36993 343567
rect 37111 343449 54993 343567
rect 55111 343449 72993 343567
rect 73111 343449 90993 343567
rect 91111 343449 108993 343567
rect 109111 343449 126993 343567
rect 127111 343449 144993 343567
rect 145111 343449 162993 343567
rect 163111 343449 180993 343567
rect 181111 343449 198993 343567
rect 199111 343449 216993 343567
rect 217111 343449 234993 343567
rect 235111 343449 252993 343567
rect 253111 343449 270993 343567
rect 271111 343449 288993 343567
rect 289111 343449 292751 343567
rect 292869 343449 293430 343567
rect -1468 343438 293430 343449
rect -998 343437 -698 343438
rect 902 343437 1202 343438
rect 18902 343437 19202 343438
rect 36902 343437 37202 343438
rect 54902 343437 55202 343438
rect 72902 343437 73202 343438
rect 90902 343437 91202 343438
rect 108902 343437 109202 343438
rect 126902 343437 127202 343438
rect 144902 343437 145202 343438
rect 162902 343437 163202 343438
rect 180902 343437 181202 343438
rect 198902 343437 199202 343438
rect 216902 343437 217202 343438
rect 234902 343437 235202 343438
rect 252902 343437 253202 343438
rect 270902 343437 271202 343438
rect 288902 343437 289202 343438
rect 292660 343437 292960 343438
rect -4288 340138 -3988 340139
rect 15302 340138 15602 340139
rect 33302 340138 33602 340139
rect 51302 340138 51602 340139
rect 69302 340138 69602 340139
rect 87302 340138 87602 340139
rect 105302 340138 105602 340139
rect 123302 340138 123602 340139
rect 141302 340138 141602 340139
rect 159302 340138 159602 340139
rect 177302 340138 177602 340139
rect 195302 340138 195602 340139
rect 213302 340138 213602 340139
rect 231302 340138 231602 340139
rect 249302 340138 249602 340139
rect 267302 340138 267602 340139
rect 285302 340138 285602 340139
rect 295950 340138 296250 340139
rect -4288 340127 296250 340138
rect -4288 340009 -4197 340127
rect -4079 340009 15393 340127
rect 15511 340009 33393 340127
rect 33511 340009 51393 340127
rect 51511 340009 69393 340127
rect 69511 340009 87393 340127
rect 87511 340009 105393 340127
rect 105511 340009 123393 340127
rect 123511 340009 141393 340127
rect 141511 340009 159393 340127
rect 159511 340009 177393 340127
rect 177511 340009 195393 340127
rect 195511 340009 213393 340127
rect 213511 340009 231393 340127
rect 231511 340009 249393 340127
rect 249511 340009 267393 340127
rect 267511 340009 285393 340127
rect 285511 340009 296041 340127
rect 296159 340009 296250 340127
rect -4288 339967 296250 340009
rect -4288 339849 -4197 339967
rect -4079 339849 15393 339967
rect 15511 339849 33393 339967
rect 33511 339849 51393 339967
rect 51511 339849 69393 339967
rect 69511 339849 87393 339967
rect 87511 339849 105393 339967
rect 105511 339849 123393 339967
rect 123511 339849 141393 339967
rect 141511 339849 159393 339967
rect 159511 339849 177393 339967
rect 177511 339849 195393 339967
rect 195511 339849 213393 339967
rect 213511 339849 231393 339967
rect 231511 339849 249393 339967
rect 249511 339849 267393 339967
rect 267511 339849 285393 339967
rect 285511 339849 296041 339967
rect 296159 339849 296250 339967
rect -4288 339838 296250 339849
rect -4288 339837 -3988 339838
rect 15302 339837 15602 339838
rect 33302 339837 33602 339838
rect 51302 339837 51602 339838
rect 69302 339837 69602 339838
rect 87302 339837 87602 339838
rect 105302 339837 105602 339838
rect 123302 339837 123602 339838
rect 141302 339837 141602 339838
rect 159302 339837 159602 339838
rect 177302 339837 177602 339838
rect 195302 339837 195602 339838
rect 213302 339837 213602 339838
rect 231302 339837 231602 339838
rect 249302 339837 249602 339838
rect 267302 339837 267602 339838
rect 285302 339837 285602 339838
rect 295950 339837 296250 339838
rect -3348 338338 -3048 338339
rect 13502 338338 13802 338339
rect 31502 338338 31802 338339
rect 49502 338338 49802 338339
rect 67502 338338 67802 338339
rect 85502 338338 85802 338339
rect 103502 338338 103802 338339
rect 121502 338338 121802 338339
rect 139502 338338 139802 338339
rect 157502 338338 157802 338339
rect 175502 338338 175802 338339
rect 193502 338338 193802 338339
rect 211502 338338 211802 338339
rect 229502 338338 229802 338339
rect 247502 338338 247802 338339
rect 265502 338338 265802 338339
rect 283502 338338 283802 338339
rect 295010 338338 295310 338339
rect -3348 338327 295310 338338
rect -3348 338209 -3257 338327
rect -3139 338209 13593 338327
rect 13711 338209 31593 338327
rect 31711 338209 49593 338327
rect 49711 338209 67593 338327
rect 67711 338209 85593 338327
rect 85711 338209 103593 338327
rect 103711 338209 121593 338327
rect 121711 338209 139593 338327
rect 139711 338209 157593 338327
rect 157711 338209 175593 338327
rect 175711 338209 193593 338327
rect 193711 338209 211593 338327
rect 211711 338209 229593 338327
rect 229711 338209 247593 338327
rect 247711 338209 265593 338327
rect 265711 338209 283593 338327
rect 283711 338209 295101 338327
rect 295219 338209 295310 338327
rect -3348 338167 295310 338209
rect -3348 338049 -3257 338167
rect -3139 338049 13593 338167
rect 13711 338049 31593 338167
rect 31711 338049 49593 338167
rect 49711 338049 67593 338167
rect 67711 338049 85593 338167
rect 85711 338049 103593 338167
rect 103711 338049 121593 338167
rect 121711 338049 139593 338167
rect 139711 338049 157593 338167
rect 157711 338049 175593 338167
rect 175711 338049 193593 338167
rect 193711 338049 211593 338167
rect 211711 338049 229593 338167
rect 229711 338049 247593 338167
rect 247711 338049 265593 338167
rect 265711 338049 283593 338167
rect 283711 338049 295101 338167
rect 295219 338049 295310 338167
rect -3348 338038 295310 338049
rect -3348 338037 -3048 338038
rect 13502 338037 13802 338038
rect 31502 338037 31802 338038
rect 49502 338037 49802 338038
rect 67502 338037 67802 338038
rect 85502 338037 85802 338038
rect 103502 338037 103802 338038
rect 121502 338037 121802 338038
rect 139502 338037 139802 338038
rect 157502 338037 157802 338038
rect 175502 338037 175802 338038
rect 193502 338037 193802 338038
rect 211502 338037 211802 338038
rect 229502 338037 229802 338038
rect 247502 338037 247802 338038
rect 265502 338037 265802 338038
rect 283502 338037 283802 338038
rect 295010 338037 295310 338038
rect -2408 336538 -2108 336539
rect 11702 336538 12002 336539
rect 29702 336538 30002 336539
rect 47702 336538 48002 336539
rect 65702 336538 66002 336539
rect 83702 336538 84002 336539
rect 101702 336538 102002 336539
rect 119702 336538 120002 336539
rect 137702 336538 138002 336539
rect 155702 336538 156002 336539
rect 173702 336538 174002 336539
rect 191702 336538 192002 336539
rect 209702 336538 210002 336539
rect 227702 336538 228002 336539
rect 245702 336538 246002 336539
rect 263702 336538 264002 336539
rect 281702 336538 282002 336539
rect 294070 336538 294370 336539
rect -2408 336527 294370 336538
rect -2408 336409 -2317 336527
rect -2199 336409 11793 336527
rect 11911 336409 29793 336527
rect 29911 336409 47793 336527
rect 47911 336409 65793 336527
rect 65911 336409 83793 336527
rect 83911 336409 101793 336527
rect 101911 336409 119793 336527
rect 119911 336409 137793 336527
rect 137911 336409 155793 336527
rect 155911 336409 173793 336527
rect 173911 336409 191793 336527
rect 191911 336409 209793 336527
rect 209911 336409 227793 336527
rect 227911 336409 245793 336527
rect 245911 336409 263793 336527
rect 263911 336409 281793 336527
rect 281911 336409 294161 336527
rect 294279 336409 294370 336527
rect -2408 336367 294370 336409
rect -2408 336249 -2317 336367
rect -2199 336249 11793 336367
rect 11911 336249 29793 336367
rect 29911 336249 47793 336367
rect 47911 336249 65793 336367
rect 65911 336249 83793 336367
rect 83911 336249 101793 336367
rect 101911 336249 119793 336367
rect 119911 336249 137793 336367
rect 137911 336249 155793 336367
rect 155911 336249 173793 336367
rect 173911 336249 191793 336367
rect 191911 336249 209793 336367
rect 209911 336249 227793 336367
rect 227911 336249 245793 336367
rect 245911 336249 263793 336367
rect 263911 336249 281793 336367
rect 281911 336249 294161 336367
rect 294279 336249 294370 336367
rect -2408 336238 294370 336249
rect -2408 336237 -2108 336238
rect 11702 336237 12002 336238
rect 29702 336237 30002 336238
rect 47702 336237 48002 336238
rect 65702 336237 66002 336238
rect 83702 336237 84002 336238
rect 101702 336237 102002 336238
rect 119702 336237 120002 336238
rect 137702 336237 138002 336238
rect 155702 336237 156002 336238
rect 173702 336237 174002 336238
rect 191702 336237 192002 336238
rect 209702 336237 210002 336238
rect 227702 336237 228002 336238
rect 245702 336237 246002 336238
rect 263702 336237 264002 336238
rect 281702 336237 282002 336238
rect 294070 336237 294370 336238
rect -1468 334738 -1168 334739
rect 9902 334738 10202 334739
rect 27902 334738 28202 334739
rect 45902 334738 46202 334739
rect 63902 334738 64202 334739
rect 81902 334738 82202 334739
rect 99902 334738 100202 334739
rect 117902 334738 118202 334739
rect 135902 334738 136202 334739
rect 153902 334738 154202 334739
rect 171902 334738 172202 334739
rect 189902 334738 190202 334739
rect 207902 334738 208202 334739
rect 225902 334738 226202 334739
rect 243902 334738 244202 334739
rect 261902 334738 262202 334739
rect 279902 334738 280202 334739
rect 293130 334738 293430 334739
rect -1468 334727 293430 334738
rect -1468 334609 -1377 334727
rect -1259 334609 9993 334727
rect 10111 334609 27993 334727
rect 28111 334609 45993 334727
rect 46111 334609 63993 334727
rect 64111 334609 81993 334727
rect 82111 334609 99993 334727
rect 100111 334609 117993 334727
rect 118111 334609 135993 334727
rect 136111 334609 153993 334727
rect 154111 334609 171993 334727
rect 172111 334609 189993 334727
rect 190111 334609 207993 334727
rect 208111 334609 225993 334727
rect 226111 334609 243993 334727
rect 244111 334609 261993 334727
rect 262111 334609 279993 334727
rect 280111 334609 293221 334727
rect 293339 334609 293430 334727
rect -1468 334567 293430 334609
rect -1468 334449 -1377 334567
rect -1259 334449 9993 334567
rect 10111 334449 27993 334567
rect 28111 334449 45993 334567
rect 46111 334449 63993 334567
rect 64111 334449 81993 334567
rect 82111 334449 99993 334567
rect 100111 334449 117993 334567
rect 118111 334449 135993 334567
rect 136111 334449 153993 334567
rect 154111 334449 171993 334567
rect 172111 334449 189993 334567
rect 190111 334449 207993 334567
rect 208111 334449 225993 334567
rect 226111 334449 243993 334567
rect 244111 334449 261993 334567
rect 262111 334449 279993 334567
rect 280111 334449 293221 334567
rect 293339 334449 293430 334567
rect -1468 334438 293430 334449
rect -1468 334437 -1168 334438
rect 9902 334437 10202 334438
rect 27902 334437 28202 334438
rect 45902 334437 46202 334438
rect 63902 334437 64202 334438
rect 81902 334437 82202 334438
rect 99902 334437 100202 334438
rect 117902 334437 118202 334438
rect 135902 334437 136202 334438
rect 153902 334437 154202 334438
rect 171902 334437 172202 334438
rect 189902 334437 190202 334438
rect 207902 334437 208202 334438
rect 225902 334437 226202 334438
rect 243902 334437 244202 334438
rect 261902 334437 262202 334438
rect 279902 334437 280202 334438
rect 293130 334437 293430 334438
rect -3818 331138 -3518 331139
rect 6302 331138 6602 331139
rect 24302 331138 24602 331139
rect 42302 331138 42602 331139
rect 60302 331138 60602 331139
rect 78302 331138 78602 331139
rect 96302 331138 96602 331139
rect 114302 331138 114602 331139
rect 132302 331138 132602 331139
rect 150302 331138 150602 331139
rect 168302 331138 168602 331139
rect 186302 331138 186602 331139
rect 204302 331138 204602 331139
rect 222302 331138 222602 331139
rect 240302 331138 240602 331139
rect 258302 331138 258602 331139
rect 276302 331138 276602 331139
rect 295480 331138 295780 331139
rect -4288 331127 296250 331138
rect -4288 331009 -3727 331127
rect -3609 331009 6393 331127
rect 6511 331009 24393 331127
rect 24511 331009 42393 331127
rect 42511 331009 60393 331127
rect 60511 331009 78393 331127
rect 78511 331009 96393 331127
rect 96511 331009 114393 331127
rect 114511 331009 132393 331127
rect 132511 331009 150393 331127
rect 150511 331009 168393 331127
rect 168511 331009 186393 331127
rect 186511 331009 204393 331127
rect 204511 331009 222393 331127
rect 222511 331009 240393 331127
rect 240511 331009 258393 331127
rect 258511 331009 276393 331127
rect 276511 331009 295571 331127
rect 295689 331009 296250 331127
rect -4288 330967 296250 331009
rect -4288 330849 -3727 330967
rect -3609 330849 6393 330967
rect 6511 330849 24393 330967
rect 24511 330849 42393 330967
rect 42511 330849 60393 330967
rect 60511 330849 78393 330967
rect 78511 330849 96393 330967
rect 96511 330849 114393 330967
rect 114511 330849 132393 330967
rect 132511 330849 150393 330967
rect 150511 330849 168393 330967
rect 168511 330849 186393 330967
rect 186511 330849 204393 330967
rect 204511 330849 222393 330967
rect 222511 330849 240393 330967
rect 240511 330849 258393 330967
rect 258511 330849 276393 330967
rect 276511 330849 295571 330967
rect 295689 330849 296250 330967
rect -4288 330838 296250 330849
rect -3818 330837 -3518 330838
rect 6302 330837 6602 330838
rect 24302 330837 24602 330838
rect 42302 330837 42602 330838
rect 60302 330837 60602 330838
rect 78302 330837 78602 330838
rect 96302 330837 96602 330838
rect 114302 330837 114602 330838
rect 132302 330837 132602 330838
rect 150302 330837 150602 330838
rect 168302 330837 168602 330838
rect 186302 330837 186602 330838
rect 204302 330837 204602 330838
rect 222302 330837 222602 330838
rect 240302 330837 240602 330838
rect 258302 330837 258602 330838
rect 276302 330837 276602 330838
rect 295480 330837 295780 330838
rect -2878 329338 -2578 329339
rect 4502 329338 4802 329339
rect 22502 329338 22802 329339
rect 40502 329338 40802 329339
rect 58502 329338 58802 329339
rect 76502 329338 76802 329339
rect 94502 329338 94802 329339
rect 112502 329338 112802 329339
rect 130502 329338 130802 329339
rect 148502 329338 148802 329339
rect 166502 329338 166802 329339
rect 184502 329338 184802 329339
rect 202502 329338 202802 329339
rect 220502 329338 220802 329339
rect 238502 329338 238802 329339
rect 256502 329338 256802 329339
rect 274502 329338 274802 329339
rect 294540 329338 294840 329339
rect -3348 329327 295310 329338
rect -3348 329209 -2787 329327
rect -2669 329209 4593 329327
rect 4711 329209 22593 329327
rect 22711 329209 40593 329327
rect 40711 329209 58593 329327
rect 58711 329209 76593 329327
rect 76711 329209 94593 329327
rect 94711 329209 112593 329327
rect 112711 329209 130593 329327
rect 130711 329209 148593 329327
rect 148711 329209 166593 329327
rect 166711 329209 184593 329327
rect 184711 329209 202593 329327
rect 202711 329209 220593 329327
rect 220711 329209 238593 329327
rect 238711 329209 256593 329327
rect 256711 329209 274593 329327
rect 274711 329209 294631 329327
rect 294749 329209 295310 329327
rect -3348 329167 295310 329209
rect -3348 329049 -2787 329167
rect -2669 329049 4593 329167
rect 4711 329049 22593 329167
rect 22711 329049 40593 329167
rect 40711 329049 58593 329167
rect 58711 329049 76593 329167
rect 76711 329049 94593 329167
rect 94711 329049 112593 329167
rect 112711 329049 130593 329167
rect 130711 329049 148593 329167
rect 148711 329049 166593 329167
rect 166711 329049 184593 329167
rect 184711 329049 202593 329167
rect 202711 329049 220593 329167
rect 220711 329049 238593 329167
rect 238711 329049 256593 329167
rect 256711 329049 274593 329167
rect 274711 329049 294631 329167
rect 294749 329049 295310 329167
rect -3348 329038 295310 329049
rect -2878 329037 -2578 329038
rect 4502 329037 4802 329038
rect 22502 329037 22802 329038
rect 40502 329037 40802 329038
rect 58502 329037 58802 329038
rect 76502 329037 76802 329038
rect 94502 329037 94802 329038
rect 112502 329037 112802 329038
rect 130502 329037 130802 329038
rect 148502 329037 148802 329038
rect 166502 329037 166802 329038
rect 184502 329037 184802 329038
rect 202502 329037 202802 329038
rect 220502 329037 220802 329038
rect 238502 329037 238802 329038
rect 256502 329037 256802 329038
rect 274502 329037 274802 329038
rect 294540 329037 294840 329038
rect -1938 327538 -1638 327539
rect 2702 327538 3002 327539
rect 20702 327538 21002 327539
rect 38702 327538 39002 327539
rect 56702 327538 57002 327539
rect 74702 327538 75002 327539
rect 92702 327538 93002 327539
rect 110702 327538 111002 327539
rect 128702 327538 129002 327539
rect 146702 327538 147002 327539
rect 164702 327538 165002 327539
rect 182702 327538 183002 327539
rect 200702 327538 201002 327539
rect 218702 327538 219002 327539
rect 236702 327538 237002 327539
rect 254702 327538 255002 327539
rect 272702 327538 273002 327539
rect 290702 327538 291002 327539
rect 293600 327538 293900 327539
rect -2408 327527 294370 327538
rect -2408 327409 -1847 327527
rect -1729 327409 2793 327527
rect 2911 327409 20793 327527
rect 20911 327409 38793 327527
rect 38911 327409 56793 327527
rect 56911 327409 74793 327527
rect 74911 327409 92793 327527
rect 92911 327409 110793 327527
rect 110911 327409 128793 327527
rect 128911 327409 146793 327527
rect 146911 327409 164793 327527
rect 164911 327409 182793 327527
rect 182911 327409 200793 327527
rect 200911 327409 218793 327527
rect 218911 327409 236793 327527
rect 236911 327409 254793 327527
rect 254911 327409 272793 327527
rect 272911 327409 290793 327527
rect 290911 327409 293691 327527
rect 293809 327409 294370 327527
rect -2408 327367 294370 327409
rect -2408 327249 -1847 327367
rect -1729 327249 2793 327367
rect 2911 327249 20793 327367
rect 20911 327249 38793 327367
rect 38911 327249 56793 327367
rect 56911 327249 74793 327367
rect 74911 327249 92793 327367
rect 92911 327249 110793 327367
rect 110911 327249 128793 327367
rect 128911 327249 146793 327367
rect 146911 327249 164793 327367
rect 164911 327249 182793 327367
rect 182911 327249 200793 327367
rect 200911 327249 218793 327367
rect 218911 327249 236793 327367
rect 236911 327249 254793 327367
rect 254911 327249 272793 327367
rect 272911 327249 290793 327367
rect 290911 327249 293691 327367
rect 293809 327249 294370 327367
rect -2408 327238 294370 327249
rect -1938 327237 -1638 327238
rect 2702 327237 3002 327238
rect 20702 327237 21002 327238
rect 38702 327237 39002 327238
rect 56702 327237 57002 327238
rect 74702 327237 75002 327238
rect 92702 327237 93002 327238
rect 110702 327237 111002 327238
rect 128702 327237 129002 327238
rect 146702 327237 147002 327238
rect 164702 327237 165002 327238
rect 182702 327237 183002 327238
rect 200702 327237 201002 327238
rect 218702 327237 219002 327238
rect 236702 327237 237002 327238
rect 254702 327237 255002 327238
rect 272702 327237 273002 327238
rect 290702 327237 291002 327238
rect 293600 327237 293900 327238
rect -998 325738 -698 325739
rect 902 325738 1202 325739
rect 18902 325738 19202 325739
rect 36902 325738 37202 325739
rect 54902 325738 55202 325739
rect 72902 325738 73202 325739
rect 90902 325738 91202 325739
rect 108902 325738 109202 325739
rect 126902 325738 127202 325739
rect 144902 325738 145202 325739
rect 162902 325738 163202 325739
rect 180902 325738 181202 325739
rect 198902 325738 199202 325739
rect 216902 325738 217202 325739
rect 234902 325738 235202 325739
rect 252902 325738 253202 325739
rect 270902 325738 271202 325739
rect 288902 325738 289202 325739
rect 292660 325738 292960 325739
rect -1468 325727 293430 325738
rect -1468 325609 -907 325727
rect -789 325609 993 325727
rect 1111 325609 18993 325727
rect 19111 325609 36993 325727
rect 37111 325609 54993 325727
rect 55111 325609 72993 325727
rect 73111 325609 90993 325727
rect 91111 325609 108993 325727
rect 109111 325609 126993 325727
rect 127111 325609 144993 325727
rect 145111 325609 162993 325727
rect 163111 325609 180993 325727
rect 181111 325609 198993 325727
rect 199111 325609 216993 325727
rect 217111 325609 234993 325727
rect 235111 325609 252993 325727
rect 253111 325609 270993 325727
rect 271111 325609 288993 325727
rect 289111 325609 292751 325727
rect 292869 325609 293430 325727
rect -1468 325567 293430 325609
rect -1468 325449 -907 325567
rect -789 325449 993 325567
rect 1111 325449 18993 325567
rect 19111 325449 36993 325567
rect 37111 325449 54993 325567
rect 55111 325449 72993 325567
rect 73111 325449 90993 325567
rect 91111 325449 108993 325567
rect 109111 325449 126993 325567
rect 127111 325449 144993 325567
rect 145111 325449 162993 325567
rect 163111 325449 180993 325567
rect 181111 325449 198993 325567
rect 199111 325449 216993 325567
rect 217111 325449 234993 325567
rect 235111 325449 252993 325567
rect 253111 325449 270993 325567
rect 271111 325449 288993 325567
rect 289111 325449 292751 325567
rect 292869 325449 293430 325567
rect -1468 325438 293430 325449
rect -998 325437 -698 325438
rect 902 325437 1202 325438
rect 18902 325437 19202 325438
rect 36902 325437 37202 325438
rect 54902 325437 55202 325438
rect 72902 325437 73202 325438
rect 90902 325437 91202 325438
rect 108902 325437 109202 325438
rect 126902 325437 127202 325438
rect 144902 325437 145202 325438
rect 162902 325437 163202 325438
rect 180902 325437 181202 325438
rect 198902 325437 199202 325438
rect 216902 325437 217202 325438
rect 234902 325437 235202 325438
rect 252902 325437 253202 325438
rect 270902 325437 271202 325438
rect 288902 325437 289202 325438
rect 292660 325437 292960 325438
rect -4288 322138 -3988 322139
rect 15302 322138 15602 322139
rect 33302 322138 33602 322139
rect 51302 322138 51602 322139
rect 69302 322138 69602 322139
rect 87302 322138 87602 322139
rect 105302 322138 105602 322139
rect 123302 322138 123602 322139
rect 141302 322138 141602 322139
rect 159302 322138 159602 322139
rect 177302 322138 177602 322139
rect 195302 322138 195602 322139
rect 213302 322138 213602 322139
rect 231302 322138 231602 322139
rect 249302 322138 249602 322139
rect 267302 322138 267602 322139
rect 285302 322138 285602 322139
rect 295950 322138 296250 322139
rect -4288 322127 296250 322138
rect -4288 322009 -4197 322127
rect -4079 322009 15393 322127
rect 15511 322009 33393 322127
rect 33511 322009 51393 322127
rect 51511 322009 69393 322127
rect 69511 322009 87393 322127
rect 87511 322009 105393 322127
rect 105511 322009 123393 322127
rect 123511 322009 141393 322127
rect 141511 322009 159393 322127
rect 159511 322009 177393 322127
rect 177511 322009 195393 322127
rect 195511 322009 213393 322127
rect 213511 322009 231393 322127
rect 231511 322009 249393 322127
rect 249511 322009 267393 322127
rect 267511 322009 285393 322127
rect 285511 322009 296041 322127
rect 296159 322009 296250 322127
rect -4288 321967 296250 322009
rect -4288 321849 -4197 321967
rect -4079 321849 15393 321967
rect 15511 321849 33393 321967
rect 33511 321849 51393 321967
rect 51511 321849 69393 321967
rect 69511 321849 87393 321967
rect 87511 321849 105393 321967
rect 105511 321849 123393 321967
rect 123511 321849 141393 321967
rect 141511 321849 159393 321967
rect 159511 321849 177393 321967
rect 177511 321849 195393 321967
rect 195511 321849 213393 321967
rect 213511 321849 231393 321967
rect 231511 321849 249393 321967
rect 249511 321849 267393 321967
rect 267511 321849 285393 321967
rect 285511 321849 296041 321967
rect 296159 321849 296250 321967
rect -4288 321838 296250 321849
rect -4288 321837 -3988 321838
rect 15302 321837 15602 321838
rect 33302 321837 33602 321838
rect 51302 321837 51602 321838
rect 69302 321837 69602 321838
rect 87302 321837 87602 321838
rect 105302 321837 105602 321838
rect 123302 321837 123602 321838
rect 141302 321837 141602 321838
rect 159302 321837 159602 321838
rect 177302 321837 177602 321838
rect 195302 321837 195602 321838
rect 213302 321837 213602 321838
rect 231302 321837 231602 321838
rect 249302 321837 249602 321838
rect 267302 321837 267602 321838
rect 285302 321837 285602 321838
rect 295950 321837 296250 321838
rect -3348 320338 -3048 320339
rect 13502 320338 13802 320339
rect 31502 320338 31802 320339
rect 49502 320338 49802 320339
rect 67502 320338 67802 320339
rect 85502 320338 85802 320339
rect 103502 320338 103802 320339
rect 121502 320338 121802 320339
rect 139502 320338 139802 320339
rect 157502 320338 157802 320339
rect 175502 320338 175802 320339
rect 193502 320338 193802 320339
rect 211502 320338 211802 320339
rect 229502 320338 229802 320339
rect 247502 320338 247802 320339
rect 265502 320338 265802 320339
rect 283502 320338 283802 320339
rect 295010 320338 295310 320339
rect -3348 320327 295310 320338
rect -3348 320209 -3257 320327
rect -3139 320209 13593 320327
rect 13711 320209 31593 320327
rect 31711 320209 49593 320327
rect 49711 320209 67593 320327
rect 67711 320209 85593 320327
rect 85711 320209 103593 320327
rect 103711 320209 121593 320327
rect 121711 320209 139593 320327
rect 139711 320209 157593 320327
rect 157711 320209 175593 320327
rect 175711 320209 193593 320327
rect 193711 320209 211593 320327
rect 211711 320209 229593 320327
rect 229711 320209 247593 320327
rect 247711 320209 265593 320327
rect 265711 320209 283593 320327
rect 283711 320209 295101 320327
rect 295219 320209 295310 320327
rect -3348 320167 295310 320209
rect -3348 320049 -3257 320167
rect -3139 320049 13593 320167
rect 13711 320049 31593 320167
rect 31711 320049 49593 320167
rect 49711 320049 67593 320167
rect 67711 320049 85593 320167
rect 85711 320049 103593 320167
rect 103711 320049 121593 320167
rect 121711 320049 139593 320167
rect 139711 320049 157593 320167
rect 157711 320049 175593 320167
rect 175711 320049 193593 320167
rect 193711 320049 211593 320167
rect 211711 320049 229593 320167
rect 229711 320049 247593 320167
rect 247711 320049 265593 320167
rect 265711 320049 283593 320167
rect 283711 320049 295101 320167
rect 295219 320049 295310 320167
rect -3348 320038 295310 320049
rect -3348 320037 -3048 320038
rect 13502 320037 13802 320038
rect 31502 320037 31802 320038
rect 49502 320037 49802 320038
rect 67502 320037 67802 320038
rect 85502 320037 85802 320038
rect 103502 320037 103802 320038
rect 121502 320037 121802 320038
rect 139502 320037 139802 320038
rect 157502 320037 157802 320038
rect 175502 320037 175802 320038
rect 193502 320037 193802 320038
rect 211502 320037 211802 320038
rect 229502 320037 229802 320038
rect 247502 320037 247802 320038
rect 265502 320037 265802 320038
rect 283502 320037 283802 320038
rect 295010 320037 295310 320038
rect -2408 318538 -2108 318539
rect 11702 318538 12002 318539
rect 29702 318538 30002 318539
rect 47702 318538 48002 318539
rect 65702 318538 66002 318539
rect 83702 318538 84002 318539
rect 101702 318538 102002 318539
rect 119702 318538 120002 318539
rect 137702 318538 138002 318539
rect 155702 318538 156002 318539
rect 173702 318538 174002 318539
rect 191702 318538 192002 318539
rect 209702 318538 210002 318539
rect 227702 318538 228002 318539
rect 245702 318538 246002 318539
rect 263702 318538 264002 318539
rect 281702 318538 282002 318539
rect 294070 318538 294370 318539
rect -2408 318527 294370 318538
rect -2408 318409 -2317 318527
rect -2199 318409 11793 318527
rect 11911 318409 29793 318527
rect 29911 318409 47793 318527
rect 47911 318409 65793 318527
rect 65911 318409 83793 318527
rect 83911 318409 101793 318527
rect 101911 318409 119793 318527
rect 119911 318409 137793 318527
rect 137911 318409 155793 318527
rect 155911 318409 173793 318527
rect 173911 318409 191793 318527
rect 191911 318409 209793 318527
rect 209911 318409 227793 318527
rect 227911 318409 245793 318527
rect 245911 318409 263793 318527
rect 263911 318409 281793 318527
rect 281911 318409 294161 318527
rect 294279 318409 294370 318527
rect -2408 318367 294370 318409
rect -2408 318249 -2317 318367
rect -2199 318249 11793 318367
rect 11911 318249 29793 318367
rect 29911 318249 47793 318367
rect 47911 318249 65793 318367
rect 65911 318249 83793 318367
rect 83911 318249 101793 318367
rect 101911 318249 119793 318367
rect 119911 318249 137793 318367
rect 137911 318249 155793 318367
rect 155911 318249 173793 318367
rect 173911 318249 191793 318367
rect 191911 318249 209793 318367
rect 209911 318249 227793 318367
rect 227911 318249 245793 318367
rect 245911 318249 263793 318367
rect 263911 318249 281793 318367
rect 281911 318249 294161 318367
rect 294279 318249 294370 318367
rect -2408 318238 294370 318249
rect -2408 318237 -2108 318238
rect 11702 318237 12002 318238
rect 29702 318237 30002 318238
rect 47702 318237 48002 318238
rect 65702 318237 66002 318238
rect 83702 318237 84002 318238
rect 101702 318237 102002 318238
rect 119702 318237 120002 318238
rect 137702 318237 138002 318238
rect 155702 318237 156002 318238
rect 173702 318237 174002 318238
rect 191702 318237 192002 318238
rect 209702 318237 210002 318238
rect 227702 318237 228002 318238
rect 245702 318237 246002 318238
rect 263702 318237 264002 318238
rect 281702 318237 282002 318238
rect 294070 318237 294370 318238
rect -1468 316738 -1168 316739
rect 9902 316738 10202 316739
rect 27902 316738 28202 316739
rect 45902 316738 46202 316739
rect 63902 316738 64202 316739
rect 81902 316738 82202 316739
rect 99902 316738 100202 316739
rect 117902 316738 118202 316739
rect 135902 316738 136202 316739
rect 153902 316738 154202 316739
rect 171902 316738 172202 316739
rect 189902 316738 190202 316739
rect 207902 316738 208202 316739
rect 225902 316738 226202 316739
rect 243902 316738 244202 316739
rect 261902 316738 262202 316739
rect 279902 316738 280202 316739
rect 293130 316738 293430 316739
rect -1468 316727 293430 316738
rect -1468 316609 -1377 316727
rect -1259 316609 9993 316727
rect 10111 316609 27993 316727
rect 28111 316609 45993 316727
rect 46111 316609 63993 316727
rect 64111 316609 81993 316727
rect 82111 316609 99993 316727
rect 100111 316609 117993 316727
rect 118111 316609 135993 316727
rect 136111 316609 153993 316727
rect 154111 316609 171993 316727
rect 172111 316609 189993 316727
rect 190111 316609 207993 316727
rect 208111 316609 225993 316727
rect 226111 316609 243993 316727
rect 244111 316609 261993 316727
rect 262111 316609 279993 316727
rect 280111 316609 293221 316727
rect 293339 316609 293430 316727
rect -1468 316567 293430 316609
rect -1468 316449 -1377 316567
rect -1259 316449 9993 316567
rect 10111 316449 27993 316567
rect 28111 316449 45993 316567
rect 46111 316449 63993 316567
rect 64111 316449 81993 316567
rect 82111 316449 99993 316567
rect 100111 316449 117993 316567
rect 118111 316449 135993 316567
rect 136111 316449 153993 316567
rect 154111 316449 171993 316567
rect 172111 316449 189993 316567
rect 190111 316449 207993 316567
rect 208111 316449 225993 316567
rect 226111 316449 243993 316567
rect 244111 316449 261993 316567
rect 262111 316449 279993 316567
rect 280111 316449 293221 316567
rect 293339 316449 293430 316567
rect -1468 316438 293430 316449
rect -1468 316437 -1168 316438
rect 9902 316437 10202 316438
rect 27902 316437 28202 316438
rect 45902 316437 46202 316438
rect 63902 316437 64202 316438
rect 81902 316437 82202 316438
rect 99902 316437 100202 316438
rect 117902 316437 118202 316438
rect 135902 316437 136202 316438
rect 153902 316437 154202 316438
rect 171902 316437 172202 316438
rect 189902 316437 190202 316438
rect 207902 316437 208202 316438
rect 225902 316437 226202 316438
rect 243902 316437 244202 316438
rect 261902 316437 262202 316438
rect 279902 316437 280202 316438
rect 293130 316437 293430 316438
rect -3818 313138 -3518 313139
rect 6302 313138 6602 313139
rect 24302 313138 24602 313139
rect 42302 313138 42602 313139
rect 60302 313138 60602 313139
rect 78302 313138 78602 313139
rect 96302 313138 96602 313139
rect 114302 313138 114602 313139
rect 132302 313138 132602 313139
rect 150302 313138 150602 313139
rect 168302 313138 168602 313139
rect 186302 313138 186602 313139
rect 204302 313138 204602 313139
rect 222302 313138 222602 313139
rect 240302 313138 240602 313139
rect 258302 313138 258602 313139
rect 276302 313138 276602 313139
rect 295480 313138 295780 313139
rect -4288 313127 296250 313138
rect -4288 313009 -3727 313127
rect -3609 313009 6393 313127
rect 6511 313009 24393 313127
rect 24511 313009 42393 313127
rect 42511 313009 60393 313127
rect 60511 313009 78393 313127
rect 78511 313009 96393 313127
rect 96511 313009 114393 313127
rect 114511 313009 132393 313127
rect 132511 313009 150393 313127
rect 150511 313009 168393 313127
rect 168511 313009 186393 313127
rect 186511 313009 204393 313127
rect 204511 313009 222393 313127
rect 222511 313009 240393 313127
rect 240511 313009 258393 313127
rect 258511 313009 276393 313127
rect 276511 313009 295571 313127
rect 295689 313009 296250 313127
rect -4288 312967 296250 313009
rect -4288 312849 -3727 312967
rect -3609 312849 6393 312967
rect 6511 312849 24393 312967
rect 24511 312849 42393 312967
rect 42511 312849 60393 312967
rect 60511 312849 78393 312967
rect 78511 312849 96393 312967
rect 96511 312849 114393 312967
rect 114511 312849 132393 312967
rect 132511 312849 150393 312967
rect 150511 312849 168393 312967
rect 168511 312849 186393 312967
rect 186511 312849 204393 312967
rect 204511 312849 222393 312967
rect 222511 312849 240393 312967
rect 240511 312849 258393 312967
rect 258511 312849 276393 312967
rect 276511 312849 295571 312967
rect 295689 312849 296250 312967
rect -4288 312838 296250 312849
rect -3818 312837 -3518 312838
rect 6302 312837 6602 312838
rect 24302 312837 24602 312838
rect 42302 312837 42602 312838
rect 60302 312837 60602 312838
rect 78302 312837 78602 312838
rect 96302 312837 96602 312838
rect 114302 312837 114602 312838
rect 132302 312837 132602 312838
rect 150302 312837 150602 312838
rect 168302 312837 168602 312838
rect 186302 312837 186602 312838
rect 204302 312837 204602 312838
rect 222302 312837 222602 312838
rect 240302 312837 240602 312838
rect 258302 312837 258602 312838
rect 276302 312837 276602 312838
rect 295480 312837 295780 312838
rect -2878 311338 -2578 311339
rect 4502 311338 4802 311339
rect 22502 311338 22802 311339
rect 40502 311338 40802 311339
rect 58502 311338 58802 311339
rect 76502 311338 76802 311339
rect 94502 311338 94802 311339
rect 112502 311338 112802 311339
rect 130502 311338 130802 311339
rect 148502 311338 148802 311339
rect 166502 311338 166802 311339
rect 184502 311338 184802 311339
rect 202502 311338 202802 311339
rect 220502 311338 220802 311339
rect 238502 311338 238802 311339
rect 256502 311338 256802 311339
rect 274502 311338 274802 311339
rect 294540 311338 294840 311339
rect -3348 311327 295310 311338
rect -3348 311209 -2787 311327
rect -2669 311209 4593 311327
rect 4711 311209 22593 311327
rect 22711 311209 40593 311327
rect 40711 311209 58593 311327
rect 58711 311209 76593 311327
rect 76711 311209 94593 311327
rect 94711 311209 112593 311327
rect 112711 311209 130593 311327
rect 130711 311209 148593 311327
rect 148711 311209 166593 311327
rect 166711 311209 184593 311327
rect 184711 311209 202593 311327
rect 202711 311209 220593 311327
rect 220711 311209 238593 311327
rect 238711 311209 256593 311327
rect 256711 311209 274593 311327
rect 274711 311209 294631 311327
rect 294749 311209 295310 311327
rect -3348 311167 295310 311209
rect -3348 311049 -2787 311167
rect -2669 311049 4593 311167
rect 4711 311049 22593 311167
rect 22711 311049 40593 311167
rect 40711 311049 58593 311167
rect 58711 311049 76593 311167
rect 76711 311049 94593 311167
rect 94711 311049 112593 311167
rect 112711 311049 130593 311167
rect 130711 311049 148593 311167
rect 148711 311049 166593 311167
rect 166711 311049 184593 311167
rect 184711 311049 202593 311167
rect 202711 311049 220593 311167
rect 220711 311049 238593 311167
rect 238711 311049 256593 311167
rect 256711 311049 274593 311167
rect 274711 311049 294631 311167
rect 294749 311049 295310 311167
rect -3348 311038 295310 311049
rect -2878 311037 -2578 311038
rect 4502 311037 4802 311038
rect 22502 311037 22802 311038
rect 40502 311037 40802 311038
rect 58502 311037 58802 311038
rect 76502 311037 76802 311038
rect 94502 311037 94802 311038
rect 112502 311037 112802 311038
rect 130502 311037 130802 311038
rect 148502 311037 148802 311038
rect 166502 311037 166802 311038
rect 184502 311037 184802 311038
rect 202502 311037 202802 311038
rect 220502 311037 220802 311038
rect 238502 311037 238802 311038
rect 256502 311037 256802 311038
rect 274502 311037 274802 311038
rect 294540 311037 294840 311038
rect -1938 309538 -1638 309539
rect 2702 309538 3002 309539
rect 20702 309538 21002 309539
rect 38702 309538 39002 309539
rect 56702 309538 57002 309539
rect 74702 309538 75002 309539
rect 92702 309538 93002 309539
rect 110702 309538 111002 309539
rect 128702 309538 129002 309539
rect 146702 309538 147002 309539
rect 164702 309538 165002 309539
rect 182702 309538 183002 309539
rect 200702 309538 201002 309539
rect 218702 309538 219002 309539
rect 236702 309538 237002 309539
rect 254702 309538 255002 309539
rect 272702 309538 273002 309539
rect 290702 309538 291002 309539
rect 293600 309538 293900 309539
rect -2408 309527 294370 309538
rect -2408 309409 -1847 309527
rect -1729 309409 2793 309527
rect 2911 309409 20793 309527
rect 20911 309409 38793 309527
rect 38911 309409 56793 309527
rect 56911 309409 74793 309527
rect 74911 309409 92793 309527
rect 92911 309409 110793 309527
rect 110911 309409 128793 309527
rect 128911 309409 146793 309527
rect 146911 309409 164793 309527
rect 164911 309409 182793 309527
rect 182911 309409 200793 309527
rect 200911 309409 218793 309527
rect 218911 309409 236793 309527
rect 236911 309409 254793 309527
rect 254911 309409 272793 309527
rect 272911 309409 290793 309527
rect 290911 309409 293691 309527
rect 293809 309409 294370 309527
rect -2408 309367 294370 309409
rect -2408 309249 -1847 309367
rect -1729 309249 2793 309367
rect 2911 309249 20793 309367
rect 20911 309249 38793 309367
rect 38911 309249 56793 309367
rect 56911 309249 74793 309367
rect 74911 309249 92793 309367
rect 92911 309249 110793 309367
rect 110911 309249 128793 309367
rect 128911 309249 146793 309367
rect 146911 309249 164793 309367
rect 164911 309249 182793 309367
rect 182911 309249 200793 309367
rect 200911 309249 218793 309367
rect 218911 309249 236793 309367
rect 236911 309249 254793 309367
rect 254911 309249 272793 309367
rect 272911 309249 290793 309367
rect 290911 309249 293691 309367
rect 293809 309249 294370 309367
rect -2408 309238 294370 309249
rect -1938 309237 -1638 309238
rect 2702 309237 3002 309238
rect 20702 309237 21002 309238
rect 38702 309237 39002 309238
rect 56702 309237 57002 309238
rect 74702 309237 75002 309238
rect 92702 309237 93002 309238
rect 110702 309237 111002 309238
rect 128702 309237 129002 309238
rect 146702 309237 147002 309238
rect 164702 309237 165002 309238
rect 182702 309237 183002 309238
rect 200702 309237 201002 309238
rect 218702 309237 219002 309238
rect 236702 309237 237002 309238
rect 254702 309237 255002 309238
rect 272702 309237 273002 309238
rect 290702 309237 291002 309238
rect 293600 309237 293900 309238
rect -998 307738 -698 307739
rect 902 307738 1202 307739
rect 18902 307738 19202 307739
rect 36902 307738 37202 307739
rect 54902 307738 55202 307739
rect 72902 307738 73202 307739
rect 90902 307738 91202 307739
rect 108902 307738 109202 307739
rect 126902 307738 127202 307739
rect 144902 307738 145202 307739
rect 162902 307738 163202 307739
rect 180902 307738 181202 307739
rect 198902 307738 199202 307739
rect 216902 307738 217202 307739
rect 234902 307738 235202 307739
rect 252902 307738 253202 307739
rect 270902 307738 271202 307739
rect 288902 307738 289202 307739
rect 292660 307738 292960 307739
rect -1468 307727 293430 307738
rect -1468 307609 -907 307727
rect -789 307609 993 307727
rect 1111 307609 18993 307727
rect 19111 307609 36993 307727
rect 37111 307609 54993 307727
rect 55111 307609 72993 307727
rect 73111 307609 90993 307727
rect 91111 307609 108993 307727
rect 109111 307609 126993 307727
rect 127111 307609 144993 307727
rect 145111 307609 162993 307727
rect 163111 307609 180993 307727
rect 181111 307609 198993 307727
rect 199111 307609 216993 307727
rect 217111 307609 234993 307727
rect 235111 307609 252993 307727
rect 253111 307609 270993 307727
rect 271111 307609 288993 307727
rect 289111 307609 292751 307727
rect 292869 307609 293430 307727
rect -1468 307567 293430 307609
rect -1468 307449 -907 307567
rect -789 307449 993 307567
rect 1111 307449 18993 307567
rect 19111 307449 36993 307567
rect 37111 307449 54993 307567
rect 55111 307449 72993 307567
rect 73111 307449 90993 307567
rect 91111 307449 108993 307567
rect 109111 307449 126993 307567
rect 127111 307449 144993 307567
rect 145111 307449 162993 307567
rect 163111 307449 180993 307567
rect 181111 307449 198993 307567
rect 199111 307449 216993 307567
rect 217111 307449 234993 307567
rect 235111 307449 252993 307567
rect 253111 307449 270993 307567
rect 271111 307449 288993 307567
rect 289111 307449 292751 307567
rect 292869 307449 293430 307567
rect -1468 307438 293430 307449
rect -998 307437 -698 307438
rect 902 307437 1202 307438
rect 18902 307437 19202 307438
rect 36902 307437 37202 307438
rect 54902 307437 55202 307438
rect 72902 307437 73202 307438
rect 90902 307437 91202 307438
rect 108902 307437 109202 307438
rect 126902 307437 127202 307438
rect 144902 307437 145202 307438
rect 162902 307437 163202 307438
rect 180902 307437 181202 307438
rect 198902 307437 199202 307438
rect 216902 307437 217202 307438
rect 234902 307437 235202 307438
rect 252902 307437 253202 307438
rect 270902 307437 271202 307438
rect 288902 307437 289202 307438
rect 292660 307437 292960 307438
rect -4288 304138 -3988 304139
rect 15302 304138 15602 304139
rect 33302 304138 33602 304139
rect 51302 304138 51602 304139
rect 69302 304138 69602 304139
rect 87302 304138 87602 304139
rect 105302 304138 105602 304139
rect 123302 304138 123602 304139
rect 141302 304138 141602 304139
rect 159302 304138 159602 304139
rect 177302 304138 177602 304139
rect 195302 304138 195602 304139
rect 213302 304138 213602 304139
rect 231302 304138 231602 304139
rect 249302 304138 249602 304139
rect 267302 304138 267602 304139
rect 285302 304138 285602 304139
rect 295950 304138 296250 304139
rect -4288 304127 296250 304138
rect -4288 304009 -4197 304127
rect -4079 304009 15393 304127
rect 15511 304009 33393 304127
rect 33511 304009 51393 304127
rect 51511 304009 69393 304127
rect 69511 304009 87393 304127
rect 87511 304009 105393 304127
rect 105511 304009 123393 304127
rect 123511 304009 141393 304127
rect 141511 304009 159393 304127
rect 159511 304009 177393 304127
rect 177511 304009 195393 304127
rect 195511 304009 213393 304127
rect 213511 304009 231393 304127
rect 231511 304009 249393 304127
rect 249511 304009 267393 304127
rect 267511 304009 285393 304127
rect 285511 304009 296041 304127
rect 296159 304009 296250 304127
rect -4288 303967 296250 304009
rect -4288 303849 -4197 303967
rect -4079 303849 15393 303967
rect 15511 303849 33393 303967
rect 33511 303849 51393 303967
rect 51511 303849 69393 303967
rect 69511 303849 87393 303967
rect 87511 303849 105393 303967
rect 105511 303849 123393 303967
rect 123511 303849 141393 303967
rect 141511 303849 159393 303967
rect 159511 303849 177393 303967
rect 177511 303849 195393 303967
rect 195511 303849 213393 303967
rect 213511 303849 231393 303967
rect 231511 303849 249393 303967
rect 249511 303849 267393 303967
rect 267511 303849 285393 303967
rect 285511 303849 296041 303967
rect 296159 303849 296250 303967
rect -4288 303838 296250 303849
rect -4288 303837 -3988 303838
rect 15302 303837 15602 303838
rect 33302 303837 33602 303838
rect 51302 303837 51602 303838
rect 69302 303837 69602 303838
rect 87302 303837 87602 303838
rect 105302 303837 105602 303838
rect 123302 303837 123602 303838
rect 141302 303837 141602 303838
rect 159302 303837 159602 303838
rect 177302 303837 177602 303838
rect 195302 303837 195602 303838
rect 213302 303837 213602 303838
rect 231302 303837 231602 303838
rect 249302 303837 249602 303838
rect 267302 303837 267602 303838
rect 285302 303837 285602 303838
rect 295950 303837 296250 303838
rect -3348 302338 -3048 302339
rect 13502 302338 13802 302339
rect 31502 302338 31802 302339
rect 49502 302338 49802 302339
rect 67502 302338 67802 302339
rect 85502 302338 85802 302339
rect 103502 302338 103802 302339
rect 121502 302338 121802 302339
rect 139502 302338 139802 302339
rect 157502 302338 157802 302339
rect 175502 302338 175802 302339
rect 193502 302338 193802 302339
rect 211502 302338 211802 302339
rect 229502 302338 229802 302339
rect 247502 302338 247802 302339
rect 265502 302338 265802 302339
rect 283502 302338 283802 302339
rect 295010 302338 295310 302339
rect -3348 302327 295310 302338
rect -3348 302209 -3257 302327
rect -3139 302209 13593 302327
rect 13711 302209 31593 302327
rect 31711 302209 49593 302327
rect 49711 302209 67593 302327
rect 67711 302209 85593 302327
rect 85711 302209 103593 302327
rect 103711 302209 121593 302327
rect 121711 302209 139593 302327
rect 139711 302209 157593 302327
rect 157711 302209 175593 302327
rect 175711 302209 193593 302327
rect 193711 302209 211593 302327
rect 211711 302209 229593 302327
rect 229711 302209 247593 302327
rect 247711 302209 265593 302327
rect 265711 302209 283593 302327
rect 283711 302209 295101 302327
rect 295219 302209 295310 302327
rect -3348 302167 295310 302209
rect -3348 302049 -3257 302167
rect -3139 302049 13593 302167
rect 13711 302049 31593 302167
rect 31711 302049 49593 302167
rect 49711 302049 67593 302167
rect 67711 302049 85593 302167
rect 85711 302049 103593 302167
rect 103711 302049 121593 302167
rect 121711 302049 139593 302167
rect 139711 302049 157593 302167
rect 157711 302049 175593 302167
rect 175711 302049 193593 302167
rect 193711 302049 211593 302167
rect 211711 302049 229593 302167
rect 229711 302049 247593 302167
rect 247711 302049 265593 302167
rect 265711 302049 283593 302167
rect 283711 302049 295101 302167
rect 295219 302049 295310 302167
rect -3348 302038 295310 302049
rect -3348 302037 -3048 302038
rect 13502 302037 13802 302038
rect 31502 302037 31802 302038
rect 49502 302037 49802 302038
rect 67502 302037 67802 302038
rect 85502 302037 85802 302038
rect 103502 302037 103802 302038
rect 121502 302037 121802 302038
rect 139502 302037 139802 302038
rect 157502 302037 157802 302038
rect 175502 302037 175802 302038
rect 193502 302037 193802 302038
rect 211502 302037 211802 302038
rect 229502 302037 229802 302038
rect 247502 302037 247802 302038
rect 265502 302037 265802 302038
rect 283502 302037 283802 302038
rect 295010 302037 295310 302038
rect -2408 300538 -2108 300539
rect 11702 300538 12002 300539
rect 29702 300538 30002 300539
rect 47702 300538 48002 300539
rect 65702 300538 66002 300539
rect 83702 300538 84002 300539
rect 101702 300538 102002 300539
rect 119702 300538 120002 300539
rect 137702 300538 138002 300539
rect 155702 300538 156002 300539
rect 173702 300538 174002 300539
rect 191702 300538 192002 300539
rect 209702 300538 210002 300539
rect 227702 300538 228002 300539
rect 245702 300538 246002 300539
rect 263702 300538 264002 300539
rect 281702 300538 282002 300539
rect 294070 300538 294370 300539
rect -2408 300527 294370 300538
rect -2408 300409 -2317 300527
rect -2199 300409 11793 300527
rect 11911 300409 29793 300527
rect 29911 300409 47793 300527
rect 47911 300409 65793 300527
rect 65911 300409 83793 300527
rect 83911 300409 101793 300527
rect 101911 300409 119793 300527
rect 119911 300409 137793 300527
rect 137911 300409 155793 300527
rect 155911 300409 173793 300527
rect 173911 300409 191793 300527
rect 191911 300409 209793 300527
rect 209911 300409 227793 300527
rect 227911 300409 245793 300527
rect 245911 300409 263793 300527
rect 263911 300409 281793 300527
rect 281911 300409 294161 300527
rect 294279 300409 294370 300527
rect -2408 300367 294370 300409
rect -2408 300249 -2317 300367
rect -2199 300249 11793 300367
rect 11911 300249 29793 300367
rect 29911 300249 47793 300367
rect 47911 300249 65793 300367
rect 65911 300249 83793 300367
rect 83911 300249 101793 300367
rect 101911 300249 119793 300367
rect 119911 300249 137793 300367
rect 137911 300249 155793 300367
rect 155911 300249 173793 300367
rect 173911 300249 191793 300367
rect 191911 300249 209793 300367
rect 209911 300249 227793 300367
rect 227911 300249 245793 300367
rect 245911 300249 263793 300367
rect 263911 300249 281793 300367
rect 281911 300249 294161 300367
rect 294279 300249 294370 300367
rect -2408 300238 294370 300249
rect -2408 300237 -2108 300238
rect 11702 300237 12002 300238
rect 29702 300237 30002 300238
rect 47702 300237 48002 300238
rect 65702 300237 66002 300238
rect 83702 300237 84002 300238
rect 101702 300237 102002 300238
rect 119702 300237 120002 300238
rect 137702 300237 138002 300238
rect 155702 300237 156002 300238
rect 173702 300237 174002 300238
rect 191702 300237 192002 300238
rect 209702 300237 210002 300238
rect 227702 300237 228002 300238
rect 245702 300237 246002 300238
rect 263702 300237 264002 300238
rect 281702 300237 282002 300238
rect 294070 300237 294370 300238
rect -1468 298738 -1168 298739
rect 9902 298738 10202 298739
rect 27902 298738 28202 298739
rect 45902 298738 46202 298739
rect 63902 298738 64202 298739
rect 81902 298738 82202 298739
rect 99902 298738 100202 298739
rect 117902 298738 118202 298739
rect 135902 298738 136202 298739
rect 153902 298738 154202 298739
rect 171902 298738 172202 298739
rect 189902 298738 190202 298739
rect 207902 298738 208202 298739
rect 225902 298738 226202 298739
rect 243902 298738 244202 298739
rect 261902 298738 262202 298739
rect 279902 298738 280202 298739
rect 293130 298738 293430 298739
rect -1468 298727 293430 298738
rect -1468 298609 -1377 298727
rect -1259 298609 9993 298727
rect 10111 298609 27993 298727
rect 28111 298609 45993 298727
rect 46111 298609 63993 298727
rect 64111 298609 81993 298727
rect 82111 298609 99993 298727
rect 100111 298609 117993 298727
rect 118111 298609 135993 298727
rect 136111 298609 153993 298727
rect 154111 298609 171993 298727
rect 172111 298609 189993 298727
rect 190111 298609 207993 298727
rect 208111 298609 225993 298727
rect 226111 298609 243993 298727
rect 244111 298609 261993 298727
rect 262111 298609 279993 298727
rect 280111 298609 293221 298727
rect 293339 298609 293430 298727
rect -1468 298567 293430 298609
rect -1468 298449 -1377 298567
rect -1259 298449 9993 298567
rect 10111 298449 27993 298567
rect 28111 298449 45993 298567
rect 46111 298449 63993 298567
rect 64111 298449 81993 298567
rect 82111 298449 99993 298567
rect 100111 298449 117993 298567
rect 118111 298449 135993 298567
rect 136111 298449 153993 298567
rect 154111 298449 171993 298567
rect 172111 298449 189993 298567
rect 190111 298449 207993 298567
rect 208111 298449 225993 298567
rect 226111 298449 243993 298567
rect 244111 298449 261993 298567
rect 262111 298449 279993 298567
rect 280111 298449 293221 298567
rect 293339 298449 293430 298567
rect -1468 298438 293430 298449
rect -1468 298437 -1168 298438
rect 9902 298437 10202 298438
rect 27902 298437 28202 298438
rect 45902 298437 46202 298438
rect 63902 298437 64202 298438
rect 81902 298437 82202 298438
rect 99902 298437 100202 298438
rect 117902 298437 118202 298438
rect 135902 298437 136202 298438
rect 153902 298437 154202 298438
rect 171902 298437 172202 298438
rect 189902 298437 190202 298438
rect 207902 298437 208202 298438
rect 225902 298437 226202 298438
rect 243902 298437 244202 298438
rect 261902 298437 262202 298438
rect 279902 298437 280202 298438
rect 293130 298437 293430 298438
rect -3818 295138 -3518 295139
rect 6302 295138 6602 295139
rect 24302 295138 24602 295139
rect 42302 295138 42602 295139
rect 60302 295138 60602 295139
rect 78302 295138 78602 295139
rect 96302 295138 96602 295139
rect 114302 295138 114602 295139
rect 132302 295138 132602 295139
rect 150302 295138 150602 295139
rect 168302 295138 168602 295139
rect 186302 295138 186602 295139
rect 204302 295138 204602 295139
rect 222302 295138 222602 295139
rect 240302 295138 240602 295139
rect 258302 295138 258602 295139
rect 276302 295138 276602 295139
rect 295480 295138 295780 295139
rect -4288 295127 296250 295138
rect -4288 295009 -3727 295127
rect -3609 295009 6393 295127
rect 6511 295009 24393 295127
rect 24511 295009 42393 295127
rect 42511 295009 60393 295127
rect 60511 295009 78393 295127
rect 78511 295009 96393 295127
rect 96511 295009 114393 295127
rect 114511 295009 132393 295127
rect 132511 295009 150393 295127
rect 150511 295009 168393 295127
rect 168511 295009 186393 295127
rect 186511 295009 204393 295127
rect 204511 295009 222393 295127
rect 222511 295009 240393 295127
rect 240511 295009 258393 295127
rect 258511 295009 276393 295127
rect 276511 295009 295571 295127
rect 295689 295009 296250 295127
rect -4288 294967 296250 295009
rect -4288 294849 -3727 294967
rect -3609 294849 6393 294967
rect 6511 294849 24393 294967
rect 24511 294849 42393 294967
rect 42511 294849 60393 294967
rect 60511 294849 78393 294967
rect 78511 294849 96393 294967
rect 96511 294849 114393 294967
rect 114511 294849 132393 294967
rect 132511 294849 150393 294967
rect 150511 294849 168393 294967
rect 168511 294849 186393 294967
rect 186511 294849 204393 294967
rect 204511 294849 222393 294967
rect 222511 294849 240393 294967
rect 240511 294849 258393 294967
rect 258511 294849 276393 294967
rect 276511 294849 295571 294967
rect 295689 294849 296250 294967
rect -4288 294838 296250 294849
rect -3818 294837 -3518 294838
rect 6302 294837 6602 294838
rect 24302 294837 24602 294838
rect 42302 294837 42602 294838
rect 60302 294837 60602 294838
rect 78302 294837 78602 294838
rect 96302 294837 96602 294838
rect 114302 294837 114602 294838
rect 132302 294837 132602 294838
rect 150302 294837 150602 294838
rect 168302 294837 168602 294838
rect 186302 294837 186602 294838
rect 204302 294837 204602 294838
rect 222302 294837 222602 294838
rect 240302 294837 240602 294838
rect 258302 294837 258602 294838
rect 276302 294837 276602 294838
rect 295480 294837 295780 294838
rect -2878 293338 -2578 293339
rect 4502 293338 4802 293339
rect 22502 293338 22802 293339
rect 40502 293338 40802 293339
rect 58502 293338 58802 293339
rect 76502 293338 76802 293339
rect 94502 293338 94802 293339
rect 112502 293338 112802 293339
rect 130502 293338 130802 293339
rect 148502 293338 148802 293339
rect 166502 293338 166802 293339
rect 184502 293338 184802 293339
rect 202502 293338 202802 293339
rect 220502 293338 220802 293339
rect 238502 293338 238802 293339
rect 256502 293338 256802 293339
rect 274502 293338 274802 293339
rect 294540 293338 294840 293339
rect -3348 293327 295310 293338
rect -3348 293209 -2787 293327
rect -2669 293209 4593 293327
rect 4711 293209 22593 293327
rect 22711 293209 40593 293327
rect 40711 293209 58593 293327
rect 58711 293209 76593 293327
rect 76711 293209 94593 293327
rect 94711 293209 112593 293327
rect 112711 293209 130593 293327
rect 130711 293209 148593 293327
rect 148711 293209 166593 293327
rect 166711 293209 184593 293327
rect 184711 293209 202593 293327
rect 202711 293209 220593 293327
rect 220711 293209 238593 293327
rect 238711 293209 256593 293327
rect 256711 293209 274593 293327
rect 274711 293209 294631 293327
rect 294749 293209 295310 293327
rect -3348 293167 295310 293209
rect -3348 293049 -2787 293167
rect -2669 293049 4593 293167
rect 4711 293049 22593 293167
rect 22711 293049 40593 293167
rect 40711 293049 58593 293167
rect 58711 293049 76593 293167
rect 76711 293049 94593 293167
rect 94711 293049 112593 293167
rect 112711 293049 130593 293167
rect 130711 293049 148593 293167
rect 148711 293049 166593 293167
rect 166711 293049 184593 293167
rect 184711 293049 202593 293167
rect 202711 293049 220593 293167
rect 220711 293049 238593 293167
rect 238711 293049 256593 293167
rect 256711 293049 274593 293167
rect 274711 293049 294631 293167
rect 294749 293049 295310 293167
rect -3348 293038 295310 293049
rect -2878 293037 -2578 293038
rect 4502 293037 4802 293038
rect 22502 293037 22802 293038
rect 40502 293037 40802 293038
rect 58502 293037 58802 293038
rect 76502 293037 76802 293038
rect 94502 293037 94802 293038
rect 112502 293037 112802 293038
rect 130502 293037 130802 293038
rect 148502 293037 148802 293038
rect 166502 293037 166802 293038
rect 184502 293037 184802 293038
rect 202502 293037 202802 293038
rect 220502 293037 220802 293038
rect 238502 293037 238802 293038
rect 256502 293037 256802 293038
rect 274502 293037 274802 293038
rect 294540 293037 294840 293038
rect -1938 291538 -1638 291539
rect 2702 291538 3002 291539
rect 20702 291538 21002 291539
rect 38702 291538 39002 291539
rect 56702 291538 57002 291539
rect 74702 291538 75002 291539
rect 92702 291538 93002 291539
rect 110702 291538 111002 291539
rect 128702 291538 129002 291539
rect 146702 291538 147002 291539
rect 164702 291538 165002 291539
rect 182702 291538 183002 291539
rect 200702 291538 201002 291539
rect 218702 291538 219002 291539
rect 236702 291538 237002 291539
rect 254702 291538 255002 291539
rect 272702 291538 273002 291539
rect 290702 291538 291002 291539
rect 293600 291538 293900 291539
rect -2408 291527 294370 291538
rect -2408 291409 -1847 291527
rect -1729 291409 2793 291527
rect 2911 291409 20793 291527
rect 20911 291409 38793 291527
rect 38911 291409 56793 291527
rect 56911 291409 74793 291527
rect 74911 291409 92793 291527
rect 92911 291409 110793 291527
rect 110911 291409 128793 291527
rect 128911 291409 146793 291527
rect 146911 291409 164793 291527
rect 164911 291409 182793 291527
rect 182911 291409 200793 291527
rect 200911 291409 218793 291527
rect 218911 291409 236793 291527
rect 236911 291409 254793 291527
rect 254911 291409 272793 291527
rect 272911 291409 290793 291527
rect 290911 291409 293691 291527
rect 293809 291409 294370 291527
rect -2408 291367 294370 291409
rect -2408 291249 -1847 291367
rect -1729 291249 2793 291367
rect 2911 291249 20793 291367
rect 20911 291249 38793 291367
rect 38911 291249 56793 291367
rect 56911 291249 74793 291367
rect 74911 291249 92793 291367
rect 92911 291249 110793 291367
rect 110911 291249 128793 291367
rect 128911 291249 146793 291367
rect 146911 291249 164793 291367
rect 164911 291249 182793 291367
rect 182911 291249 200793 291367
rect 200911 291249 218793 291367
rect 218911 291249 236793 291367
rect 236911 291249 254793 291367
rect 254911 291249 272793 291367
rect 272911 291249 290793 291367
rect 290911 291249 293691 291367
rect 293809 291249 294370 291367
rect -2408 291238 294370 291249
rect -1938 291237 -1638 291238
rect 2702 291237 3002 291238
rect 20702 291237 21002 291238
rect 38702 291237 39002 291238
rect 56702 291237 57002 291238
rect 74702 291237 75002 291238
rect 92702 291237 93002 291238
rect 110702 291237 111002 291238
rect 128702 291237 129002 291238
rect 146702 291237 147002 291238
rect 164702 291237 165002 291238
rect 182702 291237 183002 291238
rect 200702 291237 201002 291238
rect 218702 291237 219002 291238
rect 236702 291237 237002 291238
rect 254702 291237 255002 291238
rect 272702 291237 273002 291238
rect 290702 291237 291002 291238
rect 293600 291237 293900 291238
rect -998 289738 -698 289739
rect 902 289738 1202 289739
rect 18902 289738 19202 289739
rect 36902 289738 37202 289739
rect 54902 289738 55202 289739
rect 72902 289738 73202 289739
rect 90902 289738 91202 289739
rect 108902 289738 109202 289739
rect 126902 289738 127202 289739
rect 144902 289738 145202 289739
rect 162902 289738 163202 289739
rect 180902 289738 181202 289739
rect 198902 289738 199202 289739
rect 216902 289738 217202 289739
rect 234902 289738 235202 289739
rect 252902 289738 253202 289739
rect 270902 289738 271202 289739
rect 288902 289738 289202 289739
rect 292660 289738 292960 289739
rect -1468 289727 293430 289738
rect -1468 289609 -907 289727
rect -789 289609 993 289727
rect 1111 289609 18993 289727
rect 19111 289609 36993 289727
rect 37111 289609 54993 289727
rect 55111 289609 72993 289727
rect 73111 289609 90993 289727
rect 91111 289609 108993 289727
rect 109111 289609 126993 289727
rect 127111 289609 144993 289727
rect 145111 289609 162993 289727
rect 163111 289609 180993 289727
rect 181111 289609 198993 289727
rect 199111 289609 216993 289727
rect 217111 289609 234993 289727
rect 235111 289609 252993 289727
rect 253111 289609 270993 289727
rect 271111 289609 288993 289727
rect 289111 289609 292751 289727
rect 292869 289609 293430 289727
rect -1468 289567 293430 289609
rect -1468 289449 -907 289567
rect -789 289449 993 289567
rect 1111 289449 18993 289567
rect 19111 289449 36993 289567
rect 37111 289449 54993 289567
rect 55111 289449 72993 289567
rect 73111 289449 90993 289567
rect 91111 289449 108993 289567
rect 109111 289449 126993 289567
rect 127111 289449 144993 289567
rect 145111 289449 162993 289567
rect 163111 289449 180993 289567
rect 181111 289449 198993 289567
rect 199111 289449 216993 289567
rect 217111 289449 234993 289567
rect 235111 289449 252993 289567
rect 253111 289449 270993 289567
rect 271111 289449 288993 289567
rect 289111 289449 292751 289567
rect 292869 289449 293430 289567
rect -1468 289438 293430 289449
rect -998 289437 -698 289438
rect 902 289437 1202 289438
rect 18902 289437 19202 289438
rect 36902 289437 37202 289438
rect 54902 289437 55202 289438
rect 72902 289437 73202 289438
rect 90902 289437 91202 289438
rect 108902 289437 109202 289438
rect 126902 289437 127202 289438
rect 144902 289437 145202 289438
rect 162902 289437 163202 289438
rect 180902 289437 181202 289438
rect 198902 289437 199202 289438
rect 216902 289437 217202 289438
rect 234902 289437 235202 289438
rect 252902 289437 253202 289438
rect 270902 289437 271202 289438
rect 288902 289437 289202 289438
rect 292660 289437 292960 289438
rect -4288 286138 -3988 286139
rect 15302 286138 15602 286139
rect 33302 286138 33602 286139
rect 51302 286138 51602 286139
rect 69302 286138 69602 286139
rect 87302 286138 87602 286139
rect 105302 286138 105602 286139
rect 123302 286138 123602 286139
rect 141302 286138 141602 286139
rect 159302 286138 159602 286139
rect 177302 286138 177602 286139
rect 195302 286138 195602 286139
rect 213302 286138 213602 286139
rect 231302 286138 231602 286139
rect 249302 286138 249602 286139
rect 267302 286138 267602 286139
rect 285302 286138 285602 286139
rect 295950 286138 296250 286139
rect -4288 286127 296250 286138
rect -4288 286009 -4197 286127
rect -4079 286009 15393 286127
rect 15511 286009 33393 286127
rect 33511 286009 51393 286127
rect 51511 286009 69393 286127
rect 69511 286009 87393 286127
rect 87511 286009 105393 286127
rect 105511 286009 123393 286127
rect 123511 286009 141393 286127
rect 141511 286009 159393 286127
rect 159511 286009 177393 286127
rect 177511 286009 195393 286127
rect 195511 286009 213393 286127
rect 213511 286009 231393 286127
rect 231511 286009 249393 286127
rect 249511 286009 267393 286127
rect 267511 286009 285393 286127
rect 285511 286009 296041 286127
rect 296159 286009 296250 286127
rect -4288 285967 296250 286009
rect -4288 285849 -4197 285967
rect -4079 285849 15393 285967
rect 15511 285849 33393 285967
rect 33511 285849 51393 285967
rect 51511 285849 69393 285967
rect 69511 285849 87393 285967
rect 87511 285849 105393 285967
rect 105511 285849 123393 285967
rect 123511 285849 141393 285967
rect 141511 285849 159393 285967
rect 159511 285849 177393 285967
rect 177511 285849 195393 285967
rect 195511 285849 213393 285967
rect 213511 285849 231393 285967
rect 231511 285849 249393 285967
rect 249511 285849 267393 285967
rect 267511 285849 285393 285967
rect 285511 285849 296041 285967
rect 296159 285849 296250 285967
rect -4288 285838 296250 285849
rect -4288 285837 -3988 285838
rect 15302 285837 15602 285838
rect 33302 285837 33602 285838
rect 51302 285837 51602 285838
rect 69302 285837 69602 285838
rect 87302 285837 87602 285838
rect 105302 285837 105602 285838
rect 123302 285837 123602 285838
rect 141302 285837 141602 285838
rect 159302 285837 159602 285838
rect 177302 285837 177602 285838
rect 195302 285837 195602 285838
rect 213302 285837 213602 285838
rect 231302 285837 231602 285838
rect 249302 285837 249602 285838
rect 267302 285837 267602 285838
rect 285302 285837 285602 285838
rect 295950 285837 296250 285838
rect -3348 284338 -3048 284339
rect 13502 284338 13802 284339
rect 31502 284338 31802 284339
rect 49502 284338 49802 284339
rect 67502 284338 67802 284339
rect 85502 284338 85802 284339
rect 103502 284338 103802 284339
rect 121502 284338 121802 284339
rect 139502 284338 139802 284339
rect 157502 284338 157802 284339
rect 175502 284338 175802 284339
rect 193502 284338 193802 284339
rect 211502 284338 211802 284339
rect 229502 284338 229802 284339
rect 247502 284338 247802 284339
rect 265502 284338 265802 284339
rect 283502 284338 283802 284339
rect 295010 284338 295310 284339
rect -3348 284327 295310 284338
rect -3348 284209 -3257 284327
rect -3139 284209 13593 284327
rect 13711 284209 31593 284327
rect 31711 284209 49593 284327
rect 49711 284209 67593 284327
rect 67711 284209 85593 284327
rect 85711 284209 103593 284327
rect 103711 284209 121593 284327
rect 121711 284209 139593 284327
rect 139711 284209 157593 284327
rect 157711 284209 175593 284327
rect 175711 284209 193593 284327
rect 193711 284209 211593 284327
rect 211711 284209 229593 284327
rect 229711 284209 247593 284327
rect 247711 284209 265593 284327
rect 265711 284209 283593 284327
rect 283711 284209 295101 284327
rect 295219 284209 295310 284327
rect -3348 284167 295310 284209
rect -3348 284049 -3257 284167
rect -3139 284049 13593 284167
rect 13711 284049 31593 284167
rect 31711 284049 49593 284167
rect 49711 284049 67593 284167
rect 67711 284049 85593 284167
rect 85711 284049 103593 284167
rect 103711 284049 121593 284167
rect 121711 284049 139593 284167
rect 139711 284049 157593 284167
rect 157711 284049 175593 284167
rect 175711 284049 193593 284167
rect 193711 284049 211593 284167
rect 211711 284049 229593 284167
rect 229711 284049 247593 284167
rect 247711 284049 265593 284167
rect 265711 284049 283593 284167
rect 283711 284049 295101 284167
rect 295219 284049 295310 284167
rect -3348 284038 295310 284049
rect -3348 284037 -3048 284038
rect 13502 284037 13802 284038
rect 31502 284037 31802 284038
rect 49502 284037 49802 284038
rect 67502 284037 67802 284038
rect 85502 284037 85802 284038
rect 103502 284037 103802 284038
rect 121502 284037 121802 284038
rect 139502 284037 139802 284038
rect 157502 284037 157802 284038
rect 175502 284037 175802 284038
rect 193502 284037 193802 284038
rect 211502 284037 211802 284038
rect 229502 284037 229802 284038
rect 247502 284037 247802 284038
rect 265502 284037 265802 284038
rect 283502 284037 283802 284038
rect 295010 284037 295310 284038
rect -2408 282538 -2108 282539
rect 11702 282538 12002 282539
rect 29702 282538 30002 282539
rect 47702 282538 48002 282539
rect 65702 282538 66002 282539
rect 83702 282538 84002 282539
rect 101702 282538 102002 282539
rect 119702 282538 120002 282539
rect 137702 282538 138002 282539
rect 155702 282538 156002 282539
rect 173702 282538 174002 282539
rect 191702 282538 192002 282539
rect 209702 282538 210002 282539
rect 227702 282538 228002 282539
rect 245702 282538 246002 282539
rect 263702 282538 264002 282539
rect 281702 282538 282002 282539
rect 294070 282538 294370 282539
rect -2408 282527 294370 282538
rect -2408 282409 -2317 282527
rect -2199 282409 11793 282527
rect 11911 282409 29793 282527
rect 29911 282409 47793 282527
rect 47911 282409 65793 282527
rect 65911 282409 83793 282527
rect 83911 282409 101793 282527
rect 101911 282409 119793 282527
rect 119911 282409 137793 282527
rect 137911 282409 155793 282527
rect 155911 282409 173793 282527
rect 173911 282409 191793 282527
rect 191911 282409 209793 282527
rect 209911 282409 227793 282527
rect 227911 282409 245793 282527
rect 245911 282409 263793 282527
rect 263911 282409 281793 282527
rect 281911 282409 294161 282527
rect 294279 282409 294370 282527
rect -2408 282367 294370 282409
rect -2408 282249 -2317 282367
rect -2199 282249 11793 282367
rect 11911 282249 29793 282367
rect 29911 282249 47793 282367
rect 47911 282249 65793 282367
rect 65911 282249 83793 282367
rect 83911 282249 101793 282367
rect 101911 282249 119793 282367
rect 119911 282249 137793 282367
rect 137911 282249 155793 282367
rect 155911 282249 173793 282367
rect 173911 282249 191793 282367
rect 191911 282249 209793 282367
rect 209911 282249 227793 282367
rect 227911 282249 245793 282367
rect 245911 282249 263793 282367
rect 263911 282249 281793 282367
rect 281911 282249 294161 282367
rect 294279 282249 294370 282367
rect -2408 282238 294370 282249
rect -2408 282237 -2108 282238
rect 11702 282237 12002 282238
rect 29702 282237 30002 282238
rect 47702 282237 48002 282238
rect 65702 282237 66002 282238
rect 83702 282237 84002 282238
rect 101702 282237 102002 282238
rect 119702 282237 120002 282238
rect 137702 282237 138002 282238
rect 155702 282237 156002 282238
rect 173702 282237 174002 282238
rect 191702 282237 192002 282238
rect 209702 282237 210002 282238
rect 227702 282237 228002 282238
rect 245702 282237 246002 282238
rect 263702 282237 264002 282238
rect 281702 282237 282002 282238
rect 294070 282237 294370 282238
rect -1468 280738 -1168 280739
rect 9902 280738 10202 280739
rect 27902 280738 28202 280739
rect 45902 280738 46202 280739
rect 63902 280738 64202 280739
rect 81902 280738 82202 280739
rect 99902 280738 100202 280739
rect 117902 280738 118202 280739
rect 135902 280738 136202 280739
rect 153902 280738 154202 280739
rect 171902 280738 172202 280739
rect 189902 280738 190202 280739
rect 207902 280738 208202 280739
rect 225902 280738 226202 280739
rect 243902 280738 244202 280739
rect 261902 280738 262202 280739
rect 279902 280738 280202 280739
rect 293130 280738 293430 280739
rect -1468 280727 293430 280738
rect -1468 280609 -1377 280727
rect -1259 280609 9993 280727
rect 10111 280609 27993 280727
rect 28111 280609 45993 280727
rect 46111 280609 63993 280727
rect 64111 280609 81993 280727
rect 82111 280609 99993 280727
rect 100111 280609 117993 280727
rect 118111 280609 135993 280727
rect 136111 280609 153993 280727
rect 154111 280609 171993 280727
rect 172111 280609 189993 280727
rect 190111 280609 207993 280727
rect 208111 280609 225993 280727
rect 226111 280609 243993 280727
rect 244111 280609 261993 280727
rect 262111 280609 279993 280727
rect 280111 280609 293221 280727
rect 293339 280609 293430 280727
rect -1468 280567 293430 280609
rect -1468 280449 -1377 280567
rect -1259 280449 9993 280567
rect 10111 280449 27993 280567
rect 28111 280449 45993 280567
rect 46111 280449 63993 280567
rect 64111 280449 81993 280567
rect 82111 280449 99993 280567
rect 100111 280449 117993 280567
rect 118111 280449 135993 280567
rect 136111 280449 153993 280567
rect 154111 280449 171993 280567
rect 172111 280449 189993 280567
rect 190111 280449 207993 280567
rect 208111 280449 225993 280567
rect 226111 280449 243993 280567
rect 244111 280449 261993 280567
rect 262111 280449 279993 280567
rect 280111 280449 293221 280567
rect 293339 280449 293430 280567
rect -1468 280438 293430 280449
rect -1468 280437 -1168 280438
rect 9902 280437 10202 280438
rect 27902 280437 28202 280438
rect 45902 280437 46202 280438
rect 63902 280437 64202 280438
rect 81902 280437 82202 280438
rect 99902 280437 100202 280438
rect 117902 280437 118202 280438
rect 135902 280437 136202 280438
rect 153902 280437 154202 280438
rect 171902 280437 172202 280438
rect 189902 280437 190202 280438
rect 207902 280437 208202 280438
rect 225902 280437 226202 280438
rect 243902 280437 244202 280438
rect 261902 280437 262202 280438
rect 279902 280437 280202 280438
rect 293130 280437 293430 280438
rect -3818 277138 -3518 277139
rect 6302 277138 6602 277139
rect 24302 277138 24602 277139
rect 42302 277138 42602 277139
rect 60302 277138 60602 277139
rect 78302 277138 78602 277139
rect 96302 277138 96602 277139
rect 114302 277138 114602 277139
rect 132302 277138 132602 277139
rect 150302 277138 150602 277139
rect 168302 277138 168602 277139
rect 186302 277138 186602 277139
rect 204302 277138 204602 277139
rect 222302 277138 222602 277139
rect 240302 277138 240602 277139
rect 258302 277138 258602 277139
rect 276302 277138 276602 277139
rect 295480 277138 295780 277139
rect -4288 277127 296250 277138
rect -4288 277009 -3727 277127
rect -3609 277009 6393 277127
rect 6511 277009 24393 277127
rect 24511 277009 42393 277127
rect 42511 277009 60393 277127
rect 60511 277009 78393 277127
rect 78511 277009 96393 277127
rect 96511 277009 114393 277127
rect 114511 277009 132393 277127
rect 132511 277009 150393 277127
rect 150511 277009 168393 277127
rect 168511 277009 186393 277127
rect 186511 277009 204393 277127
rect 204511 277009 222393 277127
rect 222511 277009 240393 277127
rect 240511 277009 258393 277127
rect 258511 277009 276393 277127
rect 276511 277009 295571 277127
rect 295689 277009 296250 277127
rect -4288 276967 296250 277009
rect -4288 276849 -3727 276967
rect -3609 276849 6393 276967
rect 6511 276849 24393 276967
rect 24511 276849 42393 276967
rect 42511 276849 60393 276967
rect 60511 276849 78393 276967
rect 78511 276849 96393 276967
rect 96511 276849 114393 276967
rect 114511 276849 132393 276967
rect 132511 276849 150393 276967
rect 150511 276849 168393 276967
rect 168511 276849 186393 276967
rect 186511 276849 204393 276967
rect 204511 276849 222393 276967
rect 222511 276849 240393 276967
rect 240511 276849 258393 276967
rect 258511 276849 276393 276967
rect 276511 276849 295571 276967
rect 295689 276849 296250 276967
rect -4288 276838 296250 276849
rect -3818 276837 -3518 276838
rect 6302 276837 6602 276838
rect 24302 276837 24602 276838
rect 42302 276837 42602 276838
rect 60302 276837 60602 276838
rect 78302 276837 78602 276838
rect 96302 276837 96602 276838
rect 114302 276837 114602 276838
rect 132302 276837 132602 276838
rect 150302 276837 150602 276838
rect 168302 276837 168602 276838
rect 186302 276837 186602 276838
rect 204302 276837 204602 276838
rect 222302 276837 222602 276838
rect 240302 276837 240602 276838
rect 258302 276837 258602 276838
rect 276302 276837 276602 276838
rect 295480 276837 295780 276838
rect -2878 275338 -2578 275339
rect 4502 275338 4802 275339
rect 22502 275338 22802 275339
rect 40502 275338 40802 275339
rect 58502 275338 58802 275339
rect 76502 275338 76802 275339
rect 94502 275338 94802 275339
rect 112502 275338 112802 275339
rect 130502 275338 130802 275339
rect 148502 275338 148802 275339
rect 166502 275338 166802 275339
rect 184502 275338 184802 275339
rect 202502 275338 202802 275339
rect 220502 275338 220802 275339
rect 238502 275338 238802 275339
rect 256502 275338 256802 275339
rect 274502 275338 274802 275339
rect 294540 275338 294840 275339
rect -3348 275327 295310 275338
rect -3348 275209 -2787 275327
rect -2669 275209 4593 275327
rect 4711 275209 22593 275327
rect 22711 275209 40593 275327
rect 40711 275209 58593 275327
rect 58711 275209 76593 275327
rect 76711 275209 94593 275327
rect 94711 275209 112593 275327
rect 112711 275209 130593 275327
rect 130711 275209 148593 275327
rect 148711 275209 166593 275327
rect 166711 275209 184593 275327
rect 184711 275209 202593 275327
rect 202711 275209 220593 275327
rect 220711 275209 238593 275327
rect 238711 275209 256593 275327
rect 256711 275209 274593 275327
rect 274711 275209 294631 275327
rect 294749 275209 295310 275327
rect -3348 275167 295310 275209
rect -3348 275049 -2787 275167
rect -2669 275049 4593 275167
rect 4711 275049 22593 275167
rect 22711 275049 40593 275167
rect 40711 275049 58593 275167
rect 58711 275049 76593 275167
rect 76711 275049 94593 275167
rect 94711 275049 112593 275167
rect 112711 275049 130593 275167
rect 130711 275049 148593 275167
rect 148711 275049 166593 275167
rect 166711 275049 184593 275167
rect 184711 275049 202593 275167
rect 202711 275049 220593 275167
rect 220711 275049 238593 275167
rect 238711 275049 256593 275167
rect 256711 275049 274593 275167
rect 274711 275049 294631 275167
rect 294749 275049 295310 275167
rect -3348 275038 295310 275049
rect -2878 275037 -2578 275038
rect 4502 275037 4802 275038
rect 22502 275037 22802 275038
rect 40502 275037 40802 275038
rect 58502 275037 58802 275038
rect 76502 275037 76802 275038
rect 94502 275037 94802 275038
rect 112502 275037 112802 275038
rect 130502 275037 130802 275038
rect 148502 275037 148802 275038
rect 166502 275037 166802 275038
rect 184502 275037 184802 275038
rect 202502 275037 202802 275038
rect 220502 275037 220802 275038
rect 238502 275037 238802 275038
rect 256502 275037 256802 275038
rect 274502 275037 274802 275038
rect 294540 275037 294840 275038
rect -1938 273538 -1638 273539
rect 2702 273538 3002 273539
rect 20702 273538 21002 273539
rect 38702 273538 39002 273539
rect 56702 273538 57002 273539
rect 74702 273538 75002 273539
rect 92702 273538 93002 273539
rect 110702 273538 111002 273539
rect 128702 273538 129002 273539
rect 146702 273538 147002 273539
rect 164702 273538 165002 273539
rect 182702 273538 183002 273539
rect 200702 273538 201002 273539
rect 218702 273538 219002 273539
rect 236702 273538 237002 273539
rect 254702 273538 255002 273539
rect 272702 273538 273002 273539
rect 290702 273538 291002 273539
rect 293600 273538 293900 273539
rect -2408 273527 294370 273538
rect -2408 273409 -1847 273527
rect -1729 273409 2793 273527
rect 2911 273409 20793 273527
rect 20911 273409 38793 273527
rect 38911 273409 56793 273527
rect 56911 273409 74793 273527
rect 74911 273409 92793 273527
rect 92911 273409 110793 273527
rect 110911 273409 128793 273527
rect 128911 273409 146793 273527
rect 146911 273409 164793 273527
rect 164911 273409 182793 273527
rect 182911 273409 200793 273527
rect 200911 273409 218793 273527
rect 218911 273409 236793 273527
rect 236911 273409 254793 273527
rect 254911 273409 272793 273527
rect 272911 273409 290793 273527
rect 290911 273409 293691 273527
rect 293809 273409 294370 273527
rect -2408 273367 294370 273409
rect -2408 273249 -1847 273367
rect -1729 273249 2793 273367
rect 2911 273249 20793 273367
rect 20911 273249 38793 273367
rect 38911 273249 56793 273367
rect 56911 273249 74793 273367
rect 74911 273249 92793 273367
rect 92911 273249 110793 273367
rect 110911 273249 128793 273367
rect 128911 273249 146793 273367
rect 146911 273249 164793 273367
rect 164911 273249 182793 273367
rect 182911 273249 200793 273367
rect 200911 273249 218793 273367
rect 218911 273249 236793 273367
rect 236911 273249 254793 273367
rect 254911 273249 272793 273367
rect 272911 273249 290793 273367
rect 290911 273249 293691 273367
rect 293809 273249 294370 273367
rect -2408 273238 294370 273249
rect -1938 273237 -1638 273238
rect 2702 273237 3002 273238
rect 20702 273237 21002 273238
rect 38702 273237 39002 273238
rect 56702 273237 57002 273238
rect 74702 273237 75002 273238
rect 92702 273237 93002 273238
rect 110702 273237 111002 273238
rect 128702 273237 129002 273238
rect 146702 273237 147002 273238
rect 164702 273237 165002 273238
rect 182702 273237 183002 273238
rect 200702 273237 201002 273238
rect 218702 273237 219002 273238
rect 236702 273237 237002 273238
rect 254702 273237 255002 273238
rect 272702 273237 273002 273238
rect 290702 273237 291002 273238
rect 293600 273237 293900 273238
rect -998 271738 -698 271739
rect 902 271738 1202 271739
rect 18902 271738 19202 271739
rect 36902 271738 37202 271739
rect 54902 271738 55202 271739
rect 72902 271738 73202 271739
rect 90902 271738 91202 271739
rect 108902 271738 109202 271739
rect 126902 271738 127202 271739
rect 144902 271738 145202 271739
rect 162902 271738 163202 271739
rect 180902 271738 181202 271739
rect 198902 271738 199202 271739
rect 216902 271738 217202 271739
rect 234902 271738 235202 271739
rect 252902 271738 253202 271739
rect 270902 271738 271202 271739
rect 288902 271738 289202 271739
rect 292660 271738 292960 271739
rect -1468 271727 293430 271738
rect -1468 271609 -907 271727
rect -789 271609 993 271727
rect 1111 271609 18993 271727
rect 19111 271609 36993 271727
rect 37111 271609 54993 271727
rect 55111 271609 72993 271727
rect 73111 271609 90993 271727
rect 91111 271609 108993 271727
rect 109111 271609 126993 271727
rect 127111 271609 144993 271727
rect 145111 271609 162993 271727
rect 163111 271609 180993 271727
rect 181111 271609 198993 271727
rect 199111 271609 216993 271727
rect 217111 271609 234993 271727
rect 235111 271609 252993 271727
rect 253111 271609 270993 271727
rect 271111 271609 288993 271727
rect 289111 271609 292751 271727
rect 292869 271609 293430 271727
rect -1468 271567 293430 271609
rect -1468 271449 -907 271567
rect -789 271449 993 271567
rect 1111 271449 18993 271567
rect 19111 271449 36993 271567
rect 37111 271449 54993 271567
rect 55111 271449 72993 271567
rect 73111 271449 90993 271567
rect 91111 271449 108993 271567
rect 109111 271449 126993 271567
rect 127111 271449 144993 271567
rect 145111 271449 162993 271567
rect 163111 271449 180993 271567
rect 181111 271449 198993 271567
rect 199111 271449 216993 271567
rect 217111 271449 234993 271567
rect 235111 271449 252993 271567
rect 253111 271449 270993 271567
rect 271111 271449 288993 271567
rect 289111 271449 292751 271567
rect 292869 271449 293430 271567
rect -1468 271438 293430 271449
rect -998 271437 -698 271438
rect 902 271437 1202 271438
rect 18902 271437 19202 271438
rect 36902 271437 37202 271438
rect 54902 271437 55202 271438
rect 72902 271437 73202 271438
rect 90902 271437 91202 271438
rect 108902 271437 109202 271438
rect 126902 271437 127202 271438
rect 144902 271437 145202 271438
rect 162902 271437 163202 271438
rect 180902 271437 181202 271438
rect 198902 271437 199202 271438
rect 216902 271437 217202 271438
rect 234902 271437 235202 271438
rect 252902 271437 253202 271438
rect 270902 271437 271202 271438
rect 288902 271437 289202 271438
rect 292660 271437 292960 271438
rect -4288 268138 -3988 268139
rect 15302 268138 15602 268139
rect 33302 268138 33602 268139
rect 51302 268138 51602 268139
rect 69302 268138 69602 268139
rect 87302 268138 87602 268139
rect 105302 268138 105602 268139
rect 123302 268138 123602 268139
rect 141302 268138 141602 268139
rect 159302 268138 159602 268139
rect 177302 268138 177602 268139
rect 195302 268138 195602 268139
rect 213302 268138 213602 268139
rect 231302 268138 231602 268139
rect 249302 268138 249602 268139
rect 267302 268138 267602 268139
rect 285302 268138 285602 268139
rect 295950 268138 296250 268139
rect -4288 268127 296250 268138
rect -4288 268009 -4197 268127
rect -4079 268009 15393 268127
rect 15511 268009 33393 268127
rect 33511 268009 51393 268127
rect 51511 268009 69393 268127
rect 69511 268009 87393 268127
rect 87511 268009 105393 268127
rect 105511 268009 123393 268127
rect 123511 268009 141393 268127
rect 141511 268009 159393 268127
rect 159511 268009 177393 268127
rect 177511 268009 195393 268127
rect 195511 268009 213393 268127
rect 213511 268009 231393 268127
rect 231511 268009 249393 268127
rect 249511 268009 267393 268127
rect 267511 268009 285393 268127
rect 285511 268009 296041 268127
rect 296159 268009 296250 268127
rect -4288 267967 296250 268009
rect -4288 267849 -4197 267967
rect -4079 267849 15393 267967
rect 15511 267849 33393 267967
rect 33511 267849 51393 267967
rect 51511 267849 69393 267967
rect 69511 267849 87393 267967
rect 87511 267849 105393 267967
rect 105511 267849 123393 267967
rect 123511 267849 141393 267967
rect 141511 267849 159393 267967
rect 159511 267849 177393 267967
rect 177511 267849 195393 267967
rect 195511 267849 213393 267967
rect 213511 267849 231393 267967
rect 231511 267849 249393 267967
rect 249511 267849 267393 267967
rect 267511 267849 285393 267967
rect 285511 267849 296041 267967
rect 296159 267849 296250 267967
rect -4288 267838 296250 267849
rect -4288 267837 -3988 267838
rect 15302 267837 15602 267838
rect 33302 267837 33602 267838
rect 51302 267837 51602 267838
rect 69302 267837 69602 267838
rect 87302 267837 87602 267838
rect 105302 267837 105602 267838
rect 123302 267837 123602 267838
rect 141302 267837 141602 267838
rect 159302 267837 159602 267838
rect 177302 267837 177602 267838
rect 195302 267837 195602 267838
rect 213302 267837 213602 267838
rect 231302 267837 231602 267838
rect 249302 267837 249602 267838
rect 267302 267837 267602 267838
rect 285302 267837 285602 267838
rect 295950 267837 296250 267838
rect -3348 266338 -3048 266339
rect 13502 266338 13802 266339
rect 31502 266338 31802 266339
rect 49502 266338 49802 266339
rect 67502 266338 67802 266339
rect 85502 266338 85802 266339
rect 103502 266338 103802 266339
rect 121502 266338 121802 266339
rect 139502 266338 139802 266339
rect 157502 266338 157802 266339
rect 175502 266338 175802 266339
rect 193502 266338 193802 266339
rect 211502 266338 211802 266339
rect 229502 266338 229802 266339
rect 247502 266338 247802 266339
rect 265502 266338 265802 266339
rect 283502 266338 283802 266339
rect 295010 266338 295310 266339
rect -3348 266327 295310 266338
rect -3348 266209 -3257 266327
rect -3139 266209 13593 266327
rect 13711 266209 31593 266327
rect 31711 266209 49593 266327
rect 49711 266209 67593 266327
rect 67711 266209 85593 266327
rect 85711 266209 103593 266327
rect 103711 266209 121593 266327
rect 121711 266209 139593 266327
rect 139711 266209 157593 266327
rect 157711 266209 175593 266327
rect 175711 266209 193593 266327
rect 193711 266209 211593 266327
rect 211711 266209 229593 266327
rect 229711 266209 247593 266327
rect 247711 266209 265593 266327
rect 265711 266209 283593 266327
rect 283711 266209 295101 266327
rect 295219 266209 295310 266327
rect -3348 266167 295310 266209
rect -3348 266049 -3257 266167
rect -3139 266049 13593 266167
rect 13711 266049 31593 266167
rect 31711 266049 49593 266167
rect 49711 266049 67593 266167
rect 67711 266049 85593 266167
rect 85711 266049 103593 266167
rect 103711 266049 121593 266167
rect 121711 266049 139593 266167
rect 139711 266049 157593 266167
rect 157711 266049 175593 266167
rect 175711 266049 193593 266167
rect 193711 266049 211593 266167
rect 211711 266049 229593 266167
rect 229711 266049 247593 266167
rect 247711 266049 265593 266167
rect 265711 266049 283593 266167
rect 283711 266049 295101 266167
rect 295219 266049 295310 266167
rect -3348 266038 295310 266049
rect -3348 266037 -3048 266038
rect 13502 266037 13802 266038
rect 31502 266037 31802 266038
rect 49502 266037 49802 266038
rect 67502 266037 67802 266038
rect 85502 266037 85802 266038
rect 103502 266037 103802 266038
rect 121502 266037 121802 266038
rect 139502 266037 139802 266038
rect 157502 266037 157802 266038
rect 175502 266037 175802 266038
rect 193502 266037 193802 266038
rect 211502 266037 211802 266038
rect 229502 266037 229802 266038
rect 247502 266037 247802 266038
rect 265502 266037 265802 266038
rect 283502 266037 283802 266038
rect 295010 266037 295310 266038
rect -2408 264538 -2108 264539
rect 11702 264538 12002 264539
rect 29702 264538 30002 264539
rect 47702 264538 48002 264539
rect 65702 264538 66002 264539
rect 83702 264538 84002 264539
rect 101702 264538 102002 264539
rect 119702 264538 120002 264539
rect 137702 264538 138002 264539
rect 155702 264538 156002 264539
rect 173702 264538 174002 264539
rect 191702 264538 192002 264539
rect 209702 264538 210002 264539
rect 227702 264538 228002 264539
rect 245702 264538 246002 264539
rect 263702 264538 264002 264539
rect 281702 264538 282002 264539
rect 294070 264538 294370 264539
rect -2408 264527 294370 264538
rect -2408 264409 -2317 264527
rect -2199 264409 11793 264527
rect 11911 264409 29793 264527
rect 29911 264409 47793 264527
rect 47911 264409 65793 264527
rect 65911 264409 83793 264527
rect 83911 264409 101793 264527
rect 101911 264409 119793 264527
rect 119911 264409 137793 264527
rect 137911 264409 155793 264527
rect 155911 264409 173793 264527
rect 173911 264409 191793 264527
rect 191911 264409 209793 264527
rect 209911 264409 227793 264527
rect 227911 264409 245793 264527
rect 245911 264409 263793 264527
rect 263911 264409 281793 264527
rect 281911 264409 294161 264527
rect 294279 264409 294370 264527
rect -2408 264367 294370 264409
rect -2408 264249 -2317 264367
rect -2199 264249 11793 264367
rect 11911 264249 29793 264367
rect 29911 264249 47793 264367
rect 47911 264249 65793 264367
rect 65911 264249 83793 264367
rect 83911 264249 101793 264367
rect 101911 264249 119793 264367
rect 119911 264249 137793 264367
rect 137911 264249 155793 264367
rect 155911 264249 173793 264367
rect 173911 264249 191793 264367
rect 191911 264249 209793 264367
rect 209911 264249 227793 264367
rect 227911 264249 245793 264367
rect 245911 264249 263793 264367
rect 263911 264249 281793 264367
rect 281911 264249 294161 264367
rect 294279 264249 294370 264367
rect -2408 264238 294370 264249
rect -2408 264237 -2108 264238
rect 11702 264237 12002 264238
rect 29702 264237 30002 264238
rect 47702 264237 48002 264238
rect 65702 264237 66002 264238
rect 83702 264237 84002 264238
rect 101702 264237 102002 264238
rect 119702 264237 120002 264238
rect 137702 264237 138002 264238
rect 155702 264237 156002 264238
rect 173702 264237 174002 264238
rect 191702 264237 192002 264238
rect 209702 264237 210002 264238
rect 227702 264237 228002 264238
rect 245702 264237 246002 264238
rect 263702 264237 264002 264238
rect 281702 264237 282002 264238
rect 294070 264237 294370 264238
rect -1468 262738 -1168 262739
rect 9902 262738 10202 262739
rect 27902 262738 28202 262739
rect 45902 262738 46202 262739
rect 63902 262738 64202 262739
rect 81902 262738 82202 262739
rect 99902 262738 100202 262739
rect 117902 262738 118202 262739
rect 135902 262738 136202 262739
rect 153902 262738 154202 262739
rect 171902 262738 172202 262739
rect 189902 262738 190202 262739
rect 207902 262738 208202 262739
rect 225902 262738 226202 262739
rect 243902 262738 244202 262739
rect 261902 262738 262202 262739
rect 279902 262738 280202 262739
rect 293130 262738 293430 262739
rect -1468 262727 293430 262738
rect -1468 262609 -1377 262727
rect -1259 262609 9993 262727
rect 10111 262609 27993 262727
rect 28111 262609 45993 262727
rect 46111 262609 63993 262727
rect 64111 262609 81993 262727
rect 82111 262609 99993 262727
rect 100111 262609 117993 262727
rect 118111 262609 135993 262727
rect 136111 262609 153993 262727
rect 154111 262609 171993 262727
rect 172111 262609 189993 262727
rect 190111 262609 207993 262727
rect 208111 262609 225993 262727
rect 226111 262609 243993 262727
rect 244111 262609 261993 262727
rect 262111 262609 279993 262727
rect 280111 262609 293221 262727
rect 293339 262609 293430 262727
rect -1468 262567 293430 262609
rect -1468 262449 -1377 262567
rect -1259 262449 9993 262567
rect 10111 262449 27993 262567
rect 28111 262449 45993 262567
rect 46111 262449 63993 262567
rect 64111 262449 81993 262567
rect 82111 262449 99993 262567
rect 100111 262449 117993 262567
rect 118111 262449 135993 262567
rect 136111 262449 153993 262567
rect 154111 262449 171993 262567
rect 172111 262449 189993 262567
rect 190111 262449 207993 262567
rect 208111 262449 225993 262567
rect 226111 262449 243993 262567
rect 244111 262449 261993 262567
rect 262111 262449 279993 262567
rect 280111 262449 293221 262567
rect 293339 262449 293430 262567
rect -1468 262438 293430 262449
rect -1468 262437 -1168 262438
rect 9902 262437 10202 262438
rect 27902 262437 28202 262438
rect 45902 262437 46202 262438
rect 63902 262437 64202 262438
rect 81902 262437 82202 262438
rect 99902 262437 100202 262438
rect 117902 262437 118202 262438
rect 135902 262437 136202 262438
rect 153902 262437 154202 262438
rect 171902 262437 172202 262438
rect 189902 262437 190202 262438
rect 207902 262437 208202 262438
rect 225902 262437 226202 262438
rect 243902 262437 244202 262438
rect 261902 262437 262202 262438
rect 279902 262437 280202 262438
rect 293130 262437 293430 262438
rect -3818 259138 -3518 259139
rect 6302 259138 6602 259139
rect 24302 259138 24602 259139
rect 42302 259138 42602 259139
rect 60302 259138 60602 259139
rect 78302 259138 78602 259139
rect 96302 259138 96602 259139
rect 114302 259138 114602 259139
rect 132302 259138 132602 259139
rect 150302 259138 150602 259139
rect 168302 259138 168602 259139
rect 186302 259138 186602 259139
rect 204302 259138 204602 259139
rect 222302 259138 222602 259139
rect 240302 259138 240602 259139
rect 258302 259138 258602 259139
rect 276302 259138 276602 259139
rect 295480 259138 295780 259139
rect -4288 259127 296250 259138
rect -4288 259009 -3727 259127
rect -3609 259009 6393 259127
rect 6511 259009 24393 259127
rect 24511 259009 42393 259127
rect 42511 259009 60393 259127
rect 60511 259009 78393 259127
rect 78511 259009 96393 259127
rect 96511 259009 114393 259127
rect 114511 259009 132393 259127
rect 132511 259009 150393 259127
rect 150511 259009 168393 259127
rect 168511 259009 186393 259127
rect 186511 259009 204393 259127
rect 204511 259009 222393 259127
rect 222511 259009 240393 259127
rect 240511 259009 258393 259127
rect 258511 259009 276393 259127
rect 276511 259009 295571 259127
rect 295689 259009 296250 259127
rect -4288 258967 296250 259009
rect -4288 258849 -3727 258967
rect -3609 258849 6393 258967
rect 6511 258849 24393 258967
rect 24511 258849 42393 258967
rect 42511 258849 60393 258967
rect 60511 258849 78393 258967
rect 78511 258849 96393 258967
rect 96511 258849 114393 258967
rect 114511 258849 132393 258967
rect 132511 258849 150393 258967
rect 150511 258849 168393 258967
rect 168511 258849 186393 258967
rect 186511 258849 204393 258967
rect 204511 258849 222393 258967
rect 222511 258849 240393 258967
rect 240511 258849 258393 258967
rect 258511 258849 276393 258967
rect 276511 258849 295571 258967
rect 295689 258849 296250 258967
rect -4288 258838 296250 258849
rect -3818 258837 -3518 258838
rect 6302 258837 6602 258838
rect 24302 258837 24602 258838
rect 42302 258837 42602 258838
rect 60302 258837 60602 258838
rect 78302 258837 78602 258838
rect 96302 258837 96602 258838
rect 114302 258837 114602 258838
rect 132302 258837 132602 258838
rect 150302 258837 150602 258838
rect 168302 258837 168602 258838
rect 186302 258837 186602 258838
rect 204302 258837 204602 258838
rect 222302 258837 222602 258838
rect 240302 258837 240602 258838
rect 258302 258837 258602 258838
rect 276302 258837 276602 258838
rect 295480 258837 295780 258838
rect -2878 257338 -2578 257339
rect 4502 257338 4802 257339
rect 22502 257338 22802 257339
rect 40502 257338 40802 257339
rect 58502 257338 58802 257339
rect 76502 257338 76802 257339
rect 94502 257338 94802 257339
rect 112502 257338 112802 257339
rect 130502 257338 130802 257339
rect 148502 257338 148802 257339
rect 166502 257338 166802 257339
rect 184502 257338 184802 257339
rect 202502 257338 202802 257339
rect 220502 257338 220802 257339
rect 238502 257338 238802 257339
rect 256502 257338 256802 257339
rect 274502 257338 274802 257339
rect 294540 257338 294840 257339
rect -3348 257327 295310 257338
rect -3348 257209 -2787 257327
rect -2669 257209 4593 257327
rect 4711 257209 22593 257327
rect 22711 257209 40593 257327
rect 40711 257209 58593 257327
rect 58711 257209 76593 257327
rect 76711 257209 94593 257327
rect 94711 257209 112593 257327
rect 112711 257209 130593 257327
rect 130711 257209 148593 257327
rect 148711 257209 166593 257327
rect 166711 257209 184593 257327
rect 184711 257209 202593 257327
rect 202711 257209 220593 257327
rect 220711 257209 238593 257327
rect 238711 257209 256593 257327
rect 256711 257209 274593 257327
rect 274711 257209 294631 257327
rect 294749 257209 295310 257327
rect -3348 257167 295310 257209
rect -3348 257049 -2787 257167
rect -2669 257049 4593 257167
rect 4711 257049 22593 257167
rect 22711 257049 40593 257167
rect 40711 257049 58593 257167
rect 58711 257049 76593 257167
rect 76711 257049 94593 257167
rect 94711 257049 112593 257167
rect 112711 257049 130593 257167
rect 130711 257049 148593 257167
rect 148711 257049 166593 257167
rect 166711 257049 184593 257167
rect 184711 257049 202593 257167
rect 202711 257049 220593 257167
rect 220711 257049 238593 257167
rect 238711 257049 256593 257167
rect 256711 257049 274593 257167
rect 274711 257049 294631 257167
rect 294749 257049 295310 257167
rect -3348 257038 295310 257049
rect -2878 257037 -2578 257038
rect 4502 257037 4802 257038
rect 22502 257037 22802 257038
rect 40502 257037 40802 257038
rect 58502 257037 58802 257038
rect 76502 257037 76802 257038
rect 94502 257037 94802 257038
rect 112502 257037 112802 257038
rect 130502 257037 130802 257038
rect 148502 257037 148802 257038
rect 166502 257037 166802 257038
rect 184502 257037 184802 257038
rect 202502 257037 202802 257038
rect 220502 257037 220802 257038
rect 238502 257037 238802 257038
rect 256502 257037 256802 257038
rect 274502 257037 274802 257038
rect 294540 257037 294840 257038
rect -1938 255538 -1638 255539
rect 2702 255538 3002 255539
rect 20702 255538 21002 255539
rect 38702 255538 39002 255539
rect 56702 255538 57002 255539
rect 74702 255538 75002 255539
rect 92702 255538 93002 255539
rect 110702 255538 111002 255539
rect 128702 255538 129002 255539
rect 146702 255538 147002 255539
rect 164702 255538 165002 255539
rect 182702 255538 183002 255539
rect 200702 255538 201002 255539
rect 218702 255538 219002 255539
rect 236702 255538 237002 255539
rect 254702 255538 255002 255539
rect 272702 255538 273002 255539
rect 290702 255538 291002 255539
rect 293600 255538 293900 255539
rect -2408 255527 294370 255538
rect -2408 255409 -1847 255527
rect -1729 255409 2793 255527
rect 2911 255409 20793 255527
rect 20911 255409 38793 255527
rect 38911 255409 56793 255527
rect 56911 255409 74793 255527
rect 74911 255409 92793 255527
rect 92911 255409 110793 255527
rect 110911 255409 128793 255527
rect 128911 255409 146793 255527
rect 146911 255409 164793 255527
rect 164911 255409 182793 255527
rect 182911 255409 200793 255527
rect 200911 255409 218793 255527
rect 218911 255409 236793 255527
rect 236911 255409 254793 255527
rect 254911 255409 272793 255527
rect 272911 255409 290793 255527
rect 290911 255409 293691 255527
rect 293809 255409 294370 255527
rect -2408 255367 294370 255409
rect -2408 255249 -1847 255367
rect -1729 255249 2793 255367
rect 2911 255249 20793 255367
rect 20911 255249 38793 255367
rect 38911 255249 56793 255367
rect 56911 255249 74793 255367
rect 74911 255249 92793 255367
rect 92911 255249 110793 255367
rect 110911 255249 128793 255367
rect 128911 255249 146793 255367
rect 146911 255249 164793 255367
rect 164911 255249 182793 255367
rect 182911 255249 200793 255367
rect 200911 255249 218793 255367
rect 218911 255249 236793 255367
rect 236911 255249 254793 255367
rect 254911 255249 272793 255367
rect 272911 255249 290793 255367
rect 290911 255249 293691 255367
rect 293809 255249 294370 255367
rect -2408 255238 294370 255249
rect -1938 255237 -1638 255238
rect 2702 255237 3002 255238
rect 20702 255237 21002 255238
rect 38702 255237 39002 255238
rect 56702 255237 57002 255238
rect 74702 255237 75002 255238
rect 92702 255237 93002 255238
rect 110702 255237 111002 255238
rect 128702 255237 129002 255238
rect 146702 255237 147002 255238
rect 164702 255237 165002 255238
rect 182702 255237 183002 255238
rect 200702 255237 201002 255238
rect 218702 255237 219002 255238
rect 236702 255237 237002 255238
rect 254702 255237 255002 255238
rect 272702 255237 273002 255238
rect 290702 255237 291002 255238
rect 293600 255237 293900 255238
rect -998 253738 -698 253739
rect 902 253738 1202 253739
rect 18902 253738 19202 253739
rect 36902 253738 37202 253739
rect 54902 253738 55202 253739
rect 72902 253738 73202 253739
rect 90902 253738 91202 253739
rect 108902 253738 109202 253739
rect 126902 253738 127202 253739
rect 144902 253738 145202 253739
rect 162902 253738 163202 253739
rect 180902 253738 181202 253739
rect 198902 253738 199202 253739
rect 216902 253738 217202 253739
rect 234902 253738 235202 253739
rect 252902 253738 253202 253739
rect 270902 253738 271202 253739
rect 288902 253738 289202 253739
rect 292660 253738 292960 253739
rect -1468 253727 293430 253738
rect -1468 253609 -907 253727
rect -789 253609 993 253727
rect 1111 253609 18993 253727
rect 19111 253609 36993 253727
rect 37111 253609 54993 253727
rect 55111 253609 72993 253727
rect 73111 253609 90993 253727
rect 91111 253609 108993 253727
rect 109111 253609 126993 253727
rect 127111 253609 144993 253727
rect 145111 253609 162993 253727
rect 163111 253609 180993 253727
rect 181111 253609 198993 253727
rect 199111 253609 216993 253727
rect 217111 253609 234993 253727
rect 235111 253609 252993 253727
rect 253111 253609 270993 253727
rect 271111 253609 288993 253727
rect 289111 253609 292751 253727
rect 292869 253609 293430 253727
rect -1468 253567 293430 253609
rect -1468 253449 -907 253567
rect -789 253449 993 253567
rect 1111 253449 18993 253567
rect 19111 253449 36993 253567
rect 37111 253449 54993 253567
rect 55111 253449 72993 253567
rect 73111 253449 90993 253567
rect 91111 253449 108993 253567
rect 109111 253449 126993 253567
rect 127111 253449 144993 253567
rect 145111 253449 162993 253567
rect 163111 253449 180993 253567
rect 181111 253449 198993 253567
rect 199111 253449 216993 253567
rect 217111 253449 234993 253567
rect 235111 253449 252993 253567
rect 253111 253449 270993 253567
rect 271111 253449 288993 253567
rect 289111 253449 292751 253567
rect 292869 253449 293430 253567
rect -1468 253438 293430 253449
rect -998 253437 -698 253438
rect 902 253437 1202 253438
rect 18902 253437 19202 253438
rect 36902 253437 37202 253438
rect 54902 253437 55202 253438
rect 72902 253437 73202 253438
rect 90902 253437 91202 253438
rect 108902 253437 109202 253438
rect 126902 253437 127202 253438
rect 144902 253437 145202 253438
rect 162902 253437 163202 253438
rect 180902 253437 181202 253438
rect 198902 253437 199202 253438
rect 216902 253437 217202 253438
rect 234902 253437 235202 253438
rect 252902 253437 253202 253438
rect 270902 253437 271202 253438
rect 288902 253437 289202 253438
rect 292660 253437 292960 253438
rect -4288 250138 -3988 250139
rect 15302 250138 15602 250139
rect 33302 250138 33602 250139
rect 51302 250138 51602 250139
rect 69302 250138 69602 250139
rect 87302 250138 87602 250139
rect 105302 250138 105602 250139
rect 123302 250138 123602 250139
rect 141302 250138 141602 250139
rect 159302 250138 159602 250139
rect 177302 250138 177602 250139
rect 195302 250138 195602 250139
rect 213302 250138 213602 250139
rect 231302 250138 231602 250139
rect 249302 250138 249602 250139
rect 267302 250138 267602 250139
rect 285302 250138 285602 250139
rect 295950 250138 296250 250139
rect -4288 250127 296250 250138
rect -4288 250009 -4197 250127
rect -4079 250009 15393 250127
rect 15511 250009 33393 250127
rect 33511 250009 51393 250127
rect 51511 250009 69393 250127
rect 69511 250009 87393 250127
rect 87511 250009 105393 250127
rect 105511 250009 123393 250127
rect 123511 250009 141393 250127
rect 141511 250009 159393 250127
rect 159511 250009 177393 250127
rect 177511 250009 195393 250127
rect 195511 250009 213393 250127
rect 213511 250009 231393 250127
rect 231511 250009 249393 250127
rect 249511 250009 267393 250127
rect 267511 250009 285393 250127
rect 285511 250009 296041 250127
rect 296159 250009 296250 250127
rect -4288 249967 296250 250009
rect -4288 249849 -4197 249967
rect -4079 249849 15393 249967
rect 15511 249849 33393 249967
rect 33511 249849 51393 249967
rect 51511 249849 69393 249967
rect 69511 249849 87393 249967
rect 87511 249849 105393 249967
rect 105511 249849 123393 249967
rect 123511 249849 141393 249967
rect 141511 249849 159393 249967
rect 159511 249849 177393 249967
rect 177511 249849 195393 249967
rect 195511 249849 213393 249967
rect 213511 249849 231393 249967
rect 231511 249849 249393 249967
rect 249511 249849 267393 249967
rect 267511 249849 285393 249967
rect 285511 249849 296041 249967
rect 296159 249849 296250 249967
rect -4288 249838 296250 249849
rect -4288 249837 -3988 249838
rect 15302 249837 15602 249838
rect 33302 249837 33602 249838
rect 51302 249837 51602 249838
rect 69302 249837 69602 249838
rect 87302 249837 87602 249838
rect 105302 249837 105602 249838
rect 123302 249837 123602 249838
rect 141302 249837 141602 249838
rect 159302 249837 159602 249838
rect 177302 249837 177602 249838
rect 195302 249837 195602 249838
rect 213302 249837 213602 249838
rect 231302 249837 231602 249838
rect 249302 249837 249602 249838
rect 267302 249837 267602 249838
rect 285302 249837 285602 249838
rect 295950 249837 296250 249838
rect -3348 248338 -3048 248339
rect 13502 248338 13802 248339
rect 31502 248338 31802 248339
rect 49502 248338 49802 248339
rect 67502 248338 67802 248339
rect 85502 248338 85802 248339
rect 103502 248338 103802 248339
rect 121502 248338 121802 248339
rect 139502 248338 139802 248339
rect 157502 248338 157802 248339
rect 175502 248338 175802 248339
rect 193502 248338 193802 248339
rect 211502 248338 211802 248339
rect 229502 248338 229802 248339
rect 247502 248338 247802 248339
rect 265502 248338 265802 248339
rect 283502 248338 283802 248339
rect 295010 248338 295310 248339
rect -3348 248327 295310 248338
rect -3348 248209 -3257 248327
rect -3139 248209 13593 248327
rect 13711 248209 31593 248327
rect 31711 248209 49593 248327
rect 49711 248209 67593 248327
rect 67711 248209 85593 248327
rect 85711 248209 103593 248327
rect 103711 248209 121593 248327
rect 121711 248209 139593 248327
rect 139711 248209 157593 248327
rect 157711 248209 175593 248327
rect 175711 248209 193593 248327
rect 193711 248209 211593 248327
rect 211711 248209 229593 248327
rect 229711 248209 247593 248327
rect 247711 248209 265593 248327
rect 265711 248209 283593 248327
rect 283711 248209 295101 248327
rect 295219 248209 295310 248327
rect -3348 248167 295310 248209
rect -3348 248049 -3257 248167
rect -3139 248049 13593 248167
rect 13711 248049 31593 248167
rect 31711 248049 49593 248167
rect 49711 248049 67593 248167
rect 67711 248049 85593 248167
rect 85711 248049 103593 248167
rect 103711 248049 121593 248167
rect 121711 248049 139593 248167
rect 139711 248049 157593 248167
rect 157711 248049 175593 248167
rect 175711 248049 193593 248167
rect 193711 248049 211593 248167
rect 211711 248049 229593 248167
rect 229711 248049 247593 248167
rect 247711 248049 265593 248167
rect 265711 248049 283593 248167
rect 283711 248049 295101 248167
rect 295219 248049 295310 248167
rect -3348 248038 295310 248049
rect -3348 248037 -3048 248038
rect 13502 248037 13802 248038
rect 31502 248037 31802 248038
rect 49502 248037 49802 248038
rect 67502 248037 67802 248038
rect 85502 248037 85802 248038
rect 103502 248037 103802 248038
rect 121502 248037 121802 248038
rect 139502 248037 139802 248038
rect 157502 248037 157802 248038
rect 175502 248037 175802 248038
rect 193502 248037 193802 248038
rect 211502 248037 211802 248038
rect 229502 248037 229802 248038
rect 247502 248037 247802 248038
rect 265502 248037 265802 248038
rect 283502 248037 283802 248038
rect 295010 248037 295310 248038
rect -2408 246538 -2108 246539
rect 11702 246538 12002 246539
rect 29702 246538 30002 246539
rect 47702 246538 48002 246539
rect 65702 246538 66002 246539
rect 83702 246538 84002 246539
rect 101702 246538 102002 246539
rect 119702 246538 120002 246539
rect 137702 246538 138002 246539
rect 155702 246538 156002 246539
rect 173702 246538 174002 246539
rect 191702 246538 192002 246539
rect 209702 246538 210002 246539
rect 227702 246538 228002 246539
rect 245702 246538 246002 246539
rect 263702 246538 264002 246539
rect 281702 246538 282002 246539
rect 294070 246538 294370 246539
rect -2408 246527 294370 246538
rect -2408 246409 -2317 246527
rect -2199 246409 11793 246527
rect 11911 246409 29793 246527
rect 29911 246409 47793 246527
rect 47911 246409 65793 246527
rect 65911 246409 83793 246527
rect 83911 246409 101793 246527
rect 101911 246409 119793 246527
rect 119911 246409 137793 246527
rect 137911 246409 155793 246527
rect 155911 246409 173793 246527
rect 173911 246409 191793 246527
rect 191911 246409 209793 246527
rect 209911 246409 227793 246527
rect 227911 246409 245793 246527
rect 245911 246409 263793 246527
rect 263911 246409 281793 246527
rect 281911 246409 294161 246527
rect 294279 246409 294370 246527
rect -2408 246367 294370 246409
rect -2408 246249 -2317 246367
rect -2199 246249 11793 246367
rect 11911 246249 29793 246367
rect 29911 246249 47793 246367
rect 47911 246249 65793 246367
rect 65911 246249 83793 246367
rect 83911 246249 101793 246367
rect 101911 246249 119793 246367
rect 119911 246249 137793 246367
rect 137911 246249 155793 246367
rect 155911 246249 173793 246367
rect 173911 246249 191793 246367
rect 191911 246249 209793 246367
rect 209911 246249 227793 246367
rect 227911 246249 245793 246367
rect 245911 246249 263793 246367
rect 263911 246249 281793 246367
rect 281911 246249 294161 246367
rect 294279 246249 294370 246367
rect -2408 246238 294370 246249
rect -2408 246237 -2108 246238
rect 11702 246237 12002 246238
rect 29702 246237 30002 246238
rect 47702 246237 48002 246238
rect 65702 246237 66002 246238
rect 83702 246237 84002 246238
rect 101702 246237 102002 246238
rect 119702 246237 120002 246238
rect 137702 246237 138002 246238
rect 155702 246237 156002 246238
rect 173702 246237 174002 246238
rect 191702 246237 192002 246238
rect 209702 246237 210002 246238
rect 227702 246237 228002 246238
rect 245702 246237 246002 246238
rect 263702 246237 264002 246238
rect 281702 246237 282002 246238
rect 294070 246237 294370 246238
rect -1468 244738 -1168 244739
rect 9902 244738 10202 244739
rect 27902 244738 28202 244739
rect 45902 244738 46202 244739
rect 63902 244738 64202 244739
rect 81902 244738 82202 244739
rect 99902 244738 100202 244739
rect 117902 244738 118202 244739
rect 135902 244738 136202 244739
rect 153902 244738 154202 244739
rect 171902 244738 172202 244739
rect 189902 244738 190202 244739
rect 207902 244738 208202 244739
rect 225902 244738 226202 244739
rect 243902 244738 244202 244739
rect 261902 244738 262202 244739
rect 279902 244738 280202 244739
rect 293130 244738 293430 244739
rect -1468 244727 293430 244738
rect -1468 244609 -1377 244727
rect -1259 244609 9993 244727
rect 10111 244609 27993 244727
rect 28111 244609 45993 244727
rect 46111 244609 63993 244727
rect 64111 244609 81993 244727
rect 82111 244609 99993 244727
rect 100111 244609 117993 244727
rect 118111 244609 135993 244727
rect 136111 244609 153993 244727
rect 154111 244609 171993 244727
rect 172111 244609 189993 244727
rect 190111 244609 207993 244727
rect 208111 244609 225993 244727
rect 226111 244609 243993 244727
rect 244111 244609 261993 244727
rect 262111 244609 279993 244727
rect 280111 244609 293221 244727
rect 293339 244609 293430 244727
rect -1468 244567 293430 244609
rect -1468 244449 -1377 244567
rect -1259 244449 9993 244567
rect 10111 244449 27993 244567
rect 28111 244449 45993 244567
rect 46111 244449 63993 244567
rect 64111 244449 81993 244567
rect 82111 244449 99993 244567
rect 100111 244449 117993 244567
rect 118111 244449 135993 244567
rect 136111 244449 153993 244567
rect 154111 244449 171993 244567
rect 172111 244449 189993 244567
rect 190111 244449 207993 244567
rect 208111 244449 225993 244567
rect 226111 244449 243993 244567
rect 244111 244449 261993 244567
rect 262111 244449 279993 244567
rect 280111 244449 293221 244567
rect 293339 244449 293430 244567
rect -1468 244438 293430 244449
rect -1468 244437 -1168 244438
rect 9902 244437 10202 244438
rect 27902 244437 28202 244438
rect 45902 244437 46202 244438
rect 63902 244437 64202 244438
rect 81902 244437 82202 244438
rect 99902 244437 100202 244438
rect 117902 244437 118202 244438
rect 135902 244437 136202 244438
rect 153902 244437 154202 244438
rect 171902 244437 172202 244438
rect 189902 244437 190202 244438
rect 207902 244437 208202 244438
rect 225902 244437 226202 244438
rect 243902 244437 244202 244438
rect 261902 244437 262202 244438
rect 279902 244437 280202 244438
rect 293130 244437 293430 244438
rect -3818 241138 -3518 241139
rect 6302 241138 6602 241139
rect 24302 241138 24602 241139
rect 42302 241138 42602 241139
rect 60302 241138 60602 241139
rect 78302 241138 78602 241139
rect 96302 241138 96602 241139
rect 114302 241138 114602 241139
rect 132302 241138 132602 241139
rect 150302 241138 150602 241139
rect 168302 241138 168602 241139
rect 186302 241138 186602 241139
rect 204302 241138 204602 241139
rect 222302 241138 222602 241139
rect 240302 241138 240602 241139
rect 258302 241138 258602 241139
rect 276302 241138 276602 241139
rect 295480 241138 295780 241139
rect -4288 241127 296250 241138
rect -4288 241009 -3727 241127
rect -3609 241009 6393 241127
rect 6511 241009 24393 241127
rect 24511 241009 42393 241127
rect 42511 241009 60393 241127
rect 60511 241009 78393 241127
rect 78511 241009 96393 241127
rect 96511 241009 114393 241127
rect 114511 241009 132393 241127
rect 132511 241009 150393 241127
rect 150511 241009 168393 241127
rect 168511 241009 186393 241127
rect 186511 241009 204393 241127
rect 204511 241009 222393 241127
rect 222511 241009 240393 241127
rect 240511 241009 258393 241127
rect 258511 241009 276393 241127
rect 276511 241009 295571 241127
rect 295689 241009 296250 241127
rect -4288 240967 296250 241009
rect -4288 240849 -3727 240967
rect -3609 240849 6393 240967
rect 6511 240849 24393 240967
rect 24511 240849 42393 240967
rect 42511 240849 60393 240967
rect 60511 240849 78393 240967
rect 78511 240849 96393 240967
rect 96511 240849 114393 240967
rect 114511 240849 132393 240967
rect 132511 240849 150393 240967
rect 150511 240849 168393 240967
rect 168511 240849 186393 240967
rect 186511 240849 204393 240967
rect 204511 240849 222393 240967
rect 222511 240849 240393 240967
rect 240511 240849 258393 240967
rect 258511 240849 276393 240967
rect 276511 240849 295571 240967
rect 295689 240849 296250 240967
rect -4288 240838 296250 240849
rect -3818 240837 -3518 240838
rect 6302 240837 6602 240838
rect 24302 240837 24602 240838
rect 42302 240837 42602 240838
rect 60302 240837 60602 240838
rect 78302 240837 78602 240838
rect 96302 240837 96602 240838
rect 114302 240837 114602 240838
rect 132302 240837 132602 240838
rect 150302 240837 150602 240838
rect 168302 240837 168602 240838
rect 186302 240837 186602 240838
rect 204302 240837 204602 240838
rect 222302 240837 222602 240838
rect 240302 240837 240602 240838
rect 258302 240837 258602 240838
rect 276302 240837 276602 240838
rect 295480 240837 295780 240838
rect -2878 239338 -2578 239339
rect 4502 239338 4802 239339
rect 22502 239338 22802 239339
rect 40502 239338 40802 239339
rect 58502 239338 58802 239339
rect 76502 239338 76802 239339
rect 94502 239338 94802 239339
rect 112502 239338 112802 239339
rect 130502 239338 130802 239339
rect 148502 239338 148802 239339
rect 166502 239338 166802 239339
rect 184502 239338 184802 239339
rect 202502 239338 202802 239339
rect 220502 239338 220802 239339
rect 238502 239338 238802 239339
rect 256502 239338 256802 239339
rect 274502 239338 274802 239339
rect 294540 239338 294840 239339
rect -3348 239327 295310 239338
rect -3348 239209 -2787 239327
rect -2669 239209 4593 239327
rect 4711 239209 22593 239327
rect 22711 239209 40593 239327
rect 40711 239209 58593 239327
rect 58711 239209 76593 239327
rect 76711 239209 94593 239327
rect 94711 239209 112593 239327
rect 112711 239209 130593 239327
rect 130711 239209 148593 239327
rect 148711 239209 166593 239327
rect 166711 239209 184593 239327
rect 184711 239209 202593 239327
rect 202711 239209 220593 239327
rect 220711 239209 238593 239327
rect 238711 239209 256593 239327
rect 256711 239209 274593 239327
rect 274711 239209 294631 239327
rect 294749 239209 295310 239327
rect -3348 239167 295310 239209
rect -3348 239049 -2787 239167
rect -2669 239049 4593 239167
rect 4711 239049 22593 239167
rect 22711 239049 40593 239167
rect 40711 239049 58593 239167
rect 58711 239049 76593 239167
rect 76711 239049 94593 239167
rect 94711 239049 112593 239167
rect 112711 239049 130593 239167
rect 130711 239049 148593 239167
rect 148711 239049 166593 239167
rect 166711 239049 184593 239167
rect 184711 239049 202593 239167
rect 202711 239049 220593 239167
rect 220711 239049 238593 239167
rect 238711 239049 256593 239167
rect 256711 239049 274593 239167
rect 274711 239049 294631 239167
rect 294749 239049 295310 239167
rect -3348 239038 295310 239049
rect -2878 239037 -2578 239038
rect 4502 239037 4802 239038
rect 22502 239037 22802 239038
rect 40502 239037 40802 239038
rect 58502 239037 58802 239038
rect 76502 239037 76802 239038
rect 94502 239037 94802 239038
rect 112502 239037 112802 239038
rect 130502 239037 130802 239038
rect 148502 239037 148802 239038
rect 166502 239037 166802 239038
rect 184502 239037 184802 239038
rect 202502 239037 202802 239038
rect 220502 239037 220802 239038
rect 238502 239037 238802 239038
rect 256502 239037 256802 239038
rect 274502 239037 274802 239038
rect 294540 239037 294840 239038
rect -1938 237538 -1638 237539
rect 2702 237538 3002 237539
rect 20702 237538 21002 237539
rect 38702 237538 39002 237539
rect 56702 237538 57002 237539
rect 74702 237538 75002 237539
rect 92702 237538 93002 237539
rect 110702 237538 111002 237539
rect 128702 237538 129002 237539
rect 146702 237538 147002 237539
rect 164702 237538 165002 237539
rect 182702 237538 183002 237539
rect 200702 237538 201002 237539
rect 218702 237538 219002 237539
rect 236702 237538 237002 237539
rect 254702 237538 255002 237539
rect 272702 237538 273002 237539
rect 290702 237538 291002 237539
rect 293600 237538 293900 237539
rect -2408 237527 294370 237538
rect -2408 237409 -1847 237527
rect -1729 237409 2793 237527
rect 2911 237409 20793 237527
rect 20911 237409 38793 237527
rect 38911 237409 56793 237527
rect 56911 237409 74793 237527
rect 74911 237409 92793 237527
rect 92911 237409 110793 237527
rect 110911 237409 128793 237527
rect 128911 237409 146793 237527
rect 146911 237409 164793 237527
rect 164911 237409 182793 237527
rect 182911 237409 200793 237527
rect 200911 237409 218793 237527
rect 218911 237409 236793 237527
rect 236911 237409 254793 237527
rect 254911 237409 272793 237527
rect 272911 237409 290793 237527
rect 290911 237409 293691 237527
rect 293809 237409 294370 237527
rect -2408 237367 294370 237409
rect -2408 237249 -1847 237367
rect -1729 237249 2793 237367
rect 2911 237249 20793 237367
rect 20911 237249 38793 237367
rect 38911 237249 56793 237367
rect 56911 237249 74793 237367
rect 74911 237249 92793 237367
rect 92911 237249 110793 237367
rect 110911 237249 128793 237367
rect 128911 237249 146793 237367
rect 146911 237249 164793 237367
rect 164911 237249 182793 237367
rect 182911 237249 200793 237367
rect 200911 237249 218793 237367
rect 218911 237249 236793 237367
rect 236911 237249 254793 237367
rect 254911 237249 272793 237367
rect 272911 237249 290793 237367
rect 290911 237249 293691 237367
rect 293809 237249 294370 237367
rect -2408 237238 294370 237249
rect -1938 237237 -1638 237238
rect 2702 237237 3002 237238
rect 20702 237237 21002 237238
rect 38702 237237 39002 237238
rect 56702 237237 57002 237238
rect 74702 237237 75002 237238
rect 92702 237237 93002 237238
rect 110702 237237 111002 237238
rect 128702 237237 129002 237238
rect 146702 237237 147002 237238
rect 164702 237237 165002 237238
rect 182702 237237 183002 237238
rect 200702 237237 201002 237238
rect 218702 237237 219002 237238
rect 236702 237237 237002 237238
rect 254702 237237 255002 237238
rect 272702 237237 273002 237238
rect 290702 237237 291002 237238
rect 293600 237237 293900 237238
rect -998 235738 -698 235739
rect 902 235738 1202 235739
rect 18902 235738 19202 235739
rect 36902 235738 37202 235739
rect 54902 235738 55202 235739
rect 72902 235738 73202 235739
rect 90902 235738 91202 235739
rect 108902 235738 109202 235739
rect 126902 235738 127202 235739
rect 144902 235738 145202 235739
rect 162902 235738 163202 235739
rect 180902 235738 181202 235739
rect 198902 235738 199202 235739
rect 216902 235738 217202 235739
rect 234902 235738 235202 235739
rect 252902 235738 253202 235739
rect 270902 235738 271202 235739
rect 288902 235738 289202 235739
rect 292660 235738 292960 235739
rect -1468 235727 293430 235738
rect -1468 235609 -907 235727
rect -789 235609 993 235727
rect 1111 235609 18993 235727
rect 19111 235609 36993 235727
rect 37111 235609 54993 235727
rect 55111 235609 72993 235727
rect 73111 235609 90993 235727
rect 91111 235609 108993 235727
rect 109111 235609 126993 235727
rect 127111 235609 144993 235727
rect 145111 235609 162993 235727
rect 163111 235609 180993 235727
rect 181111 235609 198993 235727
rect 199111 235609 216993 235727
rect 217111 235609 234993 235727
rect 235111 235609 252993 235727
rect 253111 235609 270993 235727
rect 271111 235609 288993 235727
rect 289111 235609 292751 235727
rect 292869 235609 293430 235727
rect -1468 235567 293430 235609
rect -1468 235449 -907 235567
rect -789 235449 993 235567
rect 1111 235449 18993 235567
rect 19111 235449 36993 235567
rect 37111 235449 54993 235567
rect 55111 235449 72993 235567
rect 73111 235449 90993 235567
rect 91111 235449 108993 235567
rect 109111 235449 126993 235567
rect 127111 235449 144993 235567
rect 145111 235449 162993 235567
rect 163111 235449 180993 235567
rect 181111 235449 198993 235567
rect 199111 235449 216993 235567
rect 217111 235449 234993 235567
rect 235111 235449 252993 235567
rect 253111 235449 270993 235567
rect 271111 235449 288993 235567
rect 289111 235449 292751 235567
rect 292869 235449 293430 235567
rect -1468 235438 293430 235449
rect -998 235437 -698 235438
rect 902 235437 1202 235438
rect 18902 235437 19202 235438
rect 36902 235437 37202 235438
rect 54902 235437 55202 235438
rect 72902 235437 73202 235438
rect 90902 235437 91202 235438
rect 108902 235437 109202 235438
rect 126902 235437 127202 235438
rect 144902 235437 145202 235438
rect 162902 235437 163202 235438
rect 180902 235437 181202 235438
rect 198902 235437 199202 235438
rect 216902 235437 217202 235438
rect 234902 235437 235202 235438
rect 252902 235437 253202 235438
rect 270902 235437 271202 235438
rect 288902 235437 289202 235438
rect 292660 235437 292960 235438
rect -4288 232138 -3988 232139
rect 15302 232138 15602 232139
rect 33302 232138 33602 232139
rect 51302 232138 51602 232139
rect 69302 232138 69602 232139
rect 87302 232138 87602 232139
rect 105302 232138 105602 232139
rect 123302 232138 123602 232139
rect 141302 232138 141602 232139
rect 159302 232138 159602 232139
rect 177302 232138 177602 232139
rect 195302 232138 195602 232139
rect 213302 232138 213602 232139
rect 231302 232138 231602 232139
rect 249302 232138 249602 232139
rect 267302 232138 267602 232139
rect 285302 232138 285602 232139
rect 295950 232138 296250 232139
rect -4288 232127 296250 232138
rect -4288 232009 -4197 232127
rect -4079 232009 15393 232127
rect 15511 232009 33393 232127
rect 33511 232009 51393 232127
rect 51511 232009 69393 232127
rect 69511 232009 87393 232127
rect 87511 232009 105393 232127
rect 105511 232009 123393 232127
rect 123511 232009 141393 232127
rect 141511 232009 159393 232127
rect 159511 232009 177393 232127
rect 177511 232009 195393 232127
rect 195511 232009 213393 232127
rect 213511 232009 231393 232127
rect 231511 232009 249393 232127
rect 249511 232009 267393 232127
rect 267511 232009 285393 232127
rect 285511 232009 296041 232127
rect 296159 232009 296250 232127
rect -4288 231967 296250 232009
rect -4288 231849 -4197 231967
rect -4079 231849 15393 231967
rect 15511 231849 33393 231967
rect 33511 231849 51393 231967
rect 51511 231849 69393 231967
rect 69511 231849 87393 231967
rect 87511 231849 105393 231967
rect 105511 231849 123393 231967
rect 123511 231849 141393 231967
rect 141511 231849 159393 231967
rect 159511 231849 177393 231967
rect 177511 231849 195393 231967
rect 195511 231849 213393 231967
rect 213511 231849 231393 231967
rect 231511 231849 249393 231967
rect 249511 231849 267393 231967
rect 267511 231849 285393 231967
rect 285511 231849 296041 231967
rect 296159 231849 296250 231967
rect -4288 231838 296250 231849
rect -4288 231837 -3988 231838
rect 15302 231837 15602 231838
rect 33302 231837 33602 231838
rect 51302 231837 51602 231838
rect 69302 231837 69602 231838
rect 87302 231837 87602 231838
rect 105302 231837 105602 231838
rect 123302 231837 123602 231838
rect 141302 231837 141602 231838
rect 159302 231837 159602 231838
rect 177302 231837 177602 231838
rect 195302 231837 195602 231838
rect 213302 231837 213602 231838
rect 231302 231837 231602 231838
rect 249302 231837 249602 231838
rect 267302 231837 267602 231838
rect 285302 231837 285602 231838
rect 295950 231837 296250 231838
rect -3348 230338 -3048 230339
rect 13502 230338 13802 230339
rect 31502 230338 31802 230339
rect 49502 230338 49802 230339
rect 67502 230338 67802 230339
rect 85502 230338 85802 230339
rect 103502 230338 103802 230339
rect 121502 230338 121802 230339
rect 139502 230338 139802 230339
rect 157502 230338 157802 230339
rect 175502 230338 175802 230339
rect 193502 230338 193802 230339
rect 211502 230338 211802 230339
rect 229502 230338 229802 230339
rect 247502 230338 247802 230339
rect 265502 230338 265802 230339
rect 283502 230338 283802 230339
rect 295010 230338 295310 230339
rect -3348 230327 295310 230338
rect -3348 230209 -3257 230327
rect -3139 230209 13593 230327
rect 13711 230209 31593 230327
rect 31711 230209 49593 230327
rect 49711 230209 67593 230327
rect 67711 230209 85593 230327
rect 85711 230209 103593 230327
rect 103711 230209 121593 230327
rect 121711 230209 139593 230327
rect 139711 230209 157593 230327
rect 157711 230209 175593 230327
rect 175711 230209 193593 230327
rect 193711 230209 211593 230327
rect 211711 230209 229593 230327
rect 229711 230209 247593 230327
rect 247711 230209 265593 230327
rect 265711 230209 283593 230327
rect 283711 230209 295101 230327
rect 295219 230209 295310 230327
rect -3348 230167 295310 230209
rect -3348 230049 -3257 230167
rect -3139 230049 13593 230167
rect 13711 230049 31593 230167
rect 31711 230049 49593 230167
rect 49711 230049 67593 230167
rect 67711 230049 85593 230167
rect 85711 230049 103593 230167
rect 103711 230049 121593 230167
rect 121711 230049 139593 230167
rect 139711 230049 157593 230167
rect 157711 230049 175593 230167
rect 175711 230049 193593 230167
rect 193711 230049 211593 230167
rect 211711 230049 229593 230167
rect 229711 230049 247593 230167
rect 247711 230049 265593 230167
rect 265711 230049 283593 230167
rect 283711 230049 295101 230167
rect 295219 230049 295310 230167
rect -3348 230038 295310 230049
rect -3348 230037 -3048 230038
rect 13502 230037 13802 230038
rect 31502 230037 31802 230038
rect 49502 230037 49802 230038
rect 67502 230037 67802 230038
rect 85502 230037 85802 230038
rect 103502 230037 103802 230038
rect 121502 230037 121802 230038
rect 139502 230037 139802 230038
rect 157502 230037 157802 230038
rect 175502 230037 175802 230038
rect 193502 230037 193802 230038
rect 211502 230037 211802 230038
rect 229502 230037 229802 230038
rect 247502 230037 247802 230038
rect 265502 230037 265802 230038
rect 283502 230037 283802 230038
rect 295010 230037 295310 230038
rect -2408 228538 -2108 228539
rect 11702 228538 12002 228539
rect 29702 228538 30002 228539
rect 47702 228538 48002 228539
rect 65702 228538 66002 228539
rect 83702 228538 84002 228539
rect 101702 228538 102002 228539
rect 119702 228538 120002 228539
rect 137702 228538 138002 228539
rect 155702 228538 156002 228539
rect 173702 228538 174002 228539
rect 191702 228538 192002 228539
rect 209702 228538 210002 228539
rect 227702 228538 228002 228539
rect 245702 228538 246002 228539
rect 263702 228538 264002 228539
rect 281702 228538 282002 228539
rect 294070 228538 294370 228539
rect -2408 228527 294370 228538
rect -2408 228409 -2317 228527
rect -2199 228409 11793 228527
rect 11911 228409 29793 228527
rect 29911 228409 47793 228527
rect 47911 228409 65793 228527
rect 65911 228409 83793 228527
rect 83911 228409 101793 228527
rect 101911 228409 119793 228527
rect 119911 228409 137793 228527
rect 137911 228409 155793 228527
rect 155911 228409 173793 228527
rect 173911 228409 191793 228527
rect 191911 228409 209793 228527
rect 209911 228409 227793 228527
rect 227911 228409 245793 228527
rect 245911 228409 263793 228527
rect 263911 228409 281793 228527
rect 281911 228409 294161 228527
rect 294279 228409 294370 228527
rect -2408 228367 294370 228409
rect -2408 228249 -2317 228367
rect -2199 228249 11793 228367
rect 11911 228249 29793 228367
rect 29911 228249 47793 228367
rect 47911 228249 65793 228367
rect 65911 228249 83793 228367
rect 83911 228249 101793 228367
rect 101911 228249 119793 228367
rect 119911 228249 137793 228367
rect 137911 228249 155793 228367
rect 155911 228249 173793 228367
rect 173911 228249 191793 228367
rect 191911 228249 209793 228367
rect 209911 228249 227793 228367
rect 227911 228249 245793 228367
rect 245911 228249 263793 228367
rect 263911 228249 281793 228367
rect 281911 228249 294161 228367
rect 294279 228249 294370 228367
rect -2408 228238 294370 228249
rect -2408 228237 -2108 228238
rect 11702 228237 12002 228238
rect 29702 228237 30002 228238
rect 47702 228237 48002 228238
rect 65702 228237 66002 228238
rect 83702 228237 84002 228238
rect 101702 228237 102002 228238
rect 119702 228237 120002 228238
rect 137702 228237 138002 228238
rect 155702 228237 156002 228238
rect 173702 228237 174002 228238
rect 191702 228237 192002 228238
rect 209702 228237 210002 228238
rect 227702 228237 228002 228238
rect 245702 228237 246002 228238
rect 263702 228237 264002 228238
rect 281702 228237 282002 228238
rect 294070 228237 294370 228238
rect -1468 226738 -1168 226739
rect 9902 226738 10202 226739
rect 27902 226738 28202 226739
rect 45902 226738 46202 226739
rect 63902 226738 64202 226739
rect 81902 226738 82202 226739
rect 99902 226738 100202 226739
rect 117902 226738 118202 226739
rect 135902 226738 136202 226739
rect 153902 226738 154202 226739
rect 171902 226738 172202 226739
rect 189902 226738 190202 226739
rect 207902 226738 208202 226739
rect 225902 226738 226202 226739
rect 243902 226738 244202 226739
rect 261902 226738 262202 226739
rect 279902 226738 280202 226739
rect 293130 226738 293430 226739
rect -1468 226727 293430 226738
rect -1468 226609 -1377 226727
rect -1259 226609 9993 226727
rect 10111 226609 27993 226727
rect 28111 226609 45993 226727
rect 46111 226609 63993 226727
rect 64111 226609 81993 226727
rect 82111 226609 99993 226727
rect 100111 226609 117993 226727
rect 118111 226609 135993 226727
rect 136111 226609 153993 226727
rect 154111 226609 171993 226727
rect 172111 226609 189993 226727
rect 190111 226609 207993 226727
rect 208111 226609 225993 226727
rect 226111 226609 243993 226727
rect 244111 226609 261993 226727
rect 262111 226609 279993 226727
rect 280111 226609 293221 226727
rect 293339 226609 293430 226727
rect -1468 226567 293430 226609
rect -1468 226449 -1377 226567
rect -1259 226449 9993 226567
rect 10111 226449 27993 226567
rect 28111 226449 45993 226567
rect 46111 226449 63993 226567
rect 64111 226449 81993 226567
rect 82111 226449 99993 226567
rect 100111 226449 117993 226567
rect 118111 226449 135993 226567
rect 136111 226449 153993 226567
rect 154111 226449 171993 226567
rect 172111 226449 189993 226567
rect 190111 226449 207993 226567
rect 208111 226449 225993 226567
rect 226111 226449 243993 226567
rect 244111 226449 261993 226567
rect 262111 226449 279993 226567
rect 280111 226449 293221 226567
rect 293339 226449 293430 226567
rect -1468 226438 293430 226449
rect -1468 226437 -1168 226438
rect 9902 226437 10202 226438
rect 27902 226437 28202 226438
rect 45902 226437 46202 226438
rect 63902 226437 64202 226438
rect 81902 226437 82202 226438
rect 99902 226437 100202 226438
rect 117902 226437 118202 226438
rect 135902 226437 136202 226438
rect 153902 226437 154202 226438
rect 171902 226437 172202 226438
rect 189902 226437 190202 226438
rect 207902 226437 208202 226438
rect 225902 226437 226202 226438
rect 243902 226437 244202 226438
rect 261902 226437 262202 226438
rect 279902 226437 280202 226438
rect 293130 226437 293430 226438
rect -3818 223138 -3518 223139
rect 6302 223138 6602 223139
rect 24302 223138 24602 223139
rect 42302 223138 42602 223139
rect 60302 223138 60602 223139
rect 78302 223138 78602 223139
rect 96302 223138 96602 223139
rect 114302 223138 114602 223139
rect 132302 223138 132602 223139
rect 150302 223138 150602 223139
rect 168302 223138 168602 223139
rect 186302 223138 186602 223139
rect 204302 223138 204602 223139
rect 222302 223138 222602 223139
rect 240302 223138 240602 223139
rect 258302 223138 258602 223139
rect 276302 223138 276602 223139
rect 295480 223138 295780 223139
rect -4288 223127 296250 223138
rect -4288 223009 -3727 223127
rect -3609 223009 6393 223127
rect 6511 223009 24393 223127
rect 24511 223009 42393 223127
rect 42511 223009 60393 223127
rect 60511 223009 78393 223127
rect 78511 223009 96393 223127
rect 96511 223009 114393 223127
rect 114511 223009 132393 223127
rect 132511 223009 150393 223127
rect 150511 223009 168393 223127
rect 168511 223009 186393 223127
rect 186511 223009 204393 223127
rect 204511 223009 222393 223127
rect 222511 223009 240393 223127
rect 240511 223009 258393 223127
rect 258511 223009 276393 223127
rect 276511 223009 295571 223127
rect 295689 223009 296250 223127
rect -4288 222967 296250 223009
rect -4288 222849 -3727 222967
rect -3609 222849 6393 222967
rect 6511 222849 24393 222967
rect 24511 222849 42393 222967
rect 42511 222849 60393 222967
rect 60511 222849 78393 222967
rect 78511 222849 96393 222967
rect 96511 222849 114393 222967
rect 114511 222849 132393 222967
rect 132511 222849 150393 222967
rect 150511 222849 168393 222967
rect 168511 222849 186393 222967
rect 186511 222849 204393 222967
rect 204511 222849 222393 222967
rect 222511 222849 240393 222967
rect 240511 222849 258393 222967
rect 258511 222849 276393 222967
rect 276511 222849 295571 222967
rect 295689 222849 296250 222967
rect -4288 222838 296250 222849
rect -3818 222837 -3518 222838
rect 6302 222837 6602 222838
rect 24302 222837 24602 222838
rect 42302 222837 42602 222838
rect 60302 222837 60602 222838
rect 78302 222837 78602 222838
rect 96302 222837 96602 222838
rect 114302 222837 114602 222838
rect 132302 222837 132602 222838
rect 150302 222837 150602 222838
rect 168302 222837 168602 222838
rect 186302 222837 186602 222838
rect 204302 222837 204602 222838
rect 222302 222837 222602 222838
rect 240302 222837 240602 222838
rect 258302 222837 258602 222838
rect 276302 222837 276602 222838
rect 295480 222837 295780 222838
rect -2878 221338 -2578 221339
rect 4502 221338 4802 221339
rect 22502 221338 22802 221339
rect 40502 221338 40802 221339
rect 58502 221338 58802 221339
rect 76502 221338 76802 221339
rect 94502 221338 94802 221339
rect 112502 221338 112802 221339
rect 130502 221338 130802 221339
rect 148502 221338 148802 221339
rect 166502 221338 166802 221339
rect 184502 221338 184802 221339
rect 202502 221338 202802 221339
rect 220502 221338 220802 221339
rect 238502 221338 238802 221339
rect 256502 221338 256802 221339
rect 274502 221338 274802 221339
rect 294540 221338 294840 221339
rect -3348 221327 295310 221338
rect -3348 221209 -2787 221327
rect -2669 221209 4593 221327
rect 4711 221209 22593 221327
rect 22711 221209 40593 221327
rect 40711 221209 58593 221327
rect 58711 221209 76593 221327
rect 76711 221209 94593 221327
rect 94711 221209 112593 221327
rect 112711 221209 130593 221327
rect 130711 221209 148593 221327
rect 148711 221209 166593 221327
rect 166711 221209 184593 221327
rect 184711 221209 202593 221327
rect 202711 221209 220593 221327
rect 220711 221209 238593 221327
rect 238711 221209 256593 221327
rect 256711 221209 274593 221327
rect 274711 221209 294631 221327
rect 294749 221209 295310 221327
rect -3348 221167 295310 221209
rect -3348 221049 -2787 221167
rect -2669 221049 4593 221167
rect 4711 221049 22593 221167
rect 22711 221049 40593 221167
rect 40711 221049 58593 221167
rect 58711 221049 76593 221167
rect 76711 221049 94593 221167
rect 94711 221049 112593 221167
rect 112711 221049 130593 221167
rect 130711 221049 148593 221167
rect 148711 221049 166593 221167
rect 166711 221049 184593 221167
rect 184711 221049 202593 221167
rect 202711 221049 220593 221167
rect 220711 221049 238593 221167
rect 238711 221049 256593 221167
rect 256711 221049 274593 221167
rect 274711 221049 294631 221167
rect 294749 221049 295310 221167
rect -3348 221038 295310 221049
rect -2878 221037 -2578 221038
rect 4502 221037 4802 221038
rect 22502 221037 22802 221038
rect 40502 221037 40802 221038
rect 58502 221037 58802 221038
rect 76502 221037 76802 221038
rect 94502 221037 94802 221038
rect 112502 221037 112802 221038
rect 130502 221037 130802 221038
rect 148502 221037 148802 221038
rect 166502 221037 166802 221038
rect 184502 221037 184802 221038
rect 202502 221037 202802 221038
rect 220502 221037 220802 221038
rect 238502 221037 238802 221038
rect 256502 221037 256802 221038
rect 274502 221037 274802 221038
rect 294540 221037 294840 221038
rect -1938 219538 -1638 219539
rect 2702 219538 3002 219539
rect 20702 219538 21002 219539
rect 38702 219538 39002 219539
rect 56702 219538 57002 219539
rect 74702 219538 75002 219539
rect 92702 219538 93002 219539
rect 110702 219538 111002 219539
rect 128702 219538 129002 219539
rect 146702 219538 147002 219539
rect 164702 219538 165002 219539
rect 182702 219538 183002 219539
rect 200702 219538 201002 219539
rect 218702 219538 219002 219539
rect 236702 219538 237002 219539
rect 254702 219538 255002 219539
rect 272702 219538 273002 219539
rect 290702 219538 291002 219539
rect 293600 219538 293900 219539
rect -2408 219527 294370 219538
rect -2408 219409 -1847 219527
rect -1729 219409 2793 219527
rect 2911 219409 20793 219527
rect 20911 219409 38793 219527
rect 38911 219409 56793 219527
rect 56911 219409 74793 219527
rect 74911 219409 92793 219527
rect 92911 219409 110793 219527
rect 110911 219409 128793 219527
rect 128911 219409 146793 219527
rect 146911 219409 164793 219527
rect 164911 219409 182793 219527
rect 182911 219409 200793 219527
rect 200911 219409 218793 219527
rect 218911 219409 236793 219527
rect 236911 219409 254793 219527
rect 254911 219409 272793 219527
rect 272911 219409 290793 219527
rect 290911 219409 293691 219527
rect 293809 219409 294370 219527
rect -2408 219367 294370 219409
rect -2408 219249 -1847 219367
rect -1729 219249 2793 219367
rect 2911 219249 20793 219367
rect 20911 219249 38793 219367
rect 38911 219249 56793 219367
rect 56911 219249 74793 219367
rect 74911 219249 92793 219367
rect 92911 219249 110793 219367
rect 110911 219249 128793 219367
rect 128911 219249 146793 219367
rect 146911 219249 164793 219367
rect 164911 219249 182793 219367
rect 182911 219249 200793 219367
rect 200911 219249 218793 219367
rect 218911 219249 236793 219367
rect 236911 219249 254793 219367
rect 254911 219249 272793 219367
rect 272911 219249 290793 219367
rect 290911 219249 293691 219367
rect 293809 219249 294370 219367
rect -2408 219238 294370 219249
rect -1938 219237 -1638 219238
rect 2702 219237 3002 219238
rect 20702 219237 21002 219238
rect 38702 219237 39002 219238
rect 56702 219237 57002 219238
rect 74702 219237 75002 219238
rect 92702 219237 93002 219238
rect 110702 219237 111002 219238
rect 128702 219237 129002 219238
rect 146702 219237 147002 219238
rect 164702 219237 165002 219238
rect 182702 219237 183002 219238
rect 200702 219237 201002 219238
rect 218702 219237 219002 219238
rect 236702 219237 237002 219238
rect 254702 219237 255002 219238
rect 272702 219237 273002 219238
rect 290702 219237 291002 219238
rect 293600 219237 293900 219238
rect -998 217738 -698 217739
rect 902 217738 1202 217739
rect 18902 217738 19202 217739
rect 36902 217738 37202 217739
rect 54902 217738 55202 217739
rect 72902 217738 73202 217739
rect 90902 217738 91202 217739
rect 108902 217738 109202 217739
rect 126902 217738 127202 217739
rect 144902 217738 145202 217739
rect 162902 217738 163202 217739
rect 180902 217738 181202 217739
rect 198902 217738 199202 217739
rect 216902 217738 217202 217739
rect 234902 217738 235202 217739
rect 252902 217738 253202 217739
rect 270902 217738 271202 217739
rect 288902 217738 289202 217739
rect 292660 217738 292960 217739
rect -1468 217727 293430 217738
rect -1468 217609 -907 217727
rect -789 217609 993 217727
rect 1111 217609 18993 217727
rect 19111 217609 36993 217727
rect 37111 217609 54993 217727
rect 55111 217609 72993 217727
rect 73111 217609 90993 217727
rect 91111 217609 108993 217727
rect 109111 217609 126993 217727
rect 127111 217609 144993 217727
rect 145111 217609 162993 217727
rect 163111 217609 180993 217727
rect 181111 217609 198993 217727
rect 199111 217609 216993 217727
rect 217111 217609 234993 217727
rect 235111 217609 252993 217727
rect 253111 217609 270993 217727
rect 271111 217609 288993 217727
rect 289111 217609 292751 217727
rect 292869 217609 293430 217727
rect -1468 217567 293430 217609
rect -1468 217449 -907 217567
rect -789 217449 993 217567
rect 1111 217449 18993 217567
rect 19111 217449 36993 217567
rect 37111 217449 54993 217567
rect 55111 217449 72993 217567
rect 73111 217449 90993 217567
rect 91111 217449 108993 217567
rect 109111 217449 126993 217567
rect 127111 217449 144993 217567
rect 145111 217449 162993 217567
rect 163111 217449 180993 217567
rect 181111 217449 198993 217567
rect 199111 217449 216993 217567
rect 217111 217449 234993 217567
rect 235111 217449 252993 217567
rect 253111 217449 270993 217567
rect 271111 217449 288993 217567
rect 289111 217449 292751 217567
rect 292869 217449 293430 217567
rect -1468 217438 293430 217449
rect -998 217437 -698 217438
rect 902 217437 1202 217438
rect 18902 217437 19202 217438
rect 36902 217437 37202 217438
rect 54902 217437 55202 217438
rect 72902 217437 73202 217438
rect 90902 217437 91202 217438
rect 108902 217437 109202 217438
rect 126902 217437 127202 217438
rect 144902 217437 145202 217438
rect 162902 217437 163202 217438
rect 180902 217437 181202 217438
rect 198902 217437 199202 217438
rect 216902 217437 217202 217438
rect 234902 217437 235202 217438
rect 252902 217437 253202 217438
rect 270902 217437 271202 217438
rect 288902 217437 289202 217438
rect 292660 217437 292960 217438
rect -4288 214138 -3988 214139
rect 15302 214138 15602 214139
rect 33302 214138 33602 214139
rect 51302 214138 51602 214139
rect 69302 214138 69602 214139
rect 87302 214138 87602 214139
rect 105302 214138 105602 214139
rect 123302 214138 123602 214139
rect 141302 214138 141602 214139
rect 159302 214138 159602 214139
rect 177302 214138 177602 214139
rect 195302 214138 195602 214139
rect 213302 214138 213602 214139
rect 231302 214138 231602 214139
rect 249302 214138 249602 214139
rect 267302 214138 267602 214139
rect 285302 214138 285602 214139
rect 295950 214138 296250 214139
rect -4288 214127 296250 214138
rect -4288 214009 -4197 214127
rect -4079 214009 15393 214127
rect 15511 214009 33393 214127
rect 33511 214009 51393 214127
rect 51511 214009 69393 214127
rect 69511 214009 87393 214127
rect 87511 214009 105393 214127
rect 105511 214009 123393 214127
rect 123511 214009 141393 214127
rect 141511 214009 159393 214127
rect 159511 214009 177393 214127
rect 177511 214009 195393 214127
rect 195511 214009 213393 214127
rect 213511 214009 231393 214127
rect 231511 214009 249393 214127
rect 249511 214009 267393 214127
rect 267511 214009 285393 214127
rect 285511 214009 296041 214127
rect 296159 214009 296250 214127
rect -4288 213967 296250 214009
rect -4288 213849 -4197 213967
rect -4079 213849 15393 213967
rect 15511 213849 33393 213967
rect 33511 213849 51393 213967
rect 51511 213849 69393 213967
rect 69511 213849 87393 213967
rect 87511 213849 105393 213967
rect 105511 213849 123393 213967
rect 123511 213849 141393 213967
rect 141511 213849 159393 213967
rect 159511 213849 177393 213967
rect 177511 213849 195393 213967
rect 195511 213849 213393 213967
rect 213511 213849 231393 213967
rect 231511 213849 249393 213967
rect 249511 213849 267393 213967
rect 267511 213849 285393 213967
rect 285511 213849 296041 213967
rect 296159 213849 296250 213967
rect -4288 213838 296250 213849
rect -4288 213837 -3988 213838
rect 15302 213837 15602 213838
rect 33302 213837 33602 213838
rect 51302 213837 51602 213838
rect 69302 213837 69602 213838
rect 87302 213837 87602 213838
rect 105302 213837 105602 213838
rect 123302 213837 123602 213838
rect 141302 213837 141602 213838
rect 159302 213837 159602 213838
rect 177302 213837 177602 213838
rect 195302 213837 195602 213838
rect 213302 213837 213602 213838
rect 231302 213837 231602 213838
rect 249302 213837 249602 213838
rect 267302 213837 267602 213838
rect 285302 213837 285602 213838
rect 295950 213837 296250 213838
rect -3348 212338 -3048 212339
rect 13502 212338 13802 212339
rect 31502 212338 31802 212339
rect 49502 212338 49802 212339
rect 67502 212338 67802 212339
rect 85502 212338 85802 212339
rect 103502 212338 103802 212339
rect 121502 212338 121802 212339
rect 139502 212338 139802 212339
rect 157502 212338 157802 212339
rect 175502 212338 175802 212339
rect 193502 212338 193802 212339
rect 211502 212338 211802 212339
rect 229502 212338 229802 212339
rect 247502 212338 247802 212339
rect 265502 212338 265802 212339
rect 283502 212338 283802 212339
rect 295010 212338 295310 212339
rect -3348 212327 295310 212338
rect -3348 212209 -3257 212327
rect -3139 212209 13593 212327
rect 13711 212209 31593 212327
rect 31711 212209 49593 212327
rect 49711 212209 67593 212327
rect 67711 212209 85593 212327
rect 85711 212209 103593 212327
rect 103711 212209 121593 212327
rect 121711 212209 139593 212327
rect 139711 212209 157593 212327
rect 157711 212209 175593 212327
rect 175711 212209 193593 212327
rect 193711 212209 211593 212327
rect 211711 212209 229593 212327
rect 229711 212209 247593 212327
rect 247711 212209 265593 212327
rect 265711 212209 283593 212327
rect 283711 212209 295101 212327
rect 295219 212209 295310 212327
rect -3348 212167 295310 212209
rect -3348 212049 -3257 212167
rect -3139 212049 13593 212167
rect 13711 212049 31593 212167
rect 31711 212049 49593 212167
rect 49711 212049 67593 212167
rect 67711 212049 85593 212167
rect 85711 212049 103593 212167
rect 103711 212049 121593 212167
rect 121711 212049 139593 212167
rect 139711 212049 157593 212167
rect 157711 212049 175593 212167
rect 175711 212049 193593 212167
rect 193711 212049 211593 212167
rect 211711 212049 229593 212167
rect 229711 212049 247593 212167
rect 247711 212049 265593 212167
rect 265711 212049 283593 212167
rect 283711 212049 295101 212167
rect 295219 212049 295310 212167
rect -3348 212038 295310 212049
rect -3348 212037 -3048 212038
rect 13502 212037 13802 212038
rect 31502 212037 31802 212038
rect 49502 212037 49802 212038
rect 67502 212037 67802 212038
rect 85502 212037 85802 212038
rect 103502 212037 103802 212038
rect 121502 212037 121802 212038
rect 139502 212037 139802 212038
rect 157502 212037 157802 212038
rect 175502 212037 175802 212038
rect 193502 212037 193802 212038
rect 211502 212037 211802 212038
rect 229502 212037 229802 212038
rect 247502 212037 247802 212038
rect 265502 212037 265802 212038
rect 283502 212037 283802 212038
rect 295010 212037 295310 212038
rect -2408 210538 -2108 210539
rect 11702 210538 12002 210539
rect 29702 210538 30002 210539
rect 47702 210538 48002 210539
rect 65702 210538 66002 210539
rect 83702 210538 84002 210539
rect 101702 210538 102002 210539
rect 119702 210538 120002 210539
rect 137702 210538 138002 210539
rect 155702 210538 156002 210539
rect 173702 210538 174002 210539
rect 191702 210538 192002 210539
rect 209702 210538 210002 210539
rect 227702 210538 228002 210539
rect 245702 210538 246002 210539
rect 263702 210538 264002 210539
rect 281702 210538 282002 210539
rect 294070 210538 294370 210539
rect -2408 210527 294370 210538
rect -2408 210409 -2317 210527
rect -2199 210409 11793 210527
rect 11911 210409 29793 210527
rect 29911 210409 47793 210527
rect 47911 210409 65793 210527
rect 65911 210409 83793 210527
rect 83911 210409 101793 210527
rect 101911 210409 119793 210527
rect 119911 210409 137793 210527
rect 137911 210409 155793 210527
rect 155911 210409 173793 210527
rect 173911 210409 191793 210527
rect 191911 210409 209793 210527
rect 209911 210409 227793 210527
rect 227911 210409 245793 210527
rect 245911 210409 263793 210527
rect 263911 210409 281793 210527
rect 281911 210409 294161 210527
rect 294279 210409 294370 210527
rect -2408 210367 294370 210409
rect -2408 210249 -2317 210367
rect -2199 210249 11793 210367
rect 11911 210249 29793 210367
rect 29911 210249 47793 210367
rect 47911 210249 65793 210367
rect 65911 210249 83793 210367
rect 83911 210249 101793 210367
rect 101911 210249 119793 210367
rect 119911 210249 137793 210367
rect 137911 210249 155793 210367
rect 155911 210249 173793 210367
rect 173911 210249 191793 210367
rect 191911 210249 209793 210367
rect 209911 210249 227793 210367
rect 227911 210249 245793 210367
rect 245911 210249 263793 210367
rect 263911 210249 281793 210367
rect 281911 210249 294161 210367
rect 294279 210249 294370 210367
rect -2408 210238 294370 210249
rect -2408 210237 -2108 210238
rect 11702 210237 12002 210238
rect 29702 210237 30002 210238
rect 47702 210237 48002 210238
rect 65702 210237 66002 210238
rect 83702 210237 84002 210238
rect 101702 210237 102002 210238
rect 119702 210237 120002 210238
rect 137702 210237 138002 210238
rect 155702 210237 156002 210238
rect 173702 210237 174002 210238
rect 191702 210237 192002 210238
rect 209702 210237 210002 210238
rect 227702 210237 228002 210238
rect 245702 210237 246002 210238
rect 263702 210237 264002 210238
rect 281702 210237 282002 210238
rect 294070 210237 294370 210238
rect -1468 208738 -1168 208739
rect 9902 208738 10202 208739
rect 27902 208738 28202 208739
rect 45902 208738 46202 208739
rect 63902 208738 64202 208739
rect 81902 208738 82202 208739
rect 99902 208738 100202 208739
rect 117902 208738 118202 208739
rect 135902 208738 136202 208739
rect 153902 208738 154202 208739
rect 171902 208738 172202 208739
rect 189902 208738 190202 208739
rect 207902 208738 208202 208739
rect 225902 208738 226202 208739
rect 243902 208738 244202 208739
rect 261902 208738 262202 208739
rect 279902 208738 280202 208739
rect 293130 208738 293430 208739
rect -1468 208727 293430 208738
rect -1468 208609 -1377 208727
rect -1259 208609 9993 208727
rect 10111 208609 27993 208727
rect 28111 208609 45993 208727
rect 46111 208609 63993 208727
rect 64111 208609 81993 208727
rect 82111 208609 99993 208727
rect 100111 208609 117993 208727
rect 118111 208609 135993 208727
rect 136111 208609 153993 208727
rect 154111 208609 171993 208727
rect 172111 208609 189993 208727
rect 190111 208609 207993 208727
rect 208111 208609 225993 208727
rect 226111 208609 243993 208727
rect 244111 208609 261993 208727
rect 262111 208609 279993 208727
rect 280111 208609 293221 208727
rect 293339 208609 293430 208727
rect -1468 208567 293430 208609
rect -1468 208449 -1377 208567
rect -1259 208449 9993 208567
rect 10111 208449 27993 208567
rect 28111 208449 45993 208567
rect 46111 208449 63993 208567
rect 64111 208449 81993 208567
rect 82111 208449 99993 208567
rect 100111 208449 117993 208567
rect 118111 208449 135993 208567
rect 136111 208449 153993 208567
rect 154111 208449 171993 208567
rect 172111 208449 189993 208567
rect 190111 208449 207993 208567
rect 208111 208449 225993 208567
rect 226111 208449 243993 208567
rect 244111 208449 261993 208567
rect 262111 208449 279993 208567
rect 280111 208449 293221 208567
rect 293339 208449 293430 208567
rect -1468 208438 293430 208449
rect -1468 208437 -1168 208438
rect 9902 208437 10202 208438
rect 27902 208437 28202 208438
rect 45902 208437 46202 208438
rect 63902 208437 64202 208438
rect 81902 208437 82202 208438
rect 99902 208437 100202 208438
rect 117902 208437 118202 208438
rect 135902 208437 136202 208438
rect 153902 208437 154202 208438
rect 171902 208437 172202 208438
rect 189902 208437 190202 208438
rect 207902 208437 208202 208438
rect 225902 208437 226202 208438
rect 243902 208437 244202 208438
rect 261902 208437 262202 208438
rect 279902 208437 280202 208438
rect 293130 208437 293430 208438
rect -3818 205138 -3518 205139
rect 6302 205138 6602 205139
rect 24302 205138 24602 205139
rect 42302 205138 42602 205139
rect 60302 205138 60602 205139
rect 78302 205138 78602 205139
rect 96302 205138 96602 205139
rect 114302 205138 114602 205139
rect 132302 205138 132602 205139
rect 150302 205138 150602 205139
rect 168302 205138 168602 205139
rect 186302 205138 186602 205139
rect 204302 205138 204602 205139
rect 222302 205138 222602 205139
rect 240302 205138 240602 205139
rect 258302 205138 258602 205139
rect 276302 205138 276602 205139
rect 295480 205138 295780 205139
rect -4288 205127 296250 205138
rect -4288 205009 -3727 205127
rect -3609 205009 6393 205127
rect 6511 205009 24393 205127
rect 24511 205009 42393 205127
rect 42511 205009 60393 205127
rect 60511 205009 78393 205127
rect 78511 205009 96393 205127
rect 96511 205009 114393 205127
rect 114511 205009 132393 205127
rect 132511 205009 150393 205127
rect 150511 205009 168393 205127
rect 168511 205009 186393 205127
rect 186511 205009 204393 205127
rect 204511 205009 222393 205127
rect 222511 205009 240393 205127
rect 240511 205009 258393 205127
rect 258511 205009 276393 205127
rect 276511 205009 295571 205127
rect 295689 205009 296250 205127
rect -4288 204967 296250 205009
rect -4288 204849 -3727 204967
rect -3609 204849 6393 204967
rect 6511 204849 24393 204967
rect 24511 204849 42393 204967
rect 42511 204849 60393 204967
rect 60511 204849 78393 204967
rect 78511 204849 96393 204967
rect 96511 204849 114393 204967
rect 114511 204849 132393 204967
rect 132511 204849 150393 204967
rect 150511 204849 168393 204967
rect 168511 204849 186393 204967
rect 186511 204849 204393 204967
rect 204511 204849 222393 204967
rect 222511 204849 240393 204967
rect 240511 204849 258393 204967
rect 258511 204849 276393 204967
rect 276511 204849 295571 204967
rect 295689 204849 296250 204967
rect -4288 204838 296250 204849
rect -3818 204837 -3518 204838
rect 6302 204837 6602 204838
rect 24302 204837 24602 204838
rect 42302 204837 42602 204838
rect 60302 204837 60602 204838
rect 78302 204837 78602 204838
rect 96302 204837 96602 204838
rect 114302 204837 114602 204838
rect 132302 204837 132602 204838
rect 150302 204837 150602 204838
rect 168302 204837 168602 204838
rect 186302 204837 186602 204838
rect 204302 204837 204602 204838
rect 222302 204837 222602 204838
rect 240302 204837 240602 204838
rect 258302 204837 258602 204838
rect 276302 204837 276602 204838
rect 295480 204837 295780 204838
rect -2878 203338 -2578 203339
rect 4502 203338 4802 203339
rect 22502 203338 22802 203339
rect 40502 203338 40802 203339
rect 58502 203338 58802 203339
rect 76502 203338 76802 203339
rect 94502 203338 94802 203339
rect 112502 203338 112802 203339
rect 130502 203338 130802 203339
rect 148502 203338 148802 203339
rect 166502 203338 166802 203339
rect 184502 203338 184802 203339
rect 202502 203338 202802 203339
rect 220502 203338 220802 203339
rect 238502 203338 238802 203339
rect 256502 203338 256802 203339
rect 274502 203338 274802 203339
rect 294540 203338 294840 203339
rect -3348 203327 295310 203338
rect -3348 203209 -2787 203327
rect -2669 203209 4593 203327
rect 4711 203209 22593 203327
rect 22711 203209 40593 203327
rect 40711 203209 58593 203327
rect 58711 203209 76593 203327
rect 76711 203209 94593 203327
rect 94711 203209 112593 203327
rect 112711 203209 130593 203327
rect 130711 203209 148593 203327
rect 148711 203209 166593 203327
rect 166711 203209 184593 203327
rect 184711 203209 202593 203327
rect 202711 203209 220593 203327
rect 220711 203209 238593 203327
rect 238711 203209 256593 203327
rect 256711 203209 274593 203327
rect 274711 203209 294631 203327
rect 294749 203209 295310 203327
rect -3348 203167 295310 203209
rect -3348 203049 -2787 203167
rect -2669 203049 4593 203167
rect 4711 203049 22593 203167
rect 22711 203049 40593 203167
rect 40711 203049 58593 203167
rect 58711 203049 76593 203167
rect 76711 203049 94593 203167
rect 94711 203049 112593 203167
rect 112711 203049 130593 203167
rect 130711 203049 148593 203167
rect 148711 203049 166593 203167
rect 166711 203049 184593 203167
rect 184711 203049 202593 203167
rect 202711 203049 220593 203167
rect 220711 203049 238593 203167
rect 238711 203049 256593 203167
rect 256711 203049 274593 203167
rect 274711 203049 294631 203167
rect 294749 203049 295310 203167
rect -3348 203038 295310 203049
rect -2878 203037 -2578 203038
rect 4502 203037 4802 203038
rect 22502 203037 22802 203038
rect 40502 203037 40802 203038
rect 58502 203037 58802 203038
rect 76502 203037 76802 203038
rect 94502 203037 94802 203038
rect 112502 203037 112802 203038
rect 130502 203037 130802 203038
rect 148502 203037 148802 203038
rect 166502 203037 166802 203038
rect 184502 203037 184802 203038
rect 202502 203037 202802 203038
rect 220502 203037 220802 203038
rect 238502 203037 238802 203038
rect 256502 203037 256802 203038
rect 274502 203037 274802 203038
rect 294540 203037 294840 203038
rect -1938 201538 -1638 201539
rect 2702 201538 3002 201539
rect 20702 201538 21002 201539
rect 38702 201538 39002 201539
rect 56702 201538 57002 201539
rect 74702 201538 75002 201539
rect 92702 201538 93002 201539
rect 110702 201538 111002 201539
rect 128702 201538 129002 201539
rect 146702 201538 147002 201539
rect 164702 201538 165002 201539
rect 182702 201538 183002 201539
rect 200702 201538 201002 201539
rect 218702 201538 219002 201539
rect 236702 201538 237002 201539
rect 254702 201538 255002 201539
rect 272702 201538 273002 201539
rect 290702 201538 291002 201539
rect 293600 201538 293900 201539
rect -2408 201527 294370 201538
rect -2408 201409 -1847 201527
rect -1729 201409 2793 201527
rect 2911 201409 20793 201527
rect 20911 201409 38793 201527
rect 38911 201409 56793 201527
rect 56911 201409 74793 201527
rect 74911 201409 92793 201527
rect 92911 201409 110793 201527
rect 110911 201409 128793 201527
rect 128911 201409 146793 201527
rect 146911 201409 164793 201527
rect 164911 201409 182793 201527
rect 182911 201409 200793 201527
rect 200911 201409 218793 201527
rect 218911 201409 236793 201527
rect 236911 201409 254793 201527
rect 254911 201409 272793 201527
rect 272911 201409 290793 201527
rect 290911 201409 293691 201527
rect 293809 201409 294370 201527
rect -2408 201367 294370 201409
rect -2408 201249 -1847 201367
rect -1729 201249 2793 201367
rect 2911 201249 20793 201367
rect 20911 201249 38793 201367
rect 38911 201249 56793 201367
rect 56911 201249 74793 201367
rect 74911 201249 92793 201367
rect 92911 201249 110793 201367
rect 110911 201249 128793 201367
rect 128911 201249 146793 201367
rect 146911 201249 164793 201367
rect 164911 201249 182793 201367
rect 182911 201249 200793 201367
rect 200911 201249 218793 201367
rect 218911 201249 236793 201367
rect 236911 201249 254793 201367
rect 254911 201249 272793 201367
rect 272911 201249 290793 201367
rect 290911 201249 293691 201367
rect 293809 201249 294370 201367
rect -2408 201238 294370 201249
rect -1938 201237 -1638 201238
rect 2702 201237 3002 201238
rect 20702 201237 21002 201238
rect 38702 201237 39002 201238
rect 56702 201237 57002 201238
rect 74702 201237 75002 201238
rect 92702 201237 93002 201238
rect 110702 201237 111002 201238
rect 128702 201237 129002 201238
rect 146702 201237 147002 201238
rect 164702 201237 165002 201238
rect 182702 201237 183002 201238
rect 200702 201237 201002 201238
rect 218702 201237 219002 201238
rect 236702 201237 237002 201238
rect 254702 201237 255002 201238
rect 272702 201237 273002 201238
rect 290702 201237 291002 201238
rect 293600 201237 293900 201238
rect -998 199738 -698 199739
rect 902 199738 1202 199739
rect 18902 199738 19202 199739
rect 36902 199738 37202 199739
rect 54902 199738 55202 199739
rect 72902 199738 73202 199739
rect 90902 199738 91202 199739
rect 108902 199738 109202 199739
rect 126902 199738 127202 199739
rect 144902 199738 145202 199739
rect 162902 199738 163202 199739
rect 180902 199738 181202 199739
rect 198902 199738 199202 199739
rect 216902 199738 217202 199739
rect 234902 199738 235202 199739
rect 252902 199738 253202 199739
rect 270902 199738 271202 199739
rect 288902 199738 289202 199739
rect 292660 199738 292960 199739
rect -1468 199727 293430 199738
rect -1468 199609 -907 199727
rect -789 199609 993 199727
rect 1111 199609 18993 199727
rect 19111 199609 36993 199727
rect 37111 199609 54993 199727
rect 55111 199609 72993 199727
rect 73111 199609 90993 199727
rect 91111 199609 108993 199727
rect 109111 199609 126993 199727
rect 127111 199609 144993 199727
rect 145111 199609 162993 199727
rect 163111 199609 180993 199727
rect 181111 199609 198993 199727
rect 199111 199609 216993 199727
rect 217111 199609 234993 199727
rect 235111 199609 252993 199727
rect 253111 199609 270993 199727
rect 271111 199609 288993 199727
rect 289111 199609 292751 199727
rect 292869 199609 293430 199727
rect -1468 199567 293430 199609
rect -1468 199449 -907 199567
rect -789 199449 993 199567
rect 1111 199449 18993 199567
rect 19111 199449 36993 199567
rect 37111 199449 54993 199567
rect 55111 199449 72993 199567
rect 73111 199449 90993 199567
rect 91111 199449 108993 199567
rect 109111 199449 126993 199567
rect 127111 199449 144993 199567
rect 145111 199449 162993 199567
rect 163111 199449 180993 199567
rect 181111 199449 198993 199567
rect 199111 199449 216993 199567
rect 217111 199449 234993 199567
rect 235111 199449 252993 199567
rect 253111 199449 270993 199567
rect 271111 199449 288993 199567
rect 289111 199449 292751 199567
rect 292869 199449 293430 199567
rect -1468 199438 293430 199449
rect -998 199437 -698 199438
rect 902 199437 1202 199438
rect 18902 199437 19202 199438
rect 36902 199437 37202 199438
rect 54902 199437 55202 199438
rect 72902 199437 73202 199438
rect 90902 199437 91202 199438
rect 108902 199437 109202 199438
rect 126902 199437 127202 199438
rect 144902 199437 145202 199438
rect 162902 199437 163202 199438
rect 180902 199437 181202 199438
rect 198902 199437 199202 199438
rect 216902 199437 217202 199438
rect 234902 199437 235202 199438
rect 252902 199437 253202 199438
rect 270902 199437 271202 199438
rect 288902 199437 289202 199438
rect 292660 199437 292960 199438
rect -4288 196138 -3988 196139
rect 15302 196138 15602 196139
rect 33302 196138 33602 196139
rect 51302 196138 51602 196139
rect 69302 196138 69602 196139
rect 87302 196138 87602 196139
rect 105302 196138 105602 196139
rect 123302 196138 123602 196139
rect 141302 196138 141602 196139
rect 159302 196138 159602 196139
rect 177302 196138 177602 196139
rect 195302 196138 195602 196139
rect 213302 196138 213602 196139
rect 231302 196138 231602 196139
rect 249302 196138 249602 196139
rect 267302 196138 267602 196139
rect 285302 196138 285602 196139
rect 295950 196138 296250 196139
rect -4288 196127 296250 196138
rect -4288 196009 -4197 196127
rect -4079 196009 15393 196127
rect 15511 196009 33393 196127
rect 33511 196009 51393 196127
rect 51511 196009 69393 196127
rect 69511 196009 87393 196127
rect 87511 196009 105393 196127
rect 105511 196009 123393 196127
rect 123511 196009 141393 196127
rect 141511 196009 159393 196127
rect 159511 196009 177393 196127
rect 177511 196009 195393 196127
rect 195511 196009 213393 196127
rect 213511 196009 231393 196127
rect 231511 196009 249393 196127
rect 249511 196009 267393 196127
rect 267511 196009 285393 196127
rect 285511 196009 296041 196127
rect 296159 196009 296250 196127
rect -4288 195967 296250 196009
rect -4288 195849 -4197 195967
rect -4079 195849 15393 195967
rect 15511 195849 33393 195967
rect 33511 195849 51393 195967
rect 51511 195849 69393 195967
rect 69511 195849 87393 195967
rect 87511 195849 105393 195967
rect 105511 195849 123393 195967
rect 123511 195849 141393 195967
rect 141511 195849 159393 195967
rect 159511 195849 177393 195967
rect 177511 195849 195393 195967
rect 195511 195849 213393 195967
rect 213511 195849 231393 195967
rect 231511 195849 249393 195967
rect 249511 195849 267393 195967
rect 267511 195849 285393 195967
rect 285511 195849 296041 195967
rect 296159 195849 296250 195967
rect -4288 195838 296250 195849
rect -4288 195837 -3988 195838
rect 15302 195837 15602 195838
rect 33302 195837 33602 195838
rect 51302 195837 51602 195838
rect 69302 195837 69602 195838
rect 87302 195837 87602 195838
rect 105302 195837 105602 195838
rect 123302 195837 123602 195838
rect 141302 195837 141602 195838
rect 159302 195837 159602 195838
rect 177302 195837 177602 195838
rect 195302 195837 195602 195838
rect 213302 195837 213602 195838
rect 231302 195837 231602 195838
rect 249302 195837 249602 195838
rect 267302 195837 267602 195838
rect 285302 195837 285602 195838
rect 295950 195837 296250 195838
rect -3348 194338 -3048 194339
rect 13502 194338 13802 194339
rect 31502 194338 31802 194339
rect 49502 194338 49802 194339
rect 67502 194338 67802 194339
rect 85502 194338 85802 194339
rect 103502 194338 103802 194339
rect 121502 194338 121802 194339
rect 139502 194338 139802 194339
rect 157502 194338 157802 194339
rect 175502 194338 175802 194339
rect 193502 194338 193802 194339
rect 211502 194338 211802 194339
rect 229502 194338 229802 194339
rect 247502 194338 247802 194339
rect 265502 194338 265802 194339
rect 283502 194338 283802 194339
rect 295010 194338 295310 194339
rect -3348 194327 295310 194338
rect -3348 194209 -3257 194327
rect -3139 194209 13593 194327
rect 13711 194209 31593 194327
rect 31711 194209 49593 194327
rect 49711 194209 67593 194327
rect 67711 194209 85593 194327
rect 85711 194209 103593 194327
rect 103711 194209 121593 194327
rect 121711 194209 139593 194327
rect 139711 194209 157593 194327
rect 157711 194209 175593 194327
rect 175711 194209 193593 194327
rect 193711 194209 211593 194327
rect 211711 194209 229593 194327
rect 229711 194209 247593 194327
rect 247711 194209 265593 194327
rect 265711 194209 283593 194327
rect 283711 194209 295101 194327
rect 295219 194209 295310 194327
rect -3348 194167 295310 194209
rect -3348 194049 -3257 194167
rect -3139 194049 13593 194167
rect 13711 194049 31593 194167
rect 31711 194049 49593 194167
rect 49711 194049 67593 194167
rect 67711 194049 85593 194167
rect 85711 194049 103593 194167
rect 103711 194049 121593 194167
rect 121711 194049 139593 194167
rect 139711 194049 157593 194167
rect 157711 194049 175593 194167
rect 175711 194049 193593 194167
rect 193711 194049 211593 194167
rect 211711 194049 229593 194167
rect 229711 194049 247593 194167
rect 247711 194049 265593 194167
rect 265711 194049 283593 194167
rect 283711 194049 295101 194167
rect 295219 194049 295310 194167
rect -3348 194038 295310 194049
rect -3348 194037 -3048 194038
rect 13502 194037 13802 194038
rect 31502 194037 31802 194038
rect 49502 194037 49802 194038
rect 67502 194037 67802 194038
rect 85502 194037 85802 194038
rect 103502 194037 103802 194038
rect 121502 194037 121802 194038
rect 139502 194037 139802 194038
rect 157502 194037 157802 194038
rect 175502 194037 175802 194038
rect 193502 194037 193802 194038
rect 211502 194037 211802 194038
rect 229502 194037 229802 194038
rect 247502 194037 247802 194038
rect 265502 194037 265802 194038
rect 283502 194037 283802 194038
rect 295010 194037 295310 194038
rect -2408 192538 -2108 192539
rect 11702 192538 12002 192539
rect 29702 192538 30002 192539
rect 47702 192538 48002 192539
rect 65702 192538 66002 192539
rect 83702 192538 84002 192539
rect 101702 192538 102002 192539
rect 119702 192538 120002 192539
rect 137702 192538 138002 192539
rect 155702 192538 156002 192539
rect 173702 192538 174002 192539
rect 191702 192538 192002 192539
rect 209702 192538 210002 192539
rect 227702 192538 228002 192539
rect 245702 192538 246002 192539
rect 263702 192538 264002 192539
rect 281702 192538 282002 192539
rect 294070 192538 294370 192539
rect -2408 192527 294370 192538
rect -2408 192409 -2317 192527
rect -2199 192409 11793 192527
rect 11911 192409 29793 192527
rect 29911 192409 47793 192527
rect 47911 192409 65793 192527
rect 65911 192409 83793 192527
rect 83911 192409 101793 192527
rect 101911 192409 119793 192527
rect 119911 192409 137793 192527
rect 137911 192409 155793 192527
rect 155911 192409 173793 192527
rect 173911 192409 191793 192527
rect 191911 192409 209793 192527
rect 209911 192409 227793 192527
rect 227911 192409 245793 192527
rect 245911 192409 263793 192527
rect 263911 192409 281793 192527
rect 281911 192409 294161 192527
rect 294279 192409 294370 192527
rect -2408 192367 294370 192409
rect -2408 192249 -2317 192367
rect -2199 192249 11793 192367
rect 11911 192249 29793 192367
rect 29911 192249 47793 192367
rect 47911 192249 65793 192367
rect 65911 192249 83793 192367
rect 83911 192249 101793 192367
rect 101911 192249 119793 192367
rect 119911 192249 137793 192367
rect 137911 192249 155793 192367
rect 155911 192249 173793 192367
rect 173911 192249 191793 192367
rect 191911 192249 209793 192367
rect 209911 192249 227793 192367
rect 227911 192249 245793 192367
rect 245911 192249 263793 192367
rect 263911 192249 281793 192367
rect 281911 192249 294161 192367
rect 294279 192249 294370 192367
rect -2408 192238 294370 192249
rect -2408 192237 -2108 192238
rect 11702 192237 12002 192238
rect 29702 192237 30002 192238
rect 47702 192237 48002 192238
rect 65702 192237 66002 192238
rect 83702 192237 84002 192238
rect 101702 192237 102002 192238
rect 119702 192237 120002 192238
rect 137702 192237 138002 192238
rect 155702 192237 156002 192238
rect 173702 192237 174002 192238
rect 191702 192237 192002 192238
rect 209702 192237 210002 192238
rect 227702 192237 228002 192238
rect 245702 192237 246002 192238
rect 263702 192237 264002 192238
rect 281702 192237 282002 192238
rect 294070 192237 294370 192238
rect -1468 190738 -1168 190739
rect 9902 190738 10202 190739
rect 27902 190738 28202 190739
rect 45902 190738 46202 190739
rect 63902 190738 64202 190739
rect 81902 190738 82202 190739
rect 99902 190738 100202 190739
rect 117902 190738 118202 190739
rect 135902 190738 136202 190739
rect 153902 190738 154202 190739
rect 171902 190738 172202 190739
rect 189902 190738 190202 190739
rect 207902 190738 208202 190739
rect 225902 190738 226202 190739
rect 243902 190738 244202 190739
rect 261902 190738 262202 190739
rect 279902 190738 280202 190739
rect 293130 190738 293430 190739
rect -1468 190727 293430 190738
rect -1468 190609 -1377 190727
rect -1259 190609 9993 190727
rect 10111 190609 27993 190727
rect 28111 190609 45993 190727
rect 46111 190609 63993 190727
rect 64111 190609 81993 190727
rect 82111 190609 99993 190727
rect 100111 190609 117993 190727
rect 118111 190609 135993 190727
rect 136111 190609 153993 190727
rect 154111 190609 171993 190727
rect 172111 190609 189993 190727
rect 190111 190609 207993 190727
rect 208111 190609 225993 190727
rect 226111 190609 243993 190727
rect 244111 190609 261993 190727
rect 262111 190609 279993 190727
rect 280111 190609 293221 190727
rect 293339 190609 293430 190727
rect -1468 190567 293430 190609
rect -1468 190449 -1377 190567
rect -1259 190449 9993 190567
rect 10111 190449 27993 190567
rect 28111 190449 45993 190567
rect 46111 190449 63993 190567
rect 64111 190449 81993 190567
rect 82111 190449 99993 190567
rect 100111 190449 117993 190567
rect 118111 190449 135993 190567
rect 136111 190449 153993 190567
rect 154111 190449 171993 190567
rect 172111 190449 189993 190567
rect 190111 190449 207993 190567
rect 208111 190449 225993 190567
rect 226111 190449 243993 190567
rect 244111 190449 261993 190567
rect 262111 190449 279993 190567
rect 280111 190449 293221 190567
rect 293339 190449 293430 190567
rect -1468 190438 293430 190449
rect -1468 190437 -1168 190438
rect 9902 190437 10202 190438
rect 27902 190437 28202 190438
rect 45902 190437 46202 190438
rect 63902 190437 64202 190438
rect 81902 190437 82202 190438
rect 99902 190437 100202 190438
rect 117902 190437 118202 190438
rect 135902 190437 136202 190438
rect 153902 190437 154202 190438
rect 171902 190437 172202 190438
rect 189902 190437 190202 190438
rect 207902 190437 208202 190438
rect 225902 190437 226202 190438
rect 243902 190437 244202 190438
rect 261902 190437 262202 190438
rect 279902 190437 280202 190438
rect 293130 190437 293430 190438
rect -3818 187138 -3518 187139
rect 6302 187138 6602 187139
rect 24302 187138 24602 187139
rect 42302 187138 42602 187139
rect 60302 187138 60602 187139
rect 78302 187138 78602 187139
rect 96302 187138 96602 187139
rect 114302 187138 114602 187139
rect 132302 187138 132602 187139
rect 150302 187138 150602 187139
rect 168302 187138 168602 187139
rect 186302 187138 186602 187139
rect 204302 187138 204602 187139
rect 222302 187138 222602 187139
rect 240302 187138 240602 187139
rect 258302 187138 258602 187139
rect 276302 187138 276602 187139
rect 295480 187138 295780 187139
rect -4288 187127 296250 187138
rect -4288 187009 -3727 187127
rect -3609 187009 6393 187127
rect 6511 187009 24393 187127
rect 24511 187009 42393 187127
rect 42511 187009 60393 187127
rect 60511 187009 78393 187127
rect 78511 187009 96393 187127
rect 96511 187009 114393 187127
rect 114511 187009 132393 187127
rect 132511 187009 150393 187127
rect 150511 187009 168393 187127
rect 168511 187009 186393 187127
rect 186511 187009 204393 187127
rect 204511 187009 222393 187127
rect 222511 187009 240393 187127
rect 240511 187009 258393 187127
rect 258511 187009 276393 187127
rect 276511 187009 295571 187127
rect 295689 187009 296250 187127
rect -4288 186967 296250 187009
rect -4288 186849 -3727 186967
rect -3609 186849 6393 186967
rect 6511 186849 24393 186967
rect 24511 186849 42393 186967
rect 42511 186849 60393 186967
rect 60511 186849 78393 186967
rect 78511 186849 96393 186967
rect 96511 186849 114393 186967
rect 114511 186849 132393 186967
rect 132511 186849 150393 186967
rect 150511 186849 168393 186967
rect 168511 186849 186393 186967
rect 186511 186849 204393 186967
rect 204511 186849 222393 186967
rect 222511 186849 240393 186967
rect 240511 186849 258393 186967
rect 258511 186849 276393 186967
rect 276511 186849 295571 186967
rect 295689 186849 296250 186967
rect -4288 186838 296250 186849
rect -3818 186837 -3518 186838
rect 6302 186837 6602 186838
rect 24302 186837 24602 186838
rect 42302 186837 42602 186838
rect 60302 186837 60602 186838
rect 78302 186837 78602 186838
rect 96302 186837 96602 186838
rect 114302 186837 114602 186838
rect 132302 186837 132602 186838
rect 150302 186837 150602 186838
rect 168302 186837 168602 186838
rect 186302 186837 186602 186838
rect 204302 186837 204602 186838
rect 222302 186837 222602 186838
rect 240302 186837 240602 186838
rect 258302 186837 258602 186838
rect 276302 186837 276602 186838
rect 295480 186837 295780 186838
rect -2878 185338 -2578 185339
rect 4502 185338 4802 185339
rect 22502 185338 22802 185339
rect 40502 185338 40802 185339
rect 58502 185338 58802 185339
rect 76502 185338 76802 185339
rect 94502 185338 94802 185339
rect 112502 185338 112802 185339
rect 130502 185338 130802 185339
rect 148502 185338 148802 185339
rect 166502 185338 166802 185339
rect 184502 185338 184802 185339
rect 202502 185338 202802 185339
rect 220502 185338 220802 185339
rect 238502 185338 238802 185339
rect 256502 185338 256802 185339
rect 274502 185338 274802 185339
rect 294540 185338 294840 185339
rect -3348 185327 295310 185338
rect -3348 185209 -2787 185327
rect -2669 185209 4593 185327
rect 4711 185209 22593 185327
rect 22711 185209 40593 185327
rect 40711 185209 58593 185327
rect 58711 185209 76593 185327
rect 76711 185209 94593 185327
rect 94711 185209 112593 185327
rect 112711 185209 130593 185327
rect 130711 185209 148593 185327
rect 148711 185209 166593 185327
rect 166711 185209 184593 185327
rect 184711 185209 202593 185327
rect 202711 185209 220593 185327
rect 220711 185209 238593 185327
rect 238711 185209 256593 185327
rect 256711 185209 274593 185327
rect 274711 185209 294631 185327
rect 294749 185209 295310 185327
rect -3348 185167 295310 185209
rect -3348 185049 -2787 185167
rect -2669 185049 4593 185167
rect 4711 185049 22593 185167
rect 22711 185049 40593 185167
rect 40711 185049 58593 185167
rect 58711 185049 76593 185167
rect 76711 185049 94593 185167
rect 94711 185049 112593 185167
rect 112711 185049 130593 185167
rect 130711 185049 148593 185167
rect 148711 185049 166593 185167
rect 166711 185049 184593 185167
rect 184711 185049 202593 185167
rect 202711 185049 220593 185167
rect 220711 185049 238593 185167
rect 238711 185049 256593 185167
rect 256711 185049 274593 185167
rect 274711 185049 294631 185167
rect 294749 185049 295310 185167
rect -3348 185038 295310 185049
rect -2878 185037 -2578 185038
rect 4502 185037 4802 185038
rect 22502 185037 22802 185038
rect 40502 185037 40802 185038
rect 58502 185037 58802 185038
rect 76502 185037 76802 185038
rect 94502 185037 94802 185038
rect 112502 185037 112802 185038
rect 130502 185037 130802 185038
rect 148502 185037 148802 185038
rect 166502 185037 166802 185038
rect 184502 185037 184802 185038
rect 202502 185037 202802 185038
rect 220502 185037 220802 185038
rect 238502 185037 238802 185038
rect 256502 185037 256802 185038
rect 274502 185037 274802 185038
rect 294540 185037 294840 185038
rect -1938 183538 -1638 183539
rect 2702 183538 3002 183539
rect 20702 183538 21002 183539
rect 38702 183538 39002 183539
rect 56702 183538 57002 183539
rect 74702 183538 75002 183539
rect 92702 183538 93002 183539
rect 110702 183538 111002 183539
rect 128702 183538 129002 183539
rect 146702 183538 147002 183539
rect 164702 183538 165002 183539
rect 182702 183538 183002 183539
rect 200702 183538 201002 183539
rect 218702 183538 219002 183539
rect 236702 183538 237002 183539
rect 254702 183538 255002 183539
rect 272702 183538 273002 183539
rect 290702 183538 291002 183539
rect 293600 183538 293900 183539
rect -2408 183527 294370 183538
rect -2408 183409 -1847 183527
rect -1729 183409 2793 183527
rect 2911 183409 20793 183527
rect 20911 183409 38793 183527
rect 38911 183409 56793 183527
rect 56911 183409 74793 183527
rect 74911 183409 92793 183527
rect 92911 183409 110793 183527
rect 110911 183409 128793 183527
rect 128911 183409 146793 183527
rect 146911 183409 164793 183527
rect 164911 183409 182793 183527
rect 182911 183409 200793 183527
rect 200911 183409 218793 183527
rect 218911 183409 236793 183527
rect 236911 183409 254793 183527
rect 254911 183409 272793 183527
rect 272911 183409 290793 183527
rect 290911 183409 293691 183527
rect 293809 183409 294370 183527
rect -2408 183367 294370 183409
rect -2408 183249 -1847 183367
rect -1729 183249 2793 183367
rect 2911 183249 20793 183367
rect 20911 183249 38793 183367
rect 38911 183249 56793 183367
rect 56911 183249 74793 183367
rect 74911 183249 92793 183367
rect 92911 183249 110793 183367
rect 110911 183249 128793 183367
rect 128911 183249 146793 183367
rect 146911 183249 164793 183367
rect 164911 183249 182793 183367
rect 182911 183249 200793 183367
rect 200911 183249 218793 183367
rect 218911 183249 236793 183367
rect 236911 183249 254793 183367
rect 254911 183249 272793 183367
rect 272911 183249 290793 183367
rect 290911 183249 293691 183367
rect 293809 183249 294370 183367
rect -2408 183238 294370 183249
rect -1938 183237 -1638 183238
rect 2702 183237 3002 183238
rect 20702 183237 21002 183238
rect 38702 183237 39002 183238
rect 56702 183237 57002 183238
rect 74702 183237 75002 183238
rect 92702 183237 93002 183238
rect 110702 183237 111002 183238
rect 128702 183237 129002 183238
rect 146702 183237 147002 183238
rect 164702 183237 165002 183238
rect 182702 183237 183002 183238
rect 200702 183237 201002 183238
rect 218702 183237 219002 183238
rect 236702 183237 237002 183238
rect 254702 183237 255002 183238
rect 272702 183237 273002 183238
rect 290702 183237 291002 183238
rect 293600 183237 293900 183238
rect -998 181738 -698 181739
rect 902 181738 1202 181739
rect 18902 181738 19202 181739
rect 36902 181738 37202 181739
rect 54902 181738 55202 181739
rect 72902 181738 73202 181739
rect 90902 181738 91202 181739
rect 108902 181738 109202 181739
rect 126902 181738 127202 181739
rect 144902 181738 145202 181739
rect 162902 181738 163202 181739
rect 180902 181738 181202 181739
rect 198902 181738 199202 181739
rect 216902 181738 217202 181739
rect 234902 181738 235202 181739
rect 252902 181738 253202 181739
rect 270902 181738 271202 181739
rect 288902 181738 289202 181739
rect 292660 181738 292960 181739
rect -1468 181727 293430 181738
rect -1468 181609 -907 181727
rect -789 181609 993 181727
rect 1111 181609 18993 181727
rect 19111 181609 36993 181727
rect 37111 181609 54993 181727
rect 55111 181609 72993 181727
rect 73111 181609 90993 181727
rect 91111 181609 108993 181727
rect 109111 181609 126993 181727
rect 127111 181609 144993 181727
rect 145111 181609 162993 181727
rect 163111 181609 180993 181727
rect 181111 181609 198993 181727
rect 199111 181609 216993 181727
rect 217111 181609 234993 181727
rect 235111 181609 252993 181727
rect 253111 181609 270993 181727
rect 271111 181609 288993 181727
rect 289111 181609 292751 181727
rect 292869 181609 293430 181727
rect -1468 181567 293430 181609
rect -1468 181449 -907 181567
rect -789 181449 993 181567
rect 1111 181449 18993 181567
rect 19111 181449 36993 181567
rect 37111 181449 54993 181567
rect 55111 181449 72993 181567
rect 73111 181449 90993 181567
rect 91111 181449 108993 181567
rect 109111 181449 126993 181567
rect 127111 181449 144993 181567
rect 145111 181449 162993 181567
rect 163111 181449 180993 181567
rect 181111 181449 198993 181567
rect 199111 181449 216993 181567
rect 217111 181449 234993 181567
rect 235111 181449 252993 181567
rect 253111 181449 270993 181567
rect 271111 181449 288993 181567
rect 289111 181449 292751 181567
rect 292869 181449 293430 181567
rect -1468 181438 293430 181449
rect -998 181437 -698 181438
rect 902 181437 1202 181438
rect 18902 181437 19202 181438
rect 36902 181437 37202 181438
rect 54902 181437 55202 181438
rect 72902 181437 73202 181438
rect 90902 181437 91202 181438
rect 108902 181437 109202 181438
rect 126902 181437 127202 181438
rect 144902 181437 145202 181438
rect 162902 181437 163202 181438
rect 180902 181437 181202 181438
rect 198902 181437 199202 181438
rect 216902 181437 217202 181438
rect 234902 181437 235202 181438
rect 252902 181437 253202 181438
rect 270902 181437 271202 181438
rect 288902 181437 289202 181438
rect 292660 181437 292960 181438
rect -4288 178138 -3988 178139
rect 15302 178138 15602 178139
rect 33302 178138 33602 178139
rect 51302 178138 51602 178139
rect 69302 178138 69602 178139
rect 87302 178138 87602 178139
rect 105302 178138 105602 178139
rect 123302 178138 123602 178139
rect 141302 178138 141602 178139
rect 159302 178138 159602 178139
rect 177302 178138 177602 178139
rect 195302 178138 195602 178139
rect 213302 178138 213602 178139
rect 231302 178138 231602 178139
rect 249302 178138 249602 178139
rect 267302 178138 267602 178139
rect 285302 178138 285602 178139
rect 295950 178138 296250 178139
rect -4288 178127 296250 178138
rect -4288 178009 -4197 178127
rect -4079 178009 15393 178127
rect 15511 178009 33393 178127
rect 33511 178009 51393 178127
rect 51511 178009 69393 178127
rect 69511 178009 87393 178127
rect 87511 178009 105393 178127
rect 105511 178009 123393 178127
rect 123511 178009 141393 178127
rect 141511 178009 159393 178127
rect 159511 178009 177393 178127
rect 177511 178009 195393 178127
rect 195511 178009 213393 178127
rect 213511 178009 231393 178127
rect 231511 178009 249393 178127
rect 249511 178009 267393 178127
rect 267511 178009 285393 178127
rect 285511 178009 296041 178127
rect 296159 178009 296250 178127
rect -4288 177967 296250 178009
rect -4288 177849 -4197 177967
rect -4079 177849 15393 177967
rect 15511 177849 33393 177967
rect 33511 177849 51393 177967
rect 51511 177849 69393 177967
rect 69511 177849 87393 177967
rect 87511 177849 105393 177967
rect 105511 177849 123393 177967
rect 123511 177849 141393 177967
rect 141511 177849 159393 177967
rect 159511 177849 177393 177967
rect 177511 177849 195393 177967
rect 195511 177849 213393 177967
rect 213511 177849 231393 177967
rect 231511 177849 249393 177967
rect 249511 177849 267393 177967
rect 267511 177849 285393 177967
rect 285511 177849 296041 177967
rect 296159 177849 296250 177967
rect -4288 177838 296250 177849
rect -4288 177837 -3988 177838
rect 15302 177837 15602 177838
rect 33302 177837 33602 177838
rect 51302 177837 51602 177838
rect 69302 177837 69602 177838
rect 87302 177837 87602 177838
rect 105302 177837 105602 177838
rect 123302 177837 123602 177838
rect 141302 177837 141602 177838
rect 159302 177837 159602 177838
rect 177302 177837 177602 177838
rect 195302 177837 195602 177838
rect 213302 177837 213602 177838
rect 231302 177837 231602 177838
rect 249302 177837 249602 177838
rect 267302 177837 267602 177838
rect 285302 177837 285602 177838
rect 295950 177837 296250 177838
rect -3348 176338 -3048 176339
rect 13502 176338 13802 176339
rect 31502 176338 31802 176339
rect 49502 176338 49802 176339
rect 67502 176338 67802 176339
rect 85502 176338 85802 176339
rect 103502 176338 103802 176339
rect 121502 176338 121802 176339
rect 139502 176338 139802 176339
rect 157502 176338 157802 176339
rect 175502 176338 175802 176339
rect 193502 176338 193802 176339
rect 211502 176338 211802 176339
rect 229502 176338 229802 176339
rect 247502 176338 247802 176339
rect 265502 176338 265802 176339
rect 283502 176338 283802 176339
rect 295010 176338 295310 176339
rect -3348 176327 295310 176338
rect -3348 176209 -3257 176327
rect -3139 176209 13593 176327
rect 13711 176209 31593 176327
rect 31711 176209 49593 176327
rect 49711 176209 67593 176327
rect 67711 176209 85593 176327
rect 85711 176209 103593 176327
rect 103711 176209 121593 176327
rect 121711 176209 139593 176327
rect 139711 176209 157593 176327
rect 157711 176209 175593 176327
rect 175711 176209 193593 176327
rect 193711 176209 211593 176327
rect 211711 176209 229593 176327
rect 229711 176209 247593 176327
rect 247711 176209 265593 176327
rect 265711 176209 283593 176327
rect 283711 176209 295101 176327
rect 295219 176209 295310 176327
rect -3348 176167 295310 176209
rect -3348 176049 -3257 176167
rect -3139 176049 13593 176167
rect 13711 176049 31593 176167
rect 31711 176049 49593 176167
rect 49711 176049 67593 176167
rect 67711 176049 85593 176167
rect 85711 176049 103593 176167
rect 103711 176049 121593 176167
rect 121711 176049 139593 176167
rect 139711 176049 157593 176167
rect 157711 176049 175593 176167
rect 175711 176049 193593 176167
rect 193711 176049 211593 176167
rect 211711 176049 229593 176167
rect 229711 176049 247593 176167
rect 247711 176049 265593 176167
rect 265711 176049 283593 176167
rect 283711 176049 295101 176167
rect 295219 176049 295310 176167
rect -3348 176038 295310 176049
rect -3348 176037 -3048 176038
rect 13502 176037 13802 176038
rect 31502 176037 31802 176038
rect 49502 176037 49802 176038
rect 67502 176037 67802 176038
rect 85502 176037 85802 176038
rect 103502 176037 103802 176038
rect 121502 176037 121802 176038
rect 139502 176037 139802 176038
rect 157502 176037 157802 176038
rect 175502 176037 175802 176038
rect 193502 176037 193802 176038
rect 211502 176037 211802 176038
rect 229502 176037 229802 176038
rect 247502 176037 247802 176038
rect 265502 176037 265802 176038
rect 283502 176037 283802 176038
rect 295010 176037 295310 176038
rect -2408 174538 -2108 174539
rect 11702 174538 12002 174539
rect 29702 174538 30002 174539
rect 47702 174538 48002 174539
rect 65702 174538 66002 174539
rect 83702 174538 84002 174539
rect 101702 174538 102002 174539
rect 119702 174538 120002 174539
rect 137702 174538 138002 174539
rect 155702 174538 156002 174539
rect 173702 174538 174002 174539
rect 191702 174538 192002 174539
rect 209702 174538 210002 174539
rect 227702 174538 228002 174539
rect 245702 174538 246002 174539
rect 263702 174538 264002 174539
rect 281702 174538 282002 174539
rect 294070 174538 294370 174539
rect -2408 174527 294370 174538
rect -2408 174409 -2317 174527
rect -2199 174409 11793 174527
rect 11911 174409 29793 174527
rect 29911 174409 47793 174527
rect 47911 174409 65793 174527
rect 65911 174409 83793 174527
rect 83911 174409 101793 174527
rect 101911 174409 119793 174527
rect 119911 174409 137793 174527
rect 137911 174409 155793 174527
rect 155911 174409 173793 174527
rect 173911 174409 191793 174527
rect 191911 174409 209793 174527
rect 209911 174409 227793 174527
rect 227911 174409 245793 174527
rect 245911 174409 263793 174527
rect 263911 174409 281793 174527
rect 281911 174409 294161 174527
rect 294279 174409 294370 174527
rect -2408 174367 294370 174409
rect -2408 174249 -2317 174367
rect -2199 174249 11793 174367
rect 11911 174249 29793 174367
rect 29911 174249 47793 174367
rect 47911 174249 65793 174367
rect 65911 174249 83793 174367
rect 83911 174249 101793 174367
rect 101911 174249 119793 174367
rect 119911 174249 137793 174367
rect 137911 174249 155793 174367
rect 155911 174249 173793 174367
rect 173911 174249 191793 174367
rect 191911 174249 209793 174367
rect 209911 174249 227793 174367
rect 227911 174249 245793 174367
rect 245911 174249 263793 174367
rect 263911 174249 281793 174367
rect 281911 174249 294161 174367
rect 294279 174249 294370 174367
rect -2408 174238 294370 174249
rect -2408 174237 -2108 174238
rect 11702 174237 12002 174238
rect 29702 174237 30002 174238
rect 47702 174237 48002 174238
rect 65702 174237 66002 174238
rect 83702 174237 84002 174238
rect 101702 174237 102002 174238
rect 119702 174237 120002 174238
rect 137702 174237 138002 174238
rect 155702 174237 156002 174238
rect 173702 174237 174002 174238
rect 191702 174237 192002 174238
rect 209702 174237 210002 174238
rect 227702 174237 228002 174238
rect 245702 174237 246002 174238
rect 263702 174237 264002 174238
rect 281702 174237 282002 174238
rect 294070 174237 294370 174238
rect -1468 172738 -1168 172739
rect 9902 172738 10202 172739
rect 27902 172738 28202 172739
rect 45902 172738 46202 172739
rect 63902 172738 64202 172739
rect 81902 172738 82202 172739
rect 99902 172738 100202 172739
rect 117902 172738 118202 172739
rect 135902 172738 136202 172739
rect 153902 172738 154202 172739
rect 171902 172738 172202 172739
rect 189902 172738 190202 172739
rect 207902 172738 208202 172739
rect 225902 172738 226202 172739
rect 243902 172738 244202 172739
rect 261902 172738 262202 172739
rect 279902 172738 280202 172739
rect 293130 172738 293430 172739
rect -1468 172727 293430 172738
rect -1468 172609 -1377 172727
rect -1259 172609 9993 172727
rect 10111 172609 27993 172727
rect 28111 172609 45993 172727
rect 46111 172609 63993 172727
rect 64111 172609 81993 172727
rect 82111 172609 99993 172727
rect 100111 172609 117993 172727
rect 118111 172609 135993 172727
rect 136111 172609 153993 172727
rect 154111 172609 171993 172727
rect 172111 172609 189993 172727
rect 190111 172609 207993 172727
rect 208111 172609 225993 172727
rect 226111 172609 243993 172727
rect 244111 172609 261993 172727
rect 262111 172609 279993 172727
rect 280111 172609 293221 172727
rect 293339 172609 293430 172727
rect -1468 172567 293430 172609
rect -1468 172449 -1377 172567
rect -1259 172449 9993 172567
rect 10111 172449 27993 172567
rect 28111 172449 45993 172567
rect 46111 172449 63993 172567
rect 64111 172449 81993 172567
rect 82111 172449 99993 172567
rect 100111 172449 117993 172567
rect 118111 172449 135993 172567
rect 136111 172449 153993 172567
rect 154111 172449 171993 172567
rect 172111 172449 189993 172567
rect 190111 172449 207993 172567
rect 208111 172449 225993 172567
rect 226111 172449 243993 172567
rect 244111 172449 261993 172567
rect 262111 172449 279993 172567
rect 280111 172449 293221 172567
rect 293339 172449 293430 172567
rect -1468 172438 293430 172449
rect -1468 172437 -1168 172438
rect 9902 172437 10202 172438
rect 27902 172437 28202 172438
rect 45902 172437 46202 172438
rect 63902 172437 64202 172438
rect 81902 172437 82202 172438
rect 99902 172437 100202 172438
rect 117902 172437 118202 172438
rect 135902 172437 136202 172438
rect 153902 172437 154202 172438
rect 171902 172437 172202 172438
rect 189902 172437 190202 172438
rect 207902 172437 208202 172438
rect 225902 172437 226202 172438
rect 243902 172437 244202 172438
rect 261902 172437 262202 172438
rect 279902 172437 280202 172438
rect 293130 172437 293430 172438
rect -3818 169138 -3518 169139
rect 6302 169138 6602 169139
rect 24302 169138 24602 169139
rect 42302 169138 42602 169139
rect 60302 169138 60602 169139
rect 78302 169138 78602 169139
rect 96302 169138 96602 169139
rect 114302 169138 114602 169139
rect 132302 169138 132602 169139
rect 150302 169138 150602 169139
rect 168302 169138 168602 169139
rect 186302 169138 186602 169139
rect 204302 169138 204602 169139
rect 222302 169138 222602 169139
rect 240302 169138 240602 169139
rect 258302 169138 258602 169139
rect 276302 169138 276602 169139
rect 295480 169138 295780 169139
rect -4288 169127 296250 169138
rect -4288 169009 -3727 169127
rect -3609 169009 6393 169127
rect 6511 169009 24393 169127
rect 24511 169009 42393 169127
rect 42511 169009 60393 169127
rect 60511 169009 78393 169127
rect 78511 169009 96393 169127
rect 96511 169009 114393 169127
rect 114511 169009 132393 169127
rect 132511 169009 150393 169127
rect 150511 169009 168393 169127
rect 168511 169009 186393 169127
rect 186511 169009 204393 169127
rect 204511 169009 222393 169127
rect 222511 169009 240393 169127
rect 240511 169009 258393 169127
rect 258511 169009 276393 169127
rect 276511 169009 295571 169127
rect 295689 169009 296250 169127
rect -4288 168967 296250 169009
rect -4288 168849 -3727 168967
rect -3609 168849 6393 168967
rect 6511 168849 24393 168967
rect 24511 168849 42393 168967
rect 42511 168849 60393 168967
rect 60511 168849 78393 168967
rect 78511 168849 96393 168967
rect 96511 168849 114393 168967
rect 114511 168849 132393 168967
rect 132511 168849 150393 168967
rect 150511 168849 168393 168967
rect 168511 168849 186393 168967
rect 186511 168849 204393 168967
rect 204511 168849 222393 168967
rect 222511 168849 240393 168967
rect 240511 168849 258393 168967
rect 258511 168849 276393 168967
rect 276511 168849 295571 168967
rect 295689 168849 296250 168967
rect -4288 168838 296250 168849
rect -3818 168837 -3518 168838
rect 6302 168837 6602 168838
rect 24302 168837 24602 168838
rect 42302 168837 42602 168838
rect 60302 168837 60602 168838
rect 78302 168837 78602 168838
rect 96302 168837 96602 168838
rect 114302 168837 114602 168838
rect 132302 168837 132602 168838
rect 150302 168837 150602 168838
rect 168302 168837 168602 168838
rect 186302 168837 186602 168838
rect 204302 168837 204602 168838
rect 222302 168837 222602 168838
rect 240302 168837 240602 168838
rect 258302 168837 258602 168838
rect 276302 168837 276602 168838
rect 295480 168837 295780 168838
rect -2878 167338 -2578 167339
rect 4502 167338 4802 167339
rect 22502 167338 22802 167339
rect 40502 167338 40802 167339
rect 58502 167338 58802 167339
rect 76502 167338 76802 167339
rect 94502 167338 94802 167339
rect 112502 167338 112802 167339
rect 130502 167338 130802 167339
rect 148502 167338 148802 167339
rect 166502 167338 166802 167339
rect 184502 167338 184802 167339
rect 202502 167338 202802 167339
rect 220502 167338 220802 167339
rect 238502 167338 238802 167339
rect 256502 167338 256802 167339
rect 274502 167338 274802 167339
rect 294540 167338 294840 167339
rect -3348 167327 295310 167338
rect -3348 167209 -2787 167327
rect -2669 167209 4593 167327
rect 4711 167209 22593 167327
rect 22711 167209 40593 167327
rect 40711 167209 58593 167327
rect 58711 167209 76593 167327
rect 76711 167209 94593 167327
rect 94711 167209 112593 167327
rect 112711 167209 130593 167327
rect 130711 167209 148593 167327
rect 148711 167209 166593 167327
rect 166711 167209 184593 167327
rect 184711 167209 202593 167327
rect 202711 167209 220593 167327
rect 220711 167209 238593 167327
rect 238711 167209 256593 167327
rect 256711 167209 274593 167327
rect 274711 167209 294631 167327
rect 294749 167209 295310 167327
rect -3348 167167 295310 167209
rect -3348 167049 -2787 167167
rect -2669 167049 4593 167167
rect 4711 167049 22593 167167
rect 22711 167049 40593 167167
rect 40711 167049 58593 167167
rect 58711 167049 76593 167167
rect 76711 167049 94593 167167
rect 94711 167049 112593 167167
rect 112711 167049 130593 167167
rect 130711 167049 148593 167167
rect 148711 167049 166593 167167
rect 166711 167049 184593 167167
rect 184711 167049 202593 167167
rect 202711 167049 220593 167167
rect 220711 167049 238593 167167
rect 238711 167049 256593 167167
rect 256711 167049 274593 167167
rect 274711 167049 294631 167167
rect 294749 167049 295310 167167
rect -3348 167038 295310 167049
rect -2878 167037 -2578 167038
rect 4502 167037 4802 167038
rect 22502 167037 22802 167038
rect 40502 167037 40802 167038
rect 58502 167037 58802 167038
rect 76502 167037 76802 167038
rect 94502 167037 94802 167038
rect 112502 167037 112802 167038
rect 130502 167037 130802 167038
rect 148502 167037 148802 167038
rect 166502 167037 166802 167038
rect 184502 167037 184802 167038
rect 202502 167037 202802 167038
rect 220502 167037 220802 167038
rect 238502 167037 238802 167038
rect 256502 167037 256802 167038
rect 274502 167037 274802 167038
rect 294540 167037 294840 167038
rect -1938 165538 -1638 165539
rect 2702 165538 3002 165539
rect 20702 165538 21002 165539
rect 38702 165538 39002 165539
rect 56702 165538 57002 165539
rect 74702 165538 75002 165539
rect 92702 165538 93002 165539
rect 110702 165538 111002 165539
rect 128702 165538 129002 165539
rect 146702 165538 147002 165539
rect 164702 165538 165002 165539
rect 182702 165538 183002 165539
rect 200702 165538 201002 165539
rect 218702 165538 219002 165539
rect 236702 165538 237002 165539
rect 254702 165538 255002 165539
rect 272702 165538 273002 165539
rect 290702 165538 291002 165539
rect 293600 165538 293900 165539
rect -2408 165527 294370 165538
rect -2408 165409 -1847 165527
rect -1729 165409 2793 165527
rect 2911 165409 20793 165527
rect 20911 165409 38793 165527
rect 38911 165409 56793 165527
rect 56911 165409 74793 165527
rect 74911 165409 92793 165527
rect 92911 165409 110793 165527
rect 110911 165409 128793 165527
rect 128911 165409 146793 165527
rect 146911 165409 164793 165527
rect 164911 165409 182793 165527
rect 182911 165409 200793 165527
rect 200911 165409 218793 165527
rect 218911 165409 236793 165527
rect 236911 165409 254793 165527
rect 254911 165409 272793 165527
rect 272911 165409 290793 165527
rect 290911 165409 293691 165527
rect 293809 165409 294370 165527
rect -2408 165367 294370 165409
rect -2408 165249 -1847 165367
rect -1729 165249 2793 165367
rect 2911 165249 20793 165367
rect 20911 165249 38793 165367
rect 38911 165249 56793 165367
rect 56911 165249 74793 165367
rect 74911 165249 92793 165367
rect 92911 165249 110793 165367
rect 110911 165249 128793 165367
rect 128911 165249 146793 165367
rect 146911 165249 164793 165367
rect 164911 165249 182793 165367
rect 182911 165249 200793 165367
rect 200911 165249 218793 165367
rect 218911 165249 236793 165367
rect 236911 165249 254793 165367
rect 254911 165249 272793 165367
rect 272911 165249 290793 165367
rect 290911 165249 293691 165367
rect 293809 165249 294370 165367
rect -2408 165238 294370 165249
rect -1938 165237 -1638 165238
rect 2702 165237 3002 165238
rect 20702 165237 21002 165238
rect 38702 165237 39002 165238
rect 56702 165237 57002 165238
rect 74702 165237 75002 165238
rect 92702 165237 93002 165238
rect 110702 165237 111002 165238
rect 128702 165237 129002 165238
rect 146702 165237 147002 165238
rect 164702 165237 165002 165238
rect 182702 165237 183002 165238
rect 200702 165237 201002 165238
rect 218702 165237 219002 165238
rect 236702 165237 237002 165238
rect 254702 165237 255002 165238
rect 272702 165237 273002 165238
rect 290702 165237 291002 165238
rect 293600 165237 293900 165238
rect -998 163738 -698 163739
rect 902 163738 1202 163739
rect 18902 163738 19202 163739
rect 36902 163738 37202 163739
rect 54902 163738 55202 163739
rect 72902 163738 73202 163739
rect 90902 163738 91202 163739
rect 108902 163738 109202 163739
rect 126902 163738 127202 163739
rect 144902 163738 145202 163739
rect 162902 163738 163202 163739
rect 180902 163738 181202 163739
rect 198902 163738 199202 163739
rect 216902 163738 217202 163739
rect 234902 163738 235202 163739
rect 252902 163738 253202 163739
rect 270902 163738 271202 163739
rect 288902 163738 289202 163739
rect 292660 163738 292960 163739
rect -1468 163727 293430 163738
rect -1468 163609 -907 163727
rect -789 163609 993 163727
rect 1111 163609 18993 163727
rect 19111 163609 36993 163727
rect 37111 163609 54993 163727
rect 55111 163609 72993 163727
rect 73111 163609 90993 163727
rect 91111 163609 108993 163727
rect 109111 163609 126993 163727
rect 127111 163609 144993 163727
rect 145111 163609 162993 163727
rect 163111 163609 180993 163727
rect 181111 163609 198993 163727
rect 199111 163609 216993 163727
rect 217111 163609 234993 163727
rect 235111 163609 252993 163727
rect 253111 163609 270993 163727
rect 271111 163609 288993 163727
rect 289111 163609 292751 163727
rect 292869 163609 293430 163727
rect -1468 163567 293430 163609
rect -1468 163449 -907 163567
rect -789 163449 993 163567
rect 1111 163449 18993 163567
rect 19111 163449 36993 163567
rect 37111 163449 54993 163567
rect 55111 163449 72993 163567
rect 73111 163449 90993 163567
rect 91111 163449 108993 163567
rect 109111 163449 126993 163567
rect 127111 163449 144993 163567
rect 145111 163449 162993 163567
rect 163111 163449 180993 163567
rect 181111 163449 198993 163567
rect 199111 163449 216993 163567
rect 217111 163449 234993 163567
rect 235111 163449 252993 163567
rect 253111 163449 270993 163567
rect 271111 163449 288993 163567
rect 289111 163449 292751 163567
rect 292869 163449 293430 163567
rect -1468 163438 293430 163449
rect -998 163437 -698 163438
rect 902 163437 1202 163438
rect 18902 163437 19202 163438
rect 36902 163437 37202 163438
rect 54902 163437 55202 163438
rect 72902 163437 73202 163438
rect 90902 163437 91202 163438
rect 108902 163437 109202 163438
rect 126902 163437 127202 163438
rect 144902 163437 145202 163438
rect 162902 163437 163202 163438
rect 180902 163437 181202 163438
rect 198902 163437 199202 163438
rect 216902 163437 217202 163438
rect 234902 163437 235202 163438
rect 252902 163437 253202 163438
rect 270902 163437 271202 163438
rect 288902 163437 289202 163438
rect 292660 163437 292960 163438
rect -4288 160138 -3988 160139
rect 15302 160138 15602 160139
rect 33302 160138 33602 160139
rect 51302 160138 51602 160139
rect 69302 160138 69602 160139
rect 87302 160138 87602 160139
rect 105302 160138 105602 160139
rect 123302 160138 123602 160139
rect 141302 160138 141602 160139
rect 159302 160138 159602 160139
rect 177302 160138 177602 160139
rect 195302 160138 195602 160139
rect 213302 160138 213602 160139
rect 231302 160138 231602 160139
rect 249302 160138 249602 160139
rect 267302 160138 267602 160139
rect 285302 160138 285602 160139
rect 295950 160138 296250 160139
rect -4288 160127 296250 160138
rect -4288 160009 -4197 160127
rect -4079 160009 15393 160127
rect 15511 160009 33393 160127
rect 33511 160009 51393 160127
rect 51511 160009 69393 160127
rect 69511 160009 87393 160127
rect 87511 160009 105393 160127
rect 105511 160009 123393 160127
rect 123511 160009 141393 160127
rect 141511 160009 159393 160127
rect 159511 160009 177393 160127
rect 177511 160009 195393 160127
rect 195511 160009 213393 160127
rect 213511 160009 231393 160127
rect 231511 160009 249393 160127
rect 249511 160009 267393 160127
rect 267511 160009 285393 160127
rect 285511 160009 296041 160127
rect 296159 160009 296250 160127
rect -4288 159967 296250 160009
rect -4288 159849 -4197 159967
rect -4079 159849 15393 159967
rect 15511 159849 33393 159967
rect 33511 159849 51393 159967
rect 51511 159849 69393 159967
rect 69511 159849 87393 159967
rect 87511 159849 105393 159967
rect 105511 159849 123393 159967
rect 123511 159849 141393 159967
rect 141511 159849 159393 159967
rect 159511 159849 177393 159967
rect 177511 159849 195393 159967
rect 195511 159849 213393 159967
rect 213511 159849 231393 159967
rect 231511 159849 249393 159967
rect 249511 159849 267393 159967
rect 267511 159849 285393 159967
rect 285511 159849 296041 159967
rect 296159 159849 296250 159967
rect -4288 159838 296250 159849
rect -4288 159837 -3988 159838
rect 15302 159837 15602 159838
rect 33302 159837 33602 159838
rect 51302 159837 51602 159838
rect 69302 159837 69602 159838
rect 87302 159837 87602 159838
rect 105302 159837 105602 159838
rect 123302 159837 123602 159838
rect 141302 159837 141602 159838
rect 159302 159837 159602 159838
rect 177302 159837 177602 159838
rect 195302 159837 195602 159838
rect 213302 159837 213602 159838
rect 231302 159837 231602 159838
rect 249302 159837 249602 159838
rect 267302 159837 267602 159838
rect 285302 159837 285602 159838
rect 295950 159837 296250 159838
rect -3348 158338 -3048 158339
rect 13502 158338 13802 158339
rect 31502 158338 31802 158339
rect 49502 158338 49802 158339
rect 67502 158338 67802 158339
rect 85502 158338 85802 158339
rect 103502 158338 103802 158339
rect 121502 158338 121802 158339
rect 139502 158338 139802 158339
rect 157502 158338 157802 158339
rect 175502 158338 175802 158339
rect 193502 158338 193802 158339
rect 211502 158338 211802 158339
rect 229502 158338 229802 158339
rect 247502 158338 247802 158339
rect 265502 158338 265802 158339
rect 283502 158338 283802 158339
rect 295010 158338 295310 158339
rect -3348 158327 295310 158338
rect -3348 158209 -3257 158327
rect -3139 158209 13593 158327
rect 13711 158209 31593 158327
rect 31711 158209 49593 158327
rect 49711 158209 67593 158327
rect 67711 158209 85593 158327
rect 85711 158209 103593 158327
rect 103711 158209 121593 158327
rect 121711 158209 139593 158327
rect 139711 158209 157593 158327
rect 157711 158209 175593 158327
rect 175711 158209 193593 158327
rect 193711 158209 211593 158327
rect 211711 158209 229593 158327
rect 229711 158209 247593 158327
rect 247711 158209 265593 158327
rect 265711 158209 283593 158327
rect 283711 158209 295101 158327
rect 295219 158209 295310 158327
rect -3348 158167 295310 158209
rect -3348 158049 -3257 158167
rect -3139 158049 13593 158167
rect 13711 158049 31593 158167
rect 31711 158049 49593 158167
rect 49711 158049 67593 158167
rect 67711 158049 85593 158167
rect 85711 158049 103593 158167
rect 103711 158049 121593 158167
rect 121711 158049 139593 158167
rect 139711 158049 157593 158167
rect 157711 158049 175593 158167
rect 175711 158049 193593 158167
rect 193711 158049 211593 158167
rect 211711 158049 229593 158167
rect 229711 158049 247593 158167
rect 247711 158049 265593 158167
rect 265711 158049 283593 158167
rect 283711 158049 295101 158167
rect 295219 158049 295310 158167
rect -3348 158038 295310 158049
rect -3348 158037 -3048 158038
rect 13502 158037 13802 158038
rect 31502 158037 31802 158038
rect 49502 158037 49802 158038
rect 67502 158037 67802 158038
rect 85502 158037 85802 158038
rect 103502 158037 103802 158038
rect 121502 158037 121802 158038
rect 139502 158037 139802 158038
rect 157502 158037 157802 158038
rect 175502 158037 175802 158038
rect 193502 158037 193802 158038
rect 211502 158037 211802 158038
rect 229502 158037 229802 158038
rect 247502 158037 247802 158038
rect 265502 158037 265802 158038
rect 283502 158037 283802 158038
rect 295010 158037 295310 158038
rect -2408 156538 -2108 156539
rect 11702 156538 12002 156539
rect 29702 156538 30002 156539
rect 47702 156538 48002 156539
rect 65702 156538 66002 156539
rect 83702 156538 84002 156539
rect 101702 156538 102002 156539
rect 119702 156538 120002 156539
rect 137702 156538 138002 156539
rect 155702 156538 156002 156539
rect 173702 156538 174002 156539
rect 191702 156538 192002 156539
rect 209702 156538 210002 156539
rect 227702 156538 228002 156539
rect 245702 156538 246002 156539
rect 263702 156538 264002 156539
rect 281702 156538 282002 156539
rect 294070 156538 294370 156539
rect -2408 156527 294370 156538
rect -2408 156409 -2317 156527
rect -2199 156409 11793 156527
rect 11911 156409 29793 156527
rect 29911 156409 47793 156527
rect 47911 156409 65793 156527
rect 65911 156409 83793 156527
rect 83911 156409 101793 156527
rect 101911 156409 119793 156527
rect 119911 156409 137793 156527
rect 137911 156409 155793 156527
rect 155911 156409 173793 156527
rect 173911 156409 191793 156527
rect 191911 156409 209793 156527
rect 209911 156409 227793 156527
rect 227911 156409 245793 156527
rect 245911 156409 263793 156527
rect 263911 156409 281793 156527
rect 281911 156409 294161 156527
rect 294279 156409 294370 156527
rect -2408 156367 294370 156409
rect -2408 156249 -2317 156367
rect -2199 156249 11793 156367
rect 11911 156249 29793 156367
rect 29911 156249 47793 156367
rect 47911 156249 65793 156367
rect 65911 156249 83793 156367
rect 83911 156249 101793 156367
rect 101911 156249 119793 156367
rect 119911 156249 137793 156367
rect 137911 156249 155793 156367
rect 155911 156249 173793 156367
rect 173911 156249 191793 156367
rect 191911 156249 209793 156367
rect 209911 156249 227793 156367
rect 227911 156249 245793 156367
rect 245911 156249 263793 156367
rect 263911 156249 281793 156367
rect 281911 156249 294161 156367
rect 294279 156249 294370 156367
rect -2408 156238 294370 156249
rect -2408 156237 -2108 156238
rect 11702 156237 12002 156238
rect 29702 156237 30002 156238
rect 47702 156237 48002 156238
rect 65702 156237 66002 156238
rect 83702 156237 84002 156238
rect 101702 156237 102002 156238
rect 119702 156237 120002 156238
rect 137702 156237 138002 156238
rect 155702 156237 156002 156238
rect 173702 156237 174002 156238
rect 191702 156237 192002 156238
rect 209702 156237 210002 156238
rect 227702 156237 228002 156238
rect 245702 156237 246002 156238
rect 263702 156237 264002 156238
rect 281702 156237 282002 156238
rect 294070 156237 294370 156238
rect -1468 154738 -1168 154739
rect 9902 154738 10202 154739
rect 27902 154738 28202 154739
rect 45902 154738 46202 154739
rect 63902 154738 64202 154739
rect 81902 154738 82202 154739
rect 99902 154738 100202 154739
rect 117902 154738 118202 154739
rect 135902 154738 136202 154739
rect 153902 154738 154202 154739
rect 171902 154738 172202 154739
rect 189902 154738 190202 154739
rect 207902 154738 208202 154739
rect 225902 154738 226202 154739
rect 243902 154738 244202 154739
rect 261902 154738 262202 154739
rect 279902 154738 280202 154739
rect 293130 154738 293430 154739
rect -1468 154727 293430 154738
rect -1468 154609 -1377 154727
rect -1259 154609 9993 154727
rect 10111 154609 27993 154727
rect 28111 154609 45993 154727
rect 46111 154609 63993 154727
rect 64111 154609 81993 154727
rect 82111 154609 99993 154727
rect 100111 154609 117993 154727
rect 118111 154609 135993 154727
rect 136111 154609 153993 154727
rect 154111 154609 171993 154727
rect 172111 154609 189993 154727
rect 190111 154609 207993 154727
rect 208111 154609 225993 154727
rect 226111 154609 243993 154727
rect 244111 154609 261993 154727
rect 262111 154609 279993 154727
rect 280111 154609 293221 154727
rect 293339 154609 293430 154727
rect -1468 154567 293430 154609
rect -1468 154449 -1377 154567
rect -1259 154449 9993 154567
rect 10111 154449 27993 154567
rect 28111 154449 45993 154567
rect 46111 154449 63993 154567
rect 64111 154449 81993 154567
rect 82111 154449 99993 154567
rect 100111 154449 117993 154567
rect 118111 154449 135993 154567
rect 136111 154449 153993 154567
rect 154111 154449 171993 154567
rect 172111 154449 189993 154567
rect 190111 154449 207993 154567
rect 208111 154449 225993 154567
rect 226111 154449 243993 154567
rect 244111 154449 261993 154567
rect 262111 154449 279993 154567
rect 280111 154449 293221 154567
rect 293339 154449 293430 154567
rect -1468 154438 293430 154449
rect -1468 154437 -1168 154438
rect 9902 154437 10202 154438
rect 27902 154437 28202 154438
rect 45902 154437 46202 154438
rect 63902 154437 64202 154438
rect 81902 154437 82202 154438
rect 99902 154437 100202 154438
rect 117902 154437 118202 154438
rect 135902 154437 136202 154438
rect 153902 154437 154202 154438
rect 171902 154437 172202 154438
rect 189902 154437 190202 154438
rect 207902 154437 208202 154438
rect 225902 154437 226202 154438
rect 243902 154437 244202 154438
rect 261902 154437 262202 154438
rect 279902 154437 280202 154438
rect 293130 154437 293430 154438
rect -3818 151138 -3518 151139
rect 6302 151138 6602 151139
rect 24302 151138 24602 151139
rect 42302 151138 42602 151139
rect 60302 151138 60602 151139
rect 78302 151138 78602 151139
rect 96302 151138 96602 151139
rect 114302 151138 114602 151139
rect 132302 151138 132602 151139
rect 150302 151138 150602 151139
rect 168302 151138 168602 151139
rect 186302 151138 186602 151139
rect 204302 151138 204602 151139
rect 222302 151138 222602 151139
rect 240302 151138 240602 151139
rect 258302 151138 258602 151139
rect 276302 151138 276602 151139
rect 295480 151138 295780 151139
rect -4288 151127 296250 151138
rect -4288 151009 -3727 151127
rect -3609 151009 6393 151127
rect 6511 151009 24393 151127
rect 24511 151009 42393 151127
rect 42511 151009 60393 151127
rect 60511 151009 78393 151127
rect 78511 151009 96393 151127
rect 96511 151009 114393 151127
rect 114511 151009 132393 151127
rect 132511 151009 150393 151127
rect 150511 151009 168393 151127
rect 168511 151009 186393 151127
rect 186511 151009 204393 151127
rect 204511 151009 222393 151127
rect 222511 151009 240393 151127
rect 240511 151009 258393 151127
rect 258511 151009 276393 151127
rect 276511 151009 295571 151127
rect 295689 151009 296250 151127
rect -4288 150967 296250 151009
rect -4288 150849 -3727 150967
rect -3609 150849 6393 150967
rect 6511 150849 24393 150967
rect 24511 150849 42393 150967
rect 42511 150849 60393 150967
rect 60511 150849 78393 150967
rect 78511 150849 96393 150967
rect 96511 150849 114393 150967
rect 114511 150849 132393 150967
rect 132511 150849 150393 150967
rect 150511 150849 168393 150967
rect 168511 150849 186393 150967
rect 186511 150849 204393 150967
rect 204511 150849 222393 150967
rect 222511 150849 240393 150967
rect 240511 150849 258393 150967
rect 258511 150849 276393 150967
rect 276511 150849 295571 150967
rect 295689 150849 296250 150967
rect -4288 150838 296250 150849
rect -3818 150837 -3518 150838
rect 6302 150837 6602 150838
rect 24302 150837 24602 150838
rect 42302 150837 42602 150838
rect 60302 150837 60602 150838
rect 78302 150837 78602 150838
rect 96302 150837 96602 150838
rect 114302 150837 114602 150838
rect 132302 150837 132602 150838
rect 150302 150837 150602 150838
rect 168302 150837 168602 150838
rect 186302 150837 186602 150838
rect 204302 150837 204602 150838
rect 222302 150837 222602 150838
rect 240302 150837 240602 150838
rect 258302 150837 258602 150838
rect 276302 150837 276602 150838
rect 295480 150837 295780 150838
rect -2878 149338 -2578 149339
rect 4502 149338 4802 149339
rect 22502 149338 22802 149339
rect 40502 149338 40802 149339
rect 58502 149338 58802 149339
rect 76502 149338 76802 149339
rect 94502 149338 94802 149339
rect 112502 149338 112802 149339
rect 130502 149338 130802 149339
rect 148502 149338 148802 149339
rect 166502 149338 166802 149339
rect 184502 149338 184802 149339
rect 202502 149338 202802 149339
rect 220502 149338 220802 149339
rect 238502 149338 238802 149339
rect 256502 149338 256802 149339
rect 274502 149338 274802 149339
rect 294540 149338 294840 149339
rect -3348 149327 295310 149338
rect -3348 149209 -2787 149327
rect -2669 149209 4593 149327
rect 4711 149209 22593 149327
rect 22711 149209 40593 149327
rect 40711 149209 58593 149327
rect 58711 149209 76593 149327
rect 76711 149209 94593 149327
rect 94711 149209 112593 149327
rect 112711 149209 130593 149327
rect 130711 149209 148593 149327
rect 148711 149209 166593 149327
rect 166711 149209 184593 149327
rect 184711 149209 202593 149327
rect 202711 149209 220593 149327
rect 220711 149209 238593 149327
rect 238711 149209 256593 149327
rect 256711 149209 274593 149327
rect 274711 149209 294631 149327
rect 294749 149209 295310 149327
rect -3348 149167 295310 149209
rect -3348 149049 -2787 149167
rect -2669 149049 4593 149167
rect 4711 149049 22593 149167
rect 22711 149049 40593 149167
rect 40711 149049 58593 149167
rect 58711 149049 76593 149167
rect 76711 149049 94593 149167
rect 94711 149049 112593 149167
rect 112711 149049 130593 149167
rect 130711 149049 148593 149167
rect 148711 149049 166593 149167
rect 166711 149049 184593 149167
rect 184711 149049 202593 149167
rect 202711 149049 220593 149167
rect 220711 149049 238593 149167
rect 238711 149049 256593 149167
rect 256711 149049 274593 149167
rect 274711 149049 294631 149167
rect 294749 149049 295310 149167
rect -3348 149038 295310 149049
rect -2878 149037 -2578 149038
rect 4502 149037 4802 149038
rect 22502 149037 22802 149038
rect 40502 149037 40802 149038
rect 58502 149037 58802 149038
rect 76502 149037 76802 149038
rect 94502 149037 94802 149038
rect 112502 149037 112802 149038
rect 130502 149037 130802 149038
rect 148502 149037 148802 149038
rect 166502 149037 166802 149038
rect 184502 149037 184802 149038
rect 202502 149037 202802 149038
rect 220502 149037 220802 149038
rect 238502 149037 238802 149038
rect 256502 149037 256802 149038
rect 274502 149037 274802 149038
rect 294540 149037 294840 149038
rect -1938 147538 -1638 147539
rect 2702 147538 3002 147539
rect 20702 147538 21002 147539
rect 38702 147538 39002 147539
rect 56702 147538 57002 147539
rect 74702 147538 75002 147539
rect 92702 147538 93002 147539
rect 110702 147538 111002 147539
rect 128702 147538 129002 147539
rect 146702 147538 147002 147539
rect 164702 147538 165002 147539
rect 182702 147538 183002 147539
rect 200702 147538 201002 147539
rect 218702 147538 219002 147539
rect 236702 147538 237002 147539
rect 254702 147538 255002 147539
rect 272702 147538 273002 147539
rect 290702 147538 291002 147539
rect 293600 147538 293900 147539
rect -2408 147527 294370 147538
rect -2408 147409 -1847 147527
rect -1729 147409 2793 147527
rect 2911 147409 20793 147527
rect 20911 147409 38793 147527
rect 38911 147409 56793 147527
rect 56911 147409 74793 147527
rect 74911 147409 92793 147527
rect 92911 147409 110793 147527
rect 110911 147409 128793 147527
rect 128911 147409 146793 147527
rect 146911 147409 164793 147527
rect 164911 147409 182793 147527
rect 182911 147409 200793 147527
rect 200911 147409 218793 147527
rect 218911 147409 236793 147527
rect 236911 147409 254793 147527
rect 254911 147409 272793 147527
rect 272911 147409 290793 147527
rect 290911 147409 293691 147527
rect 293809 147409 294370 147527
rect -2408 147367 294370 147409
rect -2408 147249 -1847 147367
rect -1729 147249 2793 147367
rect 2911 147249 20793 147367
rect 20911 147249 38793 147367
rect 38911 147249 56793 147367
rect 56911 147249 74793 147367
rect 74911 147249 92793 147367
rect 92911 147249 110793 147367
rect 110911 147249 128793 147367
rect 128911 147249 146793 147367
rect 146911 147249 164793 147367
rect 164911 147249 182793 147367
rect 182911 147249 200793 147367
rect 200911 147249 218793 147367
rect 218911 147249 236793 147367
rect 236911 147249 254793 147367
rect 254911 147249 272793 147367
rect 272911 147249 290793 147367
rect 290911 147249 293691 147367
rect 293809 147249 294370 147367
rect -2408 147238 294370 147249
rect -1938 147237 -1638 147238
rect 2702 147237 3002 147238
rect 20702 147237 21002 147238
rect 38702 147237 39002 147238
rect 56702 147237 57002 147238
rect 74702 147237 75002 147238
rect 92702 147237 93002 147238
rect 110702 147237 111002 147238
rect 128702 147237 129002 147238
rect 146702 147237 147002 147238
rect 164702 147237 165002 147238
rect 182702 147237 183002 147238
rect 200702 147237 201002 147238
rect 218702 147237 219002 147238
rect 236702 147237 237002 147238
rect 254702 147237 255002 147238
rect 272702 147237 273002 147238
rect 290702 147237 291002 147238
rect 293600 147237 293900 147238
rect -998 145738 -698 145739
rect 902 145738 1202 145739
rect 18902 145738 19202 145739
rect 36902 145738 37202 145739
rect 54902 145738 55202 145739
rect 72902 145738 73202 145739
rect 90902 145738 91202 145739
rect 108902 145738 109202 145739
rect 126902 145738 127202 145739
rect 144902 145738 145202 145739
rect 162902 145738 163202 145739
rect 180902 145738 181202 145739
rect 198902 145738 199202 145739
rect 216902 145738 217202 145739
rect 234902 145738 235202 145739
rect 252902 145738 253202 145739
rect 270902 145738 271202 145739
rect 288902 145738 289202 145739
rect 292660 145738 292960 145739
rect -1468 145727 293430 145738
rect -1468 145609 -907 145727
rect -789 145609 993 145727
rect 1111 145609 18993 145727
rect 19111 145609 36993 145727
rect 37111 145609 54993 145727
rect 55111 145609 72993 145727
rect 73111 145609 90993 145727
rect 91111 145609 108993 145727
rect 109111 145609 126993 145727
rect 127111 145609 144993 145727
rect 145111 145609 162993 145727
rect 163111 145609 180993 145727
rect 181111 145609 198993 145727
rect 199111 145609 216993 145727
rect 217111 145609 234993 145727
rect 235111 145609 252993 145727
rect 253111 145609 270993 145727
rect 271111 145609 288993 145727
rect 289111 145609 292751 145727
rect 292869 145609 293430 145727
rect -1468 145567 293430 145609
rect -1468 145449 -907 145567
rect -789 145449 993 145567
rect 1111 145449 18993 145567
rect 19111 145449 36993 145567
rect 37111 145449 54993 145567
rect 55111 145449 72993 145567
rect 73111 145449 90993 145567
rect 91111 145449 108993 145567
rect 109111 145449 126993 145567
rect 127111 145449 144993 145567
rect 145111 145449 162993 145567
rect 163111 145449 180993 145567
rect 181111 145449 198993 145567
rect 199111 145449 216993 145567
rect 217111 145449 234993 145567
rect 235111 145449 252993 145567
rect 253111 145449 270993 145567
rect 271111 145449 288993 145567
rect 289111 145449 292751 145567
rect 292869 145449 293430 145567
rect -1468 145438 293430 145449
rect -998 145437 -698 145438
rect 902 145437 1202 145438
rect 18902 145437 19202 145438
rect 36902 145437 37202 145438
rect 54902 145437 55202 145438
rect 72902 145437 73202 145438
rect 90902 145437 91202 145438
rect 108902 145437 109202 145438
rect 126902 145437 127202 145438
rect 144902 145437 145202 145438
rect 162902 145437 163202 145438
rect 180902 145437 181202 145438
rect 198902 145437 199202 145438
rect 216902 145437 217202 145438
rect 234902 145437 235202 145438
rect 252902 145437 253202 145438
rect 270902 145437 271202 145438
rect 288902 145437 289202 145438
rect 292660 145437 292960 145438
rect -4288 142138 -3988 142139
rect 15302 142138 15602 142139
rect 33302 142138 33602 142139
rect 51302 142138 51602 142139
rect 69302 142138 69602 142139
rect 87302 142138 87602 142139
rect 105302 142138 105602 142139
rect 123302 142138 123602 142139
rect 141302 142138 141602 142139
rect 159302 142138 159602 142139
rect 177302 142138 177602 142139
rect 195302 142138 195602 142139
rect 213302 142138 213602 142139
rect 231302 142138 231602 142139
rect 249302 142138 249602 142139
rect 267302 142138 267602 142139
rect 285302 142138 285602 142139
rect 295950 142138 296250 142139
rect -4288 142127 296250 142138
rect -4288 142009 -4197 142127
rect -4079 142009 15393 142127
rect 15511 142009 33393 142127
rect 33511 142009 51393 142127
rect 51511 142009 69393 142127
rect 69511 142009 87393 142127
rect 87511 142009 105393 142127
rect 105511 142009 123393 142127
rect 123511 142009 141393 142127
rect 141511 142009 159393 142127
rect 159511 142009 177393 142127
rect 177511 142009 195393 142127
rect 195511 142009 213393 142127
rect 213511 142009 231393 142127
rect 231511 142009 249393 142127
rect 249511 142009 267393 142127
rect 267511 142009 285393 142127
rect 285511 142009 296041 142127
rect 296159 142009 296250 142127
rect -4288 141967 296250 142009
rect -4288 141849 -4197 141967
rect -4079 141849 15393 141967
rect 15511 141849 33393 141967
rect 33511 141849 51393 141967
rect 51511 141849 69393 141967
rect 69511 141849 87393 141967
rect 87511 141849 105393 141967
rect 105511 141849 123393 141967
rect 123511 141849 141393 141967
rect 141511 141849 159393 141967
rect 159511 141849 177393 141967
rect 177511 141849 195393 141967
rect 195511 141849 213393 141967
rect 213511 141849 231393 141967
rect 231511 141849 249393 141967
rect 249511 141849 267393 141967
rect 267511 141849 285393 141967
rect 285511 141849 296041 141967
rect 296159 141849 296250 141967
rect -4288 141838 296250 141849
rect -4288 141837 -3988 141838
rect 15302 141837 15602 141838
rect 33302 141837 33602 141838
rect 51302 141837 51602 141838
rect 69302 141837 69602 141838
rect 87302 141837 87602 141838
rect 105302 141837 105602 141838
rect 123302 141837 123602 141838
rect 141302 141837 141602 141838
rect 159302 141837 159602 141838
rect 177302 141837 177602 141838
rect 195302 141837 195602 141838
rect 213302 141837 213602 141838
rect 231302 141837 231602 141838
rect 249302 141837 249602 141838
rect 267302 141837 267602 141838
rect 285302 141837 285602 141838
rect 295950 141837 296250 141838
rect -3348 140338 -3048 140339
rect 13502 140338 13802 140339
rect 31502 140338 31802 140339
rect 49502 140338 49802 140339
rect 67502 140338 67802 140339
rect 85502 140338 85802 140339
rect 103502 140338 103802 140339
rect 121502 140338 121802 140339
rect 139502 140338 139802 140339
rect 157502 140338 157802 140339
rect 175502 140338 175802 140339
rect 193502 140338 193802 140339
rect 211502 140338 211802 140339
rect 229502 140338 229802 140339
rect 247502 140338 247802 140339
rect 265502 140338 265802 140339
rect 283502 140338 283802 140339
rect 295010 140338 295310 140339
rect -3348 140327 295310 140338
rect -3348 140209 -3257 140327
rect -3139 140209 13593 140327
rect 13711 140209 31593 140327
rect 31711 140209 49593 140327
rect 49711 140209 67593 140327
rect 67711 140209 85593 140327
rect 85711 140209 103593 140327
rect 103711 140209 121593 140327
rect 121711 140209 139593 140327
rect 139711 140209 157593 140327
rect 157711 140209 175593 140327
rect 175711 140209 193593 140327
rect 193711 140209 211593 140327
rect 211711 140209 229593 140327
rect 229711 140209 247593 140327
rect 247711 140209 265593 140327
rect 265711 140209 283593 140327
rect 283711 140209 295101 140327
rect 295219 140209 295310 140327
rect -3348 140167 295310 140209
rect -3348 140049 -3257 140167
rect -3139 140049 13593 140167
rect 13711 140049 31593 140167
rect 31711 140049 49593 140167
rect 49711 140049 67593 140167
rect 67711 140049 85593 140167
rect 85711 140049 103593 140167
rect 103711 140049 121593 140167
rect 121711 140049 139593 140167
rect 139711 140049 157593 140167
rect 157711 140049 175593 140167
rect 175711 140049 193593 140167
rect 193711 140049 211593 140167
rect 211711 140049 229593 140167
rect 229711 140049 247593 140167
rect 247711 140049 265593 140167
rect 265711 140049 283593 140167
rect 283711 140049 295101 140167
rect 295219 140049 295310 140167
rect -3348 140038 295310 140049
rect -3348 140037 -3048 140038
rect 13502 140037 13802 140038
rect 31502 140037 31802 140038
rect 49502 140037 49802 140038
rect 67502 140037 67802 140038
rect 85502 140037 85802 140038
rect 103502 140037 103802 140038
rect 121502 140037 121802 140038
rect 139502 140037 139802 140038
rect 157502 140037 157802 140038
rect 175502 140037 175802 140038
rect 193502 140037 193802 140038
rect 211502 140037 211802 140038
rect 229502 140037 229802 140038
rect 247502 140037 247802 140038
rect 265502 140037 265802 140038
rect 283502 140037 283802 140038
rect 295010 140037 295310 140038
rect -2408 138538 -2108 138539
rect 11702 138538 12002 138539
rect 29702 138538 30002 138539
rect 47702 138538 48002 138539
rect 65702 138538 66002 138539
rect 83702 138538 84002 138539
rect 101702 138538 102002 138539
rect 119702 138538 120002 138539
rect 137702 138538 138002 138539
rect 155702 138538 156002 138539
rect 173702 138538 174002 138539
rect 191702 138538 192002 138539
rect 209702 138538 210002 138539
rect 227702 138538 228002 138539
rect 245702 138538 246002 138539
rect 263702 138538 264002 138539
rect 281702 138538 282002 138539
rect 294070 138538 294370 138539
rect -2408 138527 294370 138538
rect -2408 138409 -2317 138527
rect -2199 138409 11793 138527
rect 11911 138409 29793 138527
rect 29911 138409 47793 138527
rect 47911 138409 65793 138527
rect 65911 138409 83793 138527
rect 83911 138409 101793 138527
rect 101911 138409 119793 138527
rect 119911 138409 137793 138527
rect 137911 138409 155793 138527
rect 155911 138409 173793 138527
rect 173911 138409 191793 138527
rect 191911 138409 209793 138527
rect 209911 138409 227793 138527
rect 227911 138409 245793 138527
rect 245911 138409 263793 138527
rect 263911 138409 281793 138527
rect 281911 138409 294161 138527
rect 294279 138409 294370 138527
rect -2408 138367 294370 138409
rect -2408 138249 -2317 138367
rect -2199 138249 11793 138367
rect 11911 138249 29793 138367
rect 29911 138249 47793 138367
rect 47911 138249 65793 138367
rect 65911 138249 83793 138367
rect 83911 138249 101793 138367
rect 101911 138249 119793 138367
rect 119911 138249 137793 138367
rect 137911 138249 155793 138367
rect 155911 138249 173793 138367
rect 173911 138249 191793 138367
rect 191911 138249 209793 138367
rect 209911 138249 227793 138367
rect 227911 138249 245793 138367
rect 245911 138249 263793 138367
rect 263911 138249 281793 138367
rect 281911 138249 294161 138367
rect 294279 138249 294370 138367
rect -2408 138238 294370 138249
rect -2408 138237 -2108 138238
rect 11702 138237 12002 138238
rect 29702 138237 30002 138238
rect 47702 138237 48002 138238
rect 65702 138237 66002 138238
rect 83702 138237 84002 138238
rect 101702 138237 102002 138238
rect 119702 138237 120002 138238
rect 137702 138237 138002 138238
rect 155702 138237 156002 138238
rect 173702 138237 174002 138238
rect 191702 138237 192002 138238
rect 209702 138237 210002 138238
rect 227702 138237 228002 138238
rect 245702 138237 246002 138238
rect 263702 138237 264002 138238
rect 281702 138237 282002 138238
rect 294070 138237 294370 138238
rect -1468 136738 -1168 136739
rect 9902 136738 10202 136739
rect 27902 136738 28202 136739
rect 45902 136738 46202 136739
rect 63902 136738 64202 136739
rect 81902 136738 82202 136739
rect 99902 136738 100202 136739
rect 117902 136738 118202 136739
rect 135902 136738 136202 136739
rect 153902 136738 154202 136739
rect 171902 136738 172202 136739
rect 189902 136738 190202 136739
rect 207902 136738 208202 136739
rect 225902 136738 226202 136739
rect 243902 136738 244202 136739
rect 261902 136738 262202 136739
rect 279902 136738 280202 136739
rect 293130 136738 293430 136739
rect -1468 136727 293430 136738
rect -1468 136609 -1377 136727
rect -1259 136609 9993 136727
rect 10111 136609 27993 136727
rect 28111 136609 45993 136727
rect 46111 136609 63993 136727
rect 64111 136609 81993 136727
rect 82111 136609 99993 136727
rect 100111 136609 117993 136727
rect 118111 136609 135993 136727
rect 136111 136609 153993 136727
rect 154111 136609 171993 136727
rect 172111 136609 189993 136727
rect 190111 136609 207993 136727
rect 208111 136609 225993 136727
rect 226111 136609 243993 136727
rect 244111 136609 261993 136727
rect 262111 136609 279993 136727
rect 280111 136609 293221 136727
rect 293339 136609 293430 136727
rect -1468 136567 293430 136609
rect -1468 136449 -1377 136567
rect -1259 136449 9993 136567
rect 10111 136449 27993 136567
rect 28111 136449 45993 136567
rect 46111 136449 63993 136567
rect 64111 136449 81993 136567
rect 82111 136449 99993 136567
rect 100111 136449 117993 136567
rect 118111 136449 135993 136567
rect 136111 136449 153993 136567
rect 154111 136449 171993 136567
rect 172111 136449 189993 136567
rect 190111 136449 207993 136567
rect 208111 136449 225993 136567
rect 226111 136449 243993 136567
rect 244111 136449 261993 136567
rect 262111 136449 279993 136567
rect 280111 136449 293221 136567
rect 293339 136449 293430 136567
rect -1468 136438 293430 136449
rect -1468 136437 -1168 136438
rect 9902 136437 10202 136438
rect 27902 136437 28202 136438
rect 45902 136437 46202 136438
rect 63902 136437 64202 136438
rect 81902 136437 82202 136438
rect 99902 136437 100202 136438
rect 117902 136437 118202 136438
rect 135902 136437 136202 136438
rect 153902 136437 154202 136438
rect 171902 136437 172202 136438
rect 189902 136437 190202 136438
rect 207902 136437 208202 136438
rect 225902 136437 226202 136438
rect 243902 136437 244202 136438
rect 261902 136437 262202 136438
rect 279902 136437 280202 136438
rect 293130 136437 293430 136438
rect -3818 133138 -3518 133139
rect 6302 133138 6602 133139
rect 24302 133138 24602 133139
rect 42302 133138 42602 133139
rect 60302 133138 60602 133139
rect 78302 133138 78602 133139
rect 96302 133138 96602 133139
rect 114302 133138 114602 133139
rect 132302 133138 132602 133139
rect 150302 133138 150602 133139
rect 168302 133138 168602 133139
rect 186302 133138 186602 133139
rect 204302 133138 204602 133139
rect 222302 133138 222602 133139
rect 240302 133138 240602 133139
rect 258302 133138 258602 133139
rect 276302 133138 276602 133139
rect 295480 133138 295780 133139
rect -4288 133127 296250 133138
rect -4288 133009 -3727 133127
rect -3609 133009 6393 133127
rect 6511 133009 24393 133127
rect 24511 133009 42393 133127
rect 42511 133009 60393 133127
rect 60511 133009 78393 133127
rect 78511 133009 96393 133127
rect 96511 133009 114393 133127
rect 114511 133009 132393 133127
rect 132511 133009 150393 133127
rect 150511 133009 168393 133127
rect 168511 133009 186393 133127
rect 186511 133009 204393 133127
rect 204511 133009 222393 133127
rect 222511 133009 240393 133127
rect 240511 133009 258393 133127
rect 258511 133009 276393 133127
rect 276511 133009 295571 133127
rect 295689 133009 296250 133127
rect -4288 132967 296250 133009
rect -4288 132849 -3727 132967
rect -3609 132849 6393 132967
rect 6511 132849 24393 132967
rect 24511 132849 42393 132967
rect 42511 132849 60393 132967
rect 60511 132849 78393 132967
rect 78511 132849 96393 132967
rect 96511 132849 114393 132967
rect 114511 132849 132393 132967
rect 132511 132849 150393 132967
rect 150511 132849 168393 132967
rect 168511 132849 186393 132967
rect 186511 132849 204393 132967
rect 204511 132849 222393 132967
rect 222511 132849 240393 132967
rect 240511 132849 258393 132967
rect 258511 132849 276393 132967
rect 276511 132849 295571 132967
rect 295689 132849 296250 132967
rect -4288 132838 296250 132849
rect -3818 132837 -3518 132838
rect 6302 132837 6602 132838
rect 24302 132837 24602 132838
rect 42302 132837 42602 132838
rect 60302 132837 60602 132838
rect 78302 132837 78602 132838
rect 96302 132837 96602 132838
rect 114302 132837 114602 132838
rect 132302 132837 132602 132838
rect 150302 132837 150602 132838
rect 168302 132837 168602 132838
rect 186302 132837 186602 132838
rect 204302 132837 204602 132838
rect 222302 132837 222602 132838
rect 240302 132837 240602 132838
rect 258302 132837 258602 132838
rect 276302 132837 276602 132838
rect 295480 132837 295780 132838
rect -2878 131338 -2578 131339
rect 4502 131338 4802 131339
rect 22502 131338 22802 131339
rect 40502 131338 40802 131339
rect 58502 131338 58802 131339
rect 76502 131338 76802 131339
rect 94502 131338 94802 131339
rect 112502 131338 112802 131339
rect 130502 131338 130802 131339
rect 148502 131338 148802 131339
rect 166502 131338 166802 131339
rect 184502 131338 184802 131339
rect 202502 131338 202802 131339
rect 220502 131338 220802 131339
rect 238502 131338 238802 131339
rect 256502 131338 256802 131339
rect 274502 131338 274802 131339
rect 294540 131338 294840 131339
rect -3348 131327 295310 131338
rect -3348 131209 -2787 131327
rect -2669 131209 4593 131327
rect 4711 131209 22593 131327
rect 22711 131209 40593 131327
rect 40711 131209 58593 131327
rect 58711 131209 76593 131327
rect 76711 131209 94593 131327
rect 94711 131209 112593 131327
rect 112711 131209 130593 131327
rect 130711 131209 148593 131327
rect 148711 131209 166593 131327
rect 166711 131209 184593 131327
rect 184711 131209 202593 131327
rect 202711 131209 220593 131327
rect 220711 131209 238593 131327
rect 238711 131209 256593 131327
rect 256711 131209 274593 131327
rect 274711 131209 294631 131327
rect 294749 131209 295310 131327
rect -3348 131167 295310 131209
rect -3348 131049 -2787 131167
rect -2669 131049 4593 131167
rect 4711 131049 22593 131167
rect 22711 131049 40593 131167
rect 40711 131049 58593 131167
rect 58711 131049 76593 131167
rect 76711 131049 94593 131167
rect 94711 131049 112593 131167
rect 112711 131049 130593 131167
rect 130711 131049 148593 131167
rect 148711 131049 166593 131167
rect 166711 131049 184593 131167
rect 184711 131049 202593 131167
rect 202711 131049 220593 131167
rect 220711 131049 238593 131167
rect 238711 131049 256593 131167
rect 256711 131049 274593 131167
rect 274711 131049 294631 131167
rect 294749 131049 295310 131167
rect -3348 131038 295310 131049
rect -2878 131037 -2578 131038
rect 4502 131037 4802 131038
rect 22502 131037 22802 131038
rect 40502 131037 40802 131038
rect 58502 131037 58802 131038
rect 76502 131037 76802 131038
rect 94502 131037 94802 131038
rect 112502 131037 112802 131038
rect 130502 131037 130802 131038
rect 148502 131037 148802 131038
rect 166502 131037 166802 131038
rect 184502 131037 184802 131038
rect 202502 131037 202802 131038
rect 220502 131037 220802 131038
rect 238502 131037 238802 131038
rect 256502 131037 256802 131038
rect 274502 131037 274802 131038
rect 294540 131037 294840 131038
rect -1938 129538 -1638 129539
rect 2702 129538 3002 129539
rect 20702 129538 21002 129539
rect 38702 129538 39002 129539
rect 56702 129538 57002 129539
rect 74702 129538 75002 129539
rect 92702 129538 93002 129539
rect 110702 129538 111002 129539
rect 128702 129538 129002 129539
rect 146702 129538 147002 129539
rect 164702 129538 165002 129539
rect 182702 129538 183002 129539
rect 200702 129538 201002 129539
rect 218702 129538 219002 129539
rect 236702 129538 237002 129539
rect 254702 129538 255002 129539
rect 272702 129538 273002 129539
rect 290702 129538 291002 129539
rect 293600 129538 293900 129539
rect -2408 129527 294370 129538
rect -2408 129409 -1847 129527
rect -1729 129409 2793 129527
rect 2911 129409 20793 129527
rect 20911 129409 38793 129527
rect 38911 129409 56793 129527
rect 56911 129409 74793 129527
rect 74911 129409 92793 129527
rect 92911 129409 110793 129527
rect 110911 129409 128793 129527
rect 128911 129409 146793 129527
rect 146911 129409 164793 129527
rect 164911 129409 182793 129527
rect 182911 129409 200793 129527
rect 200911 129409 218793 129527
rect 218911 129409 236793 129527
rect 236911 129409 254793 129527
rect 254911 129409 272793 129527
rect 272911 129409 290793 129527
rect 290911 129409 293691 129527
rect 293809 129409 294370 129527
rect -2408 129367 294370 129409
rect -2408 129249 -1847 129367
rect -1729 129249 2793 129367
rect 2911 129249 20793 129367
rect 20911 129249 38793 129367
rect 38911 129249 56793 129367
rect 56911 129249 74793 129367
rect 74911 129249 92793 129367
rect 92911 129249 110793 129367
rect 110911 129249 128793 129367
rect 128911 129249 146793 129367
rect 146911 129249 164793 129367
rect 164911 129249 182793 129367
rect 182911 129249 200793 129367
rect 200911 129249 218793 129367
rect 218911 129249 236793 129367
rect 236911 129249 254793 129367
rect 254911 129249 272793 129367
rect 272911 129249 290793 129367
rect 290911 129249 293691 129367
rect 293809 129249 294370 129367
rect -2408 129238 294370 129249
rect -1938 129237 -1638 129238
rect 2702 129237 3002 129238
rect 20702 129237 21002 129238
rect 38702 129237 39002 129238
rect 56702 129237 57002 129238
rect 74702 129237 75002 129238
rect 92702 129237 93002 129238
rect 110702 129237 111002 129238
rect 128702 129237 129002 129238
rect 146702 129237 147002 129238
rect 164702 129237 165002 129238
rect 182702 129237 183002 129238
rect 200702 129237 201002 129238
rect 218702 129237 219002 129238
rect 236702 129237 237002 129238
rect 254702 129237 255002 129238
rect 272702 129237 273002 129238
rect 290702 129237 291002 129238
rect 293600 129237 293900 129238
rect -998 127738 -698 127739
rect 902 127738 1202 127739
rect 18902 127738 19202 127739
rect 36902 127738 37202 127739
rect 54902 127738 55202 127739
rect 72902 127738 73202 127739
rect 90902 127738 91202 127739
rect 108902 127738 109202 127739
rect 126902 127738 127202 127739
rect 144902 127738 145202 127739
rect 162902 127738 163202 127739
rect 180902 127738 181202 127739
rect 198902 127738 199202 127739
rect 216902 127738 217202 127739
rect 234902 127738 235202 127739
rect 252902 127738 253202 127739
rect 270902 127738 271202 127739
rect 288902 127738 289202 127739
rect 292660 127738 292960 127739
rect -1468 127727 293430 127738
rect -1468 127609 -907 127727
rect -789 127609 993 127727
rect 1111 127609 18993 127727
rect 19111 127609 36993 127727
rect 37111 127609 54993 127727
rect 55111 127609 72993 127727
rect 73111 127609 90993 127727
rect 91111 127609 108993 127727
rect 109111 127609 126993 127727
rect 127111 127609 144993 127727
rect 145111 127609 162993 127727
rect 163111 127609 180993 127727
rect 181111 127609 198993 127727
rect 199111 127609 216993 127727
rect 217111 127609 234993 127727
rect 235111 127609 252993 127727
rect 253111 127609 270993 127727
rect 271111 127609 288993 127727
rect 289111 127609 292751 127727
rect 292869 127609 293430 127727
rect -1468 127567 293430 127609
rect -1468 127449 -907 127567
rect -789 127449 993 127567
rect 1111 127449 18993 127567
rect 19111 127449 36993 127567
rect 37111 127449 54993 127567
rect 55111 127449 72993 127567
rect 73111 127449 90993 127567
rect 91111 127449 108993 127567
rect 109111 127449 126993 127567
rect 127111 127449 144993 127567
rect 145111 127449 162993 127567
rect 163111 127449 180993 127567
rect 181111 127449 198993 127567
rect 199111 127449 216993 127567
rect 217111 127449 234993 127567
rect 235111 127449 252993 127567
rect 253111 127449 270993 127567
rect 271111 127449 288993 127567
rect 289111 127449 292751 127567
rect 292869 127449 293430 127567
rect -1468 127438 293430 127449
rect -998 127437 -698 127438
rect 902 127437 1202 127438
rect 18902 127437 19202 127438
rect 36902 127437 37202 127438
rect 54902 127437 55202 127438
rect 72902 127437 73202 127438
rect 90902 127437 91202 127438
rect 108902 127437 109202 127438
rect 126902 127437 127202 127438
rect 144902 127437 145202 127438
rect 162902 127437 163202 127438
rect 180902 127437 181202 127438
rect 198902 127437 199202 127438
rect 216902 127437 217202 127438
rect 234902 127437 235202 127438
rect 252902 127437 253202 127438
rect 270902 127437 271202 127438
rect 288902 127437 289202 127438
rect 292660 127437 292960 127438
rect -4288 124138 -3988 124139
rect 15302 124138 15602 124139
rect 33302 124138 33602 124139
rect 51302 124138 51602 124139
rect 69302 124138 69602 124139
rect 87302 124138 87602 124139
rect 105302 124138 105602 124139
rect 123302 124138 123602 124139
rect 141302 124138 141602 124139
rect 159302 124138 159602 124139
rect 177302 124138 177602 124139
rect 195302 124138 195602 124139
rect 213302 124138 213602 124139
rect 231302 124138 231602 124139
rect 249302 124138 249602 124139
rect 267302 124138 267602 124139
rect 285302 124138 285602 124139
rect 295950 124138 296250 124139
rect -4288 124127 296250 124138
rect -4288 124009 -4197 124127
rect -4079 124009 15393 124127
rect 15511 124009 33393 124127
rect 33511 124009 51393 124127
rect 51511 124009 69393 124127
rect 69511 124009 87393 124127
rect 87511 124009 105393 124127
rect 105511 124009 123393 124127
rect 123511 124009 141393 124127
rect 141511 124009 159393 124127
rect 159511 124009 177393 124127
rect 177511 124009 195393 124127
rect 195511 124009 213393 124127
rect 213511 124009 231393 124127
rect 231511 124009 249393 124127
rect 249511 124009 267393 124127
rect 267511 124009 285393 124127
rect 285511 124009 296041 124127
rect 296159 124009 296250 124127
rect -4288 123967 296250 124009
rect -4288 123849 -4197 123967
rect -4079 123849 15393 123967
rect 15511 123849 33393 123967
rect 33511 123849 51393 123967
rect 51511 123849 69393 123967
rect 69511 123849 87393 123967
rect 87511 123849 105393 123967
rect 105511 123849 123393 123967
rect 123511 123849 141393 123967
rect 141511 123849 159393 123967
rect 159511 123849 177393 123967
rect 177511 123849 195393 123967
rect 195511 123849 213393 123967
rect 213511 123849 231393 123967
rect 231511 123849 249393 123967
rect 249511 123849 267393 123967
rect 267511 123849 285393 123967
rect 285511 123849 296041 123967
rect 296159 123849 296250 123967
rect -4288 123838 296250 123849
rect -4288 123837 -3988 123838
rect 15302 123837 15602 123838
rect 33302 123837 33602 123838
rect 51302 123837 51602 123838
rect 69302 123837 69602 123838
rect 87302 123837 87602 123838
rect 105302 123837 105602 123838
rect 123302 123837 123602 123838
rect 141302 123837 141602 123838
rect 159302 123837 159602 123838
rect 177302 123837 177602 123838
rect 195302 123837 195602 123838
rect 213302 123837 213602 123838
rect 231302 123837 231602 123838
rect 249302 123837 249602 123838
rect 267302 123837 267602 123838
rect 285302 123837 285602 123838
rect 295950 123837 296250 123838
rect -3348 122338 -3048 122339
rect 13502 122338 13802 122339
rect 31502 122338 31802 122339
rect 49502 122338 49802 122339
rect 67502 122338 67802 122339
rect 85502 122338 85802 122339
rect 103502 122338 103802 122339
rect 121502 122338 121802 122339
rect 139502 122338 139802 122339
rect 157502 122338 157802 122339
rect 175502 122338 175802 122339
rect 193502 122338 193802 122339
rect 211502 122338 211802 122339
rect 229502 122338 229802 122339
rect 247502 122338 247802 122339
rect 265502 122338 265802 122339
rect 283502 122338 283802 122339
rect 295010 122338 295310 122339
rect -3348 122327 295310 122338
rect -3348 122209 -3257 122327
rect -3139 122209 13593 122327
rect 13711 122209 31593 122327
rect 31711 122209 49593 122327
rect 49711 122209 67593 122327
rect 67711 122209 85593 122327
rect 85711 122209 103593 122327
rect 103711 122209 121593 122327
rect 121711 122209 139593 122327
rect 139711 122209 157593 122327
rect 157711 122209 175593 122327
rect 175711 122209 193593 122327
rect 193711 122209 211593 122327
rect 211711 122209 229593 122327
rect 229711 122209 247593 122327
rect 247711 122209 265593 122327
rect 265711 122209 283593 122327
rect 283711 122209 295101 122327
rect 295219 122209 295310 122327
rect -3348 122167 295310 122209
rect -3348 122049 -3257 122167
rect -3139 122049 13593 122167
rect 13711 122049 31593 122167
rect 31711 122049 49593 122167
rect 49711 122049 67593 122167
rect 67711 122049 85593 122167
rect 85711 122049 103593 122167
rect 103711 122049 121593 122167
rect 121711 122049 139593 122167
rect 139711 122049 157593 122167
rect 157711 122049 175593 122167
rect 175711 122049 193593 122167
rect 193711 122049 211593 122167
rect 211711 122049 229593 122167
rect 229711 122049 247593 122167
rect 247711 122049 265593 122167
rect 265711 122049 283593 122167
rect 283711 122049 295101 122167
rect 295219 122049 295310 122167
rect -3348 122038 295310 122049
rect -3348 122037 -3048 122038
rect 13502 122037 13802 122038
rect 31502 122037 31802 122038
rect 49502 122037 49802 122038
rect 67502 122037 67802 122038
rect 85502 122037 85802 122038
rect 103502 122037 103802 122038
rect 121502 122037 121802 122038
rect 139502 122037 139802 122038
rect 157502 122037 157802 122038
rect 175502 122037 175802 122038
rect 193502 122037 193802 122038
rect 211502 122037 211802 122038
rect 229502 122037 229802 122038
rect 247502 122037 247802 122038
rect 265502 122037 265802 122038
rect 283502 122037 283802 122038
rect 295010 122037 295310 122038
rect -2408 120538 -2108 120539
rect 11702 120538 12002 120539
rect 29702 120538 30002 120539
rect 47702 120538 48002 120539
rect 65702 120538 66002 120539
rect 83702 120538 84002 120539
rect 101702 120538 102002 120539
rect 119702 120538 120002 120539
rect 137702 120538 138002 120539
rect 155702 120538 156002 120539
rect 173702 120538 174002 120539
rect 191702 120538 192002 120539
rect 209702 120538 210002 120539
rect 227702 120538 228002 120539
rect 245702 120538 246002 120539
rect 263702 120538 264002 120539
rect 281702 120538 282002 120539
rect 294070 120538 294370 120539
rect -2408 120527 294370 120538
rect -2408 120409 -2317 120527
rect -2199 120409 11793 120527
rect 11911 120409 29793 120527
rect 29911 120409 47793 120527
rect 47911 120409 65793 120527
rect 65911 120409 83793 120527
rect 83911 120409 101793 120527
rect 101911 120409 119793 120527
rect 119911 120409 137793 120527
rect 137911 120409 155793 120527
rect 155911 120409 173793 120527
rect 173911 120409 191793 120527
rect 191911 120409 209793 120527
rect 209911 120409 227793 120527
rect 227911 120409 245793 120527
rect 245911 120409 263793 120527
rect 263911 120409 281793 120527
rect 281911 120409 294161 120527
rect 294279 120409 294370 120527
rect -2408 120367 294370 120409
rect -2408 120249 -2317 120367
rect -2199 120249 11793 120367
rect 11911 120249 29793 120367
rect 29911 120249 47793 120367
rect 47911 120249 65793 120367
rect 65911 120249 83793 120367
rect 83911 120249 101793 120367
rect 101911 120249 119793 120367
rect 119911 120249 137793 120367
rect 137911 120249 155793 120367
rect 155911 120249 173793 120367
rect 173911 120249 191793 120367
rect 191911 120249 209793 120367
rect 209911 120249 227793 120367
rect 227911 120249 245793 120367
rect 245911 120249 263793 120367
rect 263911 120249 281793 120367
rect 281911 120249 294161 120367
rect 294279 120249 294370 120367
rect -2408 120238 294370 120249
rect -2408 120237 -2108 120238
rect 11702 120237 12002 120238
rect 29702 120237 30002 120238
rect 47702 120237 48002 120238
rect 65702 120237 66002 120238
rect 83702 120237 84002 120238
rect 101702 120237 102002 120238
rect 119702 120237 120002 120238
rect 137702 120237 138002 120238
rect 155702 120237 156002 120238
rect 173702 120237 174002 120238
rect 191702 120237 192002 120238
rect 209702 120237 210002 120238
rect 227702 120237 228002 120238
rect 245702 120237 246002 120238
rect 263702 120237 264002 120238
rect 281702 120237 282002 120238
rect 294070 120237 294370 120238
rect -1468 118738 -1168 118739
rect 9902 118738 10202 118739
rect 27902 118738 28202 118739
rect 45902 118738 46202 118739
rect 63902 118738 64202 118739
rect 81902 118738 82202 118739
rect 99902 118738 100202 118739
rect 117902 118738 118202 118739
rect 135902 118738 136202 118739
rect 153902 118738 154202 118739
rect 171902 118738 172202 118739
rect 189902 118738 190202 118739
rect 207902 118738 208202 118739
rect 225902 118738 226202 118739
rect 243902 118738 244202 118739
rect 261902 118738 262202 118739
rect 279902 118738 280202 118739
rect 293130 118738 293430 118739
rect -1468 118727 293430 118738
rect -1468 118609 -1377 118727
rect -1259 118609 9993 118727
rect 10111 118609 27993 118727
rect 28111 118609 45993 118727
rect 46111 118609 63993 118727
rect 64111 118609 81993 118727
rect 82111 118609 99993 118727
rect 100111 118609 117993 118727
rect 118111 118609 135993 118727
rect 136111 118609 153993 118727
rect 154111 118609 171993 118727
rect 172111 118609 189993 118727
rect 190111 118609 207993 118727
rect 208111 118609 225993 118727
rect 226111 118609 243993 118727
rect 244111 118609 261993 118727
rect 262111 118609 279993 118727
rect 280111 118609 293221 118727
rect 293339 118609 293430 118727
rect -1468 118567 293430 118609
rect -1468 118449 -1377 118567
rect -1259 118449 9993 118567
rect 10111 118449 27993 118567
rect 28111 118449 45993 118567
rect 46111 118449 63993 118567
rect 64111 118449 81993 118567
rect 82111 118449 99993 118567
rect 100111 118449 117993 118567
rect 118111 118449 135993 118567
rect 136111 118449 153993 118567
rect 154111 118449 171993 118567
rect 172111 118449 189993 118567
rect 190111 118449 207993 118567
rect 208111 118449 225993 118567
rect 226111 118449 243993 118567
rect 244111 118449 261993 118567
rect 262111 118449 279993 118567
rect 280111 118449 293221 118567
rect 293339 118449 293430 118567
rect -1468 118438 293430 118449
rect -1468 118437 -1168 118438
rect 9902 118437 10202 118438
rect 27902 118437 28202 118438
rect 45902 118437 46202 118438
rect 63902 118437 64202 118438
rect 81902 118437 82202 118438
rect 99902 118437 100202 118438
rect 117902 118437 118202 118438
rect 135902 118437 136202 118438
rect 153902 118437 154202 118438
rect 171902 118437 172202 118438
rect 189902 118437 190202 118438
rect 207902 118437 208202 118438
rect 225902 118437 226202 118438
rect 243902 118437 244202 118438
rect 261902 118437 262202 118438
rect 279902 118437 280202 118438
rect 293130 118437 293430 118438
rect -3818 115138 -3518 115139
rect 6302 115138 6602 115139
rect 24302 115138 24602 115139
rect 42302 115138 42602 115139
rect 60302 115138 60602 115139
rect 78302 115138 78602 115139
rect 96302 115138 96602 115139
rect 114302 115138 114602 115139
rect 132302 115138 132602 115139
rect 150302 115138 150602 115139
rect 168302 115138 168602 115139
rect 186302 115138 186602 115139
rect 204302 115138 204602 115139
rect 222302 115138 222602 115139
rect 240302 115138 240602 115139
rect 258302 115138 258602 115139
rect 276302 115138 276602 115139
rect 295480 115138 295780 115139
rect -4288 115127 296250 115138
rect -4288 115009 -3727 115127
rect -3609 115009 6393 115127
rect 6511 115009 24393 115127
rect 24511 115009 42393 115127
rect 42511 115009 60393 115127
rect 60511 115009 78393 115127
rect 78511 115009 96393 115127
rect 96511 115009 114393 115127
rect 114511 115009 132393 115127
rect 132511 115009 150393 115127
rect 150511 115009 168393 115127
rect 168511 115009 186393 115127
rect 186511 115009 204393 115127
rect 204511 115009 222393 115127
rect 222511 115009 240393 115127
rect 240511 115009 258393 115127
rect 258511 115009 276393 115127
rect 276511 115009 295571 115127
rect 295689 115009 296250 115127
rect -4288 114967 296250 115009
rect -4288 114849 -3727 114967
rect -3609 114849 6393 114967
rect 6511 114849 24393 114967
rect 24511 114849 42393 114967
rect 42511 114849 60393 114967
rect 60511 114849 78393 114967
rect 78511 114849 96393 114967
rect 96511 114849 114393 114967
rect 114511 114849 132393 114967
rect 132511 114849 150393 114967
rect 150511 114849 168393 114967
rect 168511 114849 186393 114967
rect 186511 114849 204393 114967
rect 204511 114849 222393 114967
rect 222511 114849 240393 114967
rect 240511 114849 258393 114967
rect 258511 114849 276393 114967
rect 276511 114849 295571 114967
rect 295689 114849 296250 114967
rect -4288 114838 296250 114849
rect -3818 114837 -3518 114838
rect 6302 114837 6602 114838
rect 24302 114837 24602 114838
rect 42302 114837 42602 114838
rect 60302 114837 60602 114838
rect 78302 114837 78602 114838
rect 96302 114837 96602 114838
rect 114302 114837 114602 114838
rect 132302 114837 132602 114838
rect 150302 114837 150602 114838
rect 168302 114837 168602 114838
rect 186302 114837 186602 114838
rect 204302 114837 204602 114838
rect 222302 114837 222602 114838
rect 240302 114837 240602 114838
rect 258302 114837 258602 114838
rect 276302 114837 276602 114838
rect 295480 114837 295780 114838
rect -2878 113338 -2578 113339
rect 4502 113338 4802 113339
rect 22502 113338 22802 113339
rect 40502 113338 40802 113339
rect 58502 113338 58802 113339
rect 76502 113338 76802 113339
rect 94502 113338 94802 113339
rect 112502 113338 112802 113339
rect 130502 113338 130802 113339
rect 148502 113338 148802 113339
rect 166502 113338 166802 113339
rect 184502 113338 184802 113339
rect 202502 113338 202802 113339
rect 220502 113338 220802 113339
rect 238502 113338 238802 113339
rect 256502 113338 256802 113339
rect 274502 113338 274802 113339
rect 294540 113338 294840 113339
rect -3348 113327 295310 113338
rect -3348 113209 -2787 113327
rect -2669 113209 4593 113327
rect 4711 113209 22593 113327
rect 22711 113209 40593 113327
rect 40711 113209 58593 113327
rect 58711 113209 76593 113327
rect 76711 113209 94593 113327
rect 94711 113209 112593 113327
rect 112711 113209 130593 113327
rect 130711 113209 148593 113327
rect 148711 113209 166593 113327
rect 166711 113209 184593 113327
rect 184711 113209 202593 113327
rect 202711 113209 220593 113327
rect 220711 113209 238593 113327
rect 238711 113209 256593 113327
rect 256711 113209 274593 113327
rect 274711 113209 294631 113327
rect 294749 113209 295310 113327
rect -3348 113167 295310 113209
rect -3348 113049 -2787 113167
rect -2669 113049 4593 113167
rect 4711 113049 22593 113167
rect 22711 113049 40593 113167
rect 40711 113049 58593 113167
rect 58711 113049 76593 113167
rect 76711 113049 94593 113167
rect 94711 113049 112593 113167
rect 112711 113049 130593 113167
rect 130711 113049 148593 113167
rect 148711 113049 166593 113167
rect 166711 113049 184593 113167
rect 184711 113049 202593 113167
rect 202711 113049 220593 113167
rect 220711 113049 238593 113167
rect 238711 113049 256593 113167
rect 256711 113049 274593 113167
rect 274711 113049 294631 113167
rect 294749 113049 295310 113167
rect -3348 113038 295310 113049
rect -2878 113037 -2578 113038
rect 4502 113037 4802 113038
rect 22502 113037 22802 113038
rect 40502 113037 40802 113038
rect 58502 113037 58802 113038
rect 76502 113037 76802 113038
rect 94502 113037 94802 113038
rect 112502 113037 112802 113038
rect 130502 113037 130802 113038
rect 148502 113037 148802 113038
rect 166502 113037 166802 113038
rect 184502 113037 184802 113038
rect 202502 113037 202802 113038
rect 220502 113037 220802 113038
rect 238502 113037 238802 113038
rect 256502 113037 256802 113038
rect 274502 113037 274802 113038
rect 294540 113037 294840 113038
rect -1938 111538 -1638 111539
rect 2702 111538 3002 111539
rect 20702 111538 21002 111539
rect 38702 111538 39002 111539
rect 56702 111538 57002 111539
rect 74702 111538 75002 111539
rect 92702 111538 93002 111539
rect 110702 111538 111002 111539
rect 128702 111538 129002 111539
rect 146702 111538 147002 111539
rect 164702 111538 165002 111539
rect 182702 111538 183002 111539
rect 200702 111538 201002 111539
rect 218702 111538 219002 111539
rect 236702 111538 237002 111539
rect 254702 111538 255002 111539
rect 272702 111538 273002 111539
rect 290702 111538 291002 111539
rect 293600 111538 293900 111539
rect -2408 111527 294370 111538
rect -2408 111409 -1847 111527
rect -1729 111409 2793 111527
rect 2911 111409 20793 111527
rect 20911 111409 38793 111527
rect 38911 111409 56793 111527
rect 56911 111409 74793 111527
rect 74911 111409 92793 111527
rect 92911 111409 110793 111527
rect 110911 111409 128793 111527
rect 128911 111409 146793 111527
rect 146911 111409 164793 111527
rect 164911 111409 182793 111527
rect 182911 111409 200793 111527
rect 200911 111409 218793 111527
rect 218911 111409 236793 111527
rect 236911 111409 254793 111527
rect 254911 111409 272793 111527
rect 272911 111409 290793 111527
rect 290911 111409 293691 111527
rect 293809 111409 294370 111527
rect -2408 111367 294370 111409
rect -2408 111249 -1847 111367
rect -1729 111249 2793 111367
rect 2911 111249 20793 111367
rect 20911 111249 38793 111367
rect 38911 111249 56793 111367
rect 56911 111249 74793 111367
rect 74911 111249 92793 111367
rect 92911 111249 110793 111367
rect 110911 111249 128793 111367
rect 128911 111249 146793 111367
rect 146911 111249 164793 111367
rect 164911 111249 182793 111367
rect 182911 111249 200793 111367
rect 200911 111249 218793 111367
rect 218911 111249 236793 111367
rect 236911 111249 254793 111367
rect 254911 111249 272793 111367
rect 272911 111249 290793 111367
rect 290911 111249 293691 111367
rect 293809 111249 294370 111367
rect -2408 111238 294370 111249
rect -1938 111237 -1638 111238
rect 2702 111237 3002 111238
rect 20702 111237 21002 111238
rect 38702 111237 39002 111238
rect 56702 111237 57002 111238
rect 74702 111237 75002 111238
rect 92702 111237 93002 111238
rect 110702 111237 111002 111238
rect 128702 111237 129002 111238
rect 146702 111237 147002 111238
rect 164702 111237 165002 111238
rect 182702 111237 183002 111238
rect 200702 111237 201002 111238
rect 218702 111237 219002 111238
rect 236702 111237 237002 111238
rect 254702 111237 255002 111238
rect 272702 111237 273002 111238
rect 290702 111237 291002 111238
rect 293600 111237 293900 111238
rect -998 109738 -698 109739
rect 902 109738 1202 109739
rect 18902 109738 19202 109739
rect 36902 109738 37202 109739
rect 54902 109738 55202 109739
rect 72902 109738 73202 109739
rect 90902 109738 91202 109739
rect 108902 109738 109202 109739
rect 126902 109738 127202 109739
rect 144902 109738 145202 109739
rect 162902 109738 163202 109739
rect 180902 109738 181202 109739
rect 198902 109738 199202 109739
rect 216902 109738 217202 109739
rect 234902 109738 235202 109739
rect 252902 109738 253202 109739
rect 270902 109738 271202 109739
rect 288902 109738 289202 109739
rect 292660 109738 292960 109739
rect -1468 109727 293430 109738
rect -1468 109609 -907 109727
rect -789 109609 993 109727
rect 1111 109609 18993 109727
rect 19111 109609 36993 109727
rect 37111 109609 54993 109727
rect 55111 109609 72993 109727
rect 73111 109609 90993 109727
rect 91111 109609 108993 109727
rect 109111 109609 126993 109727
rect 127111 109609 144993 109727
rect 145111 109609 162993 109727
rect 163111 109609 180993 109727
rect 181111 109609 198993 109727
rect 199111 109609 216993 109727
rect 217111 109609 234993 109727
rect 235111 109609 252993 109727
rect 253111 109609 270993 109727
rect 271111 109609 288993 109727
rect 289111 109609 292751 109727
rect 292869 109609 293430 109727
rect -1468 109567 293430 109609
rect -1468 109449 -907 109567
rect -789 109449 993 109567
rect 1111 109449 18993 109567
rect 19111 109449 36993 109567
rect 37111 109449 54993 109567
rect 55111 109449 72993 109567
rect 73111 109449 90993 109567
rect 91111 109449 108993 109567
rect 109111 109449 126993 109567
rect 127111 109449 144993 109567
rect 145111 109449 162993 109567
rect 163111 109449 180993 109567
rect 181111 109449 198993 109567
rect 199111 109449 216993 109567
rect 217111 109449 234993 109567
rect 235111 109449 252993 109567
rect 253111 109449 270993 109567
rect 271111 109449 288993 109567
rect 289111 109449 292751 109567
rect 292869 109449 293430 109567
rect -1468 109438 293430 109449
rect -998 109437 -698 109438
rect 902 109437 1202 109438
rect 18902 109437 19202 109438
rect 36902 109437 37202 109438
rect 54902 109437 55202 109438
rect 72902 109437 73202 109438
rect 90902 109437 91202 109438
rect 108902 109437 109202 109438
rect 126902 109437 127202 109438
rect 144902 109437 145202 109438
rect 162902 109437 163202 109438
rect 180902 109437 181202 109438
rect 198902 109437 199202 109438
rect 216902 109437 217202 109438
rect 234902 109437 235202 109438
rect 252902 109437 253202 109438
rect 270902 109437 271202 109438
rect 288902 109437 289202 109438
rect 292660 109437 292960 109438
rect -4288 106138 -3988 106139
rect 15302 106138 15602 106139
rect 33302 106138 33602 106139
rect 51302 106138 51602 106139
rect 69302 106138 69602 106139
rect 87302 106138 87602 106139
rect 105302 106138 105602 106139
rect 123302 106138 123602 106139
rect 141302 106138 141602 106139
rect 159302 106138 159602 106139
rect 177302 106138 177602 106139
rect 195302 106138 195602 106139
rect 213302 106138 213602 106139
rect 231302 106138 231602 106139
rect 249302 106138 249602 106139
rect 267302 106138 267602 106139
rect 285302 106138 285602 106139
rect 295950 106138 296250 106139
rect -4288 106127 296250 106138
rect -4288 106009 -4197 106127
rect -4079 106009 15393 106127
rect 15511 106009 33393 106127
rect 33511 106009 51393 106127
rect 51511 106009 69393 106127
rect 69511 106009 87393 106127
rect 87511 106009 105393 106127
rect 105511 106009 123393 106127
rect 123511 106009 141393 106127
rect 141511 106009 159393 106127
rect 159511 106009 177393 106127
rect 177511 106009 195393 106127
rect 195511 106009 213393 106127
rect 213511 106009 231393 106127
rect 231511 106009 249393 106127
rect 249511 106009 267393 106127
rect 267511 106009 285393 106127
rect 285511 106009 296041 106127
rect 296159 106009 296250 106127
rect -4288 105967 296250 106009
rect -4288 105849 -4197 105967
rect -4079 105849 15393 105967
rect 15511 105849 33393 105967
rect 33511 105849 51393 105967
rect 51511 105849 69393 105967
rect 69511 105849 87393 105967
rect 87511 105849 105393 105967
rect 105511 105849 123393 105967
rect 123511 105849 141393 105967
rect 141511 105849 159393 105967
rect 159511 105849 177393 105967
rect 177511 105849 195393 105967
rect 195511 105849 213393 105967
rect 213511 105849 231393 105967
rect 231511 105849 249393 105967
rect 249511 105849 267393 105967
rect 267511 105849 285393 105967
rect 285511 105849 296041 105967
rect 296159 105849 296250 105967
rect -4288 105838 296250 105849
rect -4288 105837 -3988 105838
rect 15302 105837 15602 105838
rect 33302 105837 33602 105838
rect 51302 105837 51602 105838
rect 69302 105837 69602 105838
rect 87302 105837 87602 105838
rect 105302 105837 105602 105838
rect 123302 105837 123602 105838
rect 141302 105837 141602 105838
rect 159302 105837 159602 105838
rect 177302 105837 177602 105838
rect 195302 105837 195602 105838
rect 213302 105837 213602 105838
rect 231302 105837 231602 105838
rect 249302 105837 249602 105838
rect 267302 105837 267602 105838
rect 285302 105837 285602 105838
rect 295950 105837 296250 105838
rect -3348 104338 -3048 104339
rect 13502 104338 13802 104339
rect 31502 104338 31802 104339
rect 49502 104338 49802 104339
rect 67502 104338 67802 104339
rect 85502 104338 85802 104339
rect 103502 104338 103802 104339
rect 121502 104338 121802 104339
rect 139502 104338 139802 104339
rect 157502 104338 157802 104339
rect 175502 104338 175802 104339
rect 193502 104338 193802 104339
rect 211502 104338 211802 104339
rect 229502 104338 229802 104339
rect 247502 104338 247802 104339
rect 265502 104338 265802 104339
rect 283502 104338 283802 104339
rect 295010 104338 295310 104339
rect -3348 104327 295310 104338
rect -3348 104209 -3257 104327
rect -3139 104209 13593 104327
rect 13711 104209 31593 104327
rect 31711 104209 49593 104327
rect 49711 104209 67593 104327
rect 67711 104209 85593 104327
rect 85711 104209 103593 104327
rect 103711 104209 121593 104327
rect 121711 104209 139593 104327
rect 139711 104209 157593 104327
rect 157711 104209 175593 104327
rect 175711 104209 193593 104327
rect 193711 104209 211593 104327
rect 211711 104209 229593 104327
rect 229711 104209 247593 104327
rect 247711 104209 265593 104327
rect 265711 104209 283593 104327
rect 283711 104209 295101 104327
rect 295219 104209 295310 104327
rect -3348 104167 295310 104209
rect -3348 104049 -3257 104167
rect -3139 104049 13593 104167
rect 13711 104049 31593 104167
rect 31711 104049 49593 104167
rect 49711 104049 67593 104167
rect 67711 104049 85593 104167
rect 85711 104049 103593 104167
rect 103711 104049 121593 104167
rect 121711 104049 139593 104167
rect 139711 104049 157593 104167
rect 157711 104049 175593 104167
rect 175711 104049 193593 104167
rect 193711 104049 211593 104167
rect 211711 104049 229593 104167
rect 229711 104049 247593 104167
rect 247711 104049 265593 104167
rect 265711 104049 283593 104167
rect 283711 104049 295101 104167
rect 295219 104049 295310 104167
rect -3348 104038 295310 104049
rect -3348 104037 -3048 104038
rect 13502 104037 13802 104038
rect 31502 104037 31802 104038
rect 49502 104037 49802 104038
rect 67502 104037 67802 104038
rect 85502 104037 85802 104038
rect 103502 104037 103802 104038
rect 121502 104037 121802 104038
rect 139502 104037 139802 104038
rect 157502 104037 157802 104038
rect 175502 104037 175802 104038
rect 193502 104037 193802 104038
rect 211502 104037 211802 104038
rect 229502 104037 229802 104038
rect 247502 104037 247802 104038
rect 265502 104037 265802 104038
rect 283502 104037 283802 104038
rect 295010 104037 295310 104038
rect -2408 102538 -2108 102539
rect 11702 102538 12002 102539
rect 29702 102538 30002 102539
rect 47702 102538 48002 102539
rect 65702 102538 66002 102539
rect 83702 102538 84002 102539
rect 101702 102538 102002 102539
rect 119702 102538 120002 102539
rect 137702 102538 138002 102539
rect 155702 102538 156002 102539
rect 173702 102538 174002 102539
rect 191702 102538 192002 102539
rect 209702 102538 210002 102539
rect 227702 102538 228002 102539
rect 245702 102538 246002 102539
rect 263702 102538 264002 102539
rect 281702 102538 282002 102539
rect 294070 102538 294370 102539
rect -2408 102527 294370 102538
rect -2408 102409 -2317 102527
rect -2199 102409 11793 102527
rect 11911 102409 29793 102527
rect 29911 102409 47793 102527
rect 47911 102409 65793 102527
rect 65911 102409 83793 102527
rect 83911 102409 101793 102527
rect 101911 102409 119793 102527
rect 119911 102409 137793 102527
rect 137911 102409 155793 102527
rect 155911 102409 173793 102527
rect 173911 102409 191793 102527
rect 191911 102409 209793 102527
rect 209911 102409 227793 102527
rect 227911 102409 245793 102527
rect 245911 102409 263793 102527
rect 263911 102409 281793 102527
rect 281911 102409 294161 102527
rect 294279 102409 294370 102527
rect -2408 102367 294370 102409
rect -2408 102249 -2317 102367
rect -2199 102249 11793 102367
rect 11911 102249 29793 102367
rect 29911 102249 47793 102367
rect 47911 102249 65793 102367
rect 65911 102249 83793 102367
rect 83911 102249 101793 102367
rect 101911 102249 119793 102367
rect 119911 102249 137793 102367
rect 137911 102249 155793 102367
rect 155911 102249 173793 102367
rect 173911 102249 191793 102367
rect 191911 102249 209793 102367
rect 209911 102249 227793 102367
rect 227911 102249 245793 102367
rect 245911 102249 263793 102367
rect 263911 102249 281793 102367
rect 281911 102249 294161 102367
rect 294279 102249 294370 102367
rect -2408 102238 294370 102249
rect -2408 102237 -2108 102238
rect 11702 102237 12002 102238
rect 29702 102237 30002 102238
rect 47702 102237 48002 102238
rect 65702 102237 66002 102238
rect 83702 102237 84002 102238
rect 101702 102237 102002 102238
rect 119702 102237 120002 102238
rect 137702 102237 138002 102238
rect 155702 102237 156002 102238
rect 173702 102237 174002 102238
rect 191702 102237 192002 102238
rect 209702 102237 210002 102238
rect 227702 102237 228002 102238
rect 245702 102237 246002 102238
rect 263702 102237 264002 102238
rect 281702 102237 282002 102238
rect 294070 102237 294370 102238
rect -1468 100738 -1168 100739
rect 9902 100738 10202 100739
rect 27902 100738 28202 100739
rect 45902 100738 46202 100739
rect 63902 100738 64202 100739
rect 81902 100738 82202 100739
rect 99902 100738 100202 100739
rect 117902 100738 118202 100739
rect 135902 100738 136202 100739
rect 153902 100738 154202 100739
rect 171902 100738 172202 100739
rect 189902 100738 190202 100739
rect 207902 100738 208202 100739
rect 225902 100738 226202 100739
rect 243902 100738 244202 100739
rect 261902 100738 262202 100739
rect 279902 100738 280202 100739
rect 293130 100738 293430 100739
rect -1468 100727 293430 100738
rect -1468 100609 -1377 100727
rect -1259 100609 9993 100727
rect 10111 100609 27993 100727
rect 28111 100609 45993 100727
rect 46111 100609 63993 100727
rect 64111 100609 81993 100727
rect 82111 100609 99993 100727
rect 100111 100609 117993 100727
rect 118111 100609 135993 100727
rect 136111 100609 153993 100727
rect 154111 100609 171993 100727
rect 172111 100609 189993 100727
rect 190111 100609 207993 100727
rect 208111 100609 225993 100727
rect 226111 100609 243993 100727
rect 244111 100609 261993 100727
rect 262111 100609 279993 100727
rect 280111 100609 293221 100727
rect 293339 100609 293430 100727
rect -1468 100567 293430 100609
rect -1468 100449 -1377 100567
rect -1259 100449 9993 100567
rect 10111 100449 27993 100567
rect 28111 100449 45993 100567
rect 46111 100449 63993 100567
rect 64111 100449 81993 100567
rect 82111 100449 99993 100567
rect 100111 100449 117993 100567
rect 118111 100449 135993 100567
rect 136111 100449 153993 100567
rect 154111 100449 171993 100567
rect 172111 100449 189993 100567
rect 190111 100449 207993 100567
rect 208111 100449 225993 100567
rect 226111 100449 243993 100567
rect 244111 100449 261993 100567
rect 262111 100449 279993 100567
rect 280111 100449 293221 100567
rect 293339 100449 293430 100567
rect -1468 100438 293430 100449
rect -1468 100437 -1168 100438
rect 9902 100437 10202 100438
rect 27902 100437 28202 100438
rect 45902 100437 46202 100438
rect 63902 100437 64202 100438
rect 81902 100437 82202 100438
rect 99902 100437 100202 100438
rect 117902 100437 118202 100438
rect 135902 100437 136202 100438
rect 153902 100437 154202 100438
rect 171902 100437 172202 100438
rect 189902 100437 190202 100438
rect 207902 100437 208202 100438
rect 225902 100437 226202 100438
rect 243902 100437 244202 100438
rect 261902 100437 262202 100438
rect 279902 100437 280202 100438
rect 293130 100437 293430 100438
rect -3818 97138 -3518 97139
rect 6302 97138 6602 97139
rect 24302 97138 24602 97139
rect 42302 97138 42602 97139
rect 60302 97138 60602 97139
rect 78302 97138 78602 97139
rect 96302 97138 96602 97139
rect 114302 97138 114602 97139
rect 132302 97138 132602 97139
rect 150302 97138 150602 97139
rect 168302 97138 168602 97139
rect 186302 97138 186602 97139
rect 204302 97138 204602 97139
rect 222302 97138 222602 97139
rect 240302 97138 240602 97139
rect 258302 97138 258602 97139
rect 276302 97138 276602 97139
rect 295480 97138 295780 97139
rect -4288 97127 296250 97138
rect -4288 97009 -3727 97127
rect -3609 97009 6393 97127
rect 6511 97009 24393 97127
rect 24511 97009 42393 97127
rect 42511 97009 60393 97127
rect 60511 97009 78393 97127
rect 78511 97009 96393 97127
rect 96511 97009 114393 97127
rect 114511 97009 132393 97127
rect 132511 97009 150393 97127
rect 150511 97009 168393 97127
rect 168511 97009 186393 97127
rect 186511 97009 204393 97127
rect 204511 97009 222393 97127
rect 222511 97009 240393 97127
rect 240511 97009 258393 97127
rect 258511 97009 276393 97127
rect 276511 97009 295571 97127
rect 295689 97009 296250 97127
rect -4288 96967 296250 97009
rect -4288 96849 -3727 96967
rect -3609 96849 6393 96967
rect 6511 96849 24393 96967
rect 24511 96849 42393 96967
rect 42511 96849 60393 96967
rect 60511 96849 78393 96967
rect 78511 96849 96393 96967
rect 96511 96849 114393 96967
rect 114511 96849 132393 96967
rect 132511 96849 150393 96967
rect 150511 96849 168393 96967
rect 168511 96849 186393 96967
rect 186511 96849 204393 96967
rect 204511 96849 222393 96967
rect 222511 96849 240393 96967
rect 240511 96849 258393 96967
rect 258511 96849 276393 96967
rect 276511 96849 295571 96967
rect 295689 96849 296250 96967
rect -4288 96838 296250 96849
rect -3818 96837 -3518 96838
rect 6302 96837 6602 96838
rect 24302 96837 24602 96838
rect 42302 96837 42602 96838
rect 60302 96837 60602 96838
rect 78302 96837 78602 96838
rect 96302 96837 96602 96838
rect 114302 96837 114602 96838
rect 132302 96837 132602 96838
rect 150302 96837 150602 96838
rect 168302 96837 168602 96838
rect 186302 96837 186602 96838
rect 204302 96837 204602 96838
rect 222302 96837 222602 96838
rect 240302 96837 240602 96838
rect 258302 96837 258602 96838
rect 276302 96837 276602 96838
rect 295480 96837 295780 96838
rect -2878 95338 -2578 95339
rect 4502 95338 4802 95339
rect 22502 95338 22802 95339
rect 40502 95338 40802 95339
rect 58502 95338 58802 95339
rect 76502 95338 76802 95339
rect 94502 95338 94802 95339
rect 112502 95338 112802 95339
rect 130502 95338 130802 95339
rect 148502 95338 148802 95339
rect 166502 95338 166802 95339
rect 184502 95338 184802 95339
rect 202502 95338 202802 95339
rect 220502 95338 220802 95339
rect 238502 95338 238802 95339
rect 256502 95338 256802 95339
rect 274502 95338 274802 95339
rect 294540 95338 294840 95339
rect -3348 95327 295310 95338
rect -3348 95209 -2787 95327
rect -2669 95209 4593 95327
rect 4711 95209 22593 95327
rect 22711 95209 40593 95327
rect 40711 95209 58593 95327
rect 58711 95209 76593 95327
rect 76711 95209 94593 95327
rect 94711 95209 112593 95327
rect 112711 95209 130593 95327
rect 130711 95209 148593 95327
rect 148711 95209 166593 95327
rect 166711 95209 184593 95327
rect 184711 95209 202593 95327
rect 202711 95209 220593 95327
rect 220711 95209 238593 95327
rect 238711 95209 256593 95327
rect 256711 95209 274593 95327
rect 274711 95209 294631 95327
rect 294749 95209 295310 95327
rect -3348 95167 295310 95209
rect -3348 95049 -2787 95167
rect -2669 95049 4593 95167
rect 4711 95049 22593 95167
rect 22711 95049 40593 95167
rect 40711 95049 58593 95167
rect 58711 95049 76593 95167
rect 76711 95049 94593 95167
rect 94711 95049 112593 95167
rect 112711 95049 130593 95167
rect 130711 95049 148593 95167
rect 148711 95049 166593 95167
rect 166711 95049 184593 95167
rect 184711 95049 202593 95167
rect 202711 95049 220593 95167
rect 220711 95049 238593 95167
rect 238711 95049 256593 95167
rect 256711 95049 274593 95167
rect 274711 95049 294631 95167
rect 294749 95049 295310 95167
rect -3348 95038 295310 95049
rect -2878 95037 -2578 95038
rect 4502 95037 4802 95038
rect 22502 95037 22802 95038
rect 40502 95037 40802 95038
rect 58502 95037 58802 95038
rect 76502 95037 76802 95038
rect 94502 95037 94802 95038
rect 112502 95037 112802 95038
rect 130502 95037 130802 95038
rect 148502 95037 148802 95038
rect 166502 95037 166802 95038
rect 184502 95037 184802 95038
rect 202502 95037 202802 95038
rect 220502 95037 220802 95038
rect 238502 95037 238802 95038
rect 256502 95037 256802 95038
rect 274502 95037 274802 95038
rect 294540 95037 294840 95038
rect -1938 93538 -1638 93539
rect 2702 93538 3002 93539
rect 20702 93538 21002 93539
rect 38702 93538 39002 93539
rect 56702 93538 57002 93539
rect 74702 93538 75002 93539
rect 92702 93538 93002 93539
rect 110702 93538 111002 93539
rect 128702 93538 129002 93539
rect 146702 93538 147002 93539
rect 164702 93538 165002 93539
rect 182702 93538 183002 93539
rect 200702 93538 201002 93539
rect 218702 93538 219002 93539
rect 236702 93538 237002 93539
rect 254702 93538 255002 93539
rect 272702 93538 273002 93539
rect 290702 93538 291002 93539
rect 293600 93538 293900 93539
rect -2408 93527 294370 93538
rect -2408 93409 -1847 93527
rect -1729 93409 2793 93527
rect 2911 93409 20793 93527
rect 20911 93409 38793 93527
rect 38911 93409 56793 93527
rect 56911 93409 74793 93527
rect 74911 93409 92793 93527
rect 92911 93409 110793 93527
rect 110911 93409 128793 93527
rect 128911 93409 146793 93527
rect 146911 93409 164793 93527
rect 164911 93409 182793 93527
rect 182911 93409 200793 93527
rect 200911 93409 218793 93527
rect 218911 93409 236793 93527
rect 236911 93409 254793 93527
rect 254911 93409 272793 93527
rect 272911 93409 290793 93527
rect 290911 93409 293691 93527
rect 293809 93409 294370 93527
rect -2408 93367 294370 93409
rect -2408 93249 -1847 93367
rect -1729 93249 2793 93367
rect 2911 93249 20793 93367
rect 20911 93249 38793 93367
rect 38911 93249 56793 93367
rect 56911 93249 74793 93367
rect 74911 93249 92793 93367
rect 92911 93249 110793 93367
rect 110911 93249 128793 93367
rect 128911 93249 146793 93367
rect 146911 93249 164793 93367
rect 164911 93249 182793 93367
rect 182911 93249 200793 93367
rect 200911 93249 218793 93367
rect 218911 93249 236793 93367
rect 236911 93249 254793 93367
rect 254911 93249 272793 93367
rect 272911 93249 290793 93367
rect 290911 93249 293691 93367
rect 293809 93249 294370 93367
rect -2408 93238 294370 93249
rect -1938 93237 -1638 93238
rect 2702 93237 3002 93238
rect 20702 93237 21002 93238
rect 38702 93237 39002 93238
rect 56702 93237 57002 93238
rect 74702 93237 75002 93238
rect 92702 93237 93002 93238
rect 110702 93237 111002 93238
rect 128702 93237 129002 93238
rect 146702 93237 147002 93238
rect 164702 93237 165002 93238
rect 182702 93237 183002 93238
rect 200702 93237 201002 93238
rect 218702 93237 219002 93238
rect 236702 93237 237002 93238
rect 254702 93237 255002 93238
rect 272702 93237 273002 93238
rect 290702 93237 291002 93238
rect 293600 93237 293900 93238
rect -998 91738 -698 91739
rect 902 91738 1202 91739
rect 18902 91738 19202 91739
rect 36902 91738 37202 91739
rect 54902 91738 55202 91739
rect 72902 91738 73202 91739
rect 90902 91738 91202 91739
rect 108902 91738 109202 91739
rect 126902 91738 127202 91739
rect 144902 91738 145202 91739
rect 162902 91738 163202 91739
rect 180902 91738 181202 91739
rect 198902 91738 199202 91739
rect 216902 91738 217202 91739
rect 234902 91738 235202 91739
rect 252902 91738 253202 91739
rect 270902 91738 271202 91739
rect 288902 91738 289202 91739
rect 292660 91738 292960 91739
rect -1468 91727 293430 91738
rect -1468 91609 -907 91727
rect -789 91609 993 91727
rect 1111 91609 18993 91727
rect 19111 91609 36993 91727
rect 37111 91609 54993 91727
rect 55111 91609 72993 91727
rect 73111 91609 90993 91727
rect 91111 91609 108993 91727
rect 109111 91609 126993 91727
rect 127111 91609 144993 91727
rect 145111 91609 162993 91727
rect 163111 91609 180993 91727
rect 181111 91609 198993 91727
rect 199111 91609 216993 91727
rect 217111 91609 234993 91727
rect 235111 91609 252993 91727
rect 253111 91609 270993 91727
rect 271111 91609 288993 91727
rect 289111 91609 292751 91727
rect 292869 91609 293430 91727
rect -1468 91567 293430 91609
rect -1468 91449 -907 91567
rect -789 91449 993 91567
rect 1111 91449 18993 91567
rect 19111 91449 36993 91567
rect 37111 91449 54993 91567
rect 55111 91449 72993 91567
rect 73111 91449 90993 91567
rect 91111 91449 108993 91567
rect 109111 91449 126993 91567
rect 127111 91449 144993 91567
rect 145111 91449 162993 91567
rect 163111 91449 180993 91567
rect 181111 91449 198993 91567
rect 199111 91449 216993 91567
rect 217111 91449 234993 91567
rect 235111 91449 252993 91567
rect 253111 91449 270993 91567
rect 271111 91449 288993 91567
rect 289111 91449 292751 91567
rect 292869 91449 293430 91567
rect -1468 91438 293430 91449
rect -998 91437 -698 91438
rect 902 91437 1202 91438
rect 18902 91437 19202 91438
rect 36902 91437 37202 91438
rect 54902 91437 55202 91438
rect 72902 91437 73202 91438
rect 90902 91437 91202 91438
rect 108902 91437 109202 91438
rect 126902 91437 127202 91438
rect 144902 91437 145202 91438
rect 162902 91437 163202 91438
rect 180902 91437 181202 91438
rect 198902 91437 199202 91438
rect 216902 91437 217202 91438
rect 234902 91437 235202 91438
rect 252902 91437 253202 91438
rect 270902 91437 271202 91438
rect 288902 91437 289202 91438
rect 292660 91437 292960 91438
rect -4288 88138 -3988 88139
rect 15302 88138 15602 88139
rect 33302 88138 33602 88139
rect 51302 88138 51602 88139
rect 69302 88138 69602 88139
rect 87302 88138 87602 88139
rect 105302 88138 105602 88139
rect 123302 88138 123602 88139
rect 141302 88138 141602 88139
rect 159302 88138 159602 88139
rect 177302 88138 177602 88139
rect 195302 88138 195602 88139
rect 213302 88138 213602 88139
rect 231302 88138 231602 88139
rect 249302 88138 249602 88139
rect 267302 88138 267602 88139
rect 285302 88138 285602 88139
rect 295950 88138 296250 88139
rect -4288 88127 296250 88138
rect -4288 88009 -4197 88127
rect -4079 88009 15393 88127
rect 15511 88009 33393 88127
rect 33511 88009 51393 88127
rect 51511 88009 69393 88127
rect 69511 88009 87393 88127
rect 87511 88009 105393 88127
rect 105511 88009 123393 88127
rect 123511 88009 141393 88127
rect 141511 88009 159393 88127
rect 159511 88009 177393 88127
rect 177511 88009 195393 88127
rect 195511 88009 213393 88127
rect 213511 88009 231393 88127
rect 231511 88009 249393 88127
rect 249511 88009 267393 88127
rect 267511 88009 285393 88127
rect 285511 88009 296041 88127
rect 296159 88009 296250 88127
rect -4288 87967 296250 88009
rect -4288 87849 -4197 87967
rect -4079 87849 15393 87967
rect 15511 87849 33393 87967
rect 33511 87849 51393 87967
rect 51511 87849 69393 87967
rect 69511 87849 87393 87967
rect 87511 87849 105393 87967
rect 105511 87849 123393 87967
rect 123511 87849 141393 87967
rect 141511 87849 159393 87967
rect 159511 87849 177393 87967
rect 177511 87849 195393 87967
rect 195511 87849 213393 87967
rect 213511 87849 231393 87967
rect 231511 87849 249393 87967
rect 249511 87849 267393 87967
rect 267511 87849 285393 87967
rect 285511 87849 296041 87967
rect 296159 87849 296250 87967
rect -4288 87838 296250 87849
rect -4288 87837 -3988 87838
rect 15302 87837 15602 87838
rect 33302 87837 33602 87838
rect 51302 87837 51602 87838
rect 69302 87837 69602 87838
rect 87302 87837 87602 87838
rect 105302 87837 105602 87838
rect 123302 87837 123602 87838
rect 141302 87837 141602 87838
rect 159302 87837 159602 87838
rect 177302 87837 177602 87838
rect 195302 87837 195602 87838
rect 213302 87837 213602 87838
rect 231302 87837 231602 87838
rect 249302 87837 249602 87838
rect 267302 87837 267602 87838
rect 285302 87837 285602 87838
rect 295950 87837 296250 87838
rect -3348 86338 -3048 86339
rect 13502 86338 13802 86339
rect 31502 86338 31802 86339
rect 49502 86338 49802 86339
rect 67502 86338 67802 86339
rect 85502 86338 85802 86339
rect 103502 86338 103802 86339
rect 121502 86338 121802 86339
rect 139502 86338 139802 86339
rect 157502 86338 157802 86339
rect 175502 86338 175802 86339
rect 193502 86338 193802 86339
rect 211502 86338 211802 86339
rect 229502 86338 229802 86339
rect 247502 86338 247802 86339
rect 265502 86338 265802 86339
rect 283502 86338 283802 86339
rect 295010 86338 295310 86339
rect -3348 86327 295310 86338
rect -3348 86209 -3257 86327
rect -3139 86209 13593 86327
rect 13711 86209 31593 86327
rect 31711 86209 49593 86327
rect 49711 86209 67593 86327
rect 67711 86209 85593 86327
rect 85711 86209 103593 86327
rect 103711 86209 121593 86327
rect 121711 86209 139593 86327
rect 139711 86209 157593 86327
rect 157711 86209 175593 86327
rect 175711 86209 193593 86327
rect 193711 86209 211593 86327
rect 211711 86209 229593 86327
rect 229711 86209 247593 86327
rect 247711 86209 265593 86327
rect 265711 86209 283593 86327
rect 283711 86209 295101 86327
rect 295219 86209 295310 86327
rect -3348 86167 295310 86209
rect -3348 86049 -3257 86167
rect -3139 86049 13593 86167
rect 13711 86049 31593 86167
rect 31711 86049 49593 86167
rect 49711 86049 67593 86167
rect 67711 86049 85593 86167
rect 85711 86049 103593 86167
rect 103711 86049 121593 86167
rect 121711 86049 139593 86167
rect 139711 86049 157593 86167
rect 157711 86049 175593 86167
rect 175711 86049 193593 86167
rect 193711 86049 211593 86167
rect 211711 86049 229593 86167
rect 229711 86049 247593 86167
rect 247711 86049 265593 86167
rect 265711 86049 283593 86167
rect 283711 86049 295101 86167
rect 295219 86049 295310 86167
rect -3348 86038 295310 86049
rect -3348 86037 -3048 86038
rect 13502 86037 13802 86038
rect 31502 86037 31802 86038
rect 49502 86037 49802 86038
rect 67502 86037 67802 86038
rect 85502 86037 85802 86038
rect 103502 86037 103802 86038
rect 121502 86037 121802 86038
rect 139502 86037 139802 86038
rect 157502 86037 157802 86038
rect 175502 86037 175802 86038
rect 193502 86037 193802 86038
rect 211502 86037 211802 86038
rect 229502 86037 229802 86038
rect 247502 86037 247802 86038
rect 265502 86037 265802 86038
rect 283502 86037 283802 86038
rect 295010 86037 295310 86038
rect -2408 84538 -2108 84539
rect 11702 84538 12002 84539
rect 29702 84538 30002 84539
rect 47702 84538 48002 84539
rect 65702 84538 66002 84539
rect 83702 84538 84002 84539
rect 101702 84538 102002 84539
rect 119702 84538 120002 84539
rect 137702 84538 138002 84539
rect 155702 84538 156002 84539
rect 173702 84538 174002 84539
rect 191702 84538 192002 84539
rect 209702 84538 210002 84539
rect 227702 84538 228002 84539
rect 245702 84538 246002 84539
rect 263702 84538 264002 84539
rect 281702 84538 282002 84539
rect 294070 84538 294370 84539
rect -2408 84527 294370 84538
rect -2408 84409 -2317 84527
rect -2199 84409 11793 84527
rect 11911 84409 29793 84527
rect 29911 84409 47793 84527
rect 47911 84409 65793 84527
rect 65911 84409 83793 84527
rect 83911 84409 101793 84527
rect 101911 84409 119793 84527
rect 119911 84409 137793 84527
rect 137911 84409 155793 84527
rect 155911 84409 173793 84527
rect 173911 84409 191793 84527
rect 191911 84409 209793 84527
rect 209911 84409 227793 84527
rect 227911 84409 245793 84527
rect 245911 84409 263793 84527
rect 263911 84409 281793 84527
rect 281911 84409 294161 84527
rect 294279 84409 294370 84527
rect -2408 84367 294370 84409
rect -2408 84249 -2317 84367
rect -2199 84249 11793 84367
rect 11911 84249 29793 84367
rect 29911 84249 47793 84367
rect 47911 84249 65793 84367
rect 65911 84249 83793 84367
rect 83911 84249 101793 84367
rect 101911 84249 119793 84367
rect 119911 84249 137793 84367
rect 137911 84249 155793 84367
rect 155911 84249 173793 84367
rect 173911 84249 191793 84367
rect 191911 84249 209793 84367
rect 209911 84249 227793 84367
rect 227911 84249 245793 84367
rect 245911 84249 263793 84367
rect 263911 84249 281793 84367
rect 281911 84249 294161 84367
rect 294279 84249 294370 84367
rect -2408 84238 294370 84249
rect -2408 84237 -2108 84238
rect 11702 84237 12002 84238
rect 29702 84237 30002 84238
rect 47702 84237 48002 84238
rect 65702 84237 66002 84238
rect 83702 84237 84002 84238
rect 101702 84237 102002 84238
rect 119702 84237 120002 84238
rect 137702 84237 138002 84238
rect 155702 84237 156002 84238
rect 173702 84237 174002 84238
rect 191702 84237 192002 84238
rect 209702 84237 210002 84238
rect 227702 84237 228002 84238
rect 245702 84237 246002 84238
rect 263702 84237 264002 84238
rect 281702 84237 282002 84238
rect 294070 84237 294370 84238
rect -1468 82738 -1168 82739
rect 9902 82738 10202 82739
rect 27902 82738 28202 82739
rect 45902 82738 46202 82739
rect 63902 82738 64202 82739
rect 81902 82738 82202 82739
rect 99902 82738 100202 82739
rect 117902 82738 118202 82739
rect 135902 82738 136202 82739
rect 153902 82738 154202 82739
rect 171902 82738 172202 82739
rect 189902 82738 190202 82739
rect 207902 82738 208202 82739
rect 225902 82738 226202 82739
rect 243902 82738 244202 82739
rect 261902 82738 262202 82739
rect 279902 82738 280202 82739
rect 293130 82738 293430 82739
rect -1468 82727 293430 82738
rect -1468 82609 -1377 82727
rect -1259 82609 9993 82727
rect 10111 82609 27993 82727
rect 28111 82609 45993 82727
rect 46111 82609 63993 82727
rect 64111 82609 81993 82727
rect 82111 82609 99993 82727
rect 100111 82609 117993 82727
rect 118111 82609 135993 82727
rect 136111 82609 153993 82727
rect 154111 82609 171993 82727
rect 172111 82609 189993 82727
rect 190111 82609 207993 82727
rect 208111 82609 225993 82727
rect 226111 82609 243993 82727
rect 244111 82609 261993 82727
rect 262111 82609 279993 82727
rect 280111 82609 293221 82727
rect 293339 82609 293430 82727
rect -1468 82567 293430 82609
rect -1468 82449 -1377 82567
rect -1259 82449 9993 82567
rect 10111 82449 27993 82567
rect 28111 82449 45993 82567
rect 46111 82449 63993 82567
rect 64111 82449 81993 82567
rect 82111 82449 99993 82567
rect 100111 82449 117993 82567
rect 118111 82449 135993 82567
rect 136111 82449 153993 82567
rect 154111 82449 171993 82567
rect 172111 82449 189993 82567
rect 190111 82449 207993 82567
rect 208111 82449 225993 82567
rect 226111 82449 243993 82567
rect 244111 82449 261993 82567
rect 262111 82449 279993 82567
rect 280111 82449 293221 82567
rect 293339 82449 293430 82567
rect -1468 82438 293430 82449
rect -1468 82437 -1168 82438
rect 9902 82437 10202 82438
rect 27902 82437 28202 82438
rect 45902 82437 46202 82438
rect 63902 82437 64202 82438
rect 81902 82437 82202 82438
rect 99902 82437 100202 82438
rect 117902 82437 118202 82438
rect 135902 82437 136202 82438
rect 153902 82437 154202 82438
rect 171902 82437 172202 82438
rect 189902 82437 190202 82438
rect 207902 82437 208202 82438
rect 225902 82437 226202 82438
rect 243902 82437 244202 82438
rect 261902 82437 262202 82438
rect 279902 82437 280202 82438
rect 293130 82437 293430 82438
rect -3818 79138 -3518 79139
rect 6302 79138 6602 79139
rect 24302 79138 24602 79139
rect 42302 79138 42602 79139
rect 60302 79138 60602 79139
rect 78302 79138 78602 79139
rect 96302 79138 96602 79139
rect 114302 79138 114602 79139
rect 132302 79138 132602 79139
rect 150302 79138 150602 79139
rect 168302 79138 168602 79139
rect 186302 79138 186602 79139
rect 204302 79138 204602 79139
rect 222302 79138 222602 79139
rect 240302 79138 240602 79139
rect 258302 79138 258602 79139
rect 276302 79138 276602 79139
rect 295480 79138 295780 79139
rect -4288 79127 296250 79138
rect -4288 79009 -3727 79127
rect -3609 79009 6393 79127
rect 6511 79009 24393 79127
rect 24511 79009 42393 79127
rect 42511 79009 60393 79127
rect 60511 79009 78393 79127
rect 78511 79009 96393 79127
rect 96511 79009 114393 79127
rect 114511 79009 132393 79127
rect 132511 79009 150393 79127
rect 150511 79009 168393 79127
rect 168511 79009 186393 79127
rect 186511 79009 204393 79127
rect 204511 79009 222393 79127
rect 222511 79009 240393 79127
rect 240511 79009 258393 79127
rect 258511 79009 276393 79127
rect 276511 79009 295571 79127
rect 295689 79009 296250 79127
rect -4288 78967 296250 79009
rect -4288 78849 -3727 78967
rect -3609 78849 6393 78967
rect 6511 78849 24393 78967
rect 24511 78849 42393 78967
rect 42511 78849 60393 78967
rect 60511 78849 78393 78967
rect 78511 78849 96393 78967
rect 96511 78849 114393 78967
rect 114511 78849 132393 78967
rect 132511 78849 150393 78967
rect 150511 78849 168393 78967
rect 168511 78849 186393 78967
rect 186511 78849 204393 78967
rect 204511 78849 222393 78967
rect 222511 78849 240393 78967
rect 240511 78849 258393 78967
rect 258511 78849 276393 78967
rect 276511 78849 295571 78967
rect 295689 78849 296250 78967
rect -4288 78838 296250 78849
rect -3818 78837 -3518 78838
rect 6302 78837 6602 78838
rect 24302 78837 24602 78838
rect 42302 78837 42602 78838
rect 60302 78837 60602 78838
rect 78302 78837 78602 78838
rect 96302 78837 96602 78838
rect 114302 78837 114602 78838
rect 132302 78837 132602 78838
rect 150302 78837 150602 78838
rect 168302 78837 168602 78838
rect 186302 78837 186602 78838
rect 204302 78837 204602 78838
rect 222302 78837 222602 78838
rect 240302 78837 240602 78838
rect 258302 78837 258602 78838
rect 276302 78837 276602 78838
rect 295480 78837 295780 78838
rect -2878 77338 -2578 77339
rect 4502 77338 4802 77339
rect 22502 77338 22802 77339
rect 40502 77338 40802 77339
rect 58502 77338 58802 77339
rect 76502 77338 76802 77339
rect 94502 77338 94802 77339
rect 112502 77338 112802 77339
rect 130502 77338 130802 77339
rect 148502 77338 148802 77339
rect 166502 77338 166802 77339
rect 184502 77338 184802 77339
rect 202502 77338 202802 77339
rect 220502 77338 220802 77339
rect 238502 77338 238802 77339
rect 256502 77338 256802 77339
rect 274502 77338 274802 77339
rect 294540 77338 294840 77339
rect -3348 77327 295310 77338
rect -3348 77209 -2787 77327
rect -2669 77209 4593 77327
rect 4711 77209 22593 77327
rect 22711 77209 40593 77327
rect 40711 77209 58593 77327
rect 58711 77209 76593 77327
rect 76711 77209 94593 77327
rect 94711 77209 112593 77327
rect 112711 77209 130593 77327
rect 130711 77209 148593 77327
rect 148711 77209 166593 77327
rect 166711 77209 184593 77327
rect 184711 77209 202593 77327
rect 202711 77209 220593 77327
rect 220711 77209 238593 77327
rect 238711 77209 256593 77327
rect 256711 77209 274593 77327
rect 274711 77209 294631 77327
rect 294749 77209 295310 77327
rect -3348 77167 295310 77209
rect -3348 77049 -2787 77167
rect -2669 77049 4593 77167
rect 4711 77049 22593 77167
rect 22711 77049 40593 77167
rect 40711 77049 58593 77167
rect 58711 77049 76593 77167
rect 76711 77049 94593 77167
rect 94711 77049 112593 77167
rect 112711 77049 130593 77167
rect 130711 77049 148593 77167
rect 148711 77049 166593 77167
rect 166711 77049 184593 77167
rect 184711 77049 202593 77167
rect 202711 77049 220593 77167
rect 220711 77049 238593 77167
rect 238711 77049 256593 77167
rect 256711 77049 274593 77167
rect 274711 77049 294631 77167
rect 294749 77049 295310 77167
rect -3348 77038 295310 77049
rect -2878 77037 -2578 77038
rect 4502 77037 4802 77038
rect 22502 77037 22802 77038
rect 40502 77037 40802 77038
rect 58502 77037 58802 77038
rect 76502 77037 76802 77038
rect 94502 77037 94802 77038
rect 112502 77037 112802 77038
rect 130502 77037 130802 77038
rect 148502 77037 148802 77038
rect 166502 77037 166802 77038
rect 184502 77037 184802 77038
rect 202502 77037 202802 77038
rect 220502 77037 220802 77038
rect 238502 77037 238802 77038
rect 256502 77037 256802 77038
rect 274502 77037 274802 77038
rect 294540 77037 294840 77038
rect -1938 75538 -1638 75539
rect 2702 75538 3002 75539
rect 20702 75538 21002 75539
rect 38702 75538 39002 75539
rect 56702 75538 57002 75539
rect 74702 75538 75002 75539
rect 92702 75538 93002 75539
rect 110702 75538 111002 75539
rect 128702 75538 129002 75539
rect 146702 75538 147002 75539
rect 164702 75538 165002 75539
rect 182702 75538 183002 75539
rect 200702 75538 201002 75539
rect 218702 75538 219002 75539
rect 236702 75538 237002 75539
rect 254702 75538 255002 75539
rect 272702 75538 273002 75539
rect 290702 75538 291002 75539
rect 293600 75538 293900 75539
rect -2408 75527 294370 75538
rect -2408 75409 -1847 75527
rect -1729 75409 2793 75527
rect 2911 75409 20793 75527
rect 20911 75409 38793 75527
rect 38911 75409 56793 75527
rect 56911 75409 74793 75527
rect 74911 75409 92793 75527
rect 92911 75409 110793 75527
rect 110911 75409 128793 75527
rect 128911 75409 146793 75527
rect 146911 75409 164793 75527
rect 164911 75409 182793 75527
rect 182911 75409 200793 75527
rect 200911 75409 218793 75527
rect 218911 75409 236793 75527
rect 236911 75409 254793 75527
rect 254911 75409 272793 75527
rect 272911 75409 290793 75527
rect 290911 75409 293691 75527
rect 293809 75409 294370 75527
rect -2408 75367 294370 75409
rect -2408 75249 -1847 75367
rect -1729 75249 2793 75367
rect 2911 75249 20793 75367
rect 20911 75249 38793 75367
rect 38911 75249 56793 75367
rect 56911 75249 74793 75367
rect 74911 75249 92793 75367
rect 92911 75249 110793 75367
rect 110911 75249 128793 75367
rect 128911 75249 146793 75367
rect 146911 75249 164793 75367
rect 164911 75249 182793 75367
rect 182911 75249 200793 75367
rect 200911 75249 218793 75367
rect 218911 75249 236793 75367
rect 236911 75249 254793 75367
rect 254911 75249 272793 75367
rect 272911 75249 290793 75367
rect 290911 75249 293691 75367
rect 293809 75249 294370 75367
rect -2408 75238 294370 75249
rect -1938 75237 -1638 75238
rect 2702 75237 3002 75238
rect 20702 75237 21002 75238
rect 38702 75237 39002 75238
rect 56702 75237 57002 75238
rect 74702 75237 75002 75238
rect 92702 75237 93002 75238
rect 110702 75237 111002 75238
rect 128702 75237 129002 75238
rect 146702 75237 147002 75238
rect 164702 75237 165002 75238
rect 182702 75237 183002 75238
rect 200702 75237 201002 75238
rect 218702 75237 219002 75238
rect 236702 75237 237002 75238
rect 254702 75237 255002 75238
rect 272702 75237 273002 75238
rect 290702 75237 291002 75238
rect 293600 75237 293900 75238
rect -998 73738 -698 73739
rect 902 73738 1202 73739
rect 18902 73738 19202 73739
rect 36902 73738 37202 73739
rect 54902 73738 55202 73739
rect 72902 73738 73202 73739
rect 90902 73738 91202 73739
rect 108902 73738 109202 73739
rect 126902 73738 127202 73739
rect 144902 73738 145202 73739
rect 162902 73738 163202 73739
rect 180902 73738 181202 73739
rect 198902 73738 199202 73739
rect 216902 73738 217202 73739
rect 234902 73738 235202 73739
rect 252902 73738 253202 73739
rect 270902 73738 271202 73739
rect 288902 73738 289202 73739
rect 292660 73738 292960 73739
rect -1468 73727 293430 73738
rect -1468 73609 -907 73727
rect -789 73609 993 73727
rect 1111 73609 18993 73727
rect 19111 73609 36993 73727
rect 37111 73609 54993 73727
rect 55111 73609 72993 73727
rect 73111 73609 90993 73727
rect 91111 73609 108993 73727
rect 109111 73609 126993 73727
rect 127111 73609 144993 73727
rect 145111 73609 162993 73727
rect 163111 73609 180993 73727
rect 181111 73609 198993 73727
rect 199111 73609 216993 73727
rect 217111 73609 234993 73727
rect 235111 73609 252993 73727
rect 253111 73609 270993 73727
rect 271111 73609 288993 73727
rect 289111 73609 292751 73727
rect 292869 73609 293430 73727
rect -1468 73567 293430 73609
rect -1468 73449 -907 73567
rect -789 73449 993 73567
rect 1111 73449 18993 73567
rect 19111 73449 36993 73567
rect 37111 73449 54993 73567
rect 55111 73449 72993 73567
rect 73111 73449 90993 73567
rect 91111 73449 108993 73567
rect 109111 73449 126993 73567
rect 127111 73449 144993 73567
rect 145111 73449 162993 73567
rect 163111 73449 180993 73567
rect 181111 73449 198993 73567
rect 199111 73449 216993 73567
rect 217111 73449 234993 73567
rect 235111 73449 252993 73567
rect 253111 73449 270993 73567
rect 271111 73449 288993 73567
rect 289111 73449 292751 73567
rect 292869 73449 293430 73567
rect -1468 73438 293430 73449
rect -998 73437 -698 73438
rect 902 73437 1202 73438
rect 18902 73437 19202 73438
rect 36902 73437 37202 73438
rect 54902 73437 55202 73438
rect 72902 73437 73202 73438
rect 90902 73437 91202 73438
rect 108902 73437 109202 73438
rect 126902 73437 127202 73438
rect 144902 73437 145202 73438
rect 162902 73437 163202 73438
rect 180902 73437 181202 73438
rect 198902 73437 199202 73438
rect 216902 73437 217202 73438
rect 234902 73437 235202 73438
rect 252902 73437 253202 73438
rect 270902 73437 271202 73438
rect 288902 73437 289202 73438
rect 292660 73437 292960 73438
rect -4288 70138 -3988 70139
rect 15302 70138 15602 70139
rect 33302 70138 33602 70139
rect 51302 70138 51602 70139
rect 69302 70138 69602 70139
rect 87302 70138 87602 70139
rect 105302 70138 105602 70139
rect 123302 70138 123602 70139
rect 141302 70138 141602 70139
rect 159302 70138 159602 70139
rect 177302 70138 177602 70139
rect 195302 70138 195602 70139
rect 213302 70138 213602 70139
rect 231302 70138 231602 70139
rect 249302 70138 249602 70139
rect 267302 70138 267602 70139
rect 285302 70138 285602 70139
rect 295950 70138 296250 70139
rect -4288 70127 296250 70138
rect -4288 70009 -4197 70127
rect -4079 70009 15393 70127
rect 15511 70009 33393 70127
rect 33511 70009 51393 70127
rect 51511 70009 69393 70127
rect 69511 70009 87393 70127
rect 87511 70009 105393 70127
rect 105511 70009 123393 70127
rect 123511 70009 141393 70127
rect 141511 70009 159393 70127
rect 159511 70009 177393 70127
rect 177511 70009 195393 70127
rect 195511 70009 213393 70127
rect 213511 70009 231393 70127
rect 231511 70009 249393 70127
rect 249511 70009 267393 70127
rect 267511 70009 285393 70127
rect 285511 70009 296041 70127
rect 296159 70009 296250 70127
rect -4288 69967 296250 70009
rect -4288 69849 -4197 69967
rect -4079 69849 15393 69967
rect 15511 69849 33393 69967
rect 33511 69849 51393 69967
rect 51511 69849 69393 69967
rect 69511 69849 87393 69967
rect 87511 69849 105393 69967
rect 105511 69849 123393 69967
rect 123511 69849 141393 69967
rect 141511 69849 159393 69967
rect 159511 69849 177393 69967
rect 177511 69849 195393 69967
rect 195511 69849 213393 69967
rect 213511 69849 231393 69967
rect 231511 69849 249393 69967
rect 249511 69849 267393 69967
rect 267511 69849 285393 69967
rect 285511 69849 296041 69967
rect 296159 69849 296250 69967
rect -4288 69838 296250 69849
rect -4288 69837 -3988 69838
rect 15302 69837 15602 69838
rect 33302 69837 33602 69838
rect 51302 69837 51602 69838
rect 69302 69837 69602 69838
rect 87302 69837 87602 69838
rect 105302 69837 105602 69838
rect 123302 69837 123602 69838
rect 141302 69837 141602 69838
rect 159302 69837 159602 69838
rect 177302 69837 177602 69838
rect 195302 69837 195602 69838
rect 213302 69837 213602 69838
rect 231302 69837 231602 69838
rect 249302 69837 249602 69838
rect 267302 69837 267602 69838
rect 285302 69837 285602 69838
rect 295950 69837 296250 69838
rect -3348 68338 -3048 68339
rect 13502 68338 13802 68339
rect 31502 68338 31802 68339
rect 49502 68338 49802 68339
rect 67502 68338 67802 68339
rect 85502 68338 85802 68339
rect 103502 68338 103802 68339
rect 121502 68338 121802 68339
rect 139502 68338 139802 68339
rect 157502 68338 157802 68339
rect 175502 68338 175802 68339
rect 193502 68338 193802 68339
rect 211502 68338 211802 68339
rect 229502 68338 229802 68339
rect 247502 68338 247802 68339
rect 265502 68338 265802 68339
rect 283502 68338 283802 68339
rect 295010 68338 295310 68339
rect -3348 68327 295310 68338
rect -3348 68209 -3257 68327
rect -3139 68209 13593 68327
rect 13711 68209 31593 68327
rect 31711 68209 49593 68327
rect 49711 68209 67593 68327
rect 67711 68209 85593 68327
rect 85711 68209 103593 68327
rect 103711 68209 121593 68327
rect 121711 68209 139593 68327
rect 139711 68209 157593 68327
rect 157711 68209 175593 68327
rect 175711 68209 193593 68327
rect 193711 68209 211593 68327
rect 211711 68209 229593 68327
rect 229711 68209 247593 68327
rect 247711 68209 265593 68327
rect 265711 68209 283593 68327
rect 283711 68209 295101 68327
rect 295219 68209 295310 68327
rect -3348 68167 295310 68209
rect -3348 68049 -3257 68167
rect -3139 68049 13593 68167
rect 13711 68049 31593 68167
rect 31711 68049 49593 68167
rect 49711 68049 67593 68167
rect 67711 68049 85593 68167
rect 85711 68049 103593 68167
rect 103711 68049 121593 68167
rect 121711 68049 139593 68167
rect 139711 68049 157593 68167
rect 157711 68049 175593 68167
rect 175711 68049 193593 68167
rect 193711 68049 211593 68167
rect 211711 68049 229593 68167
rect 229711 68049 247593 68167
rect 247711 68049 265593 68167
rect 265711 68049 283593 68167
rect 283711 68049 295101 68167
rect 295219 68049 295310 68167
rect -3348 68038 295310 68049
rect -3348 68037 -3048 68038
rect 13502 68037 13802 68038
rect 31502 68037 31802 68038
rect 49502 68037 49802 68038
rect 67502 68037 67802 68038
rect 85502 68037 85802 68038
rect 103502 68037 103802 68038
rect 121502 68037 121802 68038
rect 139502 68037 139802 68038
rect 157502 68037 157802 68038
rect 175502 68037 175802 68038
rect 193502 68037 193802 68038
rect 211502 68037 211802 68038
rect 229502 68037 229802 68038
rect 247502 68037 247802 68038
rect 265502 68037 265802 68038
rect 283502 68037 283802 68038
rect 295010 68037 295310 68038
rect -2408 66538 -2108 66539
rect 11702 66538 12002 66539
rect 29702 66538 30002 66539
rect 47702 66538 48002 66539
rect 65702 66538 66002 66539
rect 83702 66538 84002 66539
rect 101702 66538 102002 66539
rect 119702 66538 120002 66539
rect 137702 66538 138002 66539
rect 155702 66538 156002 66539
rect 173702 66538 174002 66539
rect 191702 66538 192002 66539
rect 209702 66538 210002 66539
rect 227702 66538 228002 66539
rect 245702 66538 246002 66539
rect 263702 66538 264002 66539
rect 281702 66538 282002 66539
rect 294070 66538 294370 66539
rect -2408 66527 294370 66538
rect -2408 66409 -2317 66527
rect -2199 66409 11793 66527
rect 11911 66409 29793 66527
rect 29911 66409 47793 66527
rect 47911 66409 65793 66527
rect 65911 66409 83793 66527
rect 83911 66409 101793 66527
rect 101911 66409 119793 66527
rect 119911 66409 137793 66527
rect 137911 66409 155793 66527
rect 155911 66409 173793 66527
rect 173911 66409 191793 66527
rect 191911 66409 209793 66527
rect 209911 66409 227793 66527
rect 227911 66409 245793 66527
rect 245911 66409 263793 66527
rect 263911 66409 281793 66527
rect 281911 66409 294161 66527
rect 294279 66409 294370 66527
rect -2408 66367 294370 66409
rect -2408 66249 -2317 66367
rect -2199 66249 11793 66367
rect 11911 66249 29793 66367
rect 29911 66249 47793 66367
rect 47911 66249 65793 66367
rect 65911 66249 83793 66367
rect 83911 66249 101793 66367
rect 101911 66249 119793 66367
rect 119911 66249 137793 66367
rect 137911 66249 155793 66367
rect 155911 66249 173793 66367
rect 173911 66249 191793 66367
rect 191911 66249 209793 66367
rect 209911 66249 227793 66367
rect 227911 66249 245793 66367
rect 245911 66249 263793 66367
rect 263911 66249 281793 66367
rect 281911 66249 294161 66367
rect 294279 66249 294370 66367
rect -2408 66238 294370 66249
rect -2408 66237 -2108 66238
rect 11702 66237 12002 66238
rect 29702 66237 30002 66238
rect 47702 66237 48002 66238
rect 65702 66237 66002 66238
rect 83702 66237 84002 66238
rect 101702 66237 102002 66238
rect 119702 66237 120002 66238
rect 137702 66237 138002 66238
rect 155702 66237 156002 66238
rect 173702 66237 174002 66238
rect 191702 66237 192002 66238
rect 209702 66237 210002 66238
rect 227702 66237 228002 66238
rect 245702 66237 246002 66238
rect 263702 66237 264002 66238
rect 281702 66237 282002 66238
rect 294070 66237 294370 66238
rect -1468 64738 -1168 64739
rect 9902 64738 10202 64739
rect 27902 64738 28202 64739
rect 45902 64738 46202 64739
rect 63902 64738 64202 64739
rect 81902 64738 82202 64739
rect 99902 64738 100202 64739
rect 117902 64738 118202 64739
rect 135902 64738 136202 64739
rect 153902 64738 154202 64739
rect 171902 64738 172202 64739
rect 189902 64738 190202 64739
rect 207902 64738 208202 64739
rect 225902 64738 226202 64739
rect 243902 64738 244202 64739
rect 261902 64738 262202 64739
rect 279902 64738 280202 64739
rect 293130 64738 293430 64739
rect -1468 64727 293430 64738
rect -1468 64609 -1377 64727
rect -1259 64609 9993 64727
rect 10111 64609 27993 64727
rect 28111 64609 45993 64727
rect 46111 64609 63993 64727
rect 64111 64609 81993 64727
rect 82111 64609 99993 64727
rect 100111 64609 117993 64727
rect 118111 64609 135993 64727
rect 136111 64609 153993 64727
rect 154111 64609 171993 64727
rect 172111 64609 189993 64727
rect 190111 64609 207993 64727
rect 208111 64609 225993 64727
rect 226111 64609 243993 64727
rect 244111 64609 261993 64727
rect 262111 64609 279993 64727
rect 280111 64609 293221 64727
rect 293339 64609 293430 64727
rect -1468 64567 293430 64609
rect -1468 64449 -1377 64567
rect -1259 64449 9993 64567
rect 10111 64449 27993 64567
rect 28111 64449 45993 64567
rect 46111 64449 63993 64567
rect 64111 64449 81993 64567
rect 82111 64449 99993 64567
rect 100111 64449 117993 64567
rect 118111 64449 135993 64567
rect 136111 64449 153993 64567
rect 154111 64449 171993 64567
rect 172111 64449 189993 64567
rect 190111 64449 207993 64567
rect 208111 64449 225993 64567
rect 226111 64449 243993 64567
rect 244111 64449 261993 64567
rect 262111 64449 279993 64567
rect 280111 64449 293221 64567
rect 293339 64449 293430 64567
rect -1468 64438 293430 64449
rect -1468 64437 -1168 64438
rect 9902 64437 10202 64438
rect 27902 64437 28202 64438
rect 45902 64437 46202 64438
rect 63902 64437 64202 64438
rect 81902 64437 82202 64438
rect 99902 64437 100202 64438
rect 117902 64437 118202 64438
rect 135902 64437 136202 64438
rect 153902 64437 154202 64438
rect 171902 64437 172202 64438
rect 189902 64437 190202 64438
rect 207902 64437 208202 64438
rect 225902 64437 226202 64438
rect 243902 64437 244202 64438
rect 261902 64437 262202 64438
rect 279902 64437 280202 64438
rect 293130 64437 293430 64438
rect -3818 61138 -3518 61139
rect 6302 61138 6602 61139
rect 24302 61138 24602 61139
rect 42302 61138 42602 61139
rect 60302 61138 60602 61139
rect 78302 61138 78602 61139
rect 96302 61138 96602 61139
rect 114302 61138 114602 61139
rect 132302 61138 132602 61139
rect 150302 61138 150602 61139
rect 168302 61138 168602 61139
rect 186302 61138 186602 61139
rect 204302 61138 204602 61139
rect 222302 61138 222602 61139
rect 240302 61138 240602 61139
rect 258302 61138 258602 61139
rect 276302 61138 276602 61139
rect 295480 61138 295780 61139
rect -4288 61127 296250 61138
rect -4288 61009 -3727 61127
rect -3609 61009 6393 61127
rect 6511 61009 24393 61127
rect 24511 61009 42393 61127
rect 42511 61009 60393 61127
rect 60511 61009 78393 61127
rect 78511 61009 96393 61127
rect 96511 61009 114393 61127
rect 114511 61009 132393 61127
rect 132511 61009 150393 61127
rect 150511 61009 168393 61127
rect 168511 61009 186393 61127
rect 186511 61009 204393 61127
rect 204511 61009 222393 61127
rect 222511 61009 240393 61127
rect 240511 61009 258393 61127
rect 258511 61009 276393 61127
rect 276511 61009 295571 61127
rect 295689 61009 296250 61127
rect -4288 60967 296250 61009
rect -4288 60849 -3727 60967
rect -3609 60849 6393 60967
rect 6511 60849 24393 60967
rect 24511 60849 42393 60967
rect 42511 60849 60393 60967
rect 60511 60849 78393 60967
rect 78511 60849 96393 60967
rect 96511 60849 114393 60967
rect 114511 60849 132393 60967
rect 132511 60849 150393 60967
rect 150511 60849 168393 60967
rect 168511 60849 186393 60967
rect 186511 60849 204393 60967
rect 204511 60849 222393 60967
rect 222511 60849 240393 60967
rect 240511 60849 258393 60967
rect 258511 60849 276393 60967
rect 276511 60849 295571 60967
rect 295689 60849 296250 60967
rect -4288 60838 296250 60849
rect -3818 60837 -3518 60838
rect 6302 60837 6602 60838
rect 24302 60837 24602 60838
rect 42302 60837 42602 60838
rect 60302 60837 60602 60838
rect 78302 60837 78602 60838
rect 96302 60837 96602 60838
rect 114302 60837 114602 60838
rect 132302 60837 132602 60838
rect 150302 60837 150602 60838
rect 168302 60837 168602 60838
rect 186302 60837 186602 60838
rect 204302 60837 204602 60838
rect 222302 60837 222602 60838
rect 240302 60837 240602 60838
rect 258302 60837 258602 60838
rect 276302 60837 276602 60838
rect 295480 60837 295780 60838
rect -2878 59338 -2578 59339
rect 4502 59338 4802 59339
rect 22502 59338 22802 59339
rect 40502 59338 40802 59339
rect 58502 59338 58802 59339
rect 76502 59338 76802 59339
rect 94502 59338 94802 59339
rect 112502 59338 112802 59339
rect 130502 59338 130802 59339
rect 148502 59338 148802 59339
rect 166502 59338 166802 59339
rect 184502 59338 184802 59339
rect 202502 59338 202802 59339
rect 220502 59338 220802 59339
rect 238502 59338 238802 59339
rect 256502 59338 256802 59339
rect 274502 59338 274802 59339
rect 294540 59338 294840 59339
rect -3348 59327 295310 59338
rect -3348 59209 -2787 59327
rect -2669 59209 4593 59327
rect 4711 59209 22593 59327
rect 22711 59209 40593 59327
rect 40711 59209 58593 59327
rect 58711 59209 76593 59327
rect 76711 59209 94593 59327
rect 94711 59209 112593 59327
rect 112711 59209 130593 59327
rect 130711 59209 148593 59327
rect 148711 59209 166593 59327
rect 166711 59209 184593 59327
rect 184711 59209 202593 59327
rect 202711 59209 220593 59327
rect 220711 59209 238593 59327
rect 238711 59209 256593 59327
rect 256711 59209 274593 59327
rect 274711 59209 294631 59327
rect 294749 59209 295310 59327
rect -3348 59167 295310 59209
rect -3348 59049 -2787 59167
rect -2669 59049 4593 59167
rect 4711 59049 22593 59167
rect 22711 59049 40593 59167
rect 40711 59049 58593 59167
rect 58711 59049 76593 59167
rect 76711 59049 94593 59167
rect 94711 59049 112593 59167
rect 112711 59049 130593 59167
rect 130711 59049 148593 59167
rect 148711 59049 166593 59167
rect 166711 59049 184593 59167
rect 184711 59049 202593 59167
rect 202711 59049 220593 59167
rect 220711 59049 238593 59167
rect 238711 59049 256593 59167
rect 256711 59049 274593 59167
rect 274711 59049 294631 59167
rect 294749 59049 295310 59167
rect -3348 59038 295310 59049
rect -2878 59037 -2578 59038
rect 4502 59037 4802 59038
rect 22502 59037 22802 59038
rect 40502 59037 40802 59038
rect 58502 59037 58802 59038
rect 76502 59037 76802 59038
rect 94502 59037 94802 59038
rect 112502 59037 112802 59038
rect 130502 59037 130802 59038
rect 148502 59037 148802 59038
rect 166502 59037 166802 59038
rect 184502 59037 184802 59038
rect 202502 59037 202802 59038
rect 220502 59037 220802 59038
rect 238502 59037 238802 59038
rect 256502 59037 256802 59038
rect 274502 59037 274802 59038
rect 294540 59037 294840 59038
rect -1938 57538 -1638 57539
rect 2702 57538 3002 57539
rect 20702 57538 21002 57539
rect 38702 57538 39002 57539
rect 56702 57538 57002 57539
rect 74702 57538 75002 57539
rect 92702 57538 93002 57539
rect 110702 57538 111002 57539
rect 128702 57538 129002 57539
rect 146702 57538 147002 57539
rect 164702 57538 165002 57539
rect 182702 57538 183002 57539
rect 200702 57538 201002 57539
rect 218702 57538 219002 57539
rect 236702 57538 237002 57539
rect 254702 57538 255002 57539
rect 272702 57538 273002 57539
rect 290702 57538 291002 57539
rect 293600 57538 293900 57539
rect -2408 57527 294370 57538
rect -2408 57409 -1847 57527
rect -1729 57409 2793 57527
rect 2911 57409 20793 57527
rect 20911 57409 38793 57527
rect 38911 57409 56793 57527
rect 56911 57409 74793 57527
rect 74911 57409 92793 57527
rect 92911 57409 110793 57527
rect 110911 57409 128793 57527
rect 128911 57409 146793 57527
rect 146911 57409 164793 57527
rect 164911 57409 182793 57527
rect 182911 57409 200793 57527
rect 200911 57409 218793 57527
rect 218911 57409 236793 57527
rect 236911 57409 254793 57527
rect 254911 57409 272793 57527
rect 272911 57409 290793 57527
rect 290911 57409 293691 57527
rect 293809 57409 294370 57527
rect -2408 57367 294370 57409
rect -2408 57249 -1847 57367
rect -1729 57249 2793 57367
rect 2911 57249 20793 57367
rect 20911 57249 38793 57367
rect 38911 57249 56793 57367
rect 56911 57249 74793 57367
rect 74911 57249 92793 57367
rect 92911 57249 110793 57367
rect 110911 57249 128793 57367
rect 128911 57249 146793 57367
rect 146911 57249 164793 57367
rect 164911 57249 182793 57367
rect 182911 57249 200793 57367
rect 200911 57249 218793 57367
rect 218911 57249 236793 57367
rect 236911 57249 254793 57367
rect 254911 57249 272793 57367
rect 272911 57249 290793 57367
rect 290911 57249 293691 57367
rect 293809 57249 294370 57367
rect -2408 57238 294370 57249
rect -1938 57237 -1638 57238
rect 2702 57237 3002 57238
rect 20702 57237 21002 57238
rect 38702 57237 39002 57238
rect 56702 57237 57002 57238
rect 74702 57237 75002 57238
rect 92702 57237 93002 57238
rect 110702 57237 111002 57238
rect 128702 57237 129002 57238
rect 146702 57237 147002 57238
rect 164702 57237 165002 57238
rect 182702 57237 183002 57238
rect 200702 57237 201002 57238
rect 218702 57237 219002 57238
rect 236702 57237 237002 57238
rect 254702 57237 255002 57238
rect 272702 57237 273002 57238
rect 290702 57237 291002 57238
rect 293600 57237 293900 57238
rect -998 55738 -698 55739
rect 902 55738 1202 55739
rect 18902 55738 19202 55739
rect 36902 55738 37202 55739
rect 54902 55738 55202 55739
rect 72902 55738 73202 55739
rect 90902 55738 91202 55739
rect 108902 55738 109202 55739
rect 126902 55738 127202 55739
rect 144902 55738 145202 55739
rect 162902 55738 163202 55739
rect 180902 55738 181202 55739
rect 198902 55738 199202 55739
rect 216902 55738 217202 55739
rect 234902 55738 235202 55739
rect 252902 55738 253202 55739
rect 270902 55738 271202 55739
rect 288902 55738 289202 55739
rect 292660 55738 292960 55739
rect -1468 55727 293430 55738
rect -1468 55609 -907 55727
rect -789 55609 993 55727
rect 1111 55609 18993 55727
rect 19111 55609 36993 55727
rect 37111 55609 54993 55727
rect 55111 55609 72993 55727
rect 73111 55609 90993 55727
rect 91111 55609 108993 55727
rect 109111 55609 126993 55727
rect 127111 55609 144993 55727
rect 145111 55609 162993 55727
rect 163111 55609 180993 55727
rect 181111 55609 198993 55727
rect 199111 55609 216993 55727
rect 217111 55609 234993 55727
rect 235111 55609 252993 55727
rect 253111 55609 270993 55727
rect 271111 55609 288993 55727
rect 289111 55609 292751 55727
rect 292869 55609 293430 55727
rect -1468 55567 293430 55609
rect -1468 55449 -907 55567
rect -789 55449 993 55567
rect 1111 55449 18993 55567
rect 19111 55449 36993 55567
rect 37111 55449 54993 55567
rect 55111 55449 72993 55567
rect 73111 55449 90993 55567
rect 91111 55449 108993 55567
rect 109111 55449 126993 55567
rect 127111 55449 144993 55567
rect 145111 55449 162993 55567
rect 163111 55449 180993 55567
rect 181111 55449 198993 55567
rect 199111 55449 216993 55567
rect 217111 55449 234993 55567
rect 235111 55449 252993 55567
rect 253111 55449 270993 55567
rect 271111 55449 288993 55567
rect 289111 55449 292751 55567
rect 292869 55449 293430 55567
rect -1468 55438 293430 55449
rect -998 55437 -698 55438
rect 902 55437 1202 55438
rect 18902 55437 19202 55438
rect 36902 55437 37202 55438
rect 54902 55437 55202 55438
rect 72902 55437 73202 55438
rect 90902 55437 91202 55438
rect 108902 55437 109202 55438
rect 126902 55437 127202 55438
rect 144902 55437 145202 55438
rect 162902 55437 163202 55438
rect 180902 55437 181202 55438
rect 198902 55437 199202 55438
rect 216902 55437 217202 55438
rect 234902 55437 235202 55438
rect 252902 55437 253202 55438
rect 270902 55437 271202 55438
rect 288902 55437 289202 55438
rect 292660 55437 292960 55438
rect -4288 52138 -3988 52139
rect 15302 52138 15602 52139
rect 33302 52138 33602 52139
rect 51302 52138 51602 52139
rect 69302 52138 69602 52139
rect 87302 52138 87602 52139
rect 105302 52138 105602 52139
rect 123302 52138 123602 52139
rect 141302 52138 141602 52139
rect 159302 52138 159602 52139
rect 177302 52138 177602 52139
rect 195302 52138 195602 52139
rect 213302 52138 213602 52139
rect 231302 52138 231602 52139
rect 249302 52138 249602 52139
rect 267302 52138 267602 52139
rect 285302 52138 285602 52139
rect 295950 52138 296250 52139
rect -4288 52127 296250 52138
rect -4288 52009 -4197 52127
rect -4079 52009 15393 52127
rect 15511 52009 33393 52127
rect 33511 52009 51393 52127
rect 51511 52009 69393 52127
rect 69511 52009 87393 52127
rect 87511 52009 105393 52127
rect 105511 52009 123393 52127
rect 123511 52009 141393 52127
rect 141511 52009 159393 52127
rect 159511 52009 177393 52127
rect 177511 52009 195393 52127
rect 195511 52009 213393 52127
rect 213511 52009 231393 52127
rect 231511 52009 249393 52127
rect 249511 52009 267393 52127
rect 267511 52009 285393 52127
rect 285511 52009 296041 52127
rect 296159 52009 296250 52127
rect -4288 51967 296250 52009
rect -4288 51849 -4197 51967
rect -4079 51849 15393 51967
rect 15511 51849 33393 51967
rect 33511 51849 51393 51967
rect 51511 51849 69393 51967
rect 69511 51849 87393 51967
rect 87511 51849 105393 51967
rect 105511 51849 123393 51967
rect 123511 51849 141393 51967
rect 141511 51849 159393 51967
rect 159511 51849 177393 51967
rect 177511 51849 195393 51967
rect 195511 51849 213393 51967
rect 213511 51849 231393 51967
rect 231511 51849 249393 51967
rect 249511 51849 267393 51967
rect 267511 51849 285393 51967
rect 285511 51849 296041 51967
rect 296159 51849 296250 51967
rect -4288 51838 296250 51849
rect -4288 51837 -3988 51838
rect 15302 51837 15602 51838
rect 33302 51837 33602 51838
rect 51302 51837 51602 51838
rect 69302 51837 69602 51838
rect 87302 51837 87602 51838
rect 105302 51837 105602 51838
rect 123302 51837 123602 51838
rect 141302 51837 141602 51838
rect 159302 51837 159602 51838
rect 177302 51837 177602 51838
rect 195302 51837 195602 51838
rect 213302 51837 213602 51838
rect 231302 51837 231602 51838
rect 249302 51837 249602 51838
rect 267302 51837 267602 51838
rect 285302 51837 285602 51838
rect 295950 51837 296250 51838
rect -3348 50338 -3048 50339
rect 13502 50338 13802 50339
rect 31502 50338 31802 50339
rect 49502 50338 49802 50339
rect 67502 50338 67802 50339
rect 85502 50338 85802 50339
rect 103502 50338 103802 50339
rect 121502 50338 121802 50339
rect 139502 50338 139802 50339
rect 157502 50338 157802 50339
rect 175502 50338 175802 50339
rect 193502 50338 193802 50339
rect 211502 50338 211802 50339
rect 229502 50338 229802 50339
rect 247502 50338 247802 50339
rect 265502 50338 265802 50339
rect 283502 50338 283802 50339
rect 295010 50338 295310 50339
rect -3348 50327 295310 50338
rect -3348 50209 -3257 50327
rect -3139 50209 13593 50327
rect 13711 50209 31593 50327
rect 31711 50209 49593 50327
rect 49711 50209 67593 50327
rect 67711 50209 85593 50327
rect 85711 50209 103593 50327
rect 103711 50209 121593 50327
rect 121711 50209 139593 50327
rect 139711 50209 157593 50327
rect 157711 50209 175593 50327
rect 175711 50209 193593 50327
rect 193711 50209 211593 50327
rect 211711 50209 229593 50327
rect 229711 50209 247593 50327
rect 247711 50209 265593 50327
rect 265711 50209 283593 50327
rect 283711 50209 295101 50327
rect 295219 50209 295310 50327
rect -3348 50167 295310 50209
rect -3348 50049 -3257 50167
rect -3139 50049 13593 50167
rect 13711 50049 31593 50167
rect 31711 50049 49593 50167
rect 49711 50049 67593 50167
rect 67711 50049 85593 50167
rect 85711 50049 103593 50167
rect 103711 50049 121593 50167
rect 121711 50049 139593 50167
rect 139711 50049 157593 50167
rect 157711 50049 175593 50167
rect 175711 50049 193593 50167
rect 193711 50049 211593 50167
rect 211711 50049 229593 50167
rect 229711 50049 247593 50167
rect 247711 50049 265593 50167
rect 265711 50049 283593 50167
rect 283711 50049 295101 50167
rect 295219 50049 295310 50167
rect -3348 50038 295310 50049
rect -3348 50037 -3048 50038
rect 13502 50037 13802 50038
rect 31502 50037 31802 50038
rect 49502 50037 49802 50038
rect 67502 50037 67802 50038
rect 85502 50037 85802 50038
rect 103502 50037 103802 50038
rect 121502 50037 121802 50038
rect 139502 50037 139802 50038
rect 157502 50037 157802 50038
rect 175502 50037 175802 50038
rect 193502 50037 193802 50038
rect 211502 50037 211802 50038
rect 229502 50037 229802 50038
rect 247502 50037 247802 50038
rect 265502 50037 265802 50038
rect 283502 50037 283802 50038
rect 295010 50037 295310 50038
rect -2408 48538 -2108 48539
rect 11702 48538 12002 48539
rect 29702 48538 30002 48539
rect 47702 48538 48002 48539
rect 65702 48538 66002 48539
rect 83702 48538 84002 48539
rect 101702 48538 102002 48539
rect 119702 48538 120002 48539
rect 137702 48538 138002 48539
rect 155702 48538 156002 48539
rect 173702 48538 174002 48539
rect 191702 48538 192002 48539
rect 209702 48538 210002 48539
rect 227702 48538 228002 48539
rect 245702 48538 246002 48539
rect 263702 48538 264002 48539
rect 281702 48538 282002 48539
rect 294070 48538 294370 48539
rect -2408 48527 294370 48538
rect -2408 48409 -2317 48527
rect -2199 48409 11793 48527
rect 11911 48409 29793 48527
rect 29911 48409 47793 48527
rect 47911 48409 65793 48527
rect 65911 48409 83793 48527
rect 83911 48409 101793 48527
rect 101911 48409 119793 48527
rect 119911 48409 137793 48527
rect 137911 48409 155793 48527
rect 155911 48409 173793 48527
rect 173911 48409 191793 48527
rect 191911 48409 209793 48527
rect 209911 48409 227793 48527
rect 227911 48409 245793 48527
rect 245911 48409 263793 48527
rect 263911 48409 281793 48527
rect 281911 48409 294161 48527
rect 294279 48409 294370 48527
rect -2408 48367 294370 48409
rect -2408 48249 -2317 48367
rect -2199 48249 11793 48367
rect 11911 48249 29793 48367
rect 29911 48249 47793 48367
rect 47911 48249 65793 48367
rect 65911 48249 83793 48367
rect 83911 48249 101793 48367
rect 101911 48249 119793 48367
rect 119911 48249 137793 48367
rect 137911 48249 155793 48367
rect 155911 48249 173793 48367
rect 173911 48249 191793 48367
rect 191911 48249 209793 48367
rect 209911 48249 227793 48367
rect 227911 48249 245793 48367
rect 245911 48249 263793 48367
rect 263911 48249 281793 48367
rect 281911 48249 294161 48367
rect 294279 48249 294370 48367
rect -2408 48238 294370 48249
rect -2408 48237 -2108 48238
rect 11702 48237 12002 48238
rect 29702 48237 30002 48238
rect 47702 48237 48002 48238
rect 65702 48237 66002 48238
rect 83702 48237 84002 48238
rect 101702 48237 102002 48238
rect 119702 48237 120002 48238
rect 137702 48237 138002 48238
rect 155702 48237 156002 48238
rect 173702 48237 174002 48238
rect 191702 48237 192002 48238
rect 209702 48237 210002 48238
rect 227702 48237 228002 48238
rect 245702 48237 246002 48238
rect 263702 48237 264002 48238
rect 281702 48237 282002 48238
rect 294070 48237 294370 48238
rect -1468 46738 -1168 46739
rect 9902 46738 10202 46739
rect 27902 46738 28202 46739
rect 45902 46738 46202 46739
rect 63902 46738 64202 46739
rect 81902 46738 82202 46739
rect 99902 46738 100202 46739
rect 117902 46738 118202 46739
rect 135902 46738 136202 46739
rect 153902 46738 154202 46739
rect 171902 46738 172202 46739
rect 189902 46738 190202 46739
rect 207902 46738 208202 46739
rect 225902 46738 226202 46739
rect 243902 46738 244202 46739
rect 261902 46738 262202 46739
rect 279902 46738 280202 46739
rect 293130 46738 293430 46739
rect -1468 46727 293430 46738
rect -1468 46609 -1377 46727
rect -1259 46609 9993 46727
rect 10111 46609 27993 46727
rect 28111 46609 45993 46727
rect 46111 46609 63993 46727
rect 64111 46609 81993 46727
rect 82111 46609 99993 46727
rect 100111 46609 117993 46727
rect 118111 46609 135993 46727
rect 136111 46609 153993 46727
rect 154111 46609 171993 46727
rect 172111 46609 189993 46727
rect 190111 46609 207993 46727
rect 208111 46609 225993 46727
rect 226111 46609 243993 46727
rect 244111 46609 261993 46727
rect 262111 46609 279993 46727
rect 280111 46609 293221 46727
rect 293339 46609 293430 46727
rect -1468 46567 293430 46609
rect -1468 46449 -1377 46567
rect -1259 46449 9993 46567
rect 10111 46449 27993 46567
rect 28111 46449 45993 46567
rect 46111 46449 63993 46567
rect 64111 46449 81993 46567
rect 82111 46449 99993 46567
rect 100111 46449 117993 46567
rect 118111 46449 135993 46567
rect 136111 46449 153993 46567
rect 154111 46449 171993 46567
rect 172111 46449 189993 46567
rect 190111 46449 207993 46567
rect 208111 46449 225993 46567
rect 226111 46449 243993 46567
rect 244111 46449 261993 46567
rect 262111 46449 279993 46567
rect 280111 46449 293221 46567
rect 293339 46449 293430 46567
rect -1468 46438 293430 46449
rect -1468 46437 -1168 46438
rect 9902 46437 10202 46438
rect 27902 46437 28202 46438
rect 45902 46437 46202 46438
rect 63902 46437 64202 46438
rect 81902 46437 82202 46438
rect 99902 46437 100202 46438
rect 117902 46437 118202 46438
rect 135902 46437 136202 46438
rect 153902 46437 154202 46438
rect 171902 46437 172202 46438
rect 189902 46437 190202 46438
rect 207902 46437 208202 46438
rect 225902 46437 226202 46438
rect 243902 46437 244202 46438
rect 261902 46437 262202 46438
rect 279902 46437 280202 46438
rect 293130 46437 293430 46438
rect -3818 43138 -3518 43139
rect 6302 43138 6602 43139
rect 24302 43138 24602 43139
rect 42302 43138 42602 43139
rect 60302 43138 60602 43139
rect 78302 43138 78602 43139
rect 96302 43138 96602 43139
rect 114302 43138 114602 43139
rect 132302 43138 132602 43139
rect 150302 43138 150602 43139
rect 168302 43138 168602 43139
rect 186302 43138 186602 43139
rect 204302 43138 204602 43139
rect 222302 43138 222602 43139
rect 240302 43138 240602 43139
rect 258302 43138 258602 43139
rect 276302 43138 276602 43139
rect 295480 43138 295780 43139
rect -4288 43127 296250 43138
rect -4288 43009 -3727 43127
rect -3609 43009 6393 43127
rect 6511 43009 24393 43127
rect 24511 43009 42393 43127
rect 42511 43009 60393 43127
rect 60511 43009 78393 43127
rect 78511 43009 96393 43127
rect 96511 43009 114393 43127
rect 114511 43009 132393 43127
rect 132511 43009 150393 43127
rect 150511 43009 168393 43127
rect 168511 43009 186393 43127
rect 186511 43009 204393 43127
rect 204511 43009 222393 43127
rect 222511 43009 240393 43127
rect 240511 43009 258393 43127
rect 258511 43009 276393 43127
rect 276511 43009 295571 43127
rect 295689 43009 296250 43127
rect -4288 42967 296250 43009
rect -4288 42849 -3727 42967
rect -3609 42849 6393 42967
rect 6511 42849 24393 42967
rect 24511 42849 42393 42967
rect 42511 42849 60393 42967
rect 60511 42849 78393 42967
rect 78511 42849 96393 42967
rect 96511 42849 114393 42967
rect 114511 42849 132393 42967
rect 132511 42849 150393 42967
rect 150511 42849 168393 42967
rect 168511 42849 186393 42967
rect 186511 42849 204393 42967
rect 204511 42849 222393 42967
rect 222511 42849 240393 42967
rect 240511 42849 258393 42967
rect 258511 42849 276393 42967
rect 276511 42849 295571 42967
rect 295689 42849 296250 42967
rect -4288 42838 296250 42849
rect -3818 42837 -3518 42838
rect 6302 42837 6602 42838
rect 24302 42837 24602 42838
rect 42302 42837 42602 42838
rect 60302 42837 60602 42838
rect 78302 42837 78602 42838
rect 96302 42837 96602 42838
rect 114302 42837 114602 42838
rect 132302 42837 132602 42838
rect 150302 42837 150602 42838
rect 168302 42837 168602 42838
rect 186302 42837 186602 42838
rect 204302 42837 204602 42838
rect 222302 42837 222602 42838
rect 240302 42837 240602 42838
rect 258302 42837 258602 42838
rect 276302 42837 276602 42838
rect 295480 42837 295780 42838
rect -2878 41338 -2578 41339
rect 4502 41338 4802 41339
rect 22502 41338 22802 41339
rect 40502 41338 40802 41339
rect 58502 41338 58802 41339
rect 76502 41338 76802 41339
rect 94502 41338 94802 41339
rect 112502 41338 112802 41339
rect 130502 41338 130802 41339
rect 148502 41338 148802 41339
rect 166502 41338 166802 41339
rect 184502 41338 184802 41339
rect 202502 41338 202802 41339
rect 220502 41338 220802 41339
rect 238502 41338 238802 41339
rect 256502 41338 256802 41339
rect 274502 41338 274802 41339
rect 294540 41338 294840 41339
rect -3348 41327 295310 41338
rect -3348 41209 -2787 41327
rect -2669 41209 4593 41327
rect 4711 41209 22593 41327
rect 22711 41209 40593 41327
rect 40711 41209 58593 41327
rect 58711 41209 76593 41327
rect 76711 41209 94593 41327
rect 94711 41209 112593 41327
rect 112711 41209 130593 41327
rect 130711 41209 148593 41327
rect 148711 41209 166593 41327
rect 166711 41209 184593 41327
rect 184711 41209 202593 41327
rect 202711 41209 220593 41327
rect 220711 41209 238593 41327
rect 238711 41209 256593 41327
rect 256711 41209 274593 41327
rect 274711 41209 294631 41327
rect 294749 41209 295310 41327
rect -3348 41167 295310 41209
rect -3348 41049 -2787 41167
rect -2669 41049 4593 41167
rect 4711 41049 22593 41167
rect 22711 41049 40593 41167
rect 40711 41049 58593 41167
rect 58711 41049 76593 41167
rect 76711 41049 94593 41167
rect 94711 41049 112593 41167
rect 112711 41049 130593 41167
rect 130711 41049 148593 41167
rect 148711 41049 166593 41167
rect 166711 41049 184593 41167
rect 184711 41049 202593 41167
rect 202711 41049 220593 41167
rect 220711 41049 238593 41167
rect 238711 41049 256593 41167
rect 256711 41049 274593 41167
rect 274711 41049 294631 41167
rect 294749 41049 295310 41167
rect -3348 41038 295310 41049
rect -2878 41037 -2578 41038
rect 4502 41037 4802 41038
rect 22502 41037 22802 41038
rect 40502 41037 40802 41038
rect 58502 41037 58802 41038
rect 76502 41037 76802 41038
rect 94502 41037 94802 41038
rect 112502 41037 112802 41038
rect 130502 41037 130802 41038
rect 148502 41037 148802 41038
rect 166502 41037 166802 41038
rect 184502 41037 184802 41038
rect 202502 41037 202802 41038
rect 220502 41037 220802 41038
rect 238502 41037 238802 41038
rect 256502 41037 256802 41038
rect 274502 41037 274802 41038
rect 294540 41037 294840 41038
rect -1938 39538 -1638 39539
rect 2702 39538 3002 39539
rect 20702 39538 21002 39539
rect 38702 39538 39002 39539
rect 56702 39538 57002 39539
rect 74702 39538 75002 39539
rect 92702 39538 93002 39539
rect 110702 39538 111002 39539
rect 128702 39538 129002 39539
rect 146702 39538 147002 39539
rect 164702 39538 165002 39539
rect 182702 39538 183002 39539
rect 200702 39538 201002 39539
rect 218702 39538 219002 39539
rect 236702 39538 237002 39539
rect 254702 39538 255002 39539
rect 272702 39538 273002 39539
rect 290702 39538 291002 39539
rect 293600 39538 293900 39539
rect -2408 39527 294370 39538
rect -2408 39409 -1847 39527
rect -1729 39409 2793 39527
rect 2911 39409 20793 39527
rect 20911 39409 38793 39527
rect 38911 39409 56793 39527
rect 56911 39409 74793 39527
rect 74911 39409 92793 39527
rect 92911 39409 110793 39527
rect 110911 39409 128793 39527
rect 128911 39409 146793 39527
rect 146911 39409 164793 39527
rect 164911 39409 182793 39527
rect 182911 39409 200793 39527
rect 200911 39409 218793 39527
rect 218911 39409 236793 39527
rect 236911 39409 254793 39527
rect 254911 39409 272793 39527
rect 272911 39409 290793 39527
rect 290911 39409 293691 39527
rect 293809 39409 294370 39527
rect -2408 39367 294370 39409
rect -2408 39249 -1847 39367
rect -1729 39249 2793 39367
rect 2911 39249 20793 39367
rect 20911 39249 38793 39367
rect 38911 39249 56793 39367
rect 56911 39249 74793 39367
rect 74911 39249 92793 39367
rect 92911 39249 110793 39367
rect 110911 39249 128793 39367
rect 128911 39249 146793 39367
rect 146911 39249 164793 39367
rect 164911 39249 182793 39367
rect 182911 39249 200793 39367
rect 200911 39249 218793 39367
rect 218911 39249 236793 39367
rect 236911 39249 254793 39367
rect 254911 39249 272793 39367
rect 272911 39249 290793 39367
rect 290911 39249 293691 39367
rect 293809 39249 294370 39367
rect -2408 39238 294370 39249
rect -1938 39237 -1638 39238
rect 2702 39237 3002 39238
rect 20702 39237 21002 39238
rect 38702 39237 39002 39238
rect 56702 39237 57002 39238
rect 74702 39237 75002 39238
rect 92702 39237 93002 39238
rect 110702 39237 111002 39238
rect 128702 39237 129002 39238
rect 146702 39237 147002 39238
rect 164702 39237 165002 39238
rect 182702 39237 183002 39238
rect 200702 39237 201002 39238
rect 218702 39237 219002 39238
rect 236702 39237 237002 39238
rect 254702 39237 255002 39238
rect 272702 39237 273002 39238
rect 290702 39237 291002 39238
rect 293600 39237 293900 39238
rect -998 37738 -698 37739
rect 902 37738 1202 37739
rect 18902 37738 19202 37739
rect 36902 37738 37202 37739
rect 54902 37738 55202 37739
rect 72902 37738 73202 37739
rect 90902 37738 91202 37739
rect 108902 37738 109202 37739
rect 126902 37738 127202 37739
rect 144902 37738 145202 37739
rect 162902 37738 163202 37739
rect 180902 37738 181202 37739
rect 198902 37738 199202 37739
rect 216902 37738 217202 37739
rect 234902 37738 235202 37739
rect 252902 37738 253202 37739
rect 270902 37738 271202 37739
rect 288902 37738 289202 37739
rect 292660 37738 292960 37739
rect -1468 37727 293430 37738
rect -1468 37609 -907 37727
rect -789 37609 993 37727
rect 1111 37609 18993 37727
rect 19111 37609 36993 37727
rect 37111 37609 54993 37727
rect 55111 37609 72993 37727
rect 73111 37609 90993 37727
rect 91111 37609 108993 37727
rect 109111 37609 126993 37727
rect 127111 37609 144993 37727
rect 145111 37609 162993 37727
rect 163111 37609 180993 37727
rect 181111 37609 198993 37727
rect 199111 37609 216993 37727
rect 217111 37609 234993 37727
rect 235111 37609 252993 37727
rect 253111 37609 270993 37727
rect 271111 37609 288993 37727
rect 289111 37609 292751 37727
rect 292869 37609 293430 37727
rect -1468 37567 293430 37609
rect -1468 37449 -907 37567
rect -789 37449 993 37567
rect 1111 37449 18993 37567
rect 19111 37449 36993 37567
rect 37111 37449 54993 37567
rect 55111 37449 72993 37567
rect 73111 37449 90993 37567
rect 91111 37449 108993 37567
rect 109111 37449 126993 37567
rect 127111 37449 144993 37567
rect 145111 37449 162993 37567
rect 163111 37449 180993 37567
rect 181111 37449 198993 37567
rect 199111 37449 216993 37567
rect 217111 37449 234993 37567
rect 235111 37449 252993 37567
rect 253111 37449 270993 37567
rect 271111 37449 288993 37567
rect 289111 37449 292751 37567
rect 292869 37449 293430 37567
rect -1468 37438 293430 37449
rect -998 37437 -698 37438
rect 902 37437 1202 37438
rect 18902 37437 19202 37438
rect 36902 37437 37202 37438
rect 54902 37437 55202 37438
rect 72902 37437 73202 37438
rect 90902 37437 91202 37438
rect 108902 37437 109202 37438
rect 126902 37437 127202 37438
rect 144902 37437 145202 37438
rect 162902 37437 163202 37438
rect 180902 37437 181202 37438
rect 198902 37437 199202 37438
rect 216902 37437 217202 37438
rect 234902 37437 235202 37438
rect 252902 37437 253202 37438
rect 270902 37437 271202 37438
rect 288902 37437 289202 37438
rect 292660 37437 292960 37438
rect -4288 34138 -3988 34139
rect 15302 34138 15602 34139
rect 33302 34138 33602 34139
rect 51302 34138 51602 34139
rect 69302 34138 69602 34139
rect 87302 34138 87602 34139
rect 105302 34138 105602 34139
rect 123302 34138 123602 34139
rect 141302 34138 141602 34139
rect 159302 34138 159602 34139
rect 177302 34138 177602 34139
rect 195302 34138 195602 34139
rect 213302 34138 213602 34139
rect 231302 34138 231602 34139
rect 249302 34138 249602 34139
rect 267302 34138 267602 34139
rect 285302 34138 285602 34139
rect 295950 34138 296250 34139
rect -4288 34127 296250 34138
rect -4288 34009 -4197 34127
rect -4079 34009 15393 34127
rect 15511 34009 33393 34127
rect 33511 34009 51393 34127
rect 51511 34009 69393 34127
rect 69511 34009 87393 34127
rect 87511 34009 105393 34127
rect 105511 34009 123393 34127
rect 123511 34009 141393 34127
rect 141511 34009 159393 34127
rect 159511 34009 177393 34127
rect 177511 34009 195393 34127
rect 195511 34009 213393 34127
rect 213511 34009 231393 34127
rect 231511 34009 249393 34127
rect 249511 34009 267393 34127
rect 267511 34009 285393 34127
rect 285511 34009 296041 34127
rect 296159 34009 296250 34127
rect -4288 33967 296250 34009
rect -4288 33849 -4197 33967
rect -4079 33849 15393 33967
rect 15511 33849 33393 33967
rect 33511 33849 51393 33967
rect 51511 33849 69393 33967
rect 69511 33849 87393 33967
rect 87511 33849 105393 33967
rect 105511 33849 123393 33967
rect 123511 33849 141393 33967
rect 141511 33849 159393 33967
rect 159511 33849 177393 33967
rect 177511 33849 195393 33967
rect 195511 33849 213393 33967
rect 213511 33849 231393 33967
rect 231511 33849 249393 33967
rect 249511 33849 267393 33967
rect 267511 33849 285393 33967
rect 285511 33849 296041 33967
rect 296159 33849 296250 33967
rect -4288 33838 296250 33849
rect -4288 33837 -3988 33838
rect 15302 33837 15602 33838
rect 33302 33837 33602 33838
rect 51302 33837 51602 33838
rect 69302 33837 69602 33838
rect 87302 33837 87602 33838
rect 105302 33837 105602 33838
rect 123302 33837 123602 33838
rect 141302 33837 141602 33838
rect 159302 33837 159602 33838
rect 177302 33837 177602 33838
rect 195302 33837 195602 33838
rect 213302 33837 213602 33838
rect 231302 33837 231602 33838
rect 249302 33837 249602 33838
rect 267302 33837 267602 33838
rect 285302 33837 285602 33838
rect 295950 33837 296250 33838
rect -3348 32338 -3048 32339
rect 13502 32338 13802 32339
rect 31502 32338 31802 32339
rect 49502 32338 49802 32339
rect 67502 32338 67802 32339
rect 85502 32338 85802 32339
rect 103502 32338 103802 32339
rect 121502 32338 121802 32339
rect 139502 32338 139802 32339
rect 157502 32338 157802 32339
rect 175502 32338 175802 32339
rect 193502 32338 193802 32339
rect 211502 32338 211802 32339
rect 229502 32338 229802 32339
rect 247502 32338 247802 32339
rect 265502 32338 265802 32339
rect 283502 32338 283802 32339
rect 295010 32338 295310 32339
rect -3348 32327 295310 32338
rect -3348 32209 -3257 32327
rect -3139 32209 13593 32327
rect 13711 32209 31593 32327
rect 31711 32209 49593 32327
rect 49711 32209 67593 32327
rect 67711 32209 85593 32327
rect 85711 32209 103593 32327
rect 103711 32209 121593 32327
rect 121711 32209 139593 32327
rect 139711 32209 157593 32327
rect 157711 32209 175593 32327
rect 175711 32209 193593 32327
rect 193711 32209 211593 32327
rect 211711 32209 229593 32327
rect 229711 32209 247593 32327
rect 247711 32209 265593 32327
rect 265711 32209 283593 32327
rect 283711 32209 295101 32327
rect 295219 32209 295310 32327
rect -3348 32167 295310 32209
rect -3348 32049 -3257 32167
rect -3139 32049 13593 32167
rect 13711 32049 31593 32167
rect 31711 32049 49593 32167
rect 49711 32049 67593 32167
rect 67711 32049 85593 32167
rect 85711 32049 103593 32167
rect 103711 32049 121593 32167
rect 121711 32049 139593 32167
rect 139711 32049 157593 32167
rect 157711 32049 175593 32167
rect 175711 32049 193593 32167
rect 193711 32049 211593 32167
rect 211711 32049 229593 32167
rect 229711 32049 247593 32167
rect 247711 32049 265593 32167
rect 265711 32049 283593 32167
rect 283711 32049 295101 32167
rect 295219 32049 295310 32167
rect -3348 32038 295310 32049
rect -3348 32037 -3048 32038
rect 13502 32037 13802 32038
rect 31502 32037 31802 32038
rect 49502 32037 49802 32038
rect 67502 32037 67802 32038
rect 85502 32037 85802 32038
rect 103502 32037 103802 32038
rect 121502 32037 121802 32038
rect 139502 32037 139802 32038
rect 157502 32037 157802 32038
rect 175502 32037 175802 32038
rect 193502 32037 193802 32038
rect 211502 32037 211802 32038
rect 229502 32037 229802 32038
rect 247502 32037 247802 32038
rect 265502 32037 265802 32038
rect 283502 32037 283802 32038
rect 295010 32037 295310 32038
rect -2408 30538 -2108 30539
rect 11702 30538 12002 30539
rect 29702 30538 30002 30539
rect 47702 30538 48002 30539
rect 65702 30538 66002 30539
rect 83702 30538 84002 30539
rect 101702 30538 102002 30539
rect 119702 30538 120002 30539
rect 137702 30538 138002 30539
rect 155702 30538 156002 30539
rect 173702 30538 174002 30539
rect 191702 30538 192002 30539
rect 209702 30538 210002 30539
rect 227702 30538 228002 30539
rect 245702 30538 246002 30539
rect 263702 30538 264002 30539
rect 281702 30538 282002 30539
rect 294070 30538 294370 30539
rect -2408 30527 294370 30538
rect -2408 30409 -2317 30527
rect -2199 30409 11793 30527
rect 11911 30409 29793 30527
rect 29911 30409 47793 30527
rect 47911 30409 65793 30527
rect 65911 30409 83793 30527
rect 83911 30409 101793 30527
rect 101911 30409 119793 30527
rect 119911 30409 137793 30527
rect 137911 30409 155793 30527
rect 155911 30409 173793 30527
rect 173911 30409 191793 30527
rect 191911 30409 209793 30527
rect 209911 30409 227793 30527
rect 227911 30409 245793 30527
rect 245911 30409 263793 30527
rect 263911 30409 281793 30527
rect 281911 30409 294161 30527
rect 294279 30409 294370 30527
rect -2408 30367 294370 30409
rect -2408 30249 -2317 30367
rect -2199 30249 11793 30367
rect 11911 30249 29793 30367
rect 29911 30249 47793 30367
rect 47911 30249 65793 30367
rect 65911 30249 83793 30367
rect 83911 30249 101793 30367
rect 101911 30249 119793 30367
rect 119911 30249 137793 30367
rect 137911 30249 155793 30367
rect 155911 30249 173793 30367
rect 173911 30249 191793 30367
rect 191911 30249 209793 30367
rect 209911 30249 227793 30367
rect 227911 30249 245793 30367
rect 245911 30249 263793 30367
rect 263911 30249 281793 30367
rect 281911 30249 294161 30367
rect 294279 30249 294370 30367
rect -2408 30238 294370 30249
rect -2408 30237 -2108 30238
rect 11702 30237 12002 30238
rect 29702 30237 30002 30238
rect 47702 30237 48002 30238
rect 65702 30237 66002 30238
rect 83702 30237 84002 30238
rect 101702 30237 102002 30238
rect 119702 30237 120002 30238
rect 137702 30237 138002 30238
rect 155702 30237 156002 30238
rect 173702 30237 174002 30238
rect 191702 30237 192002 30238
rect 209702 30237 210002 30238
rect 227702 30237 228002 30238
rect 245702 30237 246002 30238
rect 263702 30237 264002 30238
rect 281702 30237 282002 30238
rect 294070 30237 294370 30238
rect -1468 28738 -1168 28739
rect 9902 28738 10202 28739
rect 27902 28738 28202 28739
rect 45902 28738 46202 28739
rect 63902 28738 64202 28739
rect 81902 28738 82202 28739
rect 99902 28738 100202 28739
rect 117902 28738 118202 28739
rect 135902 28738 136202 28739
rect 153902 28738 154202 28739
rect 171902 28738 172202 28739
rect 189902 28738 190202 28739
rect 207902 28738 208202 28739
rect 225902 28738 226202 28739
rect 243902 28738 244202 28739
rect 261902 28738 262202 28739
rect 279902 28738 280202 28739
rect 293130 28738 293430 28739
rect -1468 28727 293430 28738
rect -1468 28609 -1377 28727
rect -1259 28609 9993 28727
rect 10111 28609 27993 28727
rect 28111 28609 45993 28727
rect 46111 28609 63993 28727
rect 64111 28609 81993 28727
rect 82111 28609 99993 28727
rect 100111 28609 117993 28727
rect 118111 28609 135993 28727
rect 136111 28609 153993 28727
rect 154111 28609 171993 28727
rect 172111 28609 189993 28727
rect 190111 28609 207993 28727
rect 208111 28609 225993 28727
rect 226111 28609 243993 28727
rect 244111 28609 261993 28727
rect 262111 28609 279993 28727
rect 280111 28609 293221 28727
rect 293339 28609 293430 28727
rect -1468 28567 293430 28609
rect -1468 28449 -1377 28567
rect -1259 28449 9993 28567
rect 10111 28449 27993 28567
rect 28111 28449 45993 28567
rect 46111 28449 63993 28567
rect 64111 28449 81993 28567
rect 82111 28449 99993 28567
rect 100111 28449 117993 28567
rect 118111 28449 135993 28567
rect 136111 28449 153993 28567
rect 154111 28449 171993 28567
rect 172111 28449 189993 28567
rect 190111 28449 207993 28567
rect 208111 28449 225993 28567
rect 226111 28449 243993 28567
rect 244111 28449 261993 28567
rect 262111 28449 279993 28567
rect 280111 28449 293221 28567
rect 293339 28449 293430 28567
rect -1468 28438 293430 28449
rect -1468 28437 -1168 28438
rect 9902 28437 10202 28438
rect 27902 28437 28202 28438
rect 45902 28437 46202 28438
rect 63902 28437 64202 28438
rect 81902 28437 82202 28438
rect 99902 28437 100202 28438
rect 117902 28437 118202 28438
rect 135902 28437 136202 28438
rect 153902 28437 154202 28438
rect 171902 28437 172202 28438
rect 189902 28437 190202 28438
rect 207902 28437 208202 28438
rect 225902 28437 226202 28438
rect 243902 28437 244202 28438
rect 261902 28437 262202 28438
rect 279902 28437 280202 28438
rect 293130 28437 293430 28438
rect -3818 25138 -3518 25139
rect 6302 25138 6602 25139
rect 24302 25138 24602 25139
rect 42302 25138 42602 25139
rect 60302 25138 60602 25139
rect 78302 25138 78602 25139
rect 96302 25138 96602 25139
rect 114302 25138 114602 25139
rect 132302 25138 132602 25139
rect 150302 25138 150602 25139
rect 168302 25138 168602 25139
rect 186302 25138 186602 25139
rect 204302 25138 204602 25139
rect 222302 25138 222602 25139
rect 240302 25138 240602 25139
rect 258302 25138 258602 25139
rect 276302 25138 276602 25139
rect 295480 25138 295780 25139
rect -4288 25127 296250 25138
rect -4288 25009 -3727 25127
rect -3609 25009 6393 25127
rect 6511 25009 24393 25127
rect 24511 25009 42393 25127
rect 42511 25009 60393 25127
rect 60511 25009 78393 25127
rect 78511 25009 96393 25127
rect 96511 25009 114393 25127
rect 114511 25009 132393 25127
rect 132511 25009 150393 25127
rect 150511 25009 168393 25127
rect 168511 25009 186393 25127
rect 186511 25009 204393 25127
rect 204511 25009 222393 25127
rect 222511 25009 240393 25127
rect 240511 25009 258393 25127
rect 258511 25009 276393 25127
rect 276511 25009 295571 25127
rect 295689 25009 296250 25127
rect -4288 24967 296250 25009
rect -4288 24849 -3727 24967
rect -3609 24849 6393 24967
rect 6511 24849 24393 24967
rect 24511 24849 42393 24967
rect 42511 24849 60393 24967
rect 60511 24849 78393 24967
rect 78511 24849 96393 24967
rect 96511 24849 114393 24967
rect 114511 24849 132393 24967
rect 132511 24849 150393 24967
rect 150511 24849 168393 24967
rect 168511 24849 186393 24967
rect 186511 24849 204393 24967
rect 204511 24849 222393 24967
rect 222511 24849 240393 24967
rect 240511 24849 258393 24967
rect 258511 24849 276393 24967
rect 276511 24849 295571 24967
rect 295689 24849 296250 24967
rect -4288 24838 296250 24849
rect -3818 24837 -3518 24838
rect 6302 24837 6602 24838
rect 24302 24837 24602 24838
rect 42302 24837 42602 24838
rect 60302 24837 60602 24838
rect 78302 24837 78602 24838
rect 96302 24837 96602 24838
rect 114302 24837 114602 24838
rect 132302 24837 132602 24838
rect 150302 24837 150602 24838
rect 168302 24837 168602 24838
rect 186302 24837 186602 24838
rect 204302 24837 204602 24838
rect 222302 24837 222602 24838
rect 240302 24837 240602 24838
rect 258302 24837 258602 24838
rect 276302 24837 276602 24838
rect 295480 24837 295780 24838
rect -2878 23338 -2578 23339
rect 4502 23338 4802 23339
rect 22502 23338 22802 23339
rect 40502 23338 40802 23339
rect 58502 23338 58802 23339
rect 76502 23338 76802 23339
rect 94502 23338 94802 23339
rect 112502 23338 112802 23339
rect 130502 23338 130802 23339
rect 148502 23338 148802 23339
rect 166502 23338 166802 23339
rect 184502 23338 184802 23339
rect 202502 23338 202802 23339
rect 220502 23338 220802 23339
rect 238502 23338 238802 23339
rect 256502 23338 256802 23339
rect 274502 23338 274802 23339
rect 294540 23338 294840 23339
rect -3348 23327 295310 23338
rect -3348 23209 -2787 23327
rect -2669 23209 4593 23327
rect 4711 23209 22593 23327
rect 22711 23209 40593 23327
rect 40711 23209 58593 23327
rect 58711 23209 76593 23327
rect 76711 23209 94593 23327
rect 94711 23209 112593 23327
rect 112711 23209 130593 23327
rect 130711 23209 148593 23327
rect 148711 23209 166593 23327
rect 166711 23209 184593 23327
rect 184711 23209 202593 23327
rect 202711 23209 220593 23327
rect 220711 23209 238593 23327
rect 238711 23209 256593 23327
rect 256711 23209 274593 23327
rect 274711 23209 294631 23327
rect 294749 23209 295310 23327
rect -3348 23167 295310 23209
rect -3348 23049 -2787 23167
rect -2669 23049 4593 23167
rect 4711 23049 22593 23167
rect 22711 23049 40593 23167
rect 40711 23049 58593 23167
rect 58711 23049 76593 23167
rect 76711 23049 94593 23167
rect 94711 23049 112593 23167
rect 112711 23049 130593 23167
rect 130711 23049 148593 23167
rect 148711 23049 166593 23167
rect 166711 23049 184593 23167
rect 184711 23049 202593 23167
rect 202711 23049 220593 23167
rect 220711 23049 238593 23167
rect 238711 23049 256593 23167
rect 256711 23049 274593 23167
rect 274711 23049 294631 23167
rect 294749 23049 295310 23167
rect -3348 23038 295310 23049
rect -2878 23037 -2578 23038
rect 4502 23037 4802 23038
rect 22502 23037 22802 23038
rect 40502 23037 40802 23038
rect 58502 23037 58802 23038
rect 76502 23037 76802 23038
rect 94502 23037 94802 23038
rect 112502 23037 112802 23038
rect 130502 23037 130802 23038
rect 148502 23037 148802 23038
rect 166502 23037 166802 23038
rect 184502 23037 184802 23038
rect 202502 23037 202802 23038
rect 220502 23037 220802 23038
rect 238502 23037 238802 23038
rect 256502 23037 256802 23038
rect 274502 23037 274802 23038
rect 294540 23037 294840 23038
rect -1938 21538 -1638 21539
rect 2702 21538 3002 21539
rect 20702 21538 21002 21539
rect 38702 21538 39002 21539
rect 56702 21538 57002 21539
rect 74702 21538 75002 21539
rect 92702 21538 93002 21539
rect 110702 21538 111002 21539
rect 128702 21538 129002 21539
rect 146702 21538 147002 21539
rect 164702 21538 165002 21539
rect 182702 21538 183002 21539
rect 200702 21538 201002 21539
rect 218702 21538 219002 21539
rect 236702 21538 237002 21539
rect 254702 21538 255002 21539
rect 272702 21538 273002 21539
rect 290702 21538 291002 21539
rect 293600 21538 293900 21539
rect -2408 21527 294370 21538
rect -2408 21409 -1847 21527
rect -1729 21409 2793 21527
rect 2911 21409 20793 21527
rect 20911 21409 38793 21527
rect 38911 21409 56793 21527
rect 56911 21409 74793 21527
rect 74911 21409 92793 21527
rect 92911 21409 110793 21527
rect 110911 21409 128793 21527
rect 128911 21409 146793 21527
rect 146911 21409 164793 21527
rect 164911 21409 182793 21527
rect 182911 21409 200793 21527
rect 200911 21409 218793 21527
rect 218911 21409 236793 21527
rect 236911 21409 254793 21527
rect 254911 21409 272793 21527
rect 272911 21409 290793 21527
rect 290911 21409 293691 21527
rect 293809 21409 294370 21527
rect -2408 21367 294370 21409
rect -2408 21249 -1847 21367
rect -1729 21249 2793 21367
rect 2911 21249 20793 21367
rect 20911 21249 38793 21367
rect 38911 21249 56793 21367
rect 56911 21249 74793 21367
rect 74911 21249 92793 21367
rect 92911 21249 110793 21367
rect 110911 21249 128793 21367
rect 128911 21249 146793 21367
rect 146911 21249 164793 21367
rect 164911 21249 182793 21367
rect 182911 21249 200793 21367
rect 200911 21249 218793 21367
rect 218911 21249 236793 21367
rect 236911 21249 254793 21367
rect 254911 21249 272793 21367
rect 272911 21249 290793 21367
rect 290911 21249 293691 21367
rect 293809 21249 294370 21367
rect -2408 21238 294370 21249
rect -1938 21237 -1638 21238
rect 2702 21237 3002 21238
rect 20702 21237 21002 21238
rect 38702 21237 39002 21238
rect 56702 21237 57002 21238
rect 74702 21237 75002 21238
rect 92702 21237 93002 21238
rect 110702 21237 111002 21238
rect 128702 21237 129002 21238
rect 146702 21237 147002 21238
rect 164702 21237 165002 21238
rect 182702 21237 183002 21238
rect 200702 21237 201002 21238
rect 218702 21237 219002 21238
rect 236702 21237 237002 21238
rect 254702 21237 255002 21238
rect 272702 21237 273002 21238
rect 290702 21237 291002 21238
rect 293600 21237 293900 21238
rect -998 19738 -698 19739
rect 902 19738 1202 19739
rect 18902 19738 19202 19739
rect 36902 19738 37202 19739
rect 54902 19738 55202 19739
rect 72902 19738 73202 19739
rect 90902 19738 91202 19739
rect 108902 19738 109202 19739
rect 126902 19738 127202 19739
rect 144902 19738 145202 19739
rect 162902 19738 163202 19739
rect 180902 19738 181202 19739
rect 198902 19738 199202 19739
rect 216902 19738 217202 19739
rect 234902 19738 235202 19739
rect 252902 19738 253202 19739
rect 270902 19738 271202 19739
rect 288902 19738 289202 19739
rect 292660 19738 292960 19739
rect -1468 19727 293430 19738
rect -1468 19609 -907 19727
rect -789 19609 993 19727
rect 1111 19609 18993 19727
rect 19111 19609 36993 19727
rect 37111 19609 54993 19727
rect 55111 19609 72993 19727
rect 73111 19609 90993 19727
rect 91111 19609 108993 19727
rect 109111 19609 126993 19727
rect 127111 19609 144993 19727
rect 145111 19609 162993 19727
rect 163111 19609 180993 19727
rect 181111 19609 198993 19727
rect 199111 19609 216993 19727
rect 217111 19609 234993 19727
rect 235111 19609 252993 19727
rect 253111 19609 270993 19727
rect 271111 19609 288993 19727
rect 289111 19609 292751 19727
rect 292869 19609 293430 19727
rect -1468 19567 293430 19609
rect -1468 19449 -907 19567
rect -789 19449 993 19567
rect 1111 19449 18993 19567
rect 19111 19449 36993 19567
rect 37111 19449 54993 19567
rect 55111 19449 72993 19567
rect 73111 19449 90993 19567
rect 91111 19449 108993 19567
rect 109111 19449 126993 19567
rect 127111 19449 144993 19567
rect 145111 19449 162993 19567
rect 163111 19449 180993 19567
rect 181111 19449 198993 19567
rect 199111 19449 216993 19567
rect 217111 19449 234993 19567
rect 235111 19449 252993 19567
rect 253111 19449 270993 19567
rect 271111 19449 288993 19567
rect 289111 19449 292751 19567
rect 292869 19449 293430 19567
rect -1468 19438 293430 19449
rect -998 19437 -698 19438
rect 902 19437 1202 19438
rect 18902 19437 19202 19438
rect 36902 19437 37202 19438
rect 54902 19437 55202 19438
rect 72902 19437 73202 19438
rect 90902 19437 91202 19438
rect 108902 19437 109202 19438
rect 126902 19437 127202 19438
rect 144902 19437 145202 19438
rect 162902 19437 163202 19438
rect 180902 19437 181202 19438
rect 198902 19437 199202 19438
rect 216902 19437 217202 19438
rect 234902 19437 235202 19438
rect 252902 19437 253202 19438
rect 270902 19437 271202 19438
rect 288902 19437 289202 19438
rect 292660 19437 292960 19438
rect -4288 16138 -3988 16139
rect 15302 16138 15602 16139
rect 33302 16138 33602 16139
rect 51302 16138 51602 16139
rect 69302 16138 69602 16139
rect 87302 16138 87602 16139
rect 105302 16138 105602 16139
rect 123302 16138 123602 16139
rect 141302 16138 141602 16139
rect 159302 16138 159602 16139
rect 177302 16138 177602 16139
rect 195302 16138 195602 16139
rect 213302 16138 213602 16139
rect 231302 16138 231602 16139
rect 249302 16138 249602 16139
rect 267302 16138 267602 16139
rect 285302 16138 285602 16139
rect 295950 16138 296250 16139
rect -4288 16127 296250 16138
rect -4288 16009 -4197 16127
rect -4079 16009 15393 16127
rect 15511 16009 33393 16127
rect 33511 16009 51393 16127
rect 51511 16009 69393 16127
rect 69511 16009 87393 16127
rect 87511 16009 105393 16127
rect 105511 16009 123393 16127
rect 123511 16009 141393 16127
rect 141511 16009 159393 16127
rect 159511 16009 177393 16127
rect 177511 16009 195393 16127
rect 195511 16009 213393 16127
rect 213511 16009 231393 16127
rect 231511 16009 249393 16127
rect 249511 16009 267393 16127
rect 267511 16009 285393 16127
rect 285511 16009 296041 16127
rect 296159 16009 296250 16127
rect -4288 15967 296250 16009
rect -4288 15849 -4197 15967
rect -4079 15849 15393 15967
rect 15511 15849 33393 15967
rect 33511 15849 51393 15967
rect 51511 15849 69393 15967
rect 69511 15849 87393 15967
rect 87511 15849 105393 15967
rect 105511 15849 123393 15967
rect 123511 15849 141393 15967
rect 141511 15849 159393 15967
rect 159511 15849 177393 15967
rect 177511 15849 195393 15967
rect 195511 15849 213393 15967
rect 213511 15849 231393 15967
rect 231511 15849 249393 15967
rect 249511 15849 267393 15967
rect 267511 15849 285393 15967
rect 285511 15849 296041 15967
rect 296159 15849 296250 15967
rect -4288 15838 296250 15849
rect -4288 15837 -3988 15838
rect 15302 15837 15602 15838
rect 33302 15837 33602 15838
rect 51302 15837 51602 15838
rect 69302 15837 69602 15838
rect 87302 15837 87602 15838
rect 105302 15837 105602 15838
rect 123302 15837 123602 15838
rect 141302 15837 141602 15838
rect 159302 15837 159602 15838
rect 177302 15837 177602 15838
rect 195302 15837 195602 15838
rect 213302 15837 213602 15838
rect 231302 15837 231602 15838
rect 249302 15837 249602 15838
rect 267302 15837 267602 15838
rect 285302 15837 285602 15838
rect 295950 15837 296250 15838
rect -3348 14338 -3048 14339
rect 13502 14338 13802 14339
rect 31502 14338 31802 14339
rect 49502 14338 49802 14339
rect 67502 14338 67802 14339
rect 85502 14338 85802 14339
rect 103502 14338 103802 14339
rect 121502 14338 121802 14339
rect 139502 14338 139802 14339
rect 157502 14338 157802 14339
rect 175502 14338 175802 14339
rect 193502 14338 193802 14339
rect 211502 14338 211802 14339
rect 229502 14338 229802 14339
rect 247502 14338 247802 14339
rect 265502 14338 265802 14339
rect 283502 14338 283802 14339
rect 295010 14338 295310 14339
rect -3348 14327 295310 14338
rect -3348 14209 -3257 14327
rect -3139 14209 13593 14327
rect 13711 14209 31593 14327
rect 31711 14209 49593 14327
rect 49711 14209 67593 14327
rect 67711 14209 85593 14327
rect 85711 14209 103593 14327
rect 103711 14209 121593 14327
rect 121711 14209 139593 14327
rect 139711 14209 157593 14327
rect 157711 14209 175593 14327
rect 175711 14209 193593 14327
rect 193711 14209 211593 14327
rect 211711 14209 229593 14327
rect 229711 14209 247593 14327
rect 247711 14209 265593 14327
rect 265711 14209 283593 14327
rect 283711 14209 295101 14327
rect 295219 14209 295310 14327
rect -3348 14167 295310 14209
rect -3348 14049 -3257 14167
rect -3139 14049 13593 14167
rect 13711 14049 31593 14167
rect 31711 14049 49593 14167
rect 49711 14049 67593 14167
rect 67711 14049 85593 14167
rect 85711 14049 103593 14167
rect 103711 14049 121593 14167
rect 121711 14049 139593 14167
rect 139711 14049 157593 14167
rect 157711 14049 175593 14167
rect 175711 14049 193593 14167
rect 193711 14049 211593 14167
rect 211711 14049 229593 14167
rect 229711 14049 247593 14167
rect 247711 14049 265593 14167
rect 265711 14049 283593 14167
rect 283711 14049 295101 14167
rect 295219 14049 295310 14167
rect -3348 14038 295310 14049
rect -3348 14037 -3048 14038
rect 13502 14037 13802 14038
rect 31502 14037 31802 14038
rect 49502 14037 49802 14038
rect 67502 14037 67802 14038
rect 85502 14037 85802 14038
rect 103502 14037 103802 14038
rect 121502 14037 121802 14038
rect 139502 14037 139802 14038
rect 157502 14037 157802 14038
rect 175502 14037 175802 14038
rect 193502 14037 193802 14038
rect 211502 14037 211802 14038
rect 229502 14037 229802 14038
rect 247502 14037 247802 14038
rect 265502 14037 265802 14038
rect 283502 14037 283802 14038
rect 295010 14037 295310 14038
rect -2408 12538 -2108 12539
rect 11702 12538 12002 12539
rect 29702 12538 30002 12539
rect 47702 12538 48002 12539
rect 65702 12538 66002 12539
rect 83702 12538 84002 12539
rect 101702 12538 102002 12539
rect 119702 12538 120002 12539
rect 137702 12538 138002 12539
rect 155702 12538 156002 12539
rect 173702 12538 174002 12539
rect 191702 12538 192002 12539
rect 209702 12538 210002 12539
rect 227702 12538 228002 12539
rect 245702 12538 246002 12539
rect 263702 12538 264002 12539
rect 281702 12538 282002 12539
rect 294070 12538 294370 12539
rect -2408 12527 294370 12538
rect -2408 12409 -2317 12527
rect -2199 12409 11793 12527
rect 11911 12409 29793 12527
rect 29911 12409 47793 12527
rect 47911 12409 65793 12527
rect 65911 12409 83793 12527
rect 83911 12409 101793 12527
rect 101911 12409 119793 12527
rect 119911 12409 137793 12527
rect 137911 12409 155793 12527
rect 155911 12409 173793 12527
rect 173911 12409 191793 12527
rect 191911 12409 209793 12527
rect 209911 12409 227793 12527
rect 227911 12409 245793 12527
rect 245911 12409 263793 12527
rect 263911 12409 281793 12527
rect 281911 12409 294161 12527
rect 294279 12409 294370 12527
rect -2408 12367 294370 12409
rect -2408 12249 -2317 12367
rect -2199 12249 11793 12367
rect 11911 12249 29793 12367
rect 29911 12249 47793 12367
rect 47911 12249 65793 12367
rect 65911 12249 83793 12367
rect 83911 12249 101793 12367
rect 101911 12249 119793 12367
rect 119911 12249 137793 12367
rect 137911 12249 155793 12367
rect 155911 12249 173793 12367
rect 173911 12249 191793 12367
rect 191911 12249 209793 12367
rect 209911 12249 227793 12367
rect 227911 12249 245793 12367
rect 245911 12249 263793 12367
rect 263911 12249 281793 12367
rect 281911 12249 294161 12367
rect 294279 12249 294370 12367
rect -2408 12238 294370 12249
rect -2408 12237 -2108 12238
rect 11702 12237 12002 12238
rect 29702 12237 30002 12238
rect 47702 12237 48002 12238
rect 65702 12237 66002 12238
rect 83702 12237 84002 12238
rect 101702 12237 102002 12238
rect 119702 12237 120002 12238
rect 137702 12237 138002 12238
rect 155702 12237 156002 12238
rect 173702 12237 174002 12238
rect 191702 12237 192002 12238
rect 209702 12237 210002 12238
rect 227702 12237 228002 12238
rect 245702 12237 246002 12238
rect 263702 12237 264002 12238
rect 281702 12237 282002 12238
rect 294070 12237 294370 12238
rect -1468 10738 -1168 10739
rect 9902 10738 10202 10739
rect 27902 10738 28202 10739
rect 45902 10738 46202 10739
rect 63902 10738 64202 10739
rect 81902 10738 82202 10739
rect 99902 10738 100202 10739
rect 117902 10738 118202 10739
rect 135902 10738 136202 10739
rect 153902 10738 154202 10739
rect 171902 10738 172202 10739
rect 189902 10738 190202 10739
rect 207902 10738 208202 10739
rect 225902 10738 226202 10739
rect 243902 10738 244202 10739
rect 261902 10738 262202 10739
rect 279902 10738 280202 10739
rect 293130 10738 293430 10739
rect -1468 10727 293430 10738
rect -1468 10609 -1377 10727
rect -1259 10609 9993 10727
rect 10111 10609 27993 10727
rect 28111 10609 45993 10727
rect 46111 10609 63993 10727
rect 64111 10609 81993 10727
rect 82111 10609 99993 10727
rect 100111 10609 117993 10727
rect 118111 10609 135993 10727
rect 136111 10609 153993 10727
rect 154111 10609 171993 10727
rect 172111 10609 189993 10727
rect 190111 10609 207993 10727
rect 208111 10609 225993 10727
rect 226111 10609 243993 10727
rect 244111 10609 261993 10727
rect 262111 10609 279993 10727
rect 280111 10609 293221 10727
rect 293339 10609 293430 10727
rect -1468 10567 293430 10609
rect -1468 10449 -1377 10567
rect -1259 10449 9993 10567
rect 10111 10449 27993 10567
rect 28111 10449 45993 10567
rect 46111 10449 63993 10567
rect 64111 10449 81993 10567
rect 82111 10449 99993 10567
rect 100111 10449 117993 10567
rect 118111 10449 135993 10567
rect 136111 10449 153993 10567
rect 154111 10449 171993 10567
rect 172111 10449 189993 10567
rect 190111 10449 207993 10567
rect 208111 10449 225993 10567
rect 226111 10449 243993 10567
rect 244111 10449 261993 10567
rect 262111 10449 279993 10567
rect 280111 10449 293221 10567
rect 293339 10449 293430 10567
rect -1468 10438 293430 10449
rect -1468 10437 -1168 10438
rect 9902 10437 10202 10438
rect 27902 10437 28202 10438
rect 45902 10437 46202 10438
rect 63902 10437 64202 10438
rect 81902 10437 82202 10438
rect 99902 10437 100202 10438
rect 117902 10437 118202 10438
rect 135902 10437 136202 10438
rect 153902 10437 154202 10438
rect 171902 10437 172202 10438
rect 189902 10437 190202 10438
rect 207902 10437 208202 10438
rect 225902 10437 226202 10438
rect 243902 10437 244202 10438
rect 261902 10437 262202 10438
rect 279902 10437 280202 10438
rect 293130 10437 293430 10438
rect -3818 7138 -3518 7139
rect 6302 7138 6602 7139
rect 24302 7138 24602 7139
rect 42302 7138 42602 7139
rect 60302 7138 60602 7139
rect 78302 7138 78602 7139
rect 96302 7138 96602 7139
rect 114302 7138 114602 7139
rect 132302 7138 132602 7139
rect 150302 7138 150602 7139
rect 168302 7138 168602 7139
rect 186302 7138 186602 7139
rect 204302 7138 204602 7139
rect 222302 7138 222602 7139
rect 240302 7138 240602 7139
rect 258302 7138 258602 7139
rect 276302 7138 276602 7139
rect 295480 7138 295780 7139
rect -4288 7127 296250 7138
rect -4288 7009 -3727 7127
rect -3609 7009 6393 7127
rect 6511 7009 24393 7127
rect 24511 7009 42393 7127
rect 42511 7009 60393 7127
rect 60511 7009 78393 7127
rect 78511 7009 96393 7127
rect 96511 7009 114393 7127
rect 114511 7009 132393 7127
rect 132511 7009 150393 7127
rect 150511 7009 168393 7127
rect 168511 7009 186393 7127
rect 186511 7009 204393 7127
rect 204511 7009 222393 7127
rect 222511 7009 240393 7127
rect 240511 7009 258393 7127
rect 258511 7009 276393 7127
rect 276511 7009 295571 7127
rect 295689 7009 296250 7127
rect -4288 6967 296250 7009
rect -4288 6849 -3727 6967
rect -3609 6849 6393 6967
rect 6511 6849 24393 6967
rect 24511 6849 42393 6967
rect 42511 6849 60393 6967
rect 60511 6849 78393 6967
rect 78511 6849 96393 6967
rect 96511 6849 114393 6967
rect 114511 6849 132393 6967
rect 132511 6849 150393 6967
rect 150511 6849 168393 6967
rect 168511 6849 186393 6967
rect 186511 6849 204393 6967
rect 204511 6849 222393 6967
rect 222511 6849 240393 6967
rect 240511 6849 258393 6967
rect 258511 6849 276393 6967
rect 276511 6849 295571 6967
rect 295689 6849 296250 6967
rect -4288 6838 296250 6849
rect -3818 6837 -3518 6838
rect 6302 6837 6602 6838
rect 24302 6837 24602 6838
rect 42302 6837 42602 6838
rect 60302 6837 60602 6838
rect 78302 6837 78602 6838
rect 96302 6837 96602 6838
rect 114302 6837 114602 6838
rect 132302 6837 132602 6838
rect 150302 6837 150602 6838
rect 168302 6837 168602 6838
rect 186302 6837 186602 6838
rect 204302 6837 204602 6838
rect 222302 6837 222602 6838
rect 240302 6837 240602 6838
rect 258302 6837 258602 6838
rect 276302 6837 276602 6838
rect 295480 6837 295780 6838
rect -2878 5338 -2578 5339
rect 4502 5338 4802 5339
rect 22502 5338 22802 5339
rect 40502 5338 40802 5339
rect 58502 5338 58802 5339
rect 76502 5338 76802 5339
rect 94502 5338 94802 5339
rect 112502 5338 112802 5339
rect 130502 5338 130802 5339
rect 148502 5338 148802 5339
rect 166502 5338 166802 5339
rect 184502 5338 184802 5339
rect 202502 5338 202802 5339
rect 220502 5338 220802 5339
rect 238502 5338 238802 5339
rect 256502 5338 256802 5339
rect 274502 5338 274802 5339
rect 294540 5338 294840 5339
rect -3348 5327 295310 5338
rect -3348 5209 -2787 5327
rect -2669 5209 4593 5327
rect 4711 5209 22593 5327
rect 22711 5209 40593 5327
rect 40711 5209 58593 5327
rect 58711 5209 76593 5327
rect 76711 5209 94593 5327
rect 94711 5209 112593 5327
rect 112711 5209 130593 5327
rect 130711 5209 148593 5327
rect 148711 5209 166593 5327
rect 166711 5209 184593 5327
rect 184711 5209 202593 5327
rect 202711 5209 220593 5327
rect 220711 5209 238593 5327
rect 238711 5209 256593 5327
rect 256711 5209 274593 5327
rect 274711 5209 294631 5327
rect 294749 5209 295310 5327
rect -3348 5167 295310 5209
rect -3348 5049 -2787 5167
rect -2669 5049 4593 5167
rect 4711 5049 22593 5167
rect 22711 5049 40593 5167
rect 40711 5049 58593 5167
rect 58711 5049 76593 5167
rect 76711 5049 94593 5167
rect 94711 5049 112593 5167
rect 112711 5049 130593 5167
rect 130711 5049 148593 5167
rect 148711 5049 166593 5167
rect 166711 5049 184593 5167
rect 184711 5049 202593 5167
rect 202711 5049 220593 5167
rect 220711 5049 238593 5167
rect 238711 5049 256593 5167
rect 256711 5049 274593 5167
rect 274711 5049 294631 5167
rect 294749 5049 295310 5167
rect -3348 5038 295310 5049
rect -2878 5037 -2578 5038
rect 4502 5037 4802 5038
rect 22502 5037 22802 5038
rect 40502 5037 40802 5038
rect 58502 5037 58802 5038
rect 76502 5037 76802 5038
rect 94502 5037 94802 5038
rect 112502 5037 112802 5038
rect 130502 5037 130802 5038
rect 148502 5037 148802 5038
rect 166502 5037 166802 5038
rect 184502 5037 184802 5038
rect 202502 5037 202802 5038
rect 220502 5037 220802 5038
rect 238502 5037 238802 5038
rect 256502 5037 256802 5038
rect 274502 5037 274802 5038
rect 294540 5037 294840 5038
rect -1938 3538 -1638 3539
rect 2702 3538 3002 3539
rect 20702 3538 21002 3539
rect 38702 3538 39002 3539
rect 56702 3538 57002 3539
rect 74702 3538 75002 3539
rect 92702 3538 93002 3539
rect 110702 3538 111002 3539
rect 128702 3538 129002 3539
rect 146702 3538 147002 3539
rect 164702 3538 165002 3539
rect 182702 3538 183002 3539
rect 200702 3538 201002 3539
rect 218702 3538 219002 3539
rect 236702 3538 237002 3539
rect 254702 3538 255002 3539
rect 272702 3538 273002 3539
rect 290702 3538 291002 3539
rect 293600 3538 293900 3539
rect -2408 3527 294370 3538
rect -2408 3409 -1847 3527
rect -1729 3409 2793 3527
rect 2911 3409 20793 3527
rect 20911 3409 38793 3527
rect 38911 3409 56793 3527
rect 56911 3409 74793 3527
rect 74911 3409 92793 3527
rect 92911 3409 110793 3527
rect 110911 3409 128793 3527
rect 128911 3409 146793 3527
rect 146911 3409 164793 3527
rect 164911 3409 182793 3527
rect 182911 3409 200793 3527
rect 200911 3409 218793 3527
rect 218911 3409 236793 3527
rect 236911 3409 254793 3527
rect 254911 3409 272793 3527
rect 272911 3409 290793 3527
rect 290911 3409 293691 3527
rect 293809 3409 294370 3527
rect -2408 3367 294370 3409
rect -2408 3249 -1847 3367
rect -1729 3249 2793 3367
rect 2911 3249 20793 3367
rect 20911 3249 38793 3367
rect 38911 3249 56793 3367
rect 56911 3249 74793 3367
rect 74911 3249 92793 3367
rect 92911 3249 110793 3367
rect 110911 3249 128793 3367
rect 128911 3249 146793 3367
rect 146911 3249 164793 3367
rect 164911 3249 182793 3367
rect 182911 3249 200793 3367
rect 200911 3249 218793 3367
rect 218911 3249 236793 3367
rect 236911 3249 254793 3367
rect 254911 3249 272793 3367
rect 272911 3249 290793 3367
rect 290911 3249 293691 3367
rect 293809 3249 294370 3367
rect -2408 3238 294370 3249
rect -1938 3237 -1638 3238
rect 2702 3237 3002 3238
rect 20702 3237 21002 3238
rect 38702 3237 39002 3238
rect 56702 3237 57002 3238
rect 74702 3237 75002 3238
rect 92702 3237 93002 3238
rect 110702 3237 111002 3238
rect 128702 3237 129002 3238
rect 146702 3237 147002 3238
rect 164702 3237 165002 3238
rect 182702 3237 183002 3238
rect 200702 3237 201002 3238
rect 218702 3237 219002 3238
rect 236702 3237 237002 3238
rect 254702 3237 255002 3238
rect 272702 3237 273002 3238
rect 290702 3237 291002 3238
rect 293600 3237 293900 3238
rect -998 1738 -698 1739
rect 902 1738 1202 1739
rect 18902 1738 19202 1739
rect 36902 1738 37202 1739
rect 54902 1738 55202 1739
rect 72902 1738 73202 1739
rect 90902 1738 91202 1739
rect 108902 1738 109202 1739
rect 126902 1738 127202 1739
rect 144902 1738 145202 1739
rect 162902 1738 163202 1739
rect 180902 1738 181202 1739
rect 198902 1738 199202 1739
rect 216902 1738 217202 1739
rect 234902 1738 235202 1739
rect 252902 1738 253202 1739
rect 270902 1738 271202 1739
rect 288902 1738 289202 1739
rect 292660 1738 292960 1739
rect -1468 1727 293430 1738
rect -1468 1609 -907 1727
rect -789 1609 993 1727
rect 1111 1609 18993 1727
rect 19111 1609 36993 1727
rect 37111 1609 54993 1727
rect 55111 1609 72993 1727
rect 73111 1609 90993 1727
rect 91111 1609 108993 1727
rect 109111 1609 126993 1727
rect 127111 1609 144993 1727
rect 145111 1609 162993 1727
rect 163111 1609 180993 1727
rect 181111 1609 198993 1727
rect 199111 1609 216993 1727
rect 217111 1609 234993 1727
rect 235111 1609 252993 1727
rect 253111 1609 270993 1727
rect 271111 1609 288993 1727
rect 289111 1609 292751 1727
rect 292869 1609 293430 1727
rect -1468 1567 293430 1609
rect -1468 1449 -907 1567
rect -789 1449 993 1567
rect 1111 1449 18993 1567
rect 19111 1449 36993 1567
rect 37111 1449 54993 1567
rect 55111 1449 72993 1567
rect 73111 1449 90993 1567
rect 91111 1449 108993 1567
rect 109111 1449 126993 1567
rect 127111 1449 144993 1567
rect 145111 1449 162993 1567
rect 163111 1449 180993 1567
rect 181111 1449 198993 1567
rect 199111 1449 216993 1567
rect 217111 1449 234993 1567
rect 235111 1449 252993 1567
rect 253111 1449 270993 1567
rect 271111 1449 288993 1567
rect 289111 1449 292751 1567
rect 292869 1449 293430 1567
rect -1468 1438 293430 1449
rect -998 1437 -698 1438
rect 902 1437 1202 1438
rect 18902 1437 19202 1438
rect 36902 1437 37202 1438
rect 54902 1437 55202 1438
rect 72902 1437 73202 1438
rect 90902 1437 91202 1438
rect 108902 1437 109202 1438
rect 126902 1437 127202 1438
rect 144902 1437 145202 1438
rect 162902 1437 163202 1438
rect 180902 1437 181202 1438
rect 198902 1437 199202 1438
rect 216902 1437 217202 1438
rect 234902 1437 235202 1438
rect 252902 1437 253202 1438
rect 270902 1437 271202 1438
rect 288902 1437 289202 1438
rect 292660 1437 292960 1438
rect -998 -162 -698 -161
rect 902 -162 1202 -161
rect 18902 -162 19202 -161
rect 36902 -162 37202 -161
rect 54902 -162 55202 -161
rect 72902 -162 73202 -161
rect 90902 -162 91202 -161
rect 108902 -162 109202 -161
rect 126902 -162 127202 -161
rect 144902 -162 145202 -161
rect 162902 -162 163202 -161
rect 180902 -162 181202 -161
rect 198902 -162 199202 -161
rect 216902 -162 217202 -161
rect 234902 -162 235202 -161
rect 252902 -162 253202 -161
rect 270902 -162 271202 -161
rect 288902 -162 289202 -161
rect 292660 -162 292960 -161
rect -998 -173 292960 -162
rect -998 -291 -907 -173
rect -789 -291 993 -173
rect 1111 -291 18993 -173
rect 19111 -291 36993 -173
rect 37111 -291 54993 -173
rect 55111 -291 72993 -173
rect 73111 -291 90993 -173
rect 91111 -291 108993 -173
rect 109111 -291 126993 -173
rect 127111 -291 144993 -173
rect 145111 -291 162993 -173
rect 163111 -291 180993 -173
rect 181111 -291 198993 -173
rect 199111 -291 216993 -173
rect 217111 -291 234993 -173
rect 235111 -291 252993 -173
rect 253111 -291 270993 -173
rect 271111 -291 288993 -173
rect 289111 -291 292751 -173
rect 292869 -291 292960 -173
rect -998 -333 292960 -291
rect -998 -451 -907 -333
rect -789 -451 993 -333
rect 1111 -451 18993 -333
rect 19111 -451 36993 -333
rect 37111 -451 54993 -333
rect 55111 -451 72993 -333
rect 73111 -451 90993 -333
rect 91111 -451 108993 -333
rect 109111 -451 126993 -333
rect 127111 -451 144993 -333
rect 145111 -451 162993 -333
rect 163111 -451 180993 -333
rect 181111 -451 198993 -333
rect 199111 -451 216993 -333
rect 217111 -451 234993 -333
rect 235111 -451 252993 -333
rect 253111 -451 270993 -333
rect 271111 -451 288993 -333
rect 289111 -451 292751 -333
rect 292869 -451 292960 -333
rect -998 -462 292960 -451
rect -998 -463 -698 -462
rect 902 -463 1202 -462
rect 18902 -463 19202 -462
rect 36902 -463 37202 -462
rect 54902 -463 55202 -462
rect 72902 -463 73202 -462
rect 90902 -463 91202 -462
rect 108902 -463 109202 -462
rect 126902 -463 127202 -462
rect 144902 -463 145202 -462
rect 162902 -463 163202 -462
rect 180902 -463 181202 -462
rect 198902 -463 199202 -462
rect 216902 -463 217202 -462
rect 234902 -463 235202 -462
rect 252902 -463 253202 -462
rect 270902 -463 271202 -462
rect 288902 -463 289202 -462
rect 292660 -463 292960 -462
rect -1468 -632 -1168 -631
rect 9902 -632 10202 -631
rect 27902 -632 28202 -631
rect 45902 -632 46202 -631
rect 63902 -632 64202 -631
rect 81902 -632 82202 -631
rect 99902 -632 100202 -631
rect 117902 -632 118202 -631
rect 135902 -632 136202 -631
rect 153902 -632 154202 -631
rect 171902 -632 172202 -631
rect 189902 -632 190202 -631
rect 207902 -632 208202 -631
rect 225902 -632 226202 -631
rect 243902 -632 244202 -631
rect 261902 -632 262202 -631
rect 279902 -632 280202 -631
rect 293130 -632 293430 -631
rect -1468 -643 293430 -632
rect -1468 -761 -1377 -643
rect -1259 -761 9993 -643
rect 10111 -761 27993 -643
rect 28111 -761 45993 -643
rect 46111 -761 63993 -643
rect 64111 -761 81993 -643
rect 82111 -761 99993 -643
rect 100111 -761 117993 -643
rect 118111 -761 135993 -643
rect 136111 -761 153993 -643
rect 154111 -761 171993 -643
rect 172111 -761 189993 -643
rect 190111 -761 207993 -643
rect 208111 -761 225993 -643
rect 226111 -761 243993 -643
rect 244111 -761 261993 -643
rect 262111 -761 279993 -643
rect 280111 -761 293221 -643
rect 293339 -761 293430 -643
rect -1468 -803 293430 -761
rect -1468 -921 -1377 -803
rect -1259 -921 9993 -803
rect 10111 -921 27993 -803
rect 28111 -921 45993 -803
rect 46111 -921 63993 -803
rect 64111 -921 81993 -803
rect 82111 -921 99993 -803
rect 100111 -921 117993 -803
rect 118111 -921 135993 -803
rect 136111 -921 153993 -803
rect 154111 -921 171993 -803
rect 172111 -921 189993 -803
rect 190111 -921 207993 -803
rect 208111 -921 225993 -803
rect 226111 -921 243993 -803
rect 244111 -921 261993 -803
rect 262111 -921 279993 -803
rect 280111 -921 293221 -803
rect 293339 -921 293430 -803
rect -1468 -932 293430 -921
rect -1468 -933 -1168 -932
rect 9902 -933 10202 -932
rect 27902 -933 28202 -932
rect 45902 -933 46202 -932
rect 63902 -933 64202 -932
rect 81902 -933 82202 -932
rect 99902 -933 100202 -932
rect 117902 -933 118202 -932
rect 135902 -933 136202 -932
rect 153902 -933 154202 -932
rect 171902 -933 172202 -932
rect 189902 -933 190202 -932
rect 207902 -933 208202 -932
rect 225902 -933 226202 -932
rect 243902 -933 244202 -932
rect 261902 -933 262202 -932
rect 279902 -933 280202 -932
rect 293130 -933 293430 -932
rect -1938 -1102 -1638 -1101
rect 2702 -1102 3002 -1101
rect 20702 -1102 21002 -1101
rect 38702 -1102 39002 -1101
rect 56702 -1102 57002 -1101
rect 74702 -1102 75002 -1101
rect 92702 -1102 93002 -1101
rect 110702 -1102 111002 -1101
rect 128702 -1102 129002 -1101
rect 146702 -1102 147002 -1101
rect 164702 -1102 165002 -1101
rect 182702 -1102 183002 -1101
rect 200702 -1102 201002 -1101
rect 218702 -1102 219002 -1101
rect 236702 -1102 237002 -1101
rect 254702 -1102 255002 -1101
rect 272702 -1102 273002 -1101
rect 290702 -1102 291002 -1101
rect 293600 -1102 293900 -1101
rect -1938 -1113 293900 -1102
rect -1938 -1231 -1847 -1113
rect -1729 -1231 2793 -1113
rect 2911 -1231 20793 -1113
rect 20911 -1231 38793 -1113
rect 38911 -1231 56793 -1113
rect 56911 -1231 74793 -1113
rect 74911 -1231 92793 -1113
rect 92911 -1231 110793 -1113
rect 110911 -1231 128793 -1113
rect 128911 -1231 146793 -1113
rect 146911 -1231 164793 -1113
rect 164911 -1231 182793 -1113
rect 182911 -1231 200793 -1113
rect 200911 -1231 218793 -1113
rect 218911 -1231 236793 -1113
rect 236911 -1231 254793 -1113
rect 254911 -1231 272793 -1113
rect 272911 -1231 290793 -1113
rect 290911 -1231 293691 -1113
rect 293809 -1231 293900 -1113
rect -1938 -1273 293900 -1231
rect -1938 -1391 -1847 -1273
rect -1729 -1391 2793 -1273
rect 2911 -1391 20793 -1273
rect 20911 -1391 38793 -1273
rect 38911 -1391 56793 -1273
rect 56911 -1391 74793 -1273
rect 74911 -1391 92793 -1273
rect 92911 -1391 110793 -1273
rect 110911 -1391 128793 -1273
rect 128911 -1391 146793 -1273
rect 146911 -1391 164793 -1273
rect 164911 -1391 182793 -1273
rect 182911 -1391 200793 -1273
rect 200911 -1391 218793 -1273
rect 218911 -1391 236793 -1273
rect 236911 -1391 254793 -1273
rect 254911 -1391 272793 -1273
rect 272911 -1391 290793 -1273
rect 290911 -1391 293691 -1273
rect 293809 -1391 293900 -1273
rect -1938 -1402 293900 -1391
rect -1938 -1403 -1638 -1402
rect 2702 -1403 3002 -1402
rect 20702 -1403 21002 -1402
rect 38702 -1403 39002 -1402
rect 56702 -1403 57002 -1402
rect 74702 -1403 75002 -1402
rect 92702 -1403 93002 -1402
rect 110702 -1403 111002 -1402
rect 128702 -1403 129002 -1402
rect 146702 -1403 147002 -1402
rect 164702 -1403 165002 -1402
rect 182702 -1403 183002 -1402
rect 200702 -1403 201002 -1402
rect 218702 -1403 219002 -1402
rect 236702 -1403 237002 -1402
rect 254702 -1403 255002 -1402
rect 272702 -1403 273002 -1402
rect 290702 -1403 291002 -1402
rect 293600 -1403 293900 -1402
rect -2408 -1572 -2108 -1571
rect 11702 -1572 12002 -1571
rect 29702 -1572 30002 -1571
rect 47702 -1572 48002 -1571
rect 65702 -1572 66002 -1571
rect 83702 -1572 84002 -1571
rect 101702 -1572 102002 -1571
rect 119702 -1572 120002 -1571
rect 137702 -1572 138002 -1571
rect 155702 -1572 156002 -1571
rect 173702 -1572 174002 -1571
rect 191702 -1572 192002 -1571
rect 209702 -1572 210002 -1571
rect 227702 -1572 228002 -1571
rect 245702 -1572 246002 -1571
rect 263702 -1572 264002 -1571
rect 281702 -1572 282002 -1571
rect 294070 -1572 294370 -1571
rect -2408 -1583 294370 -1572
rect -2408 -1701 -2317 -1583
rect -2199 -1701 11793 -1583
rect 11911 -1701 29793 -1583
rect 29911 -1701 47793 -1583
rect 47911 -1701 65793 -1583
rect 65911 -1701 83793 -1583
rect 83911 -1701 101793 -1583
rect 101911 -1701 119793 -1583
rect 119911 -1701 137793 -1583
rect 137911 -1701 155793 -1583
rect 155911 -1701 173793 -1583
rect 173911 -1701 191793 -1583
rect 191911 -1701 209793 -1583
rect 209911 -1701 227793 -1583
rect 227911 -1701 245793 -1583
rect 245911 -1701 263793 -1583
rect 263911 -1701 281793 -1583
rect 281911 -1701 294161 -1583
rect 294279 -1701 294370 -1583
rect -2408 -1743 294370 -1701
rect -2408 -1861 -2317 -1743
rect -2199 -1861 11793 -1743
rect 11911 -1861 29793 -1743
rect 29911 -1861 47793 -1743
rect 47911 -1861 65793 -1743
rect 65911 -1861 83793 -1743
rect 83911 -1861 101793 -1743
rect 101911 -1861 119793 -1743
rect 119911 -1861 137793 -1743
rect 137911 -1861 155793 -1743
rect 155911 -1861 173793 -1743
rect 173911 -1861 191793 -1743
rect 191911 -1861 209793 -1743
rect 209911 -1861 227793 -1743
rect 227911 -1861 245793 -1743
rect 245911 -1861 263793 -1743
rect 263911 -1861 281793 -1743
rect 281911 -1861 294161 -1743
rect 294279 -1861 294370 -1743
rect -2408 -1872 294370 -1861
rect -2408 -1873 -2108 -1872
rect 11702 -1873 12002 -1872
rect 29702 -1873 30002 -1872
rect 47702 -1873 48002 -1872
rect 65702 -1873 66002 -1872
rect 83702 -1873 84002 -1872
rect 101702 -1873 102002 -1872
rect 119702 -1873 120002 -1872
rect 137702 -1873 138002 -1872
rect 155702 -1873 156002 -1872
rect 173702 -1873 174002 -1872
rect 191702 -1873 192002 -1872
rect 209702 -1873 210002 -1872
rect 227702 -1873 228002 -1872
rect 245702 -1873 246002 -1872
rect 263702 -1873 264002 -1872
rect 281702 -1873 282002 -1872
rect 294070 -1873 294370 -1872
rect -2878 -2042 -2578 -2041
rect 4502 -2042 4802 -2041
rect 22502 -2042 22802 -2041
rect 40502 -2042 40802 -2041
rect 58502 -2042 58802 -2041
rect 76502 -2042 76802 -2041
rect 94502 -2042 94802 -2041
rect 112502 -2042 112802 -2041
rect 130502 -2042 130802 -2041
rect 148502 -2042 148802 -2041
rect 166502 -2042 166802 -2041
rect 184502 -2042 184802 -2041
rect 202502 -2042 202802 -2041
rect 220502 -2042 220802 -2041
rect 238502 -2042 238802 -2041
rect 256502 -2042 256802 -2041
rect 274502 -2042 274802 -2041
rect 294540 -2042 294840 -2041
rect -2878 -2053 294840 -2042
rect -2878 -2171 -2787 -2053
rect -2669 -2171 4593 -2053
rect 4711 -2171 22593 -2053
rect 22711 -2171 40593 -2053
rect 40711 -2171 58593 -2053
rect 58711 -2171 76593 -2053
rect 76711 -2171 94593 -2053
rect 94711 -2171 112593 -2053
rect 112711 -2171 130593 -2053
rect 130711 -2171 148593 -2053
rect 148711 -2171 166593 -2053
rect 166711 -2171 184593 -2053
rect 184711 -2171 202593 -2053
rect 202711 -2171 220593 -2053
rect 220711 -2171 238593 -2053
rect 238711 -2171 256593 -2053
rect 256711 -2171 274593 -2053
rect 274711 -2171 294631 -2053
rect 294749 -2171 294840 -2053
rect -2878 -2213 294840 -2171
rect -2878 -2331 -2787 -2213
rect -2669 -2331 4593 -2213
rect 4711 -2331 22593 -2213
rect 22711 -2331 40593 -2213
rect 40711 -2331 58593 -2213
rect 58711 -2331 76593 -2213
rect 76711 -2331 94593 -2213
rect 94711 -2331 112593 -2213
rect 112711 -2331 130593 -2213
rect 130711 -2331 148593 -2213
rect 148711 -2331 166593 -2213
rect 166711 -2331 184593 -2213
rect 184711 -2331 202593 -2213
rect 202711 -2331 220593 -2213
rect 220711 -2331 238593 -2213
rect 238711 -2331 256593 -2213
rect 256711 -2331 274593 -2213
rect 274711 -2331 294631 -2213
rect 294749 -2331 294840 -2213
rect -2878 -2342 294840 -2331
rect -2878 -2343 -2578 -2342
rect 4502 -2343 4802 -2342
rect 22502 -2343 22802 -2342
rect 40502 -2343 40802 -2342
rect 58502 -2343 58802 -2342
rect 76502 -2343 76802 -2342
rect 94502 -2343 94802 -2342
rect 112502 -2343 112802 -2342
rect 130502 -2343 130802 -2342
rect 148502 -2343 148802 -2342
rect 166502 -2343 166802 -2342
rect 184502 -2343 184802 -2342
rect 202502 -2343 202802 -2342
rect 220502 -2343 220802 -2342
rect 238502 -2343 238802 -2342
rect 256502 -2343 256802 -2342
rect 274502 -2343 274802 -2342
rect 294540 -2343 294840 -2342
rect -3348 -2512 -3048 -2511
rect 13502 -2512 13802 -2511
rect 31502 -2512 31802 -2511
rect 49502 -2512 49802 -2511
rect 67502 -2512 67802 -2511
rect 85502 -2512 85802 -2511
rect 103502 -2512 103802 -2511
rect 121502 -2512 121802 -2511
rect 139502 -2512 139802 -2511
rect 157502 -2512 157802 -2511
rect 175502 -2512 175802 -2511
rect 193502 -2512 193802 -2511
rect 211502 -2512 211802 -2511
rect 229502 -2512 229802 -2511
rect 247502 -2512 247802 -2511
rect 265502 -2512 265802 -2511
rect 283502 -2512 283802 -2511
rect 295010 -2512 295310 -2511
rect -3348 -2523 295310 -2512
rect -3348 -2641 -3257 -2523
rect -3139 -2641 13593 -2523
rect 13711 -2641 31593 -2523
rect 31711 -2641 49593 -2523
rect 49711 -2641 67593 -2523
rect 67711 -2641 85593 -2523
rect 85711 -2641 103593 -2523
rect 103711 -2641 121593 -2523
rect 121711 -2641 139593 -2523
rect 139711 -2641 157593 -2523
rect 157711 -2641 175593 -2523
rect 175711 -2641 193593 -2523
rect 193711 -2641 211593 -2523
rect 211711 -2641 229593 -2523
rect 229711 -2641 247593 -2523
rect 247711 -2641 265593 -2523
rect 265711 -2641 283593 -2523
rect 283711 -2641 295101 -2523
rect 295219 -2641 295310 -2523
rect -3348 -2683 295310 -2641
rect -3348 -2801 -3257 -2683
rect -3139 -2801 13593 -2683
rect 13711 -2801 31593 -2683
rect 31711 -2801 49593 -2683
rect 49711 -2801 67593 -2683
rect 67711 -2801 85593 -2683
rect 85711 -2801 103593 -2683
rect 103711 -2801 121593 -2683
rect 121711 -2801 139593 -2683
rect 139711 -2801 157593 -2683
rect 157711 -2801 175593 -2683
rect 175711 -2801 193593 -2683
rect 193711 -2801 211593 -2683
rect 211711 -2801 229593 -2683
rect 229711 -2801 247593 -2683
rect 247711 -2801 265593 -2683
rect 265711 -2801 283593 -2683
rect 283711 -2801 295101 -2683
rect 295219 -2801 295310 -2683
rect -3348 -2812 295310 -2801
rect -3348 -2813 -3048 -2812
rect 13502 -2813 13802 -2812
rect 31502 -2813 31802 -2812
rect 49502 -2813 49802 -2812
rect 67502 -2813 67802 -2812
rect 85502 -2813 85802 -2812
rect 103502 -2813 103802 -2812
rect 121502 -2813 121802 -2812
rect 139502 -2813 139802 -2812
rect 157502 -2813 157802 -2812
rect 175502 -2813 175802 -2812
rect 193502 -2813 193802 -2812
rect 211502 -2813 211802 -2812
rect 229502 -2813 229802 -2812
rect 247502 -2813 247802 -2812
rect 265502 -2813 265802 -2812
rect 283502 -2813 283802 -2812
rect 295010 -2813 295310 -2812
rect -3818 -2982 -3518 -2981
rect 6302 -2982 6602 -2981
rect 24302 -2982 24602 -2981
rect 42302 -2982 42602 -2981
rect 60302 -2982 60602 -2981
rect 78302 -2982 78602 -2981
rect 96302 -2982 96602 -2981
rect 114302 -2982 114602 -2981
rect 132302 -2982 132602 -2981
rect 150302 -2982 150602 -2981
rect 168302 -2982 168602 -2981
rect 186302 -2982 186602 -2981
rect 204302 -2982 204602 -2981
rect 222302 -2982 222602 -2981
rect 240302 -2982 240602 -2981
rect 258302 -2982 258602 -2981
rect 276302 -2982 276602 -2981
rect 295480 -2982 295780 -2981
rect -3818 -2993 295780 -2982
rect -3818 -3111 -3727 -2993
rect -3609 -3111 6393 -2993
rect 6511 -3111 24393 -2993
rect 24511 -3111 42393 -2993
rect 42511 -3111 60393 -2993
rect 60511 -3111 78393 -2993
rect 78511 -3111 96393 -2993
rect 96511 -3111 114393 -2993
rect 114511 -3111 132393 -2993
rect 132511 -3111 150393 -2993
rect 150511 -3111 168393 -2993
rect 168511 -3111 186393 -2993
rect 186511 -3111 204393 -2993
rect 204511 -3111 222393 -2993
rect 222511 -3111 240393 -2993
rect 240511 -3111 258393 -2993
rect 258511 -3111 276393 -2993
rect 276511 -3111 295571 -2993
rect 295689 -3111 295780 -2993
rect -3818 -3153 295780 -3111
rect -3818 -3271 -3727 -3153
rect -3609 -3271 6393 -3153
rect 6511 -3271 24393 -3153
rect 24511 -3271 42393 -3153
rect 42511 -3271 60393 -3153
rect 60511 -3271 78393 -3153
rect 78511 -3271 96393 -3153
rect 96511 -3271 114393 -3153
rect 114511 -3271 132393 -3153
rect 132511 -3271 150393 -3153
rect 150511 -3271 168393 -3153
rect 168511 -3271 186393 -3153
rect 186511 -3271 204393 -3153
rect 204511 -3271 222393 -3153
rect 222511 -3271 240393 -3153
rect 240511 -3271 258393 -3153
rect 258511 -3271 276393 -3153
rect 276511 -3271 295571 -3153
rect 295689 -3271 295780 -3153
rect -3818 -3282 295780 -3271
rect -3818 -3283 -3518 -3282
rect 6302 -3283 6602 -3282
rect 24302 -3283 24602 -3282
rect 42302 -3283 42602 -3282
rect 60302 -3283 60602 -3282
rect 78302 -3283 78602 -3282
rect 96302 -3283 96602 -3282
rect 114302 -3283 114602 -3282
rect 132302 -3283 132602 -3282
rect 150302 -3283 150602 -3282
rect 168302 -3283 168602 -3282
rect 186302 -3283 186602 -3282
rect 204302 -3283 204602 -3282
rect 222302 -3283 222602 -3282
rect 240302 -3283 240602 -3282
rect 258302 -3283 258602 -3282
rect 276302 -3283 276602 -3282
rect 295480 -3283 295780 -3282
rect -4288 -3452 -3988 -3451
rect 15302 -3452 15602 -3451
rect 33302 -3452 33602 -3451
rect 51302 -3452 51602 -3451
rect 69302 -3452 69602 -3451
rect 87302 -3452 87602 -3451
rect 105302 -3452 105602 -3451
rect 123302 -3452 123602 -3451
rect 141302 -3452 141602 -3451
rect 159302 -3452 159602 -3451
rect 177302 -3452 177602 -3451
rect 195302 -3452 195602 -3451
rect 213302 -3452 213602 -3451
rect 231302 -3452 231602 -3451
rect 249302 -3452 249602 -3451
rect 267302 -3452 267602 -3451
rect 285302 -3452 285602 -3451
rect 295950 -3452 296250 -3451
rect -4288 -3463 296250 -3452
rect -4288 -3581 -4197 -3463
rect -4079 -3581 15393 -3463
rect 15511 -3581 33393 -3463
rect 33511 -3581 51393 -3463
rect 51511 -3581 69393 -3463
rect 69511 -3581 87393 -3463
rect 87511 -3581 105393 -3463
rect 105511 -3581 123393 -3463
rect 123511 -3581 141393 -3463
rect 141511 -3581 159393 -3463
rect 159511 -3581 177393 -3463
rect 177511 -3581 195393 -3463
rect 195511 -3581 213393 -3463
rect 213511 -3581 231393 -3463
rect 231511 -3581 249393 -3463
rect 249511 -3581 267393 -3463
rect 267511 -3581 285393 -3463
rect 285511 -3581 296041 -3463
rect 296159 -3581 296250 -3463
rect -4288 -3623 296250 -3581
rect -4288 -3741 -4197 -3623
rect -4079 -3741 15393 -3623
rect 15511 -3741 33393 -3623
rect 33511 -3741 51393 -3623
rect 51511 -3741 69393 -3623
rect 69511 -3741 87393 -3623
rect 87511 -3741 105393 -3623
rect 105511 -3741 123393 -3623
rect 123511 -3741 141393 -3623
rect 141511 -3741 159393 -3623
rect 159511 -3741 177393 -3623
rect 177511 -3741 195393 -3623
rect 195511 -3741 213393 -3623
rect 213511 -3741 231393 -3623
rect 231511 -3741 249393 -3623
rect 249511 -3741 267393 -3623
rect 267511 -3741 285393 -3623
rect 285511 -3741 296041 -3623
rect 296159 -3741 296250 -3623
rect -4288 -3752 296250 -3741
rect -4288 -3753 -3988 -3752
rect 15302 -3753 15602 -3752
rect 33302 -3753 33602 -3752
rect 51302 -3753 51602 -3752
rect 69302 -3753 69602 -3752
rect 87302 -3753 87602 -3752
rect 105302 -3753 105602 -3752
rect 123302 -3753 123602 -3752
rect 141302 -3753 141602 -3752
rect 159302 -3753 159602 -3752
rect 177302 -3753 177602 -3752
rect 195302 -3753 195602 -3752
rect 213302 -3753 213602 -3752
rect 231302 -3753 231602 -3752
rect 249302 -3753 249602 -3752
rect 267302 -3753 267602 -3752
rect 285302 -3753 285602 -3752
rect 295950 -3753 296250 -3752
<< labels >>
rlabel metal3 s 291760 2898 292480 3018 6 analog_io[0]
port 0 nsew signal bidirectional
rlabel metal3 s 291760 237498 292480 237618 6 analog_io[10]
port 1 nsew signal bidirectional
rlabel metal3 s 291760 260958 292480 261078 6 analog_io[11]
port 2 nsew signal bidirectional
rlabel metal3 s 291760 284418 292480 284538 6 analog_io[12]
port 3 nsew signal bidirectional
rlabel metal3 s 291760 307878 292480 307998 6 analog_io[13]
port 4 nsew signal bidirectional
rlabel metal3 s 291760 331338 292480 331458 6 analog_io[14]
port 5 nsew signal bidirectional
rlabel metal2 s 287909 351760 287965 352480 6 analog_io[15]
port 6 nsew signal bidirectional
rlabel metal2 s 255479 351760 255535 352480 6 analog_io[16]
port 7 nsew signal bidirectional
rlabel metal2 s 223049 351760 223105 352480 6 analog_io[17]
port 8 nsew signal bidirectional
rlabel metal2 s 190573 351760 190629 352480 6 analog_io[18]
port 9 nsew signal bidirectional
rlabel metal2 s 158143 351760 158199 352480 6 analog_io[19]
port 10 nsew signal bidirectional
rlabel metal3 s 291760 26358 292480 26478 6 analog_io[1]
port 11 nsew signal bidirectional
rlabel metal2 s 125713 351760 125769 352480 6 analog_io[20]
port 12 nsew signal bidirectional
rlabel metal2 s 93237 351760 93293 352480 6 analog_io[21]
port 13 nsew signal bidirectional
rlabel metal2 s 60807 351760 60863 352480 6 analog_io[22]
port 14 nsew signal bidirectional
rlabel metal2 s 28377 351760 28433 352480 6 analog_io[23]
port 15 nsew signal bidirectional
rlabel metal3 s -480 348134 240 348254 4 analog_io[24]
port 16 nsew signal bidirectional
rlabel metal3 s -480 318214 240 318334 4 analog_io[25]
port 17 nsew signal bidirectional
rlabel metal3 s -480 288226 240 288346 4 analog_io[26]
port 18 nsew signal bidirectional
rlabel metal3 s -480 258306 240 258426 4 analog_io[27]
port 19 nsew signal bidirectional
rlabel metal3 s -480 228318 240 228438 4 analog_io[28]
port 20 nsew signal bidirectional
rlabel metal3 s 291760 49818 292480 49938 6 analog_io[2]
port 21 nsew signal bidirectional
rlabel metal3 s 291760 73278 292480 73398 6 analog_io[3]
port 22 nsew signal bidirectional
rlabel metal3 s 291760 96738 292480 96858 6 analog_io[4]
port 23 nsew signal bidirectional
rlabel metal3 s 291760 120198 292480 120318 6 analog_io[5]
port 24 nsew signal bidirectional
rlabel metal3 s 291760 143658 292480 143778 6 analog_io[6]
port 25 nsew signal bidirectional
rlabel metal3 s 291760 167118 292480 167238 6 analog_io[7]
port 26 nsew signal bidirectional
rlabel metal3 s 291760 190578 292480 190698 6 analog_io[8]
port 27 nsew signal bidirectional
rlabel metal3 s 291760 214038 292480 214158 6 analog_io[9]
port 28 nsew signal bidirectional
rlabel metal3 s 291760 8746 292480 8866 6 io_in[0]
port 29 nsew signal input
rlabel metal3 s 291760 14594 292480 14714 6 io_out[0]
port 30 nsew signal tristate
rlabel metal3 s 291760 243346 292480 243466 6 io_in[10]
port 31 nsew signal input
rlabel metal3 s 291760 249262 292480 249382 6 io_out[10]
port 32 nsew signal tristate
rlabel metal3 s 291760 266874 292480 266994 6 io_in[11]
port 33 nsew signal input
rlabel metal3 s 291760 272722 292480 272842 6 io_out[11]
port 34 nsew signal tristate
rlabel metal3 s 291760 290334 292480 290454 6 io_in[12]
port 35 nsew signal input
rlabel metal3 s 291760 296182 292480 296302 6 io_out[12]
port 36 nsew signal tristate
rlabel metal3 s 291760 313794 292480 313914 6 io_in[13]
port 37 nsew signal input
rlabel metal3 s 291760 319642 292480 319762 6 io_out[13]
port 38 nsew signal tristate
rlabel metal3 s 291760 337254 292480 337374 6 io_in[14]
port 39 nsew signal input
rlabel metal3 s 291760 343102 292480 343222 6 io_out[14]
port 40 nsew signal tristate
rlabel metal2 s 279813 351760 279869 352480 6 io_in[15]
port 41 nsew signal input
rlabel metal2 s 271717 351760 271773 352480 6 io_out[15]
port 42 nsew signal tristate
rlabel metal2 s 247383 351760 247439 352480 6 io_in[16]
port 43 nsew signal input
rlabel metal2 s 239241 351760 239297 352480 6 io_out[16]
port 44 nsew signal tristate
rlabel metal2 s 214907 351760 214963 352480 6 io_in[17]
port 45 nsew signal input
rlabel metal2 s 206811 351760 206867 352480 6 io_out[17]
port 46 nsew signal tristate
rlabel metal2 s 182477 351760 182533 352480 6 io_in[18]
port 47 nsew signal input
rlabel metal2 s 174381 351760 174437 352480 6 io_out[18]
port 48 nsew signal tristate
rlabel metal2 s 150047 351760 150103 352480 6 io_in[19]
port 49 nsew signal input
rlabel metal2 s 141905 351760 141961 352480 6 io_out[19]
port 50 nsew signal tristate
rlabel metal3 s 291760 32206 292480 32326 6 io_in[1]
port 51 nsew signal input
rlabel metal3 s 291760 38054 292480 38174 6 io_out[1]
port 52 nsew signal tristate
rlabel metal2 s 117571 351760 117627 352480 6 io_in[20]
port 53 nsew signal input
rlabel metal2 s 109475 351760 109531 352480 6 io_out[20]
port 54 nsew signal tristate
rlabel metal2 s 85141 351760 85197 352480 6 io_in[21]
port 55 nsew signal input
rlabel metal2 s 77045 351760 77101 352480 6 io_out[21]
port 56 nsew signal tristate
rlabel metal2 s 52711 351760 52767 352480 6 io_in[22]
port 57 nsew signal input
rlabel metal2 s 44569 351760 44625 352480 6 io_out[22]
port 58 nsew signal tristate
rlabel metal2 s 20235 351760 20291 352480 6 io_in[23]
port 59 nsew signal input
rlabel metal2 s 12139 351760 12195 352480 6 io_out[23]
port 60 nsew signal tristate
rlabel metal3 s -480 340654 240 340774 4 io_in[24]
port 61 nsew signal input
rlabel metal3 s -480 333174 240 333294 4 io_out[24]
port 62 nsew signal tristate
rlabel metal3 s -480 310734 240 310854 4 io_in[25]
port 63 nsew signal input
rlabel metal3 s -480 303254 240 303374 4 io_out[25]
port 64 nsew signal tristate
rlabel metal3 s -480 280746 240 280866 4 io_in[26]
port 65 nsew signal input
rlabel metal3 s -480 273266 240 273386 4 io_out[26]
port 66 nsew signal tristate
rlabel metal3 s -480 250826 240 250946 4 io_in[27]
port 67 nsew signal input
rlabel metal3 s -480 243346 240 243466 4 io_out[27]
port 68 nsew signal tristate
rlabel metal3 s -480 220838 240 220958 4 io_in[28]
port 69 nsew signal input
rlabel metal3 s -480 213358 240 213478 4 io_out[28]
port 70 nsew signal tristate
rlabel metal3 s -480 198398 240 198518 4 io_in[29]
port 71 nsew signal input
rlabel metal3 s -480 190918 240 191038 4 io_out[29]
port 72 nsew signal tristate
rlabel metal3 s 291760 55666 292480 55786 6 io_in[2]
port 73 nsew signal input
rlabel metal3 s 291760 61514 292480 61634 6 io_out[2]
port 74 nsew signal tristate
rlabel metal3 s -480 175890 240 176010 4 io_in[30]
port 75 nsew signal input
rlabel metal3 s -480 168410 240 168530 4 io_out[30]
port 76 nsew signal tristate
rlabel metal3 s -480 153450 240 153570 4 io_in[31]
port 77 nsew signal input
rlabel metal3 s -480 145970 240 146090 4 io_out[31]
port 78 nsew signal tristate
rlabel metal3 s -480 131010 240 131130 4 io_in[32]
port 79 nsew signal input
rlabel metal3 s -480 123530 240 123650 4 io_out[32]
port 80 nsew signal tristate
rlabel metal3 s -480 108502 240 108622 4 io_in[33]
port 81 nsew signal input
rlabel metal3 s -480 101022 240 101142 4 io_out[33]
port 82 nsew signal tristate
rlabel metal3 s -480 86062 240 86182 4 io_in[34]
port 83 nsew signal input
rlabel metal3 s -480 78582 240 78702 4 io_out[34]
port 84 nsew signal tristate
rlabel metal3 s -480 63622 240 63742 4 io_in[35]
port 85 nsew signal input
rlabel metal3 s -480 56074 240 56194 4 io_out[35]
port 86 nsew signal tristate
rlabel metal3 s -480 41114 240 41234 4 io_in[36]
port 87 nsew signal input
rlabel metal3 s -480 33634 240 33754 4 io_out[36]
port 88 nsew signal tristate
rlabel metal3 s -480 18674 240 18794 4 io_in[37]
port 89 nsew signal input
rlabel metal3 s -480 11194 240 11314 4 io_out[37]
port 90 nsew signal tristate
rlabel metal3 s 291760 79126 292480 79246 6 io_in[3]
port 91 nsew signal input
rlabel metal3 s 291760 84974 292480 85094 6 io_out[3]
port 92 nsew signal tristate
rlabel metal3 s 291760 102586 292480 102706 6 io_in[4]
port 93 nsew signal input
rlabel metal3 s 291760 108434 292480 108554 6 io_out[4]
port 94 nsew signal tristate
rlabel metal3 s 291760 126046 292480 126166 6 io_in[5]
port 95 nsew signal input
rlabel metal3 s 291760 131894 292480 132014 6 io_out[5]
port 96 nsew signal tristate
rlabel metal3 s 291760 149506 292480 149626 6 io_in[6]
port 97 nsew signal input
rlabel metal3 s 291760 155354 292480 155474 6 io_out[6]
port 98 nsew signal tristate
rlabel metal3 s 291760 172966 292480 173086 6 io_in[7]
port 99 nsew signal input
rlabel metal3 s 291760 178882 292480 179002 6 io_out[7]
port 100 nsew signal tristate
rlabel metal3 s 291760 196426 292480 196546 6 io_in[8]
port 101 nsew signal input
rlabel metal3 s 291760 202342 292480 202462 6 io_out[8]
port 102 nsew signal tristate
rlabel metal3 s 291760 219886 292480 220006 6 io_in[9]
port 103 nsew signal input
rlabel metal3 s 291760 225802 292480 225922 6 io_out[9]
port 104 nsew signal tristate
rlabel metal3 s 291760 20442 292480 20562 6 io_oeb[0]
port 105 nsew signal tristate
rlabel metal3 s 291760 255110 292480 255230 6 io_oeb[10]
port 106 nsew signal tristate
rlabel metal3 s 291760 278570 292480 278690 6 io_oeb[11]
port 107 nsew signal tristate
rlabel metal3 s 291760 302030 292480 302150 6 io_oeb[12]
port 108 nsew signal tristate
rlabel metal3 s 291760 325490 292480 325610 6 io_oeb[13]
port 109 nsew signal tristate
rlabel metal3 s 291760 348950 292480 349070 6 io_oeb[14]
port 110 nsew signal tristate
rlabel metal2 s 263575 351760 263631 352480 6 io_oeb[15]
port 111 nsew signal tristate
rlabel metal2 s 231145 351760 231201 352480 6 io_oeb[16]
port 112 nsew signal tristate
rlabel metal2 s 198715 351760 198771 352480 6 io_oeb[17]
port 113 nsew signal tristate
rlabel metal2 s 166239 351760 166295 352480 6 io_oeb[18]
port 114 nsew signal tristate
rlabel metal2 s 133809 351760 133865 352480 6 io_oeb[19]
port 115 nsew signal tristate
rlabel metal3 s 291760 43902 292480 44022 6 io_oeb[1]
port 116 nsew signal tristate
rlabel metal2 s 101379 351760 101435 352480 6 io_oeb[20]
port 117 nsew signal tristate
rlabel metal2 s 68903 351760 68959 352480 6 io_oeb[21]
port 118 nsew signal tristate
rlabel metal2 s 36473 351760 36529 352480 6 io_oeb[22]
port 119 nsew signal tristate
rlabel metal2 s 4043 351760 4099 352480 6 io_oeb[23]
port 120 nsew signal tristate
rlabel metal3 s -480 325694 240 325814 4 io_oeb[24]
port 121 nsew signal tristate
rlabel metal3 s -480 295706 240 295826 4 io_oeb[25]
port 122 nsew signal tristate
rlabel metal3 s -480 265786 240 265906 4 io_oeb[26]
port 123 nsew signal tristate
rlabel metal3 s -480 235798 240 235918 4 io_oeb[27]
port 124 nsew signal tristate
rlabel metal3 s -480 205878 240 205998 4 io_oeb[28]
port 125 nsew signal tristate
rlabel metal3 s -480 183438 240 183558 4 io_oeb[29]
port 126 nsew signal tristate
rlabel metal3 s 291760 67362 292480 67482 6 io_oeb[2]
port 127 nsew signal tristate
rlabel metal3 s -480 160930 240 161050 4 io_oeb[30]
port 128 nsew signal tristate
rlabel metal3 s -480 138490 240 138610 4 io_oeb[31]
port 129 nsew signal tristate
rlabel metal3 s -480 115982 240 116102 4 io_oeb[32]
port 130 nsew signal tristate
rlabel metal3 s -480 93542 240 93662 4 io_oeb[33]
port 131 nsew signal tristate
rlabel metal3 s -480 71102 240 71222 4 io_oeb[34]
port 132 nsew signal tristate
rlabel metal3 s -480 48594 240 48714 4 io_oeb[35]
port 133 nsew signal tristate
rlabel metal3 s -480 26154 240 26274 4 io_oeb[36]
port 134 nsew signal tristate
rlabel metal3 s -480 3714 240 3834 4 io_oeb[37]
port 135 nsew signal tristate
rlabel metal3 s 291760 90890 292480 91010 6 io_oeb[3]
port 136 nsew signal tristate
rlabel metal3 s 291760 114350 292480 114470 6 io_oeb[4]
port 137 nsew signal tristate
rlabel metal3 s 291760 137810 292480 137930 6 io_oeb[5]
port 138 nsew signal tristate
rlabel metal3 s 291760 161270 292480 161390 6 io_oeb[6]
port 139 nsew signal tristate
rlabel metal3 s 291760 184730 292480 184850 6 io_oeb[7]
port 140 nsew signal tristate
rlabel metal3 s 291760 208190 292480 208310 6 io_oeb[8]
port 141 nsew signal tristate
rlabel metal3 s 291760 231650 292480 231770 6 io_oeb[9]
port 142 nsew signal tristate
rlabel metal2 s 63291 -480 63347 240 8 la_data_in[0]
port 143 nsew signal input
rlabel metal2 s 241725 -480 241781 240 8 la_data_in[100]
port 144 nsew signal input
rlabel metal2 s 243473 -480 243529 240 8 la_data_in[101]
port 145 nsew signal input
rlabel metal2 s 245267 -480 245323 240 8 la_data_in[102]
port 146 nsew signal input
rlabel metal2 s 247061 -480 247117 240 8 la_data_in[103]
port 147 nsew signal input
rlabel metal2 s 248855 -480 248911 240 8 la_data_in[104]
port 148 nsew signal input
rlabel metal2 s 250603 -480 250659 240 8 la_data_in[105]
port 149 nsew signal input
rlabel metal2 s 252397 -480 252453 240 8 la_data_in[106]
port 150 nsew signal input
rlabel metal2 s 254191 -480 254247 240 8 la_data_in[107]
port 151 nsew signal input
rlabel metal2 s 255985 -480 256041 240 8 la_data_in[108]
port 152 nsew signal input
rlabel metal2 s 257779 -480 257835 240 8 la_data_in[109]
port 153 nsew signal input
rlabel metal2 s 81139 -480 81195 240 8 la_data_in[10]
port 154 nsew signal input
rlabel metal2 s 259527 -480 259583 240 8 la_data_in[110]
port 155 nsew signal input
rlabel metal2 s 261321 -480 261377 240 8 la_data_in[111]
port 156 nsew signal input
rlabel metal2 s 263115 -480 263171 240 8 la_data_in[112]
port 157 nsew signal input
rlabel metal2 s 264909 -480 264965 240 8 la_data_in[113]
port 158 nsew signal input
rlabel metal2 s 266703 -480 266759 240 8 la_data_in[114]
port 159 nsew signal input
rlabel metal2 s 268451 -480 268507 240 8 la_data_in[115]
port 160 nsew signal input
rlabel metal2 s 270245 -480 270301 240 8 la_data_in[116]
port 161 nsew signal input
rlabel metal2 s 272039 -480 272095 240 8 la_data_in[117]
port 162 nsew signal input
rlabel metal2 s 273833 -480 273889 240 8 la_data_in[118]
port 163 nsew signal input
rlabel metal2 s 275581 -480 275637 240 8 la_data_in[119]
port 164 nsew signal input
rlabel metal2 s 82933 -480 82989 240 8 la_data_in[11]
port 165 nsew signal input
rlabel metal2 s 277375 -480 277431 240 8 la_data_in[120]
port 166 nsew signal input
rlabel metal2 s 279169 -480 279225 240 8 la_data_in[121]
port 167 nsew signal input
rlabel metal2 s 280963 -480 281019 240 8 la_data_in[122]
port 168 nsew signal input
rlabel metal2 s 282757 -480 282813 240 8 la_data_in[123]
port 169 nsew signal input
rlabel metal2 s 284505 -480 284561 240 8 la_data_in[124]
port 170 nsew signal input
rlabel metal2 s 286299 -480 286355 240 8 la_data_in[125]
port 171 nsew signal input
rlabel metal2 s 288093 -480 288149 240 8 la_data_in[126]
port 172 nsew signal input
rlabel metal2 s 289887 -480 289943 240 8 la_data_in[127]
port 173 nsew signal input
rlabel metal2 s 84681 -480 84737 240 8 la_data_in[12]
port 174 nsew signal input
rlabel metal2 s 86475 -480 86531 240 8 la_data_in[13]
port 175 nsew signal input
rlabel metal2 s 88269 -480 88325 240 8 la_data_in[14]
port 176 nsew signal input
rlabel metal2 s 90063 -480 90119 240 8 la_data_in[15]
port 177 nsew signal input
rlabel metal2 s 91857 -480 91913 240 8 la_data_in[16]
port 178 nsew signal input
rlabel metal2 s 93605 -480 93661 240 8 la_data_in[17]
port 179 nsew signal input
rlabel metal2 s 95399 -480 95455 240 8 la_data_in[18]
port 180 nsew signal input
rlabel metal2 s 97193 -480 97249 240 8 la_data_in[19]
port 181 nsew signal input
rlabel metal2 s 65085 -480 65141 240 8 la_data_in[1]
port 182 nsew signal input
rlabel metal2 s 98987 -480 99043 240 8 la_data_in[20]
port 183 nsew signal input
rlabel metal2 s 100735 -480 100791 240 8 la_data_in[21]
port 184 nsew signal input
rlabel metal2 s 102529 -480 102585 240 8 la_data_in[22]
port 185 nsew signal input
rlabel metal2 s 104323 -480 104379 240 8 la_data_in[23]
port 186 nsew signal input
rlabel metal2 s 106117 -480 106173 240 8 la_data_in[24]
port 187 nsew signal input
rlabel metal2 s 107911 -480 107967 240 8 la_data_in[25]
port 188 nsew signal input
rlabel metal2 s 109659 -480 109715 240 8 la_data_in[26]
port 189 nsew signal input
rlabel metal2 s 111453 -480 111509 240 8 la_data_in[27]
port 190 nsew signal input
rlabel metal2 s 113247 -480 113303 240 8 la_data_in[28]
port 191 nsew signal input
rlabel metal2 s 115041 -480 115097 240 8 la_data_in[29]
port 192 nsew signal input
rlabel metal2 s 66879 -480 66935 240 8 la_data_in[2]
port 193 nsew signal input
rlabel metal2 s 116835 -480 116891 240 8 la_data_in[30]
port 194 nsew signal input
rlabel metal2 s 118583 -480 118639 240 8 la_data_in[31]
port 195 nsew signal input
rlabel metal2 s 120377 -480 120433 240 8 la_data_in[32]
port 196 nsew signal input
rlabel metal2 s 122171 -480 122227 240 8 la_data_in[33]
port 197 nsew signal input
rlabel metal2 s 123965 -480 124021 240 8 la_data_in[34]
port 198 nsew signal input
rlabel metal2 s 125713 -480 125769 240 8 la_data_in[35]
port 199 nsew signal input
rlabel metal2 s 127507 -480 127563 240 8 la_data_in[36]
port 200 nsew signal input
rlabel metal2 s 129301 -480 129357 240 8 la_data_in[37]
port 201 nsew signal input
rlabel metal2 s 131095 -480 131151 240 8 la_data_in[38]
port 202 nsew signal input
rlabel metal2 s 132889 -480 132945 240 8 la_data_in[39]
port 203 nsew signal input
rlabel metal2 s 68627 -480 68683 240 8 la_data_in[3]
port 204 nsew signal input
rlabel metal2 s 134637 -480 134693 240 8 la_data_in[40]
port 205 nsew signal input
rlabel metal2 s 136431 -480 136487 240 8 la_data_in[41]
port 206 nsew signal input
rlabel metal2 s 138225 -480 138281 240 8 la_data_in[42]
port 207 nsew signal input
rlabel metal2 s 140019 -480 140075 240 8 la_data_in[43]
port 208 nsew signal input
rlabel metal2 s 141813 -480 141869 240 8 la_data_in[44]
port 209 nsew signal input
rlabel metal2 s 143561 -480 143617 240 8 la_data_in[45]
port 210 nsew signal input
rlabel metal2 s 145355 -480 145411 240 8 la_data_in[46]
port 211 nsew signal input
rlabel metal2 s 147149 -480 147205 240 8 la_data_in[47]
port 212 nsew signal input
rlabel metal2 s 148943 -480 148999 240 8 la_data_in[48]
port 213 nsew signal input
rlabel metal2 s 150691 -480 150747 240 8 la_data_in[49]
port 214 nsew signal input
rlabel metal2 s 70421 -480 70477 240 8 la_data_in[4]
port 215 nsew signal input
rlabel metal2 s 152485 -480 152541 240 8 la_data_in[50]
port 216 nsew signal input
rlabel metal2 s 154279 -480 154335 240 8 la_data_in[51]
port 217 nsew signal input
rlabel metal2 s 156073 -480 156129 240 8 la_data_in[52]
port 218 nsew signal input
rlabel metal2 s 157867 -480 157923 240 8 la_data_in[53]
port 219 nsew signal input
rlabel metal2 s 159615 -480 159671 240 8 la_data_in[54]
port 220 nsew signal input
rlabel metal2 s 161409 -480 161465 240 8 la_data_in[55]
port 221 nsew signal input
rlabel metal2 s 163203 -480 163259 240 8 la_data_in[56]
port 222 nsew signal input
rlabel metal2 s 164997 -480 165053 240 8 la_data_in[57]
port 223 nsew signal input
rlabel metal2 s 166791 -480 166847 240 8 la_data_in[58]
port 224 nsew signal input
rlabel metal2 s 168539 -480 168595 240 8 la_data_in[59]
port 225 nsew signal input
rlabel metal2 s 72215 -480 72271 240 8 la_data_in[5]
port 226 nsew signal input
rlabel metal2 s 170333 -480 170389 240 8 la_data_in[60]
port 227 nsew signal input
rlabel metal2 s 172127 -480 172183 240 8 la_data_in[61]
port 228 nsew signal input
rlabel metal2 s 173921 -480 173977 240 8 la_data_in[62]
port 229 nsew signal input
rlabel metal2 s 175669 -480 175725 240 8 la_data_in[63]
port 230 nsew signal input
rlabel metal2 s 177463 -480 177519 240 8 la_data_in[64]
port 231 nsew signal input
rlabel metal2 s 179257 -480 179313 240 8 la_data_in[65]
port 232 nsew signal input
rlabel metal2 s 181051 -480 181107 240 8 la_data_in[66]
port 233 nsew signal input
rlabel metal2 s 182845 -480 182901 240 8 la_data_in[67]
port 234 nsew signal input
rlabel metal2 s 184593 -480 184649 240 8 la_data_in[68]
port 235 nsew signal input
rlabel metal2 s 186387 -480 186443 240 8 la_data_in[69]
port 236 nsew signal input
rlabel metal2 s 74009 -480 74065 240 8 la_data_in[6]
port 237 nsew signal input
rlabel metal2 s 188181 -480 188237 240 8 la_data_in[70]
port 238 nsew signal input
rlabel metal2 s 189975 -480 190031 240 8 la_data_in[71]
port 239 nsew signal input
rlabel metal2 s 191769 -480 191825 240 8 la_data_in[72]
port 240 nsew signal input
rlabel metal2 s 193517 -480 193573 240 8 la_data_in[73]
port 241 nsew signal input
rlabel metal2 s 195311 -480 195367 240 8 la_data_in[74]
port 242 nsew signal input
rlabel metal2 s 197105 -480 197161 240 8 la_data_in[75]
port 243 nsew signal input
rlabel metal2 s 198899 -480 198955 240 8 la_data_in[76]
port 244 nsew signal input
rlabel metal2 s 200647 -480 200703 240 8 la_data_in[77]
port 245 nsew signal input
rlabel metal2 s 202441 -480 202497 240 8 la_data_in[78]
port 246 nsew signal input
rlabel metal2 s 204235 -480 204291 240 8 la_data_in[79]
port 247 nsew signal input
rlabel metal2 s 75757 -480 75813 240 8 la_data_in[7]
port 248 nsew signal input
rlabel metal2 s 206029 -480 206085 240 8 la_data_in[80]
port 249 nsew signal input
rlabel metal2 s 207823 -480 207879 240 8 la_data_in[81]
port 250 nsew signal input
rlabel metal2 s 209571 -480 209627 240 8 la_data_in[82]
port 251 nsew signal input
rlabel metal2 s 211365 -480 211421 240 8 la_data_in[83]
port 252 nsew signal input
rlabel metal2 s 213159 -480 213215 240 8 la_data_in[84]
port 253 nsew signal input
rlabel metal2 s 214953 -480 215009 240 8 la_data_in[85]
port 254 nsew signal input
rlabel metal2 s 216747 -480 216803 240 8 la_data_in[86]
port 255 nsew signal input
rlabel metal2 s 218495 -480 218551 240 8 la_data_in[87]
port 256 nsew signal input
rlabel metal2 s 220289 -480 220345 240 8 la_data_in[88]
port 257 nsew signal input
rlabel metal2 s 222083 -480 222139 240 8 la_data_in[89]
port 258 nsew signal input
rlabel metal2 s 77551 -480 77607 240 8 la_data_in[8]
port 259 nsew signal input
rlabel metal2 s 223877 -480 223933 240 8 la_data_in[90]
port 260 nsew signal input
rlabel metal2 s 225625 -480 225681 240 8 la_data_in[91]
port 261 nsew signal input
rlabel metal2 s 227419 -480 227475 240 8 la_data_in[92]
port 262 nsew signal input
rlabel metal2 s 229213 -480 229269 240 8 la_data_in[93]
port 263 nsew signal input
rlabel metal2 s 231007 -480 231063 240 8 la_data_in[94]
port 264 nsew signal input
rlabel metal2 s 232801 -480 232857 240 8 la_data_in[95]
port 265 nsew signal input
rlabel metal2 s 234549 -480 234605 240 8 la_data_in[96]
port 266 nsew signal input
rlabel metal2 s 236343 -480 236399 240 8 la_data_in[97]
port 267 nsew signal input
rlabel metal2 s 238137 -480 238193 240 8 la_data_in[98]
port 268 nsew signal input
rlabel metal2 s 239931 -480 239987 240 8 la_data_in[99]
port 269 nsew signal input
rlabel metal2 s 79345 -480 79401 240 8 la_data_in[9]
port 270 nsew signal input
rlabel metal2 s 63889 -480 63945 240 8 la_data_out[0]
port 271 nsew signal tristate
rlabel metal2 s 242277 -480 242333 240 8 la_data_out[100]
port 272 nsew signal tristate
rlabel metal2 s 244071 -480 244127 240 8 la_data_out[101]
port 273 nsew signal tristate
rlabel metal2 s 245865 -480 245921 240 8 la_data_out[102]
port 274 nsew signal tristate
rlabel metal2 s 247659 -480 247715 240 8 la_data_out[103]
port 275 nsew signal tristate
rlabel metal2 s 249453 -480 249509 240 8 la_data_out[104]
port 276 nsew signal tristate
rlabel metal2 s 251201 -480 251257 240 8 la_data_out[105]
port 277 nsew signal tristate
rlabel metal2 s 252995 -480 253051 240 8 la_data_out[106]
port 278 nsew signal tristate
rlabel metal2 s 254789 -480 254845 240 8 la_data_out[107]
port 279 nsew signal tristate
rlabel metal2 s 256583 -480 256639 240 8 la_data_out[108]
port 280 nsew signal tristate
rlabel metal2 s 258377 -480 258433 240 8 la_data_out[109]
port 281 nsew signal tristate
rlabel metal2 s 81737 -480 81793 240 8 la_data_out[10]
port 282 nsew signal tristate
rlabel metal2 s 260125 -480 260181 240 8 la_data_out[110]
port 283 nsew signal tristate
rlabel metal2 s 261919 -480 261975 240 8 la_data_out[111]
port 284 nsew signal tristate
rlabel metal2 s 263713 -480 263769 240 8 la_data_out[112]
port 285 nsew signal tristate
rlabel metal2 s 265507 -480 265563 240 8 la_data_out[113]
port 286 nsew signal tristate
rlabel metal2 s 267255 -480 267311 240 8 la_data_out[114]
port 287 nsew signal tristate
rlabel metal2 s 269049 -480 269105 240 8 la_data_out[115]
port 288 nsew signal tristate
rlabel metal2 s 270843 -480 270899 240 8 la_data_out[116]
port 289 nsew signal tristate
rlabel metal2 s 272637 -480 272693 240 8 la_data_out[117]
port 290 nsew signal tristate
rlabel metal2 s 274431 -480 274487 240 8 la_data_out[118]
port 291 nsew signal tristate
rlabel metal2 s 276179 -480 276235 240 8 la_data_out[119]
port 292 nsew signal tristate
rlabel metal2 s 83531 -480 83587 240 8 la_data_out[11]
port 293 nsew signal tristate
rlabel metal2 s 277973 -480 278029 240 8 la_data_out[120]
port 294 nsew signal tristate
rlabel metal2 s 279767 -480 279823 240 8 la_data_out[121]
port 295 nsew signal tristate
rlabel metal2 s 281561 -480 281617 240 8 la_data_out[122]
port 296 nsew signal tristate
rlabel metal2 s 283355 -480 283411 240 8 la_data_out[123]
port 297 nsew signal tristate
rlabel metal2 s 285103 -480 285159 240 8 la_data_out[124]
port 298 nsew signal tristate
rlabel metal2 s 286897 -480 286953 240 8 la_data_out[125]
port 299 nsew signal tristate
rlabel metal2 s 288691 -480 288747 240 8 la_data_out[126]
port 300 nsew signal tristate
rlabel metal2 s 290485 -480 290541 240 8 la_data_out[127]
port 301 nsew signal tristate
rlabel metal2 s 85279 -480 85335 240 8 la_data_out[12]
port 302 nsew signal tristate
rlabel metal2 s 87073 -480 87129 240 8 la_data_out[13]
port 303 nsew signal tristate
rlabel metal2 s 88867 -480 88923 240 8 la_data_out[14]
port 304 nsew signal tristate
rlabel metal2 s 90661 -480 90717 240 8 la_data_out[15]
port 305 nsew signal tristate
rlabel metal2 s 92409 -480 92465 240 8 la_data_out[16]
port 306 nsew signal tristate
rlabel metal2 s 94203 -480 94259 240 8 la_data_out[17]
port 307 nsew signal tristate
rlabel metal2 s 95997 -480 96053 240 8 la_data_out[18]
port 308 nsew signal tristate
rlabel metal2 s 97791 -480 97847 240 8 la_data_out[19]
port 309 nsew signal tristate
rlabel metal2 s 65683 -480 65739 240 8 la_data_out[1]
port 310 nsew signal tristate
rlabel metal2 s 99585 -480 99641 240 8 la_data_out[20]
port 311 nsew signal tristate
rlabel metal2 s 101333 -480 101389 240 8 la_data_out[21]
port 312 nsew signal tristate
rlabel metal2 s 103127 -480 103183 240 8 la_data_out[22]
port 313 nsew signal tristate
rlabel metal2 s 104921 -480 104977 240 8 la_data_out[23]
port 314 nsew signal tristate
rlabel metal2 s 106715 -480 106771 240 8 la_data_out[24]
port 315 nsew signal tristate
rlabel metal2 s 108509 -480 108565 240 8 la_data_out[25]
port 316 nsew signal tristate
rlabel metal2 s 110257 -480 110313 240 8 la_data_out[26]
port 317 nsew signal tristate
rlabel metal2 s 112051 -480 112107 240 8 la_data_out[27]
port 318 nsew signal tristate
rlabel metal2 s 113845 -480 113901 240 8 la_data_out[28]
port 319 nsew signal tristate
rlabel metal2 s 115639 -480 115695 240 8 la_data_out[29]
port 320 nsew signal tristate
rlabel metal2 s 67431 -480 67487 240 8 la_data_out[2]
port 321 nsew signal tristate
rlabel metal2 s 117387 -480 117443 240 8 la_data_out[30]
port 322 nsew signal tristate
rlabel metal2 s 119181 -480 119237 240 8 la_data_out[31]
port 323 nsew signal tristate
rlabel metal2 s 120975 -480 121031 240 8 la_data_out[32]
port 324 nsew signal tristate
rlabel metal2 s 122769 -480 122825 240 8 la_data_out[33]
port 325 nsew signal tristate
rlabel metal2 s 124563 -480 124619 240 8 la_data_out[34]
port 326 nsew signal tristate
rlabel metal2 s 126311 -480 126367 240 8 la_data_out[35]
port 327 nsew signal tristate
rlabel metal2 s 128105 -480 128161 240 8 la_data_out[36]
port 328 nsew signal tristate
rlabel metal2 s 129899 -480 129955 240 8 la_data_out[37]
port 329 nsew signal tristate
rlabel metal2 s 131693 -480 131749 240 8 la_data_out[38]
port 330 nsew signal tristate
rlabel metal2 s 133487 -480 133543 240 8 la_data_out[39]
port 331 nsew signal tristate
rlabel metal2 s 69225 -480 69281 240 8 la_data_out[3]
port 332 nsew signal tristate
rlabel metal2 s 135235 -480 135291 240 8 la_data_out[40]
port 333 nsew signal tristate
rlabel metal2 s 137029 -480 137085 240 8 la_data_out[41]
port 334 nsew signal tristate
rlabel metal2 s 138823 -480 138879 240 8 la_data_out[42]
port 335 nsew signal tristate
rlabel metal2 s 140617 -480 140673 240 8 la_data_out[43]
port 336 nsew signal tristate
rlabel metal2 s 142365 -480 142421 240 8 la_data_out[44]
port 337 nsew signal tristate
rlabel metal2 s 144159 -480 144215 240 8 la_data_out[45]
port 338 nsew signal tristate
rlabel metal2 s 145953 -480 146009 240 8 la_data_out[46]
port 339 nsew signal tristate
rlabel metal2 s 147747 -480 147803 240 8 la_data_out[47]
port 340 nsew signal tristate
rlabel metal2 s 149541 -480 149597 240 8 la_data_out[48]
port 341 nsew signal tristate
rlabel metal2 s 151289 -480 151345 240 8 la_data_out[49]
port 342 nsew signal tristate
rlabel metal2 s 71019 -480 71075 240 8 la_data_out[4]
port 343 nsew signal tristate
rlabel metal2 s 153083 -480 153139 240 8 la_data_out[50]
port 344 nsew signal tristate
rlabel metal2 s 154877 -480 154933 240 8 la_data_out[51]
port 345 nsew signal tristate
rlabel metal2 s 156671 -480 156727 240 8 la_data_out[52]
port 346 nsew signal tristate
rlabel metal2 s 158465 -480 158521 240 8 la_data_out[53]
port 347 nsew signal tristate
rlabel metal2 s 160213 -480 160269 240 8 la_data_out[54]
port 348 nsew signal tristate
rlabel metal2 s 162007 -480 162063 240 8 la_data_out[55]
port 349 nsew signal tristate
rlabel metal2 s 163801 -480 163857 240 8 la_data_out[56]
port 350 nsew signal tristate
rlabel metal2 s 165595 -480 165651 240 8 la_data_out[57]
port 351 nsew signal tristate
rlabel metal2 s 167343 -480 167399 240 8 la_data_out[58]
port 352 nsew signal tristate
rlabel metal2 s 169137 -480 169193 240 8 la_data_out[59]
port 353 nsew signal tristate
rlabel metal2 s 72813 -480 72869 240 8 la_data_out[5]
port 354 nsew signal tristate
rlabel metal2 s 170931 -480 170987 240 8 la_data_out[60]
port 355 nsew signal tristate
rlabel metal2 s 172725 -480 172781 240 8 la_data_out[61]
port 356 nsew signal tristate
rlabel metal2 s 174519 -480 174575 240 8 la_data_out[62]
port 357 nsew signal tristate
rlabel metal2 s 176267 -480 176323 240 8 la_data_out[63]
port 358 nsew signal tristate
rlabel metal2 s 178061 -480 178117 240 8 la_data_out[64]
port 359 nsew signal tristate
rlabel metal2 s 179855 -480 179911 240 8 la_data_out[65]
port 360 nsew signal tristate
rlabel metal2 s 181649 -480 181705 240 8 la_data_out[66]
port 361 nsew signal tristate
rlabel metal2 s 183443 -480 183499 240 8 la_data_out[67]
port 362 nsew signal tristate
rlabel metal2 s 185191 -480 185247 240 8 la_data_out[68]
port 363 nsew signal tristate
rlabel metal2 s 186985 -480 187041 240 8 la_data_out[69]
port 364 nsew signal tristate
rlabel metal2 s 74607 -480 74663 240 8 la_data_out[6]
port 365 nsew signal tristate
rlabel metal2 s 188779 -480 188835 240 8 la_data_out[70]
port 366 nsew signal tristate
rlabel metal2 s 190573 -480 190629 240 8 la_data_out[71]
port 367 nsew signal tristate
rlabel metal2 s 192321 -480 192377 240 8 la_data_out[72]
port 368 nsew signal tristate
rlabel metal2 s 194115 -480 194171 240 8 la_data_out[73]
port 369 nsew signal tristate
rlabel metal2 s 195909 -480 195965 240 8 la_data_out[74]
port 370 nsew signal tristate
rlabel metal2 s 197703 -480 197759 240 8 la_data_out[75]
port 371 nsew signal tristate
rlabel metal2 s 199497 -480 199553 240 8 la_data_out[76]
port 372 nsew signal tristate
rlabel metal2 s 201245 -480 201301 240 8 la_data_out[77]
port 373 nsew signal tristate
rlabel metal2 s 203039 -480 203095 240 8 la_data_out[78]
port 374 nsew signal tristate
rlabel metal2 s 204833 -480 204889 240 8 la_data_out[79]
port 375 nsew signal tristate
rlabel metal2 s 76355 -480 76411 240 8 la_data_out[7]
port 376 nsew signal tristate
rlabel metal2 s 206627 -480 206683 240 8 la_data_out[80]
port 377 nsew signal tristate
rlabel metal2 s 208421 -480 208477 240 8 la_data_out[81]
port 378 nsew signal tristate
rlabel metal2 s 210169 -480 210225 240 8 la_data_out[82]
port 379 nsew signal tristate
rlabel metal2 s 211963 -480 212019 240 8 la_data_out[83]
port 380 nsew signal tristate
rlabel metal2 s 213757 -480 213813 240 8 la_data_out[84]
port 381 nsew signal tristate
rlabel metal2 s 215551 -480 215607 240 8 la_data_out[85]
port 382 nsew signal tristate
rlabel metal2 s 217299 -480 217355 240 8 la_data_out[86]
port 383 nsew signal tristate
rlabel metal2 s 219093 -480 219149 240 8 la_data_out[87]
port 384 nsew signal tristate
rlabel metal2 s 220887 -480 220943 240 8 la_data_out[88]
port 385 nsew signal tristate
rlabel metal2 s 222681 -480 222737 240 8 la_data_out[89]
port 386 nsew signal tristate
rlabel metal2 s 78149 -480 78205 240 8 la_data_out[8]
port 387 nsew signal tristate
rlabel metal2 s 224475 -480 224531 240 8 la_data_out[90]
port 388 nsew signal tristate
rlabel metal2 s 226223 -480 226279 240 8 la_data_out[91]
port 389 nsew signal tristate
rlabel metal2 s 228017 -480 228073 240 8 la_data_out[92]
port 390 nsew signal tristate
rlabel metal2 s 229811 -480 229867 240 8 la_data_out[93]
port 391 nsew signal tristate
rlabel metal2 s 231605 -480 231661 240 8 la_data_out[94]
port 392 nsew signal tristate
rlabel metal2 s 233399 -480 233455 240 8 la_data_out[95]
port 393 nsew signal tristate
rlabel metal2 s 235147 -480 235203 240 8 la_data_out[96]
port 394 nsew signal tristate
rlabel metal2 s 236941 -480 236997 240 8 la_data_out[97]
port 395 nsew signal tristate
rlabel metal2 s 238735 -480 238791 240 8 la_data_out[98]
port 396 nsew signal tristate
rlabel metal2 s 240529 -480 240585 240 8 la_data_out[99]
port 397 nsew signal tristate
rlabel metal2 s 79943 -480 79999 240 8 la_data_out[9]
port 398 nsew signal tristate
rlabel metal2 s 64487 -480 64543 240 8 la_oen[0]
port 399 nsew signal input
rlabel metal2 s 242875 -480 242931 240 8 la_oen[100]
port 400 nsew signal input
rlabel metal2 s 244669 -480 244725 240 8 la_oen[101]
port 401 nsew signal input
rlabel metal2 s 246463 -480 246519 240 8 la_oen[102]
port 402 nsew signal input
rlabel metal2 s 248257 -480 248313 240 8 la_oen[103]
port 403 nsew signal input
rlabel metal2 s 250051 -480 250107 240 8 la_oen[104]
port 404 nsew signal input
rlabel metal2 s 251799 -480 251855 240 8 la_oen[105]
port 405 nsew signal input
rlabel metal2 s 253593 -480 253649 240 8 la_oen[106]
port 406 nsew signal input
rlabel metal2 s 255387 -480 255443 240 8 la_oen[107]
port 407 nsew signal input
rlabel metal2 s 257181 -480 257237 240 8 la_oen[108]
port 408 nsew signal input
rlabel metal2 s 258929 -480 258985 240 8 la_oen[109]
port 409 nsew signal input
rlabel metal2 s 82335 -480 82391 240 8 la_oen[10]
port 410 nsew signal input
rlabel metal2 s 260723 -480 260779 240 8 la_oen[110]
port 411 nsew signal input
rlabel metal2 s 262517 -480 262573 240 8 la_oen[111]
port 412 nsew signal input
rlabel metal2 s 264311 -480 264367 240 8 la_oen[112]
port 413 nsew signal input
rlabel metal2 s 266105 -480 266161 240 8 la_oen[113]
port 414 nsew signal input
rlabel metal2 s 267853 -480 267909 240 8 la_oen[114]
port 415 nsew signal input
rlabel metal2 s 269647 -480 269703 240 8 la_oen[115]
port 416 nsew signal input
rlabel metal2 s 271441 -480 271497 240 8 la_oen[116]
port 417 nsew signal input
rlabel metal2 s 273235 -480 273291 240 8 la_oen[117]
port 418 nsew signal input
rlabel metal2 s 275029 -480 275085 240 8 la_oen[118]
port 419 nsew signal input
rlabel metal2 s 276777 -480 276833 240 8 la_oen[119]
port 420 nsew signal input
rlabel metal2 s 84083 -480 84139 240 8 la_oen[11]
port 421 nsew signal input
rlabel metal2 s 278571 -480 278627 240 8 la_oen[120]
port 422 nsew signal input
rlabel metal2 s 280365 -480 280421 240 8 la_oen[121]
port 423 nsew signal input
rlabel metal2 s 282159 -480 282215 240 8 la_oen[122]
port 424 nsew signal input
rlabel metal2 s 283907 -480 283963 240 8 la_oen[123]
port 425 nsew signal input
rlabel metal2 s 285701 -480 285757 240 8 la_oen[124]
port 426 nsew signal input
rlabel metal2 s 287495 -480 287551 240 8 la_oen[125]
port 427 nsew signal input
rlabel metal2 s 289289 -480 289345 240 8 la_oen[126]
port 428 nsew signal input
rlabel metal2 s 291083 -480 291139 240 8 la_oen[127]
port 429 nsew signal input
rlabel metal2 s 85877 -480 85933 240 8 la_oen[12]
port 430 nsew signal input
rlabel metal2 s 87671 -480 87727 240 8 la_oen[13]
port 431 nsew signal input
rlabel metal2 s 89465 -480 89521 240 8 la_oen[14]
port 432 nsew signal input
rlabel metal2 s 91259 -480 91315 240 8 la_oen[15]
port 433 nsew signal input
rlabel metal2 s 93007 -480 93063 240 8 la_oen[16]
port 434 nsew signal input
rlabel metal2 s 94801 -480 94857 240 8 la_oen[17]
port 435 nsew signal input
rlabel metal2 s 96595 -480 96651 240 8 la_oen[18]
port 436 nsew signal input
rlabel metal2 s 98389 -480 98445 240 8 la_oen[19]
port 437 nsew signal input
rlabel metal2 s 66281 -480 66337 240 8 la_oen[1]
port 438 nsew signal input
rlabel metal2 s 100183 -480 100239 240 8 la_oen[20]
port 439 nsew signal input
rlabel metal2 s 101931 -480 101987 240 8 la_oen[21]
port 440 nsew signal input
rlabel metal2 s 103725 -480 103781 240 8 la_oen[22]
port 441 nsew signal input
rlabel metal2 s 105519 -480 105575 240 8 la_oen[23]
port 442 nsew signal input
rlabel metal2 s 107313 -480 107369 240 8 la_oen[24]
port 443 nsew signal input
rlabel metal2 s 109061 -480 109117 240 8 la_oen[25]
port 444 nsew signal input
rlabel metal2 s 110855 -480 110911 240 8 la_oen[26]
port 445 nsew signal input
rlabel metal2 s 112649 -480 112705 240 8 la_oen[27]
port 446 nsew signal input
rlabel metal2 s 114443 -480 114499 240 8 la_oen[28]
port 447 nsew signal input
rlabel metal2 s 116237 -480 116293 240 8 la_oen[29]
port 448 nsew signal input
rlabel metal2 s 68029 -480 68085 240 8 la_oen[2]
port 449 nsew signal input
rlabel metal2 s 117985 -480 118041 240 8 la_oen[30]
port 450 nsew signal input
rlabel metal2 s 119779 -480 119835 240 8 la_oen[31]
port 451 nsew signal input
rlabel metal2 s 121573 -480 121629 240 8 la_oen[32]
port 452 nsew signal input
rlabel metal2 s 123367 -480 123423 240 8 la_oen[33]
port 453 nsew signal input
rlabel metal2 s 125161 -480 125217 240 8 la_oen[34]
port 454 nsew signal input
rlabel metal2 s 126909 -480 126965 240 8 la_oen[35]
port 455 nsew signal input
rlabel metal2 s 128703 -480 128759 240 8 la_oen[36]
port 456 nsew signal input
rlabel metal2 s 130497 -480 130553 240 8 la_oen[37]
port 457 nsew signal input
rlabel metal2 s 132291 -480 132347 240 8 la_oen[38]
port 458 nsew signal input
rlabel metal2 s 134039 -480 134095 240 8 la_oen[39]
port 459 nsew signal input
rlabel metal2 s 69823 -480 69879 240 8 la_oen[3]
port 460 nsew signal input
rlabel metal2 s 135833 -480 135889 240 8 la_oen[40]
port 461 nsew signal input
rlabel metal2 s 137627 -480 137683 240 8 la_oen[41]
port 462 nsew signal input
rlabel metal2 s 139421 -480 139477 240 8 la_oen[42]
port 463 nsew signal input
rlabel metal2 s 141215 -480 141271 240 8 la_oen[43]
port 464 nsew signal input
rlabel metal2 s 142963 -480 143019 240 8 la_oen[44]
port 465 nsew signal input
rlabel metal2 s 144757 -480 144813 240 8 la_oen[45]
port 466 nsew signal input
rlabel metal2 s 146551 -480 146607 240 8 la_oen[46]
port 467 nsew signal input
rlabel metal2 s 148345 -480 148401 240 8 la_oen[47]
port 468 nsew signal input
rlabel metal2 s 150139 -480 150195 240 8 la_oen[48]
port 469 nsew signal input
rlabel metal2 s 151887 -480 151943 240 8 la_oen[49]
port 470 nsew signal input
rlabel metal2 s 71617 -480 71673 240 8 la_oen[4]
port 471 nsew signal input
rlabel metal2 s 153681 -480 153737 240 8 la_oen[50]
port 472 nsew signal input
rlabel metal2 s 155475 -480 155531 240 8 la_oen[51]
port 473 nsew signal input
rlabel metal2 s 157269 -480 157325 240 8 la_oen[52]
port 474 nsew signal input
rlabel metal2 s 159017 -480 159073 240 8 la_oen[53]
port 475 nsew signal input
rlabel metal2 s 160811 -480 160867 240 8 la_oen[54]
port 476 nsew signal input
rlabel metal2 s 162605 -480 162661 240 8 la_oen[55]
port 477 nsew signal input
rlabel metal2 s 164399 -480 164455 240 8 la_oen[56]
port 478 nsew signal input
rlabel metal2 s 166193 -480 166249 240 8 la_oen[57]
port 479 nsew signal input
rlabel metal2 s 167941 -480 167997 240 8 la_oen[58]
port 480 nsew signal input
rlabel metal2 s 169735 -480 169791 240 8 la_oen[59]
port 481 nsew signal input
rlabel metal2 s 73411 -480 73467 240 8 la_oen[5]
port 482 nsew signal input
rlabel metal2 s 171529 -480 171585 240 8 la_oen[60]
port 483 nsew signal input
rlabel metal2 s 173323 -480 173379 240 8 la_oen[61]
port 484 nsew signal input
rlabel metal2 s 175117 -480 175173 240 8 la_oen[62]
port 485 nsew signal input
rlabel metal2 s 176865 -480 176921 240 8 la_oen[63]
port 486 nsew signal input
rlabel metal2 s 178659 -480 178715 240 8 la_oen[64]
port 487 nsew signal input
rlabel metal2 s 180453 -480 180509 240 8 la_oen[65]
port 488 nsew signal input
rlabel metal2 s 182247 -480 182303 240 8 la_oen[66]
port 489 nsew signal input
rlabel metal2 s 183995 -480 184051 240 8 la_oen[67]
port 490 nsew signal input
rlabel metal2 s 185789 -480 185845 240 8 la_oen[68]
port 491 nsew signal input
rlabel metal2 s 187583 -480 187639 240 8 la_oen[69]
port 492 nsew signal input
rlabel metal2 s 75205 -480 75261 240 8 la_oen[6]
port 493 nsew signal input
rlabel metal2 s 189377 -480 189433 240 8 la_oen[70]
port 494 nsew signal input
rlabel metal2 s 191171 -480 191227 240 8 la_oen[71]
port 495 nsew signal input
rlabel metal2 s 192919 -480 192975 240 8 la_oen[72]
port 496 nsew signal input
rlabel metal2 s 194713 -480 194769 240 8 la_oen[73]
port 497 nsew signal input
rlabel metal2 s 196507 -480 196563 240 8 la_oen[74]
port 498 nsew signal input
rlabel metal2 s 198301 -480 198357 240 8 la_oen[75]
port 499 nsew signal input
rlabel metal2 s 200095 -480 200151 240 8 la_oen[76]
port 500 nsew signal input
rlabel metal2 s 201843 -480 201899 240 8 la_oen[77]
port 501 nsew signal input
rlabel metal2 s 203637 -480 203693 240 8 la_oen[78]
port 502 nsew signal input
rlabel metal2 s 205431 -480 205487 240 8 la_oen[79]
port 503 nsew signal input
rlabel metal2 s 76953 -480 77009 240 8 la_oen[7]
port 504 nsew signal input
rlabel metal2 s 207225 -480 207281 240 8 la_oen[80]
port 505 nsew signal input
rlabel metal2 s 208973 -480 209029 240 8 la_oen[81]
port 506 nsew signal input
rlabel metal2 s 210767 -480 210823 240 8 la_oen[82]
port 507 nsew signal input
rlabel metal2 s 212561 -480 212617 240 8 la_oen[83]
port 508 nsew signal input
rlabel metal2 s 214355 -480 214411 240 8 la_oen[84]
port 509 nsew signal input
rlabel metal2 s 216149 -480 216205 240 8 la_oen[85]
port 510 nsew signal input
rlabel metal2 s 217897 -480 217953 240 8 la_oen[86]
port 511 nsew signal input
rlabel metal2 s 219691 -480 219747 240 8 la_oen[87]
port 512 nsew signal input
rlabel metal2 s 221485 -480 221541 240 8 la_oen[88]
port 513 nsew signal input
rlabel metal2 s 223279 -480 223335 240 8 la_oen[89]
port 514 nsew signal input
rlabel metal2 s 78747 -480 78803 240 8 la_oen[8]
port 515 nsew signal input
rlabel metal2 s 225073 -480 225129 240 8 la_oen[90]
port 516 nsew signal input
rlabel metal2 s 226821 -480 226877 240 8 la_oen[91]
port 517 nsew signal input
rlabel metal2 s 228615 -480 228671 240 8 la_oen[92]
port 518 nsew signal input
rlabel metal2 s 230409 -480 230465 240 8 la_oen[93]
port 519 nsew signal input
rlabel metal2 s 232203 -480 232259 240 8 la_oen[94]
port 520 nsew signal input
rlabel metal2 s 233951 -480 234007 240 8 la_oen[95]
port 521 nsew signal input
rlabel metal2 s 235745 -480 235801 240 8 la_oen[96]
port 522 nsew signal input
rlabel metal2 s 237539 -480 237595 240 8 la_oen[97]
port 523 nsew signal input
rlabel metal2 s 239333 -480 239389 240 8 la_oen[98]
port 524 nsew signal input
rlabel metal2 s 241127 -480 241183 240 8 la_oen[99]
port 525 nsew signal input
rlabel metal2 s 80541 -480 80597 240 8 la_oen[9]
port 526 nsew signal input
rlabel metal2 s 291681 -480 291737 240 8 user_clock2
port 527 nsew signal input
rlabel metal2 s 271 -480 327 240 8 wb_clk_i
port 528 nsew signal input
rlabel metal2 s 823 -480 879 240 8 wb_rst_i
port 529 nsew signal input
rlabel metal2 s 1421 -480 1477 240 8 wbs_ack_o
port 530 nsew signal tristate
rlabel metal2 s 3813 -480 3869 240 8 wbs_adr_i[0]
port 531 nsew signal input
rlabel metal2 s 24053 -480 24109 240 8 wbs_adr_i[10]
port 532 nsew signal input
rlabel metal2 s 25801 -480 25857 240 8 wbs_adr_i[11]
port 533 nsew signal input
rlabel metal2 s 27595 -480 27651 240 8 wbs_adr_i[12]
port 534 nsew signal input
rlabel metal2 s 29389 -480 29445 240 8 wbs_adr_i[13]
port 535 nsew signal input
rlabel metal2 s 31183 -480 31239 240 8 wbs_adr_i[14]
port 536 nsew signal input
rlabel metal2 s 32977 -480 33033 240 8 wbs_adr_i[15]
port 537 nsew signal input
rlabel metal2 s 34725 -480 34781 240 8 wbs_adr_i[16]
port 538 nsew signal input
rlabel metal2 s 36519 -480 36575 240 8 wbs_adr_i[17]
port 539 nsew signal input
rlabel metal2 s 38313 -480 38369 240 8 wbs_adr_i[18]
port 540 nsew signal input
rlabel metal2 s 40107 -480 40163 240 8 wbs_adr_i[19]
port 541 nsew signal input
rlabel metal2 s 6205 -480 6261 240 8 wbs_adr_i[1]
port 542 nsew signal input
rlabel metal2 s 41901 -480 41957 240 8 wbs_adr_i[20]
port 543 nsew signal input
rlabel metal2 s 43649 -480 43705 240 8 wbs_adr_i[21]
port 544 nsew signal input
rlabel metal2 s 45443 -480 45499 240 8 wbs_adr_i[22]
port 545 nsew signal input
rlabel metal2 s 47237 -480 47293 240 8 wbs_adr_i[23]
port 546 nsew signal input
rlabel metal2 s 49031 -480 49087 240 8 wbs_adr_i[24]
port 547 nsew signal input
rlabel metal2 s 50779 -480 50835 240 8 wbs_adr_i[25]
port 548 nsew signal input
rlabel metal2 s 52573 -480 52629 240 8 wbs_adr_i[26]
port 549 nsew signal input
rlabel metal2 s 54367 -480 54423 240 8 wbs_adr_i[27]
port 550 nsew signal input
rlabel metal2 s 56161 -480 56217 240 8 wbs_adr_i[28]
port 551 nsew signal input
rlabel metal2 s 57955 -480 58011 240 8 wbs_adr_i[29]
port 552 nsew signal input
rlabel metal2 s 8597 -480 8653 240 8 wbs_adr_i[2]
port 553 nsew signal input
rlabel metal2 s 59703 -480 59759 240 8 wbs_adr_i[30]
port 554 nsew signal input
rlabel metal2 s 61497 -480 61553 240 8 wbs_adr_i[31]
port 555 nsew signal input
rlabel metal2 s 10943 -480 10999 240 8 wbs_adr_i[3]
port 556 nsew signal input
rlabel metal2 s 13335 -480 13391 240 8 wbs_adr_i[4]
port 557 nsew signal input
rlabel metal2 s 15129 -480 15185 240 8 wbs_adr_i[5]
port 558 nsew signal input
rlabel metal2 s 16923 -480 16979 240 8 wbs_adr_i[6]
port 559 nsew signal input
rlabel metal2 s 18671 -480 18727 240 8 wbs_adr_i[7]
port 560 nsew signal input
rlabel metal2 s 20465 -480 20521 240 8 wbs_adr_i[8]
port 561 nsew signal input
rlabel metal2 s 22259 -480 22315 240 8 wbs_adr_i[9]
port 562 nsew signal input
rlabel metal2 s 2019 -480 2075 240 8 wbs_cyc_i
port 563 nsew signal input
rlabel metal2 s 4411 -480 4467 240 8 wbs_dat_i[0]
port 564 nsew signal input
rlabel metal2 s 24651 -480 24707 240 8 wbs_dat_i[10]
port 565 nsew signal input
rlabel metal2 s 26399 -480 26455 240 8 wbs_dat_i[11]
port 566 nsew signal input
rlabel metal2 s 28193 -480 28249 240 8 wbs_dat_i[12]
port 567 nsew signal input
rlabel metal2 s 29987 -480 30043 240 8 wbs_dat_i[13]
port 568 nsew signal input
rlabel metal2 s 31781 -480 31837 240 8 wbs_dat_i[14]
port 569 nsew signal input
rlabel metal2 s 33575 -480 33631 240 8 wbs_dat_i[15]
port 570 nsew signal input
rlabel metal2 s 35323 -480 35379 240 8 wbs_dat_i[16]
port 571 nsew signal input
rlabel metal2 s 37117 -480 37173 240 8 wbs_dat_i[17]
port 572 nsew signal input
rlabel metal2 s 38911 -480 38967 240 8 wbs_dat_i[18]
port 573 nsew signal input
rlabel metal2 s 40705 -480 40761 240 8 wbs_dat_i[19]
port 574 nsew signal input
rlabel metal2 s 6803 -480 6859 240 8 wbs_dat_i[1]
port 575 nsew signal input
rlabel metal2 s 42453 -480 42509 240 8 wbs_dat_i[20]
port 576 nsew signal input
rlabel metal2 s 44247 -480 44303 240 8 wbs_dat_i[21]
port 577 nsew signal input
rlabel metal2 s 46041 -480 46097 240 8 wbs_dat_i[22]
port 578 nsew signal input
rlabel metal2 s 47835 -480 47891 240 8 wbs_dat_i[23]
port 579 nsew signal input
rlabel metal2 s 49629 -480 49685 240 8 wbs_dat_i[24]
port 580 nsew signal input
rlabel metal2 s 51377 -480 51433 240 8 wbs_dat_i[25]
port 581 nsew signal input
rlabel metal2 s 53171 -480 53227 240 8 wbs_dat_i[26]
port 582 nsew signal input
rlabel metal2 s 54965 -480 55021 240 8 wbs_dat_i[27]
port 583 nsew signal input
rlabel metal2 s 56759 -480 56815 240 8 wbs_dat_i[28]
port 584 nsew signal input
rlabel metal2 s 58553 -480 58609 240 8 wbs_dat_i[29]
port 585 nsew signal input
rlabel metal2 s 9149 -480 9205 240 8 wbs_dat_i[2]
port 586 nsew signal input
rlabel metal2 s 60301 -480 60357 240 8 wbs_dat_i[30]
port 587 nsew signal input
rlabel metal2 s 62095 -480 62151 240 8 wbs_dat_i[31]
port 588 nsew signal input
rlabel metal2 s 11541 -480 11597 240 8 wbs_dat_i[3]
port 589 nsew signal input
rlabel metal2 s 13933 -480 13989 240 8 wbs_dat_i[4]
port 590 nsew signal input
rlabel metal2 s 15727 -480 15783 240 8 wbs_dat_i[5]
port 591 nsew signal input
rlabel metal2 s 17475 -480 17531 240 8 wbs_dat_i[6]
port 592 nsew signal input
rlabel metal2 s 19269 -480 19325 240 8 wbs_dat_i[7]
port 593 nsew signal input
rlabel metal2 s 21063 -480 21119 240 8 wbs_dat_i[8]
port 594 nsew signal input
rlabel metal2 s 22857 -480 22913 240 8 wbs_dat_i[9]
port 595 nsew signal input
rlabel metal2 s 5009 -480 5065 240 8 wbs_dat_o[0]
port 596 nsew signal tristate
rlabel metal2 s 25249 -480 25305 240 8 wbs_dat_o[10]
port 597 nsew signal tristate
rlabel metal2 s 26997 -480 27053 240 8 wbs_dat_o[11]
port 598 nsew signal tristate
rlabel metal2 s 28791 -480 28847 240 8 wbs_dat_o[12]
port 599 nsew signal tristate
rlabel metal2 s 30585 -480 30641 240 8 wbs_dat_o[13]
port 600 nsew signal tristate
rlabel metal2 s 32379 -480 32435 240 8 wbs_dat_o[14]
port 601 nsew signal tristate
rlabel metal2 s 34127 -480 34183 240 8 wbs_dat_o[15]
port 602 nsew signal tristate
rlabel metal2 s 35921 -480 35977 240 8 wbs_dat_o[16]
port 603 nsew signal tristate
rlabel metal2 s 37715 -480 37771 240 8 wbs_dat_o[17]
port 604 nsew signal tristate
rlabel metal2 s 39509 -480 39565 240 8 wbs_dat_o[18]
port 605 nsew signal tristate
rlabel metal2 s 41303 -480 41359 240 8 wbs_dat_o[19]
port 606 nsew signal tristate
rlabel metal2 s 7401 -480 7457 240 8 wbs_dat_o[1]
port 607 nsew signal tristate
rlabel metal2 s 43051 -480 43107 240 8 wbs_dat_o[20]
port 608 nsew signal tristate
rlabel metal2 s 44845 -480 44901 240 8 wbs_dat_o[21]
port 609 nsew signal tristate
rlabel metal2 s 46639 -480 46695 240 8 wbs_dat_o[22]
port 610 nsew signal tristate
rlabel metal2 s 48433 -480 48489 240 8 wbs_dat_o[23]
port 611 nsew signal tristate
rlabel metal2 s 50227 -480 50283 240 8 wbs_dat_o[24]
port 612 nsew signal tristate
rlabel metal2 s 51975 -480 52031 240 8 wbs_dat_o[25]
port 613 nsew signal tristate
rlabel metal2 s 53769 -480 53825 240 8 wbs_dat_o[26]
port 614 nsew signal tristate
rlabel metal2 s 55563 -480 55619 240 8 wbs_dat_o[27]
port 615 nsew signal tristate
rlabel metal2 s 57357 -480 57413 240 8 wbs_dat_o[28]
port 616 nsew signal tristate
rlabel metal2 s 59105 -480 59161 240 8 wbs_dat_o[29]
port 617 nsew signal tristate
rlabel metal2 s 9747 -480 9803 240 8 wbs_dat_o[2]
port 618 nsew signal tristate
rlabel metal2 s 60899 -480 60955 240 8 wbs_dat_o[30]
port 619 nsew signal tristate
rlabel metal2 s 62693 -480 62749 240 8 wbs_dat_o[31]
port 620 nsew signal tristate
rlabel metal2 s 12139 -480 12195 240 8 wbs_dat_o[3]
port 621 nsew signal tristate
rlabel metal2 s 14531 -480 14587 240 8 wbs_dat_o[4]
port 622 nsew signal tristate
rlabel metal2 s 16325 -480 16381 240 8 wbs_dat_o[5]
port 623 nsew signal tristate
rlabel metal2 s 18073 -480 18129 240 8 wbs_dat_o[6]
port 624 nsew signal tristate
rlabel metal2 s 19867 -480 19923 240 8 wbs_dat_o[7]
port 625 nsew signal tristate
rlabel metal2 s 21661 -480 21717 240 8 wbs_dat_o[8]
port 626 nsew signal tristate
rlabel metal2 s 23455 -480 23511 240 8 wbs_dat_o[9]
port 627 nsew signal tristate
rlabel metal2 s 5607 -480 5663 240 8 wbs_sel_i[0]
port 628 nsew signal input
rlabel metal2 s 7999 -480 8055 240 8 wbs_sel_i[1]
port 629 nsew signal input
rlabel metal2 s 10345 -480 10401 240 8 wbs_sel_i[2]
port 630 nsew signal input
rlabel metal2 s 12737 -480 12793 240 8 wbs_sel_i[3]
port 631 nsew signal input
rlabel metal2 s 2617 -480 2673 240 8 wbs_stb_i
port 632 nsew signal input
rlabel metal2 s 3215 -480 3271 240 8 wbs_we_i
port 633 nsew signal input
rlabel metal4 s 288902 -932 289202 352900 6 vccd1
port 634 nsew power bidirectional
rlabel metal4 s 270902 -932 271202 352900 6 vccd1.extra1
port 635 nsew power bidirectional
rlabel metal4 s 252902 -932 253202 352900 6 vccd1.extra2
port 636 nsew power bidirectional
rlabel metal4 s 234902 -932 235202 352900 6 vccd1.extra3
port 637 nsew power bidirectional
rlabel metal4 s 216902 -932 217202 352900 6 vccd1.extra4
port 638 nsew power bidirectional
rlabel metal4 s 198902 -932 199202 352900 6 vccd1.extra5
port 639 nsew power bidirectional
rlabel metal4 s 180902 -932 181202 352900 6 vccd1.extra6
port 640 nsew power bidirectional
rlabel metal4 s 162902 -932 163202 352900 6 vccd1.extra7
port 641 nsew power bidirectional
rlabel metal4 s 144902 -932 145202 352900 6 vccd1.extra8
port 642 nsew power bidirectional
rlabel metal4 s 126902 -932 127202 352900 6 vccd1.extra9
port 643 nsew power bidirectional
rlabel metal4 s 108902 -932 109202 352900 6 vccd1.extra10
port 644 nsew power bidirectional
rlabel metal4 s 90902 -932 91202 352900 6 vccd1.extra11
port 645 nsew power bidirectional
rlabel metal4 s 72902 -932 73202 352900 6 vccd1.extra12
port 646 nsew power bidirectional
rlabel metal4 s 54902 -932 55202 352900 6 vccd1.extra13
port 647 nsew power bidirectional
rlabel metal4 s 36902 -932 37202 352900 6 vccd1.extra14
port 648 nsew power bidirectional
rlabel metal4 s 18902 -932 19202 352900 6 vccd1.extra15
port 649 nsew power bidirectional
rlabel metal4 s 902 -932 1202 352900 6 vccd1.extra16
port 650 nsew power bidirectional
rlabel metal4 s 292660 -462 292960 352430 6 vccd1.extra17
port 651 nsew power bidirectional
rlabel metal4 s -998 -462 -698 352430 4 vccd1.extra18
port 652 nsew power bidirectional
rlabel metal5 s -998 352130 292960 352430 6 vccd1.extra19
port 653 nsew power bidirectional
rlabel metal5 s -1468 343438 293430 343738 6 vccd1.extra20
port 654 nsew power bidirectional
rlabel metal5 s -1468 325438 293430 325738 6 vccd1.extra21
port 655 nsew power bidirectional
rlabel metal5 s -1468 307438 293430 307738 6 vccd1.extra22
port 656 nsew power bidirectional
rlabel metal5 s -1468 289438 293430 289738 6 vccd1.extra23
port 657 nsew power bidirectional
rlabel metal5 s -1468 271438 293430 271738 6 vccd1.extra24
port 658 nsew power bidirectional
rlabel metal5 s -1468 253438 293430 253738 6 vccd1.extra25
port 659 nsew power bidirectional
rlabel metal5 s -1468 235438 293430 235738 6 vccd1.extra26
port 660 nsew power bidirectional
rlabel metal5 s -1468 217438 293430 217738 6 vccd1.extra27
port 661 nsew power bidirectional
rlabel metal5 s -1468 199438 293430 199738 6 vccd1.extra28
port 662 nsew power bidirectional
rlabel metal5 s -1468 181438 293430 181738 6 vccd1.extra29
port 663 nsew power bidirectional
rlabel metal5 s -1468 163438 293430 163738 6 vccd1.extra30
port 664 nsew power bidirectional
rlabel metal5 s -1468 145438 293430 145738 6 vccd1.extra31
port 665 nsew power bidirectional
rlabel metal5 s -1468 127438 293430 127738 6 vccd1.extra32
port 666 nsew power bidirectional
rlabel metal5 s -1468 109438 293430 109738 6 vccd1.extra33
port 667 nsew power bidirectional
rlabel metal5 s -1468 91438 293430 91738 6 vccd1.extra34
port 668 nsew power bidirectional
rlabel metal5 s -1468 73438 293430 73738 6 vccd1.extra35
port 669 nsew power bidirectional
rlabel metal5 s -1468 55438 293430 55738 6 vccd1.extra36
port 670 nsew power bidirectional
rlabel metal5 s -1468 37438 293430 37738 6 vccd1.extra37
port 671 nsew power bidirectional
rlabel metal5 s -1468 19438 293430 19738 6 vccd1.extra38
port 672 nsew power bidirectional
rlabel metal5 s -1468 1438 293430 1738 6 vccd1.extra39
port 673 nsew power bidirectional
rlabel metal5 s -998 -462 292960 -162 8 vccd1.extra40
port 674 nsew power bidirectional
rlabel metal4 s 293130 -932 293430 352900 6 vssd1
port 675 nsew ground bidirectional
rlabel metal4 s 279902 -932 280202 352900 6 vssd1.extra1
port 676 nsew ground bidirectional
rlabel metal4 s 261902 -932 262202 352900 6 vssd1.extra2
port 677 nsew ground bidirectional
rlabel metal4 s 243902 -932 244202 352900 6 vssd1.extra3
port 678 nsew ground bidirectional
rlabel metal4 s 225902 -932 226202 352900 6 vssd1.extra4
port 679 nsew ground bidirectional
rlabel metal4 s 207902 -932 208202 352900 6 vssd1.extra5
port 680 nsew ground bidirectional
rlabel metal4 s 189902 -932 190202 352900 6 vssd1.extra6
port 681 nsew ground bidirectional
rlabel metal4 s 171902 -932 172202 352900 6 vssd1.extra7
port 682 nsew ground bidirectional
rlabel metal4 s 153902 -932 154202 352900 6 vssd1.extra8
port 683 nsew ground bidirectional
rlabel metal4 s 135902 -932 136202 352900 6 vssd1.extra9
port 684 nsew ground bidirectional
rlabel metal4 s 117902 -932 118202 352900 6 vssd1.extra10
port 685 nsew ground bidirectional
rlabel metal4 s 99902 -932 100202 352900 6 vssd1.extra11
port 686 nsew ground bidirectional
rlabel metal4 s 81902 -932 82202 352900 6 vssd1.extra12
port 687 nsew ground bidirectional
rlabel metal4 s 63902 -932 64202 352900 6 vssd1.extra13
port 688 nsew ground bidirectional
rlabel metal4 s 45902 -932 46202 352900 6 vssd1.extra14
port 689 nsew ground bidirectional
rlabel metal4 s 27902 -932 28202 352900 6 vssd1.extra15
port 690 nsew ground bidirectional
rlabel metal4 s 9902 -932 10202 352900 6 vssd1.extra16
port 691 nsew ground bidirectional
rlabel metal4 s -1468 -932 -1168 352900 4 vssd1.extra17
port 692 nsew ground bidirectional
rlabel metal5 s -1468 352600 293430 352900 6 vssd1.extra18
port 693 nsew ground bidirectional
rlabel metal5 s -1468 334438 293430 334738 6 vssd1.extra19
port 694 nsew ground bidirectional
rlabel metal5 s -1468 316438 293430 316738 6 vssd1.extra20
port 695 nsew ground bidirectional
rlabel metal5 s -1468 298438 293430 298738 6 vssd1.extra21
port 696 nsew ground bidirectional
rlabel metal5 s -1468 280438 293430 280738 6 vssd1.extra22
port 697 nsew ground bidirectional
rlabel metal5 s -1468 262438 293430 262738 6 vssd1.extra23
port 698 nsew ground bidirectional
rlabel metal5 s -1468 244438 293430 244738 6 vssd1.extra24
port 699 nsew ground bidirectional
rlabel metal5 s -1468 226438 293430 226738 6 vssd1.extra25
port 700 nsew ground bidirectional
rlabel metal5 s -1468 208438 293430 208738 6 vssd1.extra26
port 701 nsew ground bidirectional
rlabel metal5 s -1468 190438 293430 190738 6 vssd1.extra27
port 702 nsew ground bidirectional
rlabel metal5 s -1468 172438 293430 172738 6 vssd1.extra28
port 703 nsew ground bidirectional
rlabel metal5 s -1468 154438 293430 154738 6 vssd1.extra29
port 704 nsew ground bidirectional
rlabel metal5 s -1468 136438 293430 136738 6 vssd1.extra30
port 705 nsew ground bidirectional
rlabel metal5 s -1468 118438 293430 118738 6 vssd1.extra31
port 706 nsew ground bidirectional
rlabel metal5 s -1468 100438 293430 100738 6 vssd1.extra32
port 707 nsew ground bidirectional
rlabel metal5 s -1468 82438 293430 82738 6 vssd1.extra33
port 708 nsew ground bidirectional
rlabel metal5 s -1468 64438 293430 64738 6 vssd1.extra34
port 709 nsew ground bidirectional
rlabel metal5 s -1468 46438 293430 46738 6 vssd1.extra35
port 710 nsew ground bidirectional
rlabel metal5 s -1468 28438 293430 28738 6 vssd1.extra36
port 711 nsew ground bidirectional
rlabel metal5 s -1468 10438 293430 10738 6 vssd1.extra37
port 712 nsew ground bidirectional
rlabel metal5 s -1468 -932 293430 -632 8 vssd1.extra38
port 713 nsew ground bidirectional
rlabel metal4 s 290702 -1872 291002 353840 6 vccd2
port 714 nsew power bidirectional
rlabel metal4 s 272702 -1872 273002 353840 6 vccd2.extra1
port 715 nsew power bidirectional
rlabel metal4 s 254702 -1872 255002 353840 6 vccd2.extra2
port 716 nsew power bidirectional
rlabel metal4 s 236702 -1872 237002 353840 6 vccd2.extra3
port 717 nsew power bidirectional
rlabel metal4 s 218702 -1872 219002 353840 6 vccd2.extra4
port 718 nsew power bidirectional
rlabel metal4 s 200702 -1872 201002 353840 6 vccd2.extra5
port 719 nsew power bidirectional
rlabel metal4 s 182702 -1872 183002 353840 6 vccd2.extra6
port 720 nsew power bidirectional
rlabel metal4 s 164702 -1872 165002 353840 6 vccd2.extra7
port 721 nsew power bidirectional
rlabel metal4 s 146702 -1872 147002 353840 6 vccd2.extra8
port 722 nsew power bidirectional
rlabel metal4 s 128702 -1872 129002 353840 6 vccd2.extra9
port 723 nsew power bidirectional
rlabel metal4 s 110702 -1872 111002 353840 6 vccd2.extra10
port 724 nsew power bidirectional
rlabel metal4 s 92702 -1872 93002 353840 6 vccd2.extra11
port 725 nsew power bidirectional
rlabel metal4 s 74702 -1872 75002 353840 6 vccd2.extra12
port 726 nsew power bidirectional
rlabel metal4 s 56702 -1872 57002 353840 6 vccd2.extra13
port 727 nsew power bidirectional
rlabel metal4 s 38702 -1872 39002 353840 6 vccd2.extra14
port 728 nsew power bidirectional
rlabel metal4 s 20702 -1872 21002 353840 6 vccd2.extra15
port 729 nsew power bidirectional
rlabel metal4 s 2702 -1872 3002 353840 6 vccd2.extra16
port 730 nsew power bidirectional
rlabel metal4 s 293600 -1402 293900 353370 6 vccd2.extra17
port 731 nsew power bidirectional
rlabel metal4 s -1938 -1402 -1638 353370 4 vccd2.extra18
port 732 nsew power bidirectional
rlabel metal5 s -1938 353070 293900 353370 6 vccd2.extra19
port 733 nsew power bidirectional
rlabel metal5 s -2408 345238 294370 345538 6 vccd2.extra20
port 734 nsew power bidirectional
rlabel metal5 s -2408 327238 294370 327538 6 vccd2.extra21
port 735 nsew power bidirectional
rlabel metal5 s -2408 309238 294370 309538 6 vccd2.extra22
port 736 nsew power bidirectional
rlabel metal5 s -2408 291238 294370 291538 6 vccd2.extra23
port 737 nsew power bidirectional
rlabel metal5 s -2408 273238 294370 273538 6 vccd2.extra24
port 738 nsew power bidirectional
rlabel metal5 s -2408 255238 294370 255538 6 vccd2.extra25
port 739 nsew power bidirectional
rlabel metal5 s -2408 237238 294370 237538 6 vccd2.extra26
port 740 nsew power bidirectional
rlabel metal5 s -2408 219238 294370 219538 6 vccd2.extra27
port 741 nsew power bidirectional
rlabel metal5 s -2408 201238 294370 201538 6 vccd2.extra28
port 742 nsew power bidirectional
rlabel metal5 s -2408 183238 294370 183538 6 vccd2.extra29
port 743 nsew power bidirectional
rlabel metal5 s -2408 165238 294370 165538 6 vccd2.extra30
port 744 nsew power bidirectional
rlabel metal5 s -2408 147238 294370 147538 6 vccd2.extra31
port 745 nsew power bidirectional
rlabel metal5 s -2408 129238 294370 129538 6 vccd2.extra32
port 746 nsew power bidirectional
rlabel metal5 s -2408 111238 294370 111538 6 vccd2.extra33
port 747 nsew power bidirectional
rlabel metal5 s -2408 93238 294370 93538 6 vccd2.extra34
port 748 nsew power bidirectional
rlabel metal5 s -2408 75238 294370 75538 6 vccd2.extra35
port 749 nsew power bidirectional
rlabel metal5 s -2408 57238 294370 57538 6 vccd2.extra36
port 750 nsew power bidirectional
rlabel metal5 s -2408 39238 294370 39538 6 vccd2.extra37
port 751 nsew power bidirectional
rlabel metal5 s -2408 21238 294370 21538 6 vccd2.extra38
port 752 nsew power bidirectional
rlabel metal5 s -2408 3238 294370 3538 6 vccd2.extra39
port 753 nsew power bidirectional
rlabel metal5 s -1938 -1402 293900 -1102 8 vccd2.extra40
port 754 nsew power bidirectional
rlabel metal4 s 294070 -1872 294370 353840 6 vssd2
port 755 nsew ground bidirectional
rlabel metal4 s 281702 -1872 282002 353840 6 vssd2.extra1
port 756 nsew ground bidirectional
rlabel metal4 s 263702 -1872 264002 353840 6 vssd2.extra2
port 757 nsew ground bidirectional
rlabel metal4 s 245702 -1872 246002 353840 6 vssd2.extra3
port 758 nsew ground bidirectional
rlabel metal4 s 227702 -1872 228002 353840 6 vssd2.extra4
port 759 nsew ground bidirectional
rlabel metal4 s 209702 -1872 210002 353840 6 vssd2.extra5
port 760 nsew ground bidirectional
rlabel metal4 s 191702 -1872 192002 353840 6 vssd2.extra6
port 761 nsew ground bidirectional
rlabel metal4 s 173702 -1872 174002 353840 6 vssd2.extra7
port 762 nsew ground bidirectional
rlabel metal4 s 155702 -1872 156002 353840 6 vssd2.extra8
port 763 nsew ground bidirectional
rlabel metal4 s 137702 -1872 138002 353840 6 vssd2.extra9
port 764 nsew ground bidirectional
rlabel metal4 s 119702 -1872 120002 353840 6 vssd2.extra10
port 765 nsew ground bidirectional
rlabel metal4 s 101702 -1872 102002 353840 6 vssd2.extra11
port 766 nsew ground bidirectional
rlabel metal4 s 83702 -1872 84002 353840 6 vssd2.extra12
port 767 nsew ground bidirectional
rlabel metal4 s 65702 -1872 66002 353840 6 vssd2.extra13
port 768 nsew ground bidirectional
rlabel metal4 s 47702 -1872 48002 353840 6 vssd2.extra14
port 769 nsew ground bidirectional
rlabel metal4 s 29702 -1872 30002 353840 6 vssd2.extra15
port 770 nsew ground bidirectional
rlabel metal4 s 11702 -1872 12002 353840 6 vssd2.extra16
port 771 nsew ground bidirectional
rlabel metal4 s -2408 -1872 -2108 353840 4 vssd2.extra17
port 772 nsew ground bidirectional
rlabel metal5 s -2408 353540 294370 353840 6 vssd2.extra18
port 773 nsew ground bidirectional
rlabel metal5 s -2408 336238 294370 336538 6 vssd2.extra19
port 774 nsew ground bidirectional
rlabel metal5 s -2408 318238 294370 318538 6 vssd2.extra20
port 775 nsew ground bidirectional
rlabel metal5 s -2408 300238 294370 300538 6 vssd2.extra21
port 776 nsew ground bidirectional
rlabel metal5 s -2408 282238 294370 282538 6 vssd2.extra22
port 777 nsew ground bidirectional
rlabel metal5 s -2408 264238 294370 264538 6 vssd2.extra23
port 778 nsew ground bidirectional
rlabel metal5 s -2408 246238 294370 246538 6 vssd2.extra24
port 779 nsew ground bidirectional
rlabel metal5 s -2408 228238 294370 228538 6 vssd2.extra25
port 780 nsew ground bidirectional
rlabel metal5 s -2408 210238 294370 210538 6 vssd2.extra26
port 781 nsew ground bidirectional
rlabel metal5 s -2408 192238 294370 192538 6 vssd2.extra27
port 782 nsew ground bidirectional
rlabel metal5 s -2408 174238 294370 174538 6 vssd2.extra28
port 783 nsew ground bidirectional
rlabel metal5 s -2408 156238 294370 156538 6 vssd2.extra29
port 784 nsew ground bidirectional
rlabel metal5 s -2408 138238 294370 138538 6 vssd2.extra30
port 785 nsew ground bidirectional
rlabel metal5 s -2408 120238 294370 120538 6 vssd2.extra31
port 786 nsew ground bidirectional
rlabel metal5 s -2408 102238 294370 102538 6 vssd2.extra32
port 787 nsew ground bidirectional
rlabel metal5 s -2408 84238 294370 84538 6 vssd2.extra33
port 788 nsew ground bidirectional
rlabel metal5 s -2408 66238 294370 66538 6 vssd2.extra34
port 789 nsew ground bidirectional
rlabel metal5 s -2408 48238 294370 48538 6 vssd2.extra35
port 790 nsew ground bidirectional
rlabel metal5 s -2408 30238 294370 30538 6 vssd2.extra36
port 791 nsew ground bidirectional
rlabel metal5 s -2408 12238 294370 12538 6 vssd2.extra37
port 792 nsew ground bidirectional
rlabel metal5 s -2408 -1872 294370 -1572 8 vssd2.extra38
port 793 nsew ground bidirectional
rlabel metal4 s 274502 -2812 274802 354780 6 vdda1
port 794 nsew power bidirectional
rlabel metal4 s 256502 -2812 256802 354780 6 vdda1.extra1
port 795 nsew power bidirectional
rlabel metal4 s 238502 -2812 238802 354780 6 vdda1.extra2
port 796 nsew power bidirectional
rlabel metal4 s 220502 -2812 220802 354780 6 vdda1.extra3
port 797 nsew power bidirectional
rlabel metal4 s 202502 -2812 202802 354780 6 vdda1.extra4
port 798 nsew power bidirectional
rlabel metal4 s 184502 -2812 184802 354780 6 vdda1.extra5
port 799 nsew power bidirectional
rlabel metal4 s 166502 -2812 166802 354780 6 vdda1.extra6
port 800 nsew power bidirectional
rlabel metal4 s 148502 -2812 148802 354780 6 vdda1.extra7
port 801 nsew power bidirectional
rlabel metal4 s 130502 -2812 130802 354780 6 vdda1.extra8
port 802 nsew power bidirectional
rlabel metal4 s 112502 -2812 112802 354780 6 vdda1.extra9
port 803 nsew power bidirectional
rlabel metal4 s 94502 -2812 94802 354780 6 vdda1.extra10
port 804 nsew power bidirectional
rlabel metal4 s 76502 -2812 76802 354780 6 vdda1.extra11
port 805 nsew power bidirectional
rlabel metal4 s 58502 -2812 58802 354780 6 vdda1.extra12
port 806 nsew power bidirectional
rlabel metal4 s 40502 -2812 40802 354780 6 vdda1.extra13
port 807 nsew power bidirectional
rlabel metal4 s 22502 -2812 22802 354780 6 vdda1.extra14
port 808 nsew power bidirectional
rlabel metal4 s 4502 -2812 4802 354780 6 vdda1.extra15
port 809 nsew power bidirectional
rlabel metal4 s 294540 -2342 294840 354310 6 vdda1.extra16
port 810 nsew power bidirectional
rlabel metal4 s -2878 -2342 -2578 354310 4 vdda1.extra17
port 811 nsew power bidirectional
rlabel metal5 s -2878 354010 294840 354310 6 vdda1.extra18
port 812 nsew power bidirectional
rlabel metal5 s -3348 347038 295310 347338 6 vdda1.extra19
port 813 nsew power bidirectional
rlabel metal5 s -3348 329038 295310 329338 6 vdda1.extra20
port 814 nsew power bidirectional
rlabel metal5 s -3348 311038 295310 311338 6 vdda1.extra21
port 815 nsew power bidirectional
rlabel metal5 s -3348 293038 295310 293338 6 vdda1.extra22
port 816 nsew power bidirectional
rlabel metal5 s -3348 275038 295310 275338 6 vdda1.extra23
port 817 nsew power bidirectional
rlabel metal5 s -3348 257038 295310 257338 6 vdda1.extra24
port 818 nsew power bidirectional
rlabel metal5 s -3348 239038 295310 239338 6 vdda1.extra25
port 819 nsew power bidirectional
rlabel metal5 s -3348 221038 295310 221338 6 vdda1.extra26
port 820 nsew power bidirectional
rlabel metal5 s -3348 203038 295310 203338 6 vdda1.extra27
port 821 nsew power bidirectional
rlabel metal5 s -3348 185038 295310 185338 6 vdda1.extra28
port 822 nsew power bidirectional
rlabel metal5 s -3348 167038 295310 167338 6 vdda1.extra29
port 823 nsew power bidirectional
rlabel metal5 s -3348 149038 295310 149338 6 vdda1.extra30
port 824 nsew power bidirectional
rlabel metal5 s -3348 131038 295310 131338 6 vdda1.extra31
port 825 nsew power bidirectional
rlabel metal5 s -3348 113038 295310 113338 6 vdda1.extra32
port 826 nsew power bidirectional
rlabel metal5 s -3348 95038 295310 95338 6 vdda1.extra33
port 827 nsew power bidirectional
rlabel metal5 s -3348 77038 295310 77338 6 vdda1.extra34
port 828 nsew power bidirectional
rlabel metal5 s -3348 59038 295310 59338 6 vdda1.extra35
port 829 nsew power bidirectional
rlabel metal5 s -3348 41038 295310 41338 6 vdda1.extra36
port 830 nsew power bidirectional
rlabel metal5 s -3348 23038 295310 23338 6 vdda1.extra37
port 831 nsew power bidirectional
rlabel metal5 s -3348 5038 295310 5338 6 vdda1.extra38
port 832 nsew power bidirectional
rlabel metal5 s -2878 -2342 294840 -2042 8 vdda1.extra39
port 833 nsew power bidirectional
rlabel metal4 s 295010 -2812 295310 354780 6 vssa1
port 834 nsew ground bidirectional
rlabel metal4 s 283502 -2812 283802 354780 6 vssa1.extra1
port 835 nsew ground bidirectional
rlabel metal4 s 265502 -2812 265802 354780 6 vssa1.extra2
port 836 nsew ground bidirectional
rlabel metal4 s 247502 -2812 247802 354780 6 vssa1.extra3
port 837 nsew ground bidirectional
rlabel metal4 s 229502 -2812 229802 354780 6 vssa1.extra4
port 838 nsew ground bidirectional
rlabel metal4 s 211502 -2812 211802 354780 6 vssa1.extra5
port 839 nsew ground bidirectional
rlabel metal4 s 193502 -2812 193802 354780 6 vssa1.extra6
port 840 nsew ground bidirectional
rlabel metal4 s 175502 -2812 175802 354780 6 vssa1.extra7
port 841 nsew ground bidirectional
rlabel metal4 s 157502 -2812 157802 354780 6 vssa1.extra8
port 842 nsew ground bidirectional
rlabel metal4 s 139502 -2812 139802 354780 6 vssa1.extra9
port 843 nsew ground bidirectional
rlabel metal4 s 121502 -2812 121802 354780 6 vssa1.extra10
port 844 nsew ground bidirectional
rlabel metal4 s 103502 -2812 103802 354780 6 vssa1.extra11
port 845 nsew ground bidirectional
rlabel metal4 s 85502 -2812 85802 354780 6 vssa1.extra12
port 846 nsew ground bidirectional
rlabel metal4 s 67502 -2812 67802 354780 6 vssa1.extra13
port 847 nsew ground bidirectional
rlabel metal4 s 49502 -2812 49802 354780 6 vssa1.extra14
port 848 nsew ground bidirectional
rlabel metal4 s 31502 -2812 31802 354780 6 vssa1.extra15
port 849 nsew ground bidirectional
rlabel metal4 s 13502 -2812 13802 354780 6 vssa1.extra16
port 850 nsew ground bidirectional
rlabel metal4 s -3348 -2812 -3048 354780 4 vssa1.extra17
port 851 nsew ground bidirectional
rlabel metal5 s -3348 354480 295310 354780 6 vssa1.extra18
port 852 nsew ground bidirectional
rlabel metal5 s -3348 338038 295310 338338 6 vssa1.extra19
port 853 nsew ground bidirectional
rlabel metal5 s -3348 320038 295310 320338 6 vssa1.extra20
port 854 nsew ground bidirectional
rlabel metal5 s -3348 302038 295310 302338 6 vssa1.extra21
port 855 nsew ground bidirectional
rlabel metal5 s -3348 284038 295310 284338 6 vssa1.extra22
port 856 nsew ground bidirectional
rlabel metal5 s -3348 266038 295310 266338 6 vssa1.extra23
port 857 nsew ground bidirectional
rlabel metal5 s -3348 248038 295310 248338 6 vssa1.extra24
port 858 nsew ground bidirectional
rlabel metal5 s -3348 230038 295310 230338 6 vssa1.extra25
port 859 nsew ground bidirectional
rlabel metal5 s -3348 212038 295310 212338 6 vssa1.extra26
port 860 nsew ground bidirectional
rlabel metal5 s -3348 194038 295310 194338 6 vssa1.extra27
port 861 nsew ground bidirectional
rlabel metal5 s -3348 176038 295310 176338 6 vssa1.extra28
port 862 nsew ground bidirectional
rlabel metal5 s -3348 158038 295310 158338 6 vssa1.extra29
port 863 nsew ground bidirectional
rlabel metal5 s -3348 140038 295310 140338 6 vssa1.extra30
port 864 nsew ground bidirectional
rlabel metal5 s -3348 122038 295310 122338 6 vssa1.extra31
port 865 nsew ground bidirectional
rlabel metal5 s -3348 104038 295310 104338 6 vssa1.extra32
port 866 nsew ground bidirectional
rlabel metal5 s -3348 86038 295310 86338 6 vssa1.extra33
port 867 nsew ground bidirectional
rlabel metal5 s -3348 68038 295310 68338 6 vssa1.extra34
port 868 nsew ground bidirectional
rlabel metal5 s -3348 50038 295310 50338 6 vssa1.extra35
port 869 nsew ground bidirectional
rlabel metal5 s -3348 32038 295310 32338 6 vssa1.extra36
port 870 nsew ground bidirectional
rlabel metal5 s -3348 14038 295310 14338 6 vssa1.extra37
port 871 nsew ground bidirectional
rlabel metal5 s -3348 -2812 295310 -2512 8 vssa1.extra38
port 872 nsew ground bidirectional
rlabel metal4 s 276302 -3752 276602 355720 6 vdda2
port 873 nsew power bidirectional
rlabel metal4 s 258302 -3752 258602 355720 6 vdda2.extra1
port 874 nsew power bidirectional
rlabel metal4 s 240302 -3752 240602 355720 6 vdda2.extra2
port 875 nsew power bidirectional
rlabel metal4 s 222302 -3752 222602 355720 6 vdda2.extra3
port 876 nsew power bidirectional
rlabel metal4 s 204302 -3752 204602 355720 6 vdda2.extra4
port 877 nsew power bidirectional
rlabel metal4 s 186302 -3752 186602 355720 6 vdda2.extra5
port 878 nsew power bidirectional
rlabel metal4 s 168302 -3752 168602 355720 6 vdda2.extra6
port 879 nsew power bidirectional
rlabel metal4 s 150302 -3752 150602 355720 6 vdda2.extra7
port 880 nsew power bidirectional
rlabel metal4 s 132302 -3752 132602 355720 6 vdda2.extra8
port 881 nsew power bidirectional
rlabel metal4 s 114302 -3752 114602 355720 6 vdda2.extra9
port 882 nsew power bidirectional
rlabel metal4 s 96302 -3752 96602 355720 6 vdda2.extra10
port 883 nsew power bidirectional
rlabel metal4 s 78302 -3752 78602 355720 6 vdda2.extra11
port 884 nsew power bidirectional
rlabel metal4 s 60302 -3752 60602 355720 6 vdda2.extra12
port 885 nsew power bidirectional
rlabel metal4 s 42302 -3752 42602 355720 6 vdda2.extra13
port 886 nsew power bidirectional
rlabel metal4 s 24302 -3752 24602 355720 6 vdda2.extra14
port 887 nsew power bidirectional
rlabel metal4 s 6302 -3752 6602 355720 6 vdda2.extra15
port 888 nsew power bidirectional
rlabel metal4 s 295480 -3282 295780 355250 6 vdda2.extra16
port 889 nsew power bidirectional
rlabel metal4 s -3818 -3282 -3518 355250 4 vdda2.extra17
port 890 nsew power bidirectional
rlabel metal5 s -3818 354950 295780 355250 6 vdda2.extra18
port 891 nsew power bidirectional
rlabel metal5 s -4288 348838 296250 349138 6 vdda2.extra19
port 892 nsew power bidirectional
rlabel metal5 s -4288 330838 296250 331138 6 vdda2.extra20
port 893 nsew power bidirectional
rlabel metal5 s -4288 312838 296250 313138 6 vdda2.extra21
port 894 nsew power bidirectional
rlabel metal5 s -4288 294838 296250 295138 6 vdda2.extra22
port 895 nsew power bidirectional
rlabel metal5 s -4288 276838 296250 277138 6 vdda2.extra23
port 896 nsew power bidirectional
rlabel metal5 s -4288 258838 296250 259138 6 vdda2.extra24
port 897 nsew power bidirectional
rlabel metal5 s -4288 240838 296250 241138 6 vdda2.extra25
port 898 nsew power bidirectional
rlabel metal5 s -4288 222838 296250 223138 6 vdda2.extra26
port 899 nsew power bidirectional
rlabel metal5 s -4288 204838 296250 205138 6 vdda2.extra27
port 900 nsew power bidirectional
rlabel metal5 s -4288 186838 296250 187138 6 vdda2.extra28
port 901 nsew power bidirectional
rlabel metal5 s -4288 168838 296250 169138 6 vdda2.extra29
port 902 nsew power bidirectional
rlabel metal5 s -4288 150838 296250 151138 6 vdda2.extra30
port 903 nsew power bidirectional
rlabel metal5 s -4288 132838 296250 133138 6 vdda2.extra31
port 904 nsew power bidirectional
rlabel metal5 s -4288 114838 296250 115138 6 vdda2.extra32
port 905 nsew power bidirectional
rlabel metal5 s -4288 96838 296250 97138 6 vdda2.extra33
port 906 nsew power bidirectional
rlabel metal5 s -4288 78838 296250 79138 6 vdda2.extra34
port 907 nsew power bidirectional
rlabel metal5 s -4288 60838 296250 61138 6 vdda2.extra35
port 908 nsew power bidirectional
rlabel metal5 s -4288 42838 296250 43138 6 vdda2.extra36
port 909 nsew power bidirectional
rlabel metal5 s -4288 24838 296250 25138 6 vdda2.extra37
port 910 nsew power bidirectional
rlabel metal5 s -4288 6838 296250 7138 6 vdda2.extra38
port 911 nsew power bidirectional
rlabel metal5 s -3818 -3282 295780 -2982 8 vdda2.extra39
port 912 nsew power bidirectional
rlabel metal4 s 295950 -3752 296250 355720 6 vssa2
port 913 nsew ground bidirectional
rlabel metal4 s 285302 -3752 285602 355720 6 vssa2.extra1
port 914 nsew ground bidirectional
rlabel metal4 s 267302 -3752 267602 355720 6 vssa2.extra2
port 915 nsew ground bidirectional
rlabel metal4 s 249302 -3752 249602 355720 6 vssa2.extra3
port 916 nsew ground bidirectional
rlabel metal4 s 231302 -3752 231602 355720 6 vssa2.extra4
port 917 nsew ground bidirectional
rlabel metal4 s 213302 -3752 213602 355720 6 vssa2.extra5
port 918 nsew ground bidirectional
rlabel metal4 s 195302 -3752 195602 355720 6 vssa2.extra6
port 919 nsew ground bidirectional
rlabel metal4 s 177302 -3752 177602 355720 6 vssa2.extra7
port 920 nsew ground bidirectional
rlabel metal4 s 159302 -3752 159602 355720 6 vssa2.extra8
port 921 nsew ground bidirectional
rlabel metal4 s 141302 -3752 141602 355720 6 vssa2.extra9
port 922 nsew ground bidirectional
rlabel metal4 s 123302 -3752 123602 355720 6 vssa2.extra10
port 923 nsew ground bidirectional
rlabel metal4 s 105302 -3752 105602 355720 6 vssa2.extra11
port 924 nsew ground bidirectional
rlabel metal4 s 87302 -3752 87602 355720 6 vssa2.extra12
port 925 nsew ground bidirectional
rlabel metal4 s 69302 -3752 69602 355720 6 vssa2.extra13
port 926 nsew ground bidirectional
rlabel metal4 s 51302 -3752 51602 355720 6 vssa2.extra14
port 927 nsew ground bidirectional
rlabel metal4 s 33302 -3752 33602 355720 6 vssa2.extra15
port 928 nsew ground bidirectional
rlabel metal4 s 15302 -3752 15602 355720 6 vssa2.extra16
port 929 nsew ground bidirectional
rlabel metal4 s -4288 -3752 -3988 355720 4 vssa2.extra17
port 930 nsew ground bidirectional
rlabel metal5 s -4288 355420 296250 355720 6 vssa2.extra18
port 931 nsew ground bidirectional
rlabel metal5 s -4288 339838 296250 340138 6 vssa2.extra19
port 932 nsew ground bidirectional
rlabel metal5 s -4288 321838 296250 322138 6 vssa2.extra20
port 933 nsew ground bidirectional
rlabel metal5 s -4288 303838 296250 304138 6 vssa2.extra21
port 934 nsew ground bidirectional
rlabel metal5 s -4288 285838 296250 286138 6 vssa2.extra22
port 935 nsew ground bidirectional
rlabel metal5 s -4288 267838 296250 268138 6 vssa2.extra23
port 936 nsew ground bidirectional
rlabel metal5 s -4288 249838 296250 250138 6 vssa2.extra24
port 937 nsew ground bidirectional
rlabel metal5 s -4288 231838 296250 232138 6 vssa2.extra25
port 938 nsew ground bidirectional
rlabel metal5 s -4288 213838 296250 214138 6 vssa2.extra26
port 939 nsew ground bidirectional
rlabel metal5 s -4288 195838 296250 196138 6 vssa2.extra27
port 940 nsew ground bidirectional
rlabel metal5 s -4288 177838 296250 178138 6 vssa2.extra28
port 941 nsew ground bidirectional
rlabel metal5 s -4288 159838 296250 160138 6 vssa2.extra29
port 942 nsew ground bidirectional
rlabel metal5 s -4288 141838 296250 142138 6 vssa2.extra30
port 943 nsew ground bidirectional
rlabel metal5 s -4288 123838 296250 124138 6 vssa2.extra31
port 944 nsew ground bidirectional
rlabel metal5 s -4288 105838 296250 106138 6 vssa2.extra32
port 945 nsew ground bidirectional
rlabel metal5 s -4288 87838 296250 88138 6 vssa2.extra33
port 946 nsew ground bidirectional
rlabel metal5 s -4288 69838 296250 70138 6 vssa2.extra34
port 947 nsew ground bidirectional
rlabel metal5 s -4288 51838 296250 52138 6 vssa2.extra35
port 948 nsew ground bidirectional
rlabel metal5 s -4288 33838 296250 34138 6 vssa2.extra36
port 949 nsew ground bidirectional
rlabel metal5 s -4288 15838 296250 16138 6 vssa2.extra37
port 950 nsew ground bidirectional
rlabel metal5 s -4288 -3752 296250 -3452 8 vssa2.extra38
port 951 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 292000 352000
<< end >>
