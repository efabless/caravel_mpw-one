DFFRAM.cdl