magic
tech sky130A
magscale 1 2
timestamp 1611263055
<< obsli1 >>
rect 920 2159 10367 11441
<< obsm1 >>
rect 920 1164 26574 12504
<< obsm2 >>
rect 1216 167 26570 13705
<< metal3 >>
rect 14000 13608 34000 13728
rect 14000 13064 34000 13184
rect 14000 12520 34000 12640
rect 14000 11976 34000 12096
rect 14000 11432 34000 11552
rect 14000 10888 34000 11008
rect 14000 10344 34000 10464
rect 14000 9800 34000 9920
rect 14000 9256 34000 9376
rect 14000 8712 34000 8832
rect 14000 8168 34000 8288
rect 14000 7624 34000 7744
rect 14000 7080 34000 7200
rect 14000 6536 34000 6656
rect 14000 5992 34000 6112
rect 14000 5448 34000 5568
rect 14000 4904 34000 5024
rect 14000 4360 34000 4480
rect 14000 3816 34000 3936
rect 14000 3272 34000 3392
rect 14000 2728 34000 2848
rect 14000 2184 34000 2304
rect 14000 1640 34000 1760
rect 14000 1096 34000 1216
rect 14000 552 34000 672
rect 14000 144 34000 264
<< obsm3 >>
rect 2060 2143 5380 11457
<< metal4 >>
rect -1620 -364 -1300 13964
rect -960 296 -640 13304
rect -300 956 20 12644
rect 360 1616 680 11984
rect 2060 956 2380 12644
rect 2960 -364 3280 13964
rect 3560 956 3880 12644
rect 4460 -364 4780 13964
rect 5060 956 5380 12644
rect 5960 -364 6280 13964
rect 7324 1616 7644 11984
rect 7984 956 8304 12644
rect 8644 296 8964 13304
rect 9304 -364 9624 13964
<< metal5 >>
rect -1620 13644 9624 13964
rect -960 12984 8964 13304
rect -300 12324 8304 12644
rect 360 11664 7644 11984
rect -300 10116 8304 10436
rect -1620 9416 9624 9736
rect -300 8516 8304 8836
rect -1620 7816 9624 8136
rect -300 6916 8304 7236
rect -1620 6216 9624 6536
rect -300 5316 8304 5636
rect -1620 4616 9624 4936
rect -300 3716 8304 4036
rect 360 1616 7644 1936
rect -300 956 8304 1276
rect -960 296 8964 616
rect -1620 -364 9624 -44
<< labels >>
rlabel metal3 s 14000 1096 34000 1216 6 mgmt_gpio_in
port 1 nsew signal output
rlabel metal3 s 14000 1640 34000 1760 6 mgmt_gpio_oeb
port 2 nsew signal input
rlabel metal3 s 14000 2184 34000 2304 6 mgmt_gpio_out
port 3 nsew signal input
rlabel metal3 s 14000 552 34000 672 6 one
port 4 nsew signal output
rlabel metal3 s 14000 2728 34000 2848 6 pad_gpio_ana_en
port 5 nsew signal output
rlabel metal3 s 14000 3272 34000 3392 6 pad_gpio_ana_pol
port 6 nsew signal output
rlabel metal3 s 14000 3816 34000 3936 6 pad_gpio_ana_sel
port 7 nsew signal output
rlabel metal3 s 14000 4360 34000 4480 6 pad_gpio_dm[0]
port 8 nsew signal output
rlabel metal3 s 14000 4904 34000 5024 6 pad_gpio_dm[1]
port 9 nsew signal output
rlabel metal3 s 14000 5448 34000 5568 6 pad_gpio_dm[2]
port 10 nsew signal output
rlabel metal3 s 14000 5992 34000 6112 6 pad_gpio_holdover
port 11 nsew signal output
rlabel metal3 s 14000 6536 34000 6656 6 pad_gpio_ib_mode_sel
port 12 nsew signal output
rlabel metal3 s 14000 7080 34000 7200 6 pad_gpio_in
port 13 nsew signal input
rlabel metal3 s 14000 7624 34000 7744 6 pad_gpio_inenb
port 14 nsew signal output
rlabel metal3 s 14000 8168 34000 8288 6 pad_gpio_out
port 15 nsew signal output
rlabel metal3 s 14000 8712 34000 8832 6 pad_gpio_outenb
port 16 nsew signal output
rlabel metal3 s 14000 9256 34000 9376 6 pad_gpio_slow_sel
port 17 nsew signal output
rlabel metal3 s 14000 9800 34000 9920 6 pad_gpio_vtrip_sel
port 18 nsew signal output
rlabel metal3 s 14000 10344 34000 10464 6 resetn
port 19 nsew signal input
rlabel metal3 s 14000 10888 34000 11008 6 serial_clock
port 20 nsew signal input
rlabel metal3 s 14000 11432 34000 11552 6 serial_data_in
port 21 nsew signal input
rlabel metal3 s 14000 11976 34000 12096 6 serial_data_out
port 22 nsew signal output
rlabel metal3 s 14000 12520 34000 12640 6 user_gpio_in
port 23 nsew signal output
rlabel metal3 s 14000 13064 34000 13184 6 user_gpio_oeb
port 24 nsew signal input
rlabel metal3 s 14000 13608 34000 13728 6 user_gpio_out
port 25 nsew signal input
rlabel metal3 s 14000 144 34000 264 6 zero
port 26 nsew signal output
rlabel metal4 s 5060 956 5380 12644 6 vccd
port 27 nsew power bidirectional
rlabel metal4 s 2060 956 2380 12644 6 vccd
port 28 nsew power bidirectional
rlabel metal4 s 7324 1616 7644 11984 6 vccd
port 29 nsew power bidirectional
rlabel metal4 s 360 1616 680 11984 6 vccd
port 30 nsew power bidirectional
rlabel metal5 s 360 11664 7644 11984 6 vccd
port 31 nsew power bidirectional
rlabel metal5 s -300 10116 8304 10436 6 vccd
port 32 nsew power bidirectional
rlabel metal5 s -300 6916 8304 7236 6 vccd
port 33 nsew power bidirectional
rlabel metal5 s -300 3716 8304 4036 6 vccd
port 34 nsew power bidirectional
rlabel metal5 s 360 1616 7644 1936 6 vccd
port 35 nsew power bidirectional
rlabel metal4 s 7984 956 8304 12644 6 vssd
port 36 nsew ground bidirectional
rlabel metal4 s 3560 956 3880 12644 6 vssd
port 37 nsew ground bidirectional
rlabel metal4 s -300 956 20 12644 4 vssd
port 38 nsew ground bidirectional
rlabel metal5 s -300 12324 8304 12644 6 vssd
port 39 nsew ground bidirectional
rlabel metal5 s -300 8516 8304 8836 6 vssd
port 40 nsew ground bidirectional
rlabel metal5 s -300 5316 8304 5636 6 vssd
port 41 nsew ground bidirectional
rlabel metal5 s -300 956 8304 1276 6 vssd
port 42 nsew ground bidirectional
rlabel metal4 s 5960 -364 6280 13964 6 vccd1
port 43 nsew power bidirectional
rlabel metal4 s 2960 -364 3280 13964 6 vccd1
port 44 nsew power bidirectional
rlabel metal4 s 8644 296 8964 13304 6 vccd1
port 45 nsew power bidirectional
rlabel metal4 s -960 296 -640 13304 4 vccd1
port 46 nsew power bidirectional
rlabel metal5 s -960 12984 8964 13304 6 vccd1
port 47 nsew power bidirectional
rlabel metal5 s -1620 7816 9624 8136 6 vccd1
port 48 nsew power bidirectional
rlabel metal5 s -1620 4616 9624 4936 6 vccd1
port 49 nsew power bidirectional
rlabel metal5 s -960 296 8964 616 6 vccd1
port 50 nsew power bidirectional
rlabel metal4 s 9304 -364 9624 13964 6 vssd1
port 51 nsew ground bidirectional
rlabel metal4 s 4460 -364 4780 13964 6 vssd1
port 52 nsew ground bidirectional
rlabel metal4 s -1620 -364 -1300 13964 4 vssd1
port 53 nsew ground bidirectional
rlabel metal5 s -1620 13644 9624 13964 6 vssd1
port 54 nsew ground bidirectional
rlabel metal5 s -1620 9416 9624 9736 6 vssd1
port 55 nsew ground bidirectional
rlabel metal5 s -1620 6216 9624 6536 6 vssd1
port 56 nsew ground bidirectional
rlabel metal5 s -1620 -364 9624 -44 8 vssd1
port 57 nsew ground bidirectional
<< properties >>
string LEFclass BLOCK
string FIXED_BBOX 0 0 34000 14000
string LEFview TRUE
string GDS_FILE ../gds/gpio_control_block.gds
string GDS_END 348020
string GDS_START 146164
<< end >>

