magic
tech sky130A
magscale 1 2
timestamp 1606424343
<< metal3 >>
rect -5178 3222 -1806 3250
rect -5178 78 -1890 3222
rect -1826 78 -1806 3222
rect -5178 50 -1806 78
rect -1686 3222 1686 3250
rect -1686 78 1602 3222
rect 1666 78 1686 3222
rect -1686 50 1686 78
rect 1806 3222 5178 3250
rect 1806 78 5094 3222
rect 5158 78 5178 3222
rect 1806 50 5178 78
rect -5178 -78 -1806 -50
rect -5178 -3222 -1890 -78
rect -1826 -3222 -1806 -78
rect -5178 -3250 -1806 -3222
rect -1686 -78 1686 -50
rect -1686 -3222 1602 -78
rect 1666 -3222 1686 -78
rect -1686 -3250 1686 -3222
rect 1806 -78 5178 -50
rect 1806 -3222 5094 -78
rect 5158 -3222 5178 -78
rect 1806 -3250 5178 -3222
<< via3 >>
rect -1890 78 -1826 3222
rect 1602 78 1666 3222
rect 5094 78 5158 3222
rect -1890 -3222 -1826 -78
rect 1602 -3222 1666 -78
rect 5094 -3222 5158 -78
<< mimcap >>
rect -5078 3110 -2078 3150
rect -5078 190 -5038 3110
rect -2118 190 -2078 3110
rect -5078 150 -2078 190
rect -1586 3110 1414 3150
rect -1586 190 -1546 3110
rect 1374 190 1414 3110
rect -1586 150 1414 190
rect 1906 3110 4906 3150
rect 1906 190 1946 3110
rect 4866 190 4906 3110
rect 1906 150 4906 190
rect -5078 -190 -2078 -150
rect -5078 -3110 -5038 -190
rect -2118 -3110 -2078 -190
rect -5078 -3150 -2078 -3110
rect -1586 -190 1414 -150
rect -1586 -3110 -1546 -190
rect 1374 -3110 1414 -190
rect -1586 -3150 1414 -3110
rect 1906 -190 4906 -150
rect 1906 -3110 1946 -190
rect 4866 -3110 4906 -190
rect 1906 -3150 4906 -3110
<< mimcapcontact >>
rect -5038 190 -2118 3110
rect -1546 190 1374 3110
rect 1946 190 4866 3110
rect -5038 -3110 -2118 -190
rect -1546 -3110 1374 -190
rect 1946 -3110 4866 -190
<< metal4 >>
rect -3630 3111 -3526 3300
rect -1910 3222 -1806 3300
rect -5039 3110 -2117 3111
rect -5039 190 -5038 3110
rect -2118 190 -2117 3110
rect -5039 189 -2117 190
rect -3630 -189 -3526 189
rect -1910 78 -1890 3222
rect -1826 78 -1806 3222
rect -138 3111 -34 3300
rect 1582 3222 1686 3300
rect -1547 3110 1375 3111
rect -1547 190 -1546 3110
rect 1374 190 1375 3110
rect -1547 189 1375 190
rect -1910 -78 -1806 78
rect -5039 -190 -2117 -189
rect -5039 -3110 -5038 -190
rect -2118 -3110 -2117 -190
rect -5039 -3111 -2117 -3110
rect -3630 -3300 -3526 -3111
rect -1910 -3222 -1890 -78
rect -1826 -3222 -1806 -78
rect -138 -189 -34 189
rect 1582 78 1602 3222
rect 1666 78 1686 3222
rect 3354 3111 3458 3300
rect 5074 3222 5178 3300
rect 1945 3110 4867 3111
rect 1945 190 1946 3110
rect 4866 190 4867 3110
rect 1945 189 4867 190
rect 1582 -78 1686 78
rect -1547 -190 1375 -189
rect -1547 -3110 -1546 -190
rect 1374 -3110 1375 -190
rect -1547 -3111 1375 -3110
rect -1910 -3300 -1806 -3222
rect -138 -3300 -34 -3111
rect 1582 -3222 1602 -78
rect 1666 -3222 1686 -78
rect 3354 -189 3458 189
rect 5074 78 5094 3222
rect 5158 78 5178 3222
rect 5074 -78 5178 78
rect 1945 -190 4867 -189
rect 1945 -3110 1946 -190
rect 4866 -3110 4867 -190
rect 1945 -3111 4867 -3110
rect 1582 -3300 1686 -3222
rect 3354 -3300 3458 -3111
rect 5074 -3222 5094 -78
rect 5158 -3222 5178 -78
rect 5074 -3300 5178 -3222
<< properties >>
string gencell sky130_fd_pr__cap_mim_m3_1
string FIXED_BBOX 1806 50 5006 3250
string parameters w 15.0 l 15.0 val 235.2 carea 1.00 cperi 0.17 nx 3 ny 2 dummy 0 square 1 lmin 2.00 wmin 2.00 lmax 30.0 wmax 30.0 dc 0 bconnect 1 tconnect 1
string library sky130
<< end >>
