* SPICE NETLIST
***************************************

.SUBCKT MN g s d b
.ENDS
***************************************
.SUBCKT MP g s d b
.ENDS
***************************************
.SUBCKT condiode pin0 pin1
.ENDS
***************************************
.SUBCKT condiodeHvPsub pin0 pin1
.ENDS
***************************************
.SUBCKT nvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20nativevhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT n20vhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT n20nativevhviso1 pin0 pin1 pin2 pin3 pin4
.ENDS
***************************************
.SUBCKT pvhv pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT p20vhv1 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcnwvc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcnwvc2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xchvnwc pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT Dpar d0 d1
.ENDS
***************************************
.SUBCKT xcmvpp pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_nhvnative10x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp2_phv5x4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap2_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_wafflecap1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l40 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l20 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l10 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_atlas_fingercap_l5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1_met5pullin pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_5x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_4x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_3x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_2x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp_hd5_1x1 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvppx4_2xnhvnative10x4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym50p4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_lim5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_lim4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp6p8x6p1_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_polym4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m4shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3_lishield pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp8p6x7p9_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp1p8x1p8_m3shield c0 c1 b term4
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4m5shield pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp11p5x11p7_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4p4x4p6_m1m2 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp5 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp4 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT xcmvpp3 pin0 pin1 pin2
.ENDS
***************************************
.SUBCKT balun pin0 pin1 pin2 pin3 pin4 pin5
.ENDS
***************************************
.SUBCKT ind4 pin0 pin1 pin2 pin3
.ENDS
***************************************
.SUBCKT xhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p35 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_0p69 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_1p41 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_2p85 POS NEG SUB
.ENDS
***************************************
.SUBCKT xhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT xuhrpoly_5p73 POS NEG SUB
.ENDS
***************************************
.SUBCKT Probe probe conductor
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808671
** N=117 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808672
** N=175 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808673
** N=26 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808663
** N=118 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_2 2 3 4
** N=27 EP=3 IP=48 FDC=22
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
M18 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=41400 $Y=0 $D=49
M19 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=43410 $Y=0 $D=49
M20 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=46000 $Y=0 $D=49
M21 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=48010 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_3 2 3 4
** N=26 EP=3 IP=48 FDC=22
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
M18 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=41400 $Y=0 $D=49
M19 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=43410 $Y=0 $D=49
M20 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=46000 $Y=0 $D=49
M21 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=48010 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_pr__nfet_01v8__example_55959141808670
** N=21 EP=0 IP=10 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_4 2 3 4
** N=22 EP=3 IP=39 FDC=18
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_5 2 3 4
** N=23 EP=3 IP=39 FDC=18
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_6 2 3 4
** N=22 EP=3 IP=39 FDC=18
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_7 2 3 4
** N=30 EP=3 IP=48 FDC=22
*.SEEDPROM
M0 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250001 sb=250020 a=10 p=41 mult=1 $X=0 $Y=0 $D=49
M1 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250003 sb=250020 a=10 p=41 mult=1 $X=2010 $Y=0 $D=49
M2 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250006 sb=250020 a=10 p=41 mult=1 $X=4600 $Y=0 $D=49
M3 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250008 sb=250020 a=10 p=41 mult=1 $X=6610 $Y=0 $D=49
M4 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250010 sb=250020 a=10 p=41 mult=1 $X=9200 $Y=0 $D=49
M5 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250012 sb=250020 a=10 p=41 mult=1 $X=11210 $Y=0 $D=49
M6 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250015 sb=250020 a=10 p=41 mult=1 $X=13800 $Y=0 $D=49
M7 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250017 sb=250020 a=10 p=41 mult=1 $X=15810 $Y=0 $D=49
M8 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=18400 $Y=0 $D=49
M9 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=20410 $Y=0 $D=49
M10 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=23000 $Y=0 $D=49
M11 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=25010 $Y=0 $D=49
M12 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=27600 $Y=0 $D=49
M13 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250020 a=10 p=41 mult=1 $X=29610 $Y=0 $D=49
M14 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250017 a=10 p=41 mult=1 $X=32200 $Y=0 $D=49
M15 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250015 a=10 p=41 mult=1 $X=34210 $Y=0 $D=49
M16 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250012 a=10 p=41 mult=1 $X=36800 $Y=0 $D=49
M17 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250010 a=10 p=41 mult=1 $X=38810 $Y=0 $D=49
M18 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250008 a=10 p=41 mult=1 $X=41400 $Y=0 $D=49
M19 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250006 a=10 p=41 mult=1 $X=43410 $Y=0 $D=49
M20 4 3 2 2 nhv L=0.5 W=20 AD=15.1 AS=13.9 PD=21.51 PS=41.39 NRD=2.5308 NRS=2.2458 m=1 r=40 sa=250020 sb=250003 a=10 p=41 mult=1 $X=46000 $Y=0 $D=49
M21 2 3 4 2 nhv L=0.5 W=20 AD=13.9 AS=15.1 PD=41.39 PS=21.51 NRD=2.2458 NRS=2.5308 m=1 r=40 sa=250020 sb=250001 a=10 p=41 mult=1 $X=48010 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT ICV_8
** N=486 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_9
** N=280 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_10
** N=513 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_11
** N=316 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_12
** N=244 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_13
** N=273 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_14
** N=198 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s2__example_55959141808676
** N=88 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdftpl1s__example_55959141808675
** N=59 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1__example_55959141808662
** N=58 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_15
** N=567 EP=0 IP=4 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_16
** N=398 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_17
** N=259 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__hvdfl1sd__example_5595914180851
** N=15 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 1 2
** N=7 EP=2 IP=2 FDC=1
M0 1 2 1 1 nhv L=4 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 r=1.25 sa=2e+06 sb=2e+06 a=20 p=18 mult=1 $X=0 $Y=0 $D=49
.ENDS
***************************************
.SUBCKT sky130_fd_io__sio_clamp_pcap_4x5 1 2
** N=81 EP=2 IP=4 FDC=1
X0 1 2 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=1145 720 0 0 $X=700 $Y=540
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808679
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808678
** N=22 EP=0 IP=0 FDC=0
.ENDS
***************************************
.SUBCKT ICV_18 2 4
** N=702 EP=2 IP=88 FDC=1
*.SEEDPROM
X0 2 4 sky130_fd_io__sio_clamp_pcap_4x5 $T=25830 -68720 0 90 $X=19080 $Y=-68720
.ENDS
***************************************
.SUBCKT sky130_fd_io__esd_rcclamp_nfetcap 2 3
** N=122 EP=2 IP=2 FDC=1
*.SEEDPROM
M0 2 3 2 2 nhv L=8 W=5 AD=1.325 AS=1.325 PD=10.53 PS=10.53 NRD=0 NRS=0 m=1 r=0.625 sa=4e+06 sb=4e+06 a=40 p=26 mult=1 $X=895 $Y=630 $D=49
.ENDS
***************************************
.SUBCKT ICV_19 2 4
** N=308 EP=2 IP=282 FDC=3
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=7080 -68470 0 90 $X=420 $Y=-68720
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=13300 -68470 0 90 $X=6640 $Y=-68720
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=19520 -68470 0 90 $X=12860 $Y=-68720
.ENDS
***************************************
.SUBCKT ICV_20
** N=258 EP=0 IP=8 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_21
** N=1121 EP=0 IP=12 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_22 2 4
** N=308 EP=2 IP=282 FDC=3
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=7080 -58710 0 90 $X=420 $Y=-58960
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=13300 -58710 0 90 $X=6640 $Y=-58960
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=19520 -58710 0 90 $X=12860 $Y=-58960
.ENDS
***************************************
.SUBCKT ICV_23
** N=241 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_24
** N=1237 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_25 2 4
** N=305 EP=2 IP=282 FDC=3
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=7080 -48950 0 90 $X=420 $Y=-49200
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=13300 -48950 0 90 $X=6640 $Y=-49200
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=19520 -48950 0 90 $X=12860 $Y=-49200
.ENDS
***************************************
.SUBCKT ICV_26
** N=594 EP=0 IP=15 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_27
** N=981 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_28
** N=610 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_29
** N=2681 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_30 2 4
** N=588 EP=2 IP=564 FDC=6
*.SEEDPROM
X0 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=29430 7080 0 180 $X=19390 $Y=420
X1 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=29430 13300 0 180 $X=19390 $Y=6640
X2 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=29430 19520 0 180 $X=19390 $Y=12860
X3 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=39190 7080 0 180 $X=29150 $Y=420
X4 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=39190 13300 0 180 $X=29150 $Y=6640
X5 2 4 sky130_fd_io__esd_rcclamp_nfetcap $T=39190 19520 0 180 $X=29150 $Y=12860
.ENDS
***************************************
.SUBCKT ICV_31
** N=953 EP=0 IP=1 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_32
** N=502 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_33
** N=164 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_34
** N=221 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_35
** N=416 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_36
** N=1602 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_37
** N=1538 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd__example_55959141808336
** N=22 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT sky130_fd_pr__dfl1sd2__example_55959141808666
** N=23 EP=0 IP=0 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_38
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_39
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_40
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_41
** N=3 EP=0 IP=6 FDC=0
*.SEEDPROM
.ENDS
***************************************
.SUBCKT ICV_1 2 3 4
** N=257 EP=3 IP=16 FDC=50
*.SEEDPROM
M0 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=14 sa=250000 sb=250020 a=3.5 p=15 mult=1 $X=0 $Y=0 $D=109
M1 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250001 sb=250020 a=3.5 p=15 mult=1 $X=780 $Y=0 $D=109
M2 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250020 a=3.5 p=15 mult=1 $X=1560 $Y=0 $D=109
M3 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250020 a=3.5 p=15 mult=1 $X=2340 $Y=0 $D=109
M4 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250003 sb=250020 a=3.5 p=15 mult=1 $X=3120 $Y=0 $D=109
M5 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250004 sb=250020 a=3.5 p=15 mult=1 $X=3900 $Y=0 $D=109
M6 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250020 a=3.5 p=15 mult=1 $X=4680 $Y=0 $D=109
M7 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250020 a=3.5 p=15 mult=1 $X=5460 $Y=0 $D=109
M8 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250006 sb=250020 a=3.5 p=15 mult=1 $X=6240 $Y=0 $D=109
M9 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250007 sb=250020 a=3.5 p=15 mult=1 $X=7020 $Y=0 $D=109
M10 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250008 sb=250020 a=3.5 p=15 mult=1 $X=7800 $Y=0 $D=109
M11 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250020 a=3.5 p=15 mult=1 $X=8580 $Y=0 $D=109
M12 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250020 a=3.5 p=15 mult=1 $X=9360 $Y=0 $D=109
M13 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250010 sb=250020 a=3.5 p=15 mult=1 $X=10140 $Y=0 $D=109
M14 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250011 sb=250020 a=3.5 p=15 mult=1 $X=10920 $Y=0 $D=109
M15 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250012 sb=250020 a=3.5 p=15 mult=1 $X=11700 $Y=0 $D=109
M16 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250012 sb=250020 a=3.5 p=15 mult=1 $X=12480 $Y=0 $D=109
M17 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250013 sb=250020 a=3.5 p=15 mult=1 $X=13260 $Y=0 $D=109
M18 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250014 sb=250020 a=3.5 p=15 mult=1 $X=14040 $Y=0 $D=109
M19 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250015 sb=250020 a=3.5 p=15 mult=1 $X=14820 $Y=0 $D=109
M20 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250016 sb=250020 a=3.5 p=15 mult=1 $X=15600 $Y=0 $D=109
M21 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250016 sb=250020 a=3.5 p=15 mult=1 $X=16380 $Y=0 $D=109
M22 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250017 sb=250020 a=3.5 p=15 mult=1 $X=17160 $Y=0 $D=109
M23 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250018 sb=250020 a=3.5 p=15 mult=1 $X=17940 $Y=0 $D=109
M24 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250019 sb=250020 a=3.5 p=15 mult=1 $X=18720 $Y=0 $D=109
M25 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250019 a=3.5 p=15 mult=1 $X=19500 $Y=0 $D=109
M26 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250018 a=3.5 p=15 mult=1 $X=20280 $Y=0 $D=109
M27 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250017 a=3.5 p=15 mult=1 $X=21060 $Y=0 $D=109
M28 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250016 a=3.5 p=15 mult=1 $X=21840 $Y=0 $D=109
M29 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250016 a=3.5 p=15 mult=1 $X=22620 $Y=0 $D=109
M30 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250015 a=3.5 p=15 mult=1 $X=23400 $Y=0 $D=109
M31 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250014 a=3.5 p=15 mult=1 $X=24180 $Y=0 $D=109
M32 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250013 a=3.5 p=15 mult=1 $X=24960 $Y=0 $D=109
M33 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250012 a=3.5 p=15 mult=1 $X=25740 $Y=0 $D=109
M34 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250012 a=3.5 p=15 mult=1 $X=26520 $Y=0 $D=109
M35 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250011 a=3.5 p=15 mult=1 $X=27300 $Y=0 $D=109
M36 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250010 a=3.5 p=15 mult=1 $X=28080 $Y=0 $D=109
M37 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250009 a=3.5 p=15 mult=1 $X=28860 $Y=0 $D=109
M38 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250009 a=3.5 p=15 mult=1 $X=29640 $Y=0 $D=109
M39 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250008 a=3.5 p=15 mult=1 $X=30420 $Y=0 $D=109
M40 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250007 a=3.5 p=15 mult=1 $X=31200 $Y=0 $D=109
M41 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250006 a=3.5 p=15 mult=1 $X=31980 $Y=0 $D=109
M42 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250005 a=3.5 p=15 mult=1 $X=32760 $Y=0 $D=109
M43 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250005 a=3.5 p=15 mult=1 $X=33540 $Y=0 $D=109
M44 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250004 a=3.5 p=15 mult=1 $X=34320 $Y=0 $D=109
M45 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250003 a=3.5 p=15 mult=1 $X=35100 $Y=0 $D=109
M46 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250002 a=3.5 p=15 mult=1 $X=35880 $Y=0 $D=109
M47 2 3 4 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250002 a=3.5 p=15 mult=1 $X=36660 $Y=0 $D=109
M48 4 3 2 2 phv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250001 a=3.5 p=15 mult=1 $X=37440 $Y=0 $D=109
M49 2 3 4 2 phv L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250020 sb=250000 a=3.5 p=15 mult=1 $X=38220 $Y=0 $D=109
.ENDS
***************************************
.SUBCKT sky130_ef_io__vddio_hvc_clamped_pad VSSD VSSIO VDDIO VSSA AMUXBUS_B AMUXBUS_A VSSIO_Q VSWITCH VCCHIB VCCD VDDA
** N=1179 EP=11 IP=1295 FDC=241
M0 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250001 sb=250020 a=5 p=21 mult=1 $X=15885 $Y=183145 $D=49
M1 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250003 sb=250020 a=5 p=21 mult=1 $X=17895 $Y=183145 $D=49
M2 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250006 sb=250020 a=5 p=21 mult=1 $X=20485 $Y=183145 $D=49
M3 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250008 sb=250020 a=5 p=21 mult=1 $X=22495 $Y=183145 $D=49
M4 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250010 sb=250020 a=5 p=21 mult=1 $X=25085 $Y=183145 $D=49
M5 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250012 sb=250020 a=5 p=21 mult=1 $X=27095 $Y=183145 $D=49
M6 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250015 sb=250020 a=5 p=21 mult=1 $X=29685 $Y=183145 $D=49
M7 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250017 sb=250020 a=5 p=21 mult=1 $X=31695 $Y=183145 $D=49
M8 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=34285 $Y=183145 $D=49
M9 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=36295 $Y=183145 $D=49
M10 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=38885 $Y=183145 $D=49
M11 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=40895 $Y=183145 $D=49
M12 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=43485 $Y=183145 $D=49
M13 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250020 a=5 p=21 mult=1 $X=45495 $Y=183145 $D=49
M14 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250017 a=5 p=21 mult=1 $X=48085 $Y=183145 $D=49
M15 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250015 a=5 p=21 mult=1 $X=50095 $Y=183145 $D=49
M16 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250012 a=5 p=21 mult=1 $X=52685 $Y=183145 $D=49
M17 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250010 a=5 p=21 mult=1 $X=54695 $Y=183145 $D=49
M18 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=1.855 PD=7.28 PS=14.53 NRD=0 NRS=0 m=1 r=14 sa=250000 sb=250011 a=3.5 p=15 mult=1 $X=54915 $Y=30545 $D=49
M19 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250001 sb=250010 a=3.5 p=15 mult=1 $X=55695 $Y=30545 $D=49
M20 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250009 a=3.5 p=15 mult=1 $X=56475 $Y=30545 $D=49
M21 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250002 sb=250009 a=3.5 p=15 mult=1 $X=57255 $Y=30545 $D=49
M22 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250008 a=5 p=21 mult=1 $X=57285 $Y=183145 $D=49
M23 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250003 sb=250008 a=3.5 p=15 mult=1 $X=58035 $Y=30545 $D=49
M24 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250004 sb=250007 a=3.5 p=15 mult=1 $X=58815 $Y=30545 $D=49
M25 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250006 a=5 p=21 mult=1 $X=59295 $Y=183145 $D=49
M26 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250006 a=3.5 p=15 mult=1 $X=59595 $Y=30545 $D=49
M27 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250005 sb=250005 a=3.5 p=15 mult=1 $X=60375 $Y=30545 $D=49
M28 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250006 sb=250005 a=3.5 p=15 mult=1 $X=61155 $Y=30545 $D=49
M29 VDDIO 4 VSSIO VSSIO nhv L=0.5 W=10 AD=7.55 AS=6.95 PD=11.51 PS=21.39 NRD=5.073 NRS=4.503 m=1 r=20 sa=250020 sb=250003 a=5 p=21 mult=1 $X=61885 $Y=183145 $D=49
M30 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250007 sb=250004 a=3.5 p=15 mult=1 $X=61935 $Y=30545 $D=49
M31 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250008 sb=250003 a=3.5 p=15 mult=1 $X=62715 $Y=30545 $D=49
M32 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250002 a=3.5 p=15 mult=1 $X=63495 $Y=30545 $D=49
M33 VSSIO 4 VDDIO VSSIO nhv L=0.5 W=10 AD=6.95 AS=7.55 PD=21.39 PS=11.51 NRD=4.503 NRS=5.073 m=1 r=20 sa=250020 sb=250001 a=5 p=21 mult=1 $X=63895 $Y=183145 $D=49
M34 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250009 sb=250002 a=3.5 p=15 mult=1 $X=64275 $Y=30545 $D=49
M35 VSSIO 5 4 VSSIO nhv L=0.5 W=7 AD=0.98 AS=0.98 PD=7.28 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250010 sb=250001 a=3.5 p=15 mult=1 $X=65055 $Y=30545 $D=49
M36 4 5 VSSIO VSSIO nhv L=0.5 W=7 AD=1.855 AS=0.98 PD=14.53 PS=7.28 NRD=0 NRS=0 m=1 r=14 sa=250011 sb=250000 a=3.5 p=15 mult=1 $X=65835 $Y=30545 $D=49
X37 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=19700 $D=150
X38 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=51225 $Y=43275 $D=150
X39 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=64770 $Y=38800 $D=150
X40 VSSIO VDDIO condiode a=1e-06 p=0.004 m=1 ahftempperim=0.004 $X=68375 $Y=195640 $D=150
X41 VSSD VDDIO Dpar a=126.766 p=0 m=1 $[nwdiode] $X=8835 $Y=41140 $D=189
X42 VSSD VDDIO Dpar a=369.745 p=100.13 m=1 $[nwdiode] $X=5200 $Y=26890 $D=191
X43 VSSD VDDIO Dpar a=10358.7 p=619.08 m=1 $[dnwdiode_psub] $X=9500 $Y=131800 $D=193
X44 VSSIO VDDIO Dpar a=137.463 p=47.72 m=1 $[dnwdiode_pw] $X=53530 $Y=29360 $D=194
X45 VSSIO VDDIO Dpar a=8184.99 p=443.22 m=1 $[dnwdiode_pw] $X=10695 $Y=43000 $D=194
X46 VSSIO VDDIO Dpar a=1172.63 p=163 m=1 $[dnwdiode_pw] $X=13380 $Y=170 $D=194
R47 7 6 L=1550 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=1070 $Y=41405 $D=257
R48 7 VDDIO L=700 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=9500 $Y=72320 $D=257
R49 6 5 L=470 W=0.33 m=1 mult=1 model="mrp1" $[mrp1] $X=70725 $Y=39980 $D=257
R50 VDDIO VDDIO 0.01 m=1 $[short] $X=6670 $Y=103310 $D=286
X51 VSSIO 4 VDDIO ICV_2 $T=15885 160145 0 0 $X=14310 $Y=159965
X52 VSSIO 4 VDDIO ICV_3 $T=15885 137145 0 0 $X=14310 $Y=136965
X53 VSSIO 4 VDDIO ICV_4 $T=25085 114145 0 0 $X=23510 $Y=113965
X54 VSSIO 4 VDDIO ICV_5 $T=25085 91145 0 0 $X=23510 $Y=90965
X55 VSSIO 4 VDDIO ICV_6 $T=25085 68145 0 0 $X=23510 $Y=67965
X56 VSSIO 4 VDDIO ICV_7 $T=15885 45145 0 0 $X=14310 $Y=44965
X67 VSSIO 5 sky130_fd_pr__model__nfet_highvoltage__example_55959141808664 $T=61815 25110 0 180 $X=57370 $Y=19930
X68 VSSIO 5 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 7170 0 180 $X=13630 $Y=420
X69 VSSIO 5 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 13390 0 180 $X=13630 $Y=6640
X70 VSSIO 5 sky130_fd_io__sio_clamp_pcap_4x5 $T=19920 19610 0 180 $X=13630 $Y=12860
X71 VSSIO 5 ICV_18 $T=0 0 0 90 $X=59000 $Y=19080
X72 VSSIO 5 ICV_19 $T=0 0 0 90 $X=58430 $Y=-2035
X75 VSSIO 5 ICV_22 $T=0 0 0 90 $X=48670 $Y=-2035
X78 VSSIO 5 ICV_25 $T=0 0 0 90 $X=38910 $Y=-2035
X83 VSSIO 5 ICV_30 $T=0 0 0 0 $X=16700 $Y=-2035
X91 VDDIO 5 4 ICV_1 $T=6340 27765 0 0 $X=5745 $Y=27435
*.CALIBRE WARNING SHORT Short circuit(s) detected by extraction in this cell. See extraction report for details.
.ENDS
***************************************
