magic
tech sky130A
magscale 1 2
timestamp 1608238675
<< metal1 >>
rect 452176 1008113 452182 1008165
rect 452234 1008153 452240 1008165
rect 472144 1008153 472150 1008165
rect 452234 1008125 472150 1008153
rect 452234 1008113 452240 1008125
rect 472144 1008113 472150 1008125
rect 472202 1008113 472208 1008165
rect 434992 1008039 434998 1008091
rect 435050 1008079 435056 1008091
rect 471568 1008079 471574 1008091
rect 435050 1008051 471574 1008079
rect 435050 1008039 435056 1008051
rect 471568 1008039 471574 1008051
rect 471626 1008039 471632 1008091
rect 434704 1007965 434710 1008017
rect 434762 1008005 434768 1008017
rect 452176 1008005 452182 1008017
rect 434762 1007977 452182 1008005
rect 434762 1007965 434768 1007977
rect 452176 1007965 452182 1007977
rect 452234 1007965 452240 1008017
rect 367216 1005449 367222 1005501
rect 367274 1005489 367280 1005501
rect 383632 1005489 383638 1005501
rect 367274 1005461 383638 1005489
rect 367274 1005449 367280 1005461
rect 383632 1005449 383638 1005461
rect 383690 1005449 383696 1005501
rect 434608 1005449 434614 1005501
rect 434666 1005489 434672 1005501
rect 471856 1005489 471862 1005501
rect 434666 1005461 471862 1005489
rect 434666 1005449 434672 1005461
rect 471856 1005449 471862 1005461
rect 471914 1005449 471920 1005501
rect 434896 1005301 434902 1005353
rect 434954 1005341 434960 1005353
rect 469360 1005341 469366 1005353
rect 434954 1005313 469366 1005341
rect 434954 1005301 434960 1005313
rect 469360 1005301 469366 1005313
rect 469418 1005301 469424 1005353
rect 164272 1005227 164278 1005279
rect 164330 1005267 164336 1005279
rect 172816 1005267 172822 1005279
rect 164330 1005239 172822 1005267
rect 164330 1005227 164336 1005239
rect 172816 1005227 172822 1005239
rect 172874 1005227 172880 1005279
rect 437488 1005227 437494 1005279
rect 437546 1005267 437552 1005279
rect 470128 1005267 470134 1005279
rect 437546 1005239 470134 1005267
rect 437546 1005227 437552 1005239
rect 470128 1005227 470134 1005239
rect 470186 1005227 470192 1005279
rect 218800 1005153 218806 1005205
rect 218858 1005193 218864 1005205
rect 222640 1005193 222646 1005205
rect 218858 1005165 222646 1005193
rect 218858 1005153 218864 1005165
rect 222640 1005153 222646 1005165
rect 222698 1005153 222704 1005205
rect 316816 1005153 316822 1005205
rect 316874 1005193 316880 1005205
rect 331216 1005193 331222 1005205
rect 316874 1005165 331222 1005193
rect 316874 1005153 316880 1005165
rect 331216 1005153 331222 1005165
rect 331274 1005153 331280 1005205
rect 195280 1003229 195286 1003281
rect 195338 1003269 195344 1003281
rect 377296 1003269 377302 1003281
rect 195338 1003241 209150 1003269
rect 195338 1003229 195344 1003241
rect 209122 1003207 209150 1003241
rect 357442 1003241 377302 1003269
rect 357442 1003207 357470 1003241
rect 377296 1003229 377302 1003241
rect 377354 1003229 377360 1003281
rect 434608 1003269 434614 1003281
rect 428674 1003241 434614 1003269
rect 428674 1003207 428702 1003241
rect 434608 1003229 434614 1003241
rect 434666 1003229 434672 1003281
rect 439120 1003229 439126 1003281
rect 439178 1003269 439184 1003281
rect 466480 1003269 466486 1003281
rect 439178 1003241 466486 1003269
rect 439178 1003229 439184 1003241
rect 466480 1003229 466486 1003241
rect 466538 1003229 466544 1003281
rect 519664 1003269 519670 1003281
rect 502402 1003241 519670 1003269
rect 502402 1003207 502430 1003241
rect 519664 1003229 519670 1003241
rect 519722 1003229 519728 1003281
rect 160432 1003155 160438 1003207
rect 160490 1003195 160496 1003207
rect 164272 1003195 164278 1003207
rect 160490 1003167 164278 1003195
rect 160490 1003155 160496 1003167
rect 164272 1003155 164278 1003167
rect 164330 1003155 164336 1003207
rect 209104 1003155 209110 1003207
rect 209162 1003155 209168 1003207
rect 211792 1003155 211798 1003207
rect 211850 1003195 211856 1003207
rect 213808 1003195 213814 1003207
rect 211850 1003167 213814 1003195
rect 211850 1003155 211856 1003167
rect 213808 1003155 213814 1003167
rect 213866 1003155 213872 1003207
rect 357424 1003155 357430 1003207
rect 357482 1003155 357488 1003207
rect 362512 1003155 362518 1003207
rect 362570 1003195 362576 1003207
rect 367216 1003195 367222 1003207
rect 362570 1003167 367222 1003195
rect 362570 1003155 362576 1003167
rect 367216 1003155 367222 1003167
rect 367274 1003155 367280 1003207
rect 428656 1003155 428662 1003207
rect 428714 1003155 428720 1003207
rect 429520 1003155 429526 1003207
rect 429578 1003195 429584 1003207
rect 466384 1003195 466390 1003207
rect 429578 1003167 466390 1003195
rect 429578 1003155 429584 1003167
rect 466384 1003155 466390 1003167
rect 466442 1003155 466448 1003207
rect 502384 1003155 502390 1003207
rect 502442 1003155 502448 1003207
rect 519760 1003195 519766 1003207
rect 502882 1003167 519766 1003195
rect 425392 1003081 425398 1003133
rect 425450 1003121 425456 1003133
rect 466288 1003121 466294 1003133
rect 425450 1003093 466294 1003121
rect 425450 1003081 425456 1003093
rect 466288 1003081 466294 1003093
rect 466346 1003081 466352 1003133
rect 428272 1003007 428278 1003059
rect 428330 1003047 428336 1003059
rect 429136 1003047 429142 1003059
rect 428330 1003019 429142 1003047
rect 428330 1003007 428336 1003019
rect 429136 1003007 429142 1003019
rect 429194 1003007 429200 1003059
rect 430288 1003007 430294 1003059
rect 430346 1003047 430352 1003059
rect 434896 1003047 434902 1003059
rect 430346 1003019 434902 1003047
rect 430346 1003007 430352 1003019
rect 434896 1003007 434902 1003019
rect 434954 1003007 434960 1003059
rect 435376 1003007 435382 1003059
rect 435434 1003047 435440 1003059
rect 466192 1003047 466198 1003059
rect 435434 1003019 466198 1003047
rect 435434 1003007 435440 1003019
rect 466192 1003007 466198 1003019
rect 466250 1003007 466256 1003059
rect 501328 1003007 501334 1003059
rect 501386 1003047 501392 1003059
rect 502882 1003047 502910 1003167
rect 519760 1003155 519766 1003167
rect 519818 1003155 519824 1003207
rect 501386 1003019 502910 1003047
rect 501386 1003007 501392 1003019
rect 502960 1003007 502966 1003059
rect 503018 1003047 503024 1003059
rect 519856 1003047 519862 1003059
rect 503018 1003019 519862 1003047
rect 503018 1003007 503024 1003019
rect 519856 1003007 519862 1003019
rect 519914 1003007 519920 1003059
rect 555376 1003007 555382 1003059
rect 555434 1003047 555440 1003059
rect 572752 1003047 572758 1003059
rect 555434 1003019 572758 1003047
rect 555434 1003007 555440 1003019
rect 572752 1003007 572758 1003019
rect 572810 1003007 572816 1003059
rect 161488 1002933 161494 1002985
rect 161546 1002973 161552 1002985
rect 169936 1002973 169942 1002985
rect 161546 1002945 169942 1002973
rect 161546 1002933 161552 1002945
rect 169936 1002933 169942 1002945
rect 169994 1002933 170000 1002985
rect 298288 1002933 298294 1002985
rect 298346 1002973 298352 1002985
rect 312112 1002973 312118 1002985
rect 298346 1002945 312118 1002973
rect 298346 1002933 298352 1002945
rect 312112 1002933 312118 1002945
rect 312170 1002933 312176 1002985
rect 426064 1002933 426070 1002985
rect 426122 1002973 426128 1002985
rect 426122 1002945 439070 1002973
rect 426122 1002933 426128 1002945
rect 299344 1002859 299350 1002911
rect 299402 1002899 299408 1002911
rect 308848 1002899 308854 1002911
rect 299402 1002871 308854 1002899
rect 299402 1002859 299408 1002871
rect 308848 1002859 308854 1002871
rect 308906 1002859 308912 1002911
rect 423856 1002859 423862 1002911
rect 423914 1002899 423920 1002911
rect 435376 1002899 435382 1002911
rect 423914 1002871 435382 1002899
rect 423914 1002859 423920 1002871
rect 435376 1002859 435382 1002871
rect 435434 1002859 435440 1002911
rect 299440 1002785 299446 1002837
rect 299498 1002825 299504 1002837
rect 309328 1002825 309334 1002837
rect 299498 1002797 309334 1002825
rect 299498 1002785 299504 1002797
rect 309328 1002785 309334 1002797
rect 309386 1002785 309392 1002837
rect 424336 1002785 424342 1002837
rect 424394 1002825 424400 1002837
rect 429520 1002825 429526 1002837
rect 424394 1002797 429526 1002825
rect 424394 1002785 424400 1002797
rect 429520 1002785 429526 1002797
rect 429578 1002785 429584 1002837
rect 432016 1002785 432022 1002837
rect 432074 1002825 432080 1002837
rect 434992 1002825 434998 1002837
rect 432074 1002797 434998 1002825
rect 432074 1002785 432080 1002797
rect 434992 1002785 434998 1002797
rect 435050 1002785 435056 1002837
rect 439042 1002825 439070 1002945
rect 439216 1002933 439222 1002985
rect 439274 1002973 439280 1002985
rect 465520 1002973 465526 1002985
rect 439274 1002945 465526 1002973
rect 439274 1002933 439280 1002945
rect 465520 1002933 465526 1002945
rect 465578 1002933 465584 1002985
rect 554320 1002933 554326 1002985
rect 554378 1002973 554384 1002985
rect 573040 1002973 573046 1002985
rect 554378 1002945 573046 1002973
rect 554378 1002933 554384 1002945
rect 573040 1002933 573046 1002945
rect 573098 1002933 573104 1002985
rect 553744 1002859 553750 1002911
rect 553802 1002899 553808 1002911
rect 570736 1002899 570742 1002911
rect 553802 1002871 570742 1002899
rect 553802 1002859 553808 1002871
rect 570736 1002859 570742 1002871
rect 570794 1002859 570800 1002911
rect 439216 1002825 439222 1002837
rect 439042 1002797 439222 1002825
rect 439216 1002785 439222 1002797
rect 439274 1002785 439280 1002837
rect 299248 1002711 299254 1002763
rect 299306 1002751 299312 1002763
rect 308272 1002751 308278 1002763
rect 299306 1002723 308278 1002751
rect 299306 1002711 299312 1002723
rect 308272 1002711 308278 1002723
rect 308330 1002711 308336 1002763
rect 358576 1002711 358582 1002763
rect 358634 1002751 358640 1002763
rect 373360 1002751 373366 1002763
rect 358634 1002723 373366 1002751
rect 358634 1002711 358640 1002723
rect 373360 1002711 373366 1002723
rect 373418 1002711 373424 1002763
rect 424816 1002711 424822 1002763
rect 424874 1002751 424880 1002763
rect 439120 1002751 439126 1002763
rect 424874 1002723 439126 1002751
rect 424874 1002711 424880 1002723
rect 439120 1002711 439126 1002723
rect 439178 1002711 439184 1002763
rect 554896 1002711 554902 1002763
rect 554954 1002751 554960 1002763
rect 571216 1002751 571222 1002763
rect 554954 1002723 571222 1002751
rect 554954 1002711 554960 1002723
rect 571216 1002711 571222 1002723
rect 571274 1002711 571280 1002763
rect 358000 1002637 358006 1002689
rect 358058 1002677 358064 1002689
rect 372496 1002677 372502 1002689
rect 358058 1002649 372502 1002677
rect 358058 1002637 358064 1002649
rect 372496 1002637 372502 1002649
rect 372554 1002637 372560 1002689
rect 427600 1002637 427606 1002689
rect 427658 1002677 427664 1002689
rect 435088 1002677 435094 1002689
rect 427658 1002649 435094 1002677
rect 427658 1002637 427664 1002649
rect 435088 1002637 435094 1002649
rect 435146 1002637 435152 1002689
rect 143920 1002563 143926 1002615
rect 143978 1002603 143984 1002615
rect 153328 1002603 153334 1002615
rect 143978 1002575 153334 1002603
rect 143978 1002563 143984 1002575
rect 153328 1002563 153334 1002575
rect 153386 1002563 153392 1002615
rect 429232 1002563 429238 1002615
rect 429290 1002603 429296 1002615
rect 434704 1002603 434710 1002615
rect 429290 1002575 434710 1002603
rect 429290 1002563 429296 1002575
rect 434704 1002563 434710 1002575
rect 434762 1002563 434768 1002615
rect 553264 1002563 553270 1002615
rect 553322 1002603 553328 1002615
rect 572944 1002603 572950 1002615
rect 553322 1002575 572950 1002603
rect 553322 1002563 553328 1002575
rect 572944 1002563 572950 1002575
rect 573002 1002563 573008 1002615
rect 143728 1002489 143734 1002541
rect 143786 1002529 143792 1002541
rect 152656 1002529 152662 1002541
rect 143786 1002501 152662 1002529
rect 143786 1002489 143792 1002501
rect 152656 1002489 152662 1002501
rect 152714 1002489 152720 1002541
rect 361840 1002489 361846 1002541
rect 361898 1002529 361904 1002541
rect 371536 1002529 371542 1002541
rect 361898 1002501 371542 1002529
rect 361898 1002489 361904 1002501
rect 371536 1002489 371542 1002501
rect 371594 1002489 371600 1002541
rect 426640 1002489 426646 1002541
rect 426698 1002529 426704 1002541
rect 435184 1002529 435190 1002541
rect 426698 1002501 435190 1002529
rect 426698 1002489 426704 1002501
rect 435184 1002489 435190 1002501
rect 435242 1002489 435248 1002541
rect 144016 1002415 144022 1002467
rect 144074 1002455 144080 1002467
rect 151600 1002455 151606 1002467
rect 144074 1002427 151606 1002455
rect 144074 1002415 144080 1002427
rect 151600 1002415 151606 1002427
rect 151658 1002415 151664 1002467
rect 427120 1002415 427126 1002467
rect 427178 1002455 427184 1002467
rect 435280 1002455 435286 1002467
rect 427178 1002427 435286 1002455
rect 427178 1002415 427184 1002427
rect 435280 1002415 435286 1002427
rect 435338 1002415 435344 1002467
rect 143824 1002341 143830 1002393
rect 143882 1002381 143888 1002393
rect 151024 1002381 151030 1002393
rect 143882 1002353 151030 1002381
rect 143882 1002341 143888 1002353
rect 151024 1002341 151030 1002353
rect 151082 1002341 151088 1002393
rect 362896 1002341 362902 1002393
rect 362954 1002381 362960 1002393
rect 371632 1002381 371638 1002393
rect 362954 1002353 371638 1002381
rect 362954 1002341 362960 1002353
rect 371632 1002341 371638 1002353
rect 371690 1002341 371696 1002393
rect 429136 1002341 429142 1002393
rect 429194 1002381 429200 1002393
rect 443536 1002381 443542 1002393
rect 429194 1002353 443542 1002381
rect 429194 1002341 429200 1002353
rect 443536 1002341 443542 1002353
rect 443594 1002341 443600 1002393
rect 144112 1002267 144118 1002319
rect 144170 1002307 144176 1002319
rect 175696 1002307 175702 1002319
rect 144170 1002279 175702 1002307
rect 144170 1002267 144176 1002279
rect 175696 1002267 175702 1002279
rect 175754 1002267 175760 1002319
rect 359056 1002267 359062 1002319
rect 359114 1002307 359120 1002319
rect 365776 1002307 365782 1002319
rect 359114 1002279 365782 1002307
rect 359114 1002267 359120 1002279
rect 365776 1002267 365782 1002279
rect 365834 1002267 365840 1002319
rect 489136 1002267 489142 1002319
rect 489194 1002307 489200 1002319
rect 519088 1002307 519094 1002319
rect 489194 1002279 519094 1002307
rect 489194 1002267 489200 1002279
rect 519088 1002267 519094 1002279
rect 519146 1002267 519152 1002319
rect 361360 1002193 361366 1002245
rect 361418 1002233 361424 1002245
rect 379984 1002233 379990 1002245
rect 361418 1002205 379990 1002233
rect 361418 1002193 361424 1002205
rect 379984 1002193 379990 1002205
rect 380042 1002193 380048 1002245
rect 356368 1001231 356374 1001283
rect 356426 1001271 356432 1001283
rect 379792 1001271 379798 1001283
rect 356426 1001243 379798 1001271
rect 356426 1001231 356432 1001243
rect 379792 1001231 379798 1001243
rect 379850 1001231 379856 1001283
rect 357136 1001083 357142 1001135
rect 357194 1001123 357200 1001135
rect 380080 1001123 380086 1001135
rect 357194 1001095 380086 1001123
rect 357194 1001083 357200 1001095
rect 380080 1001083 380086 1001095
rect 380138 1001083 380144 1001135
rect 465232 1001009 465238 1001061
rect 465290 1001049 465296 1001061
rect 472528 1001049 472534 1001061
rect 465290 1001021 472534 1001049
rect 465290 1001009 465296 1001021
rect 472528 1001009 472534 1001021
rect 472586 1001009 472592 1001061
rect 365776 1000935 365782 1000987
rect 365834 1000975 365840 1000987
rect 383152 1000975 383158 1000987
rect 365834 1000947 383158 1000975
rect 365834 1000935 365840 1000947
rect 383152 1000935 383158 1000947
rect 383210 1000935 383216 1000987
rect 506320 1000935 506326 1000987
rect 506378 1000975 506384 1000987
rect 515536 1000975 515542 1000987
rect 506378 1000947 515542 1000975
rect 506378 1000935 506384 1000947
rect 515536 1000935 515542 1000947
rect 515594 1000935 515600 1000987
rect 360208 1000861 360214 1000913
rect 360266 1000901 360272 1000913
rect 383440 1000901 383446 1000913
rect 360266 1000873 383446 1000901
rect 360266 1000861 360272 1000873
rect 383440 1000861 383446 1000873
rect 383498 1000861 383504 1000913
rect 430960 1000861 430966 1000913
rect 431018 1000901 431024 1000913
rect 472432 1000901 472438 1000913
rect 431018 1000873 472438 1000901
rect 431018 1000861 431024 1000873
rect 472432 1000861 472438 1000873
rect 472490 1000861 472496 1000913
rect 359632 1000787 359638 1000839
rect 359690 1000827 359696 1000839
rect 383248 1000827 383254 1000839
rect 359690 1000799 383254 1000827
rect 359690 1000787 359696 1000799
rect 383248 1000787 383254 1000799
rect 383306 1000787 383312 1000839
rect 429904 1000787 429910 1000839
rect 429962 1000827 429968 1000839
rect 472624 1000827 472630 1000839
rect 429962 1000799 472630 1000827
rect 429962 1000787 429968 1000799
rect 472624 1000787 472630 1000799
rect 472682 1000787 472688 1000839
rect 507856 1000787 507862 1000839
rect 507914 1000827 507920 1000839
rect 512656 1000827 512662 1000839
rect 507914 1000799 512662 1000827
rect 507914 1000787 507920 1000799
rect 512656 1000787 512662 1000799
rect 512714 1000787 512720 1000839
rect 552304 1000787 552310 1000839
rect 552362 1000827 552368 1000839
rect 573136 1000827 573142 1000839
rect 552362 1000799 573142 1000827
rect 552362 1000787 552368 1000799
rect 573136 1000787 573142 1000799
rect 573194 1000787 573200 1000839
rect 506896 1000639 506902 1000691
rect 506954 1000679 506960 1000691
rect 512176 1000679 512182 1000691
rect 506954 1000651 512182 1000679
rect 506954 1000639 506960 1000651
rect 512176 1000639 512182 1000651
rect 512234 1000639 512240 1000691
rect 377296 999825 377302 999877
rect 377354 999865 377360 999877
rect 383344 999865 383350 999877
rect 377354 999837 383350 999865
rect 377354 999825 377360 999837
rect 383344 999825 383350 999837
rect 383402 999825 383408 999877
rect 504688 999825 504694 999877
rect 504746 999865 504752 999877
rect 512080 999865 512086 999877
rect 504746 999837 512086 999865
rect 504746 999825 504752 999837
rect 512080 999825 512086 999837
rect 512138 999825 512144 999877
rect 509680 999751 509686 999803
rect 509738 999791 509744 999803
rect 519952 999791 519958 999803
rect 509738 999763 519958 999791
rect 509738 999751 509744 999763
rect 519952 999751 519958 999763
rect 520010 999751 520016 999803
rect 613456 999751 613462 999803
rect 613514 999791 613520 999803
rect 625840 999791 625846 999803
rect 613514 999763 625846 999791
rect 613514 999751 613520 999763
rect 625840 999751 625846 999763
rect 625898 999751 625904 999803
rect 503632 999677 503638 999729
rect 503690 999717 503696 999729
rect 512272 999717 512278 999729
rect 503690 999689 512278 999717
rect 503690 999677 503696 999689
rect 512272 999677 512278 999689
rect 512330 999677 512336 999729
rect 610576 999677 610582 999729
rect 610634 999717 610640 999729
rect 625552 999717 625558 999729
rect 610634 999689 625558 999717
rect 610634 999677 610640 999689
rect 625552 999677 625558 999689
rect 625610 999677 625616 999729
rect 195472 999603 195478 999655
rect 195530 999643 195536 999655
rect 195530 999615 207134 999643
rect 195530 999603 195536 999615
rect 195184 999455 195190 999507
rect 195242 999495 195248 999507
rect 207106 999495 207134 999615
rect 500752 999603 500758 999655
rect 500810 999643 500816 999655
rect 511984 999643 511990 999655
rect 500810 999615 511990 999643
rect 500810 999603 500816 999615
rect 511984 999603 511990 999615
rect 512042 999603 512048 999655
rect 512080 999603 512086 999655
rect 512138 999603 512144 999655
rect 604240 999603 604246 999655
rect 604298 999643 604304 999655
rect 625648 999643 625654 999655
rect 604298 999615 625654 999643
rect 604298 999603 604304 999615
rect 625648 999603 625654 999615
rect 625706 999603 625712 999655
rect 503632 999529 503638 999581
rect 503690 999569 503696 999581
rect 512098 999569 512126 999603
rect 503690 999541 512126 999569
rect 503690 999529 503696 999541
rect 609040 999529 609046 999581
rect 609098 999569 609104 999581
rect 625456 999569 625462 999581
rect 609098 999541 625462 999569
rect 609098 999529 609104 999541
rect 625456 999529 625462 999541
rect 625514 999529 625520 999581
rect 226000 999495 226006 999507
rect 195242 999467 207038 999495
rect 207106 999467 226006 999495
rect 195242 999455 195248 999467
rect 92656 999381 92662 999433
rect 92714 999421 92720 999433
rect 126640 999421 126646 999433
rect 92714 999393 126646 999421
rect 92714 999381 92720 999393
rect 126640 999381 126646 999393
rect 126698 999381 126704 999433
rect 143728 999381 143734 999433
rect 143786 999421 143792 999433
rect 155536 999421 155542 999433
rect 143786 999393 155542 999421
rect 143786 999381 143792 999393
rect 155536 999381 155542 999393
rect 155594 999381 155600 999433
rect 195088 999381 195094 999433
rect 195146 999421 195152 999433
rect 206896 999421 206902 999433
rect 195146 999393 206902 999421
rect 195146 999381 195152 999393
rect 206896 999381 206902 999393
rect 206954 999381 206960 999433
rect 207010 999421 207038 999467
rect 226000 999455 226006 999467
rect 226058 999455 226064 999507
rect 371536 999455 371542 999507
rect 371594 999495 371600 999507
rect 371594 999467 380030 999495
rect 371594 999455 371600 999467
rect 222928 999421 222934 999433
rect 207010 999393 222934 999421
rect 222928 999381 222934 999393
rect 222986 999381 222992 999433
rect 246544 999381 246550 999433
rect 246602 999421 246608 999433
rect 258352 999421 258358 999433
rect 246602 999393 258358 999421
rect 246602 999381 246608 999393
rect 258352 999381 258358 999393
rect 258410 999381 258416 999433
rect 298192 999381 298198 999433
rect 298250 999421 298256 999433
rect 309904 999421 309910 999433
rect 298250 999393 309910 999421
rect 298250 999381 298256 999393
rect 309904 999381 309910 999393
rect 309962 999381 309968 999433
rect 371632 999381 371638 999433
rect 371690 999421 371696 999433
rect 379888 999421 379894 999433
rect 371690 999393 379894 999421
rect 371690 999381 371696 999393
rect 379888 999381 379894 999393
rect 379946 999381 379952 999433
rect 380002 999421 380030 999467
rect 502000 999455 502006 999507
rect 502058 999495 502064 999507
rect 512080 999495 512086 999507
rect 502058 999467 512086 999495
rect 502058 999455 502064 999467
rect 512080 999455 512086 999467
rect 512138 999455 512144 999507
rect 596176 999455 596182 999507
rect 596234 999495 596240 999507
rect 625840 999495 625846 999507
rect 596234 999467 625846 999495
rect 596234 999455 596240 999467
rect 625840 999455 625846 999467
rect 625898 999455 625904 999507
rect 380002 999393 380510 999421
rect 313744 999307 313750 999359
rect 313802 999347 313808 999359
rect 328336 999347 328342 999359
rect 313802 999319 328342 999347
rect 313802 999307 313808 999319
rect 328336 999307 328342 999319
rect 328394 999307 328400 999359
rect 364528 999307 364534 999359
rect 364586 999347 364592 999359
rect 380368 999347 380374 999359
rect 364586 999319 380374 999347
rect 364586 999307 364592 999319
rect 380368 999307 380374 999319
rect 380426 999307 380432 999359
rect 380482 999347 380510 999393
rect 488944 999381 488950 999433
rect 489002 999421 489008 999433
rect 509680 999421 509686 999433
rect 489002 999393 509686 999421
rect 489002 999381 489008 999393
rect 509680 999381 509686 999393
rect 509738 999381 509744 999433
rect 552976 999381 552982 999433
rect 553034 999421 553040 999433
rect 553034 999393 561566 999421
rect 553034 999381 553040 999393
rect 383536 999347 383542 999359
rect 380482 999319 383542 999347
rect 383536 999307 383542 999319
rect 383594 999307 383600 999359
rect 561538 999347 561566 999393
rect 593296 999381 593302 999433
rect 593354 999421 593360 999433
rect 625744 999421 625750 999433
rect 593354 999393 625750 999421
rect 593354 999381 593360 999393
rect 625744 999381 625750 999393
rect 625802 999381 625808 999433
rect 567376 999347 567382 999359
rect 561538 999319 567382 999347
rect 567376 999307 567382 999319
rect 567434 999307 567440 999359
rect 466288 999233 466294 999285
rect 466346 999273 466352 999285
rect 472048 999273 472054 999285
rect 466346 999245 472054 999273
rect 466346 999233 466352 999245
rect 472048 999233 472054 999245
rect 472106 999233 472112 999285
rect 558832 999233 558838 999285
rect 558890 999273 558896 999285
rect 573712 999273 573718 999285
rect 558890 999245 573718 999273
rect 558890 999233 558896 999245
rect 573712 999233 573718 999245
rect 573770 999233 573776 999285
rect 466480 999011 466486 999063
rect 466538 999051 466544 999063
rect 472240 999051 472246 999063
rect 466538 999023 472246 999051
rect 466538 999011 466544 999023
rect 472240 999011 472246 999023
rect 472298 999011 472304 999063
rect 465520 998937 465526 998989
rect 465578 998977 465584 998989
rect 471952 998977 471958 998989
rect 465578 998949 471958 998977
rect 465578 998937 465584 998949
rect 471952 998937 471958 998949
rect 472010 998937 472016 998989
rect 379984 998863 379990 998915
rect 380042 998903 380048 998915
rect 383056 998903 383062 998915
rect 380042 998875 383062 998903
rect 380042 998863 380048 998875
rect 383056 998863 383062 998875
rect 383114 998863 383120 998915
rect 557200 998789 557206 998841
rect 557258 998829 557264 998841
rect 573904 998829 573910 998841
rect 557258 998801 573910 998829
rect 557258 998789 557264 998801
rect 573904 998789 573910 998801
rect 573962 998789 573968 998841
rect 298384 997901 298390 997953
rect 298442 997941 298448 997953
rect 348880 997941 348886 997953
rect 298442 997913 348886 997941
rect 298442 997901 298448 997913
rect 348880 997901 348886 997913
rect 348938 997901 348944 997953
rect 572752 997901 572758 997953
rect 572810 997941 572816 997953
rect 604240 997941 604246 997953
rect 572810 997913 604246 997941
rect 572810 997901 572816 997913
rect 604240 997901 604246 997913
rect 604298 997901 604304 997953
rect 314800 997827 314806 997879
rect 314858 997867 314864 997879
rect 365200 997867 365206 997879
rect 314858 997839 365206 997867
rect 314858 997827 314864 997839
rect 365200 997827 365206 997839
rect 365258 997827 365264 997879
rect 555952 997827 555958 997879
rect 556010 997867 556016 997879
rect 593296 997867 593302 997879
rect 556010 997839 593302 997867
rect 556010 997827 556016 997839
rect 593296 997827 593302 997839
rect 593354 997827 593360 997879
rect 328336 997753 328342 997805
rect 328394 997793 328400 997805
rect 364528 997793 364534 997805
rect 328394 997765 364534 997793
rect 328394 997753 328400 997765
rect 364528 997753 364534 997765
rect 364586 997753 364592 997805
rect 558160 997753 558166 997805
rect 558218 997793 558224 997805
rect 596176 997793 596182 997805
rect 558218 997765 596182 997793
rect 558218 997753 558224 997765
rect 596176 997753 596182 997765
rect 596234 997753 596240 997805
rect 571216 997679 571222 997731
rect 571274 997719 571280 997731
rect 610576 997719 610582 997731
rect 571274 997691 610582 997719
rect 571274 997679 571280 997691
rect 610576 997679 610582 997691
rect 610634 997679 610640 997731
rect 557776 997605 557782 997657
rect 557834 997645 557840 997657
rect 613456 997645 613462 997657
rect 557834 997617 613462 997645
rect 557834 997605 557840 997617
rect 613456 997605 613462 997617
rect 613514 997605 613520 997657
rect 559408 997531 559414 997583
rect 559466 997571 559472 997583
rect 622000 997571 622006 997583
rect 559466 997543 622006 997571
rect 559466 997531 559472 997543
rect 622000 997531 622006 997543
rect 622058 997531 622064 997583
rect 573136 997457 573142 997509
rect 573194 997497 573200 997509
rect 609040 997497 609046 997509
rect 573194 997469 609046 997497
rect 573194 997457 573200 997469
rect 609040 997457 609046 997469
rect 609098 997457 609104 997509
rect 572944 997383 572950 997435
rect 573002 997423 573008 997435
rect 621904 997423 621910 997435
rect 573002 997395 621910 997423
rect 573002 997383 573008 997395
rect 621904 997383 621910 997395
rect 621962 997383 621968 997435
rect 298096 997087 298102 997139
rect 298154 997127 298160 997139
rect 313744 997127 313750 997139
rect 298154 997099 313750 997127
rect 298154 997087 298160 997099
rect 313744 997087 313750 997099
rect 313802 997087 313808 997139
rect 511984 996717 511990 996769
rect 512042 996757 512048 996769
rect 518320 996757 518326 996769
rect 512042 996729 518326 996757
rect 512042 996717 512048 996729
rect 518320 996717 518326 996729
rect 518378 996717 518384 996769
rect 196816 996643 196822 996695
rect 196874 996683 196880 996695
rect 196874 996655 205310 996683
rect 196874 996643 196880 996655
rect 97936 996495 97942 996547
rect 97994 996535 98000 996547
rect 104656 996535 104662 996547
rect 97994 996507 104662 996535
rect 97994 996495 98000 996507
rect 104656 996495 104662 996507
rect 104714 996495 104720 996547
rect 195760 996495 195766 996547
rect 195818 996535 195824 996547
rect 205168 996535 205174 996547
rect 195818 996507 205174 996535
rect 195818 996495 195824 996507
rect 205168 996495 205174 996507
rect 205226 996495 205232 996547
rect 205282 996535 205310 996655
rect 507472 996569 507478 996621
rect 507530 996609 507536 996621
rect 521296 996609 521302 996621
rect 507530 996581 521302 996609
rect 507530 996569 507536 996581
rect 521296 996569 521302 996581
rect 521354 996569 521360 996621
rect 207952 996535 207958 996547
rect 205282 996507 207958 996535
rect 207952 996495 207958 996507
rect 208010 996495 208016 996547
rect 309904 996495 309910 996547
rect 309962 996535 309968 996547
rect 311536 996535 311542 996547
rect 309962 996507 311542 996535
rect 309962 996495 309968 996507
rect 311536 996495 311542 996507
rect 311594 996495 311600 996547
rect 379888 996495 379894 996547
rect 379946 996535 379952 996547
rect 382960 996535 382966 996547
rect 379946 996507 382966 996535
rect 379946 996495 379952 996507
rect 382960 996495 382966 996507
rect 383018 996495 383024 996547
rect 505744 996495 505750 996547
rect 505802 996535 505808 996547
rect 519184 996535 519190 996547
rect 505802 996507 519190 996535
rect 505802 996495 505808 996507
rect 519184 996495 519190 996507
rect 519242 996495 519248 996547
rect 313168 996421 313174 996473
rect 313226 996461 313232 996473
rect 363952 996461 363958 996473
rect 313226 996433 363958 996461
rect 313226 996421 313232 996433
rect 363952 996421 363958 996433
rect 364010 996421 364016 996473
rect 225232 996387 225238 996399
rect 210178 996359 225238 996387
rect 107536 996273 107542 996325
rect 107594 996313 107600 996325
rect 126736 996313 126742 996325
rect 107594 996285 126742 996313
rect 107594 996273 107600 996285
rect 126736 996273 126742 996285
rect 126794 996273 126800 996325
rect 144208 996273 144214 996325
rect 144266 996313 144272 996325
rect 144266 996285 159230 996313
rect 144266 996273 144272 996285
rect 159202 996251 159230 996285
rect 159184 996199 159190 996251
rect 159242 996239 159248 996251
rect 159242 996211 160670 996239
rect 159242 996199 159248 996211
rect 107920 996051 107926 996103
rect 107978 996091 107984 996103
rect 159760 996091 159766 996103
rect 107978 996063 159766 996091
rect 107978 996051 107984 996063
rect 159760 996051 159766 996063
rect 159818 996091 159824 996103
rect 160642 996091 160670 996211
rect 210178 996103 210206 996359
rect 225232 996347 225238 996359
rect 225290 996347 225296 996399
rect 262480 996347 262486 996399
rect 262538 996387 262544 996399
rect 270640 996387 270646 996399
rect 262538 996359 270646 996387
rect 262538 996347 262544 996359
rect 270640 996347 270646 996359
rect 270698 996347 270704 996399
rect 262498 996239 262526 996347
rect 246466 996211 262526 996239
rect 246466 996165 246494 996211
rect 210658 996137 246494 996165
rect 246562 996137 262046 996165
rect 210160 996091 210166 996103
rect 159818 996063 160574 996091
rect 160642 996063 210166 996091
rect 159818 996051 159824 996063
rect 108976 995977 108982 996029
rect 109034 996017 109040 996029
rect 160432 996017 160438 996029
rect 109034 995989 160438 996017
rect 109034 995977 109040 995989
rect 160432 995977 160438 995989
rect 160490 995977 160496 996029
rect 160546 996017 160574 996063
rect 210160 996051 210166 996063
rect 210218 996051 210224 996103
rect 210658 996029 210686 996137
rect 225232 996051 225238 996103
rect 225290 996091 225296 996103
rect 246562 996091 246590 996137
rect 262018 996103 262046 996137
rect 263056 996125 263062 996177
rect 263114 996165 263120 996177
rect 314800 996165 314806 996177
rect 263114 996137 314806 996165
rect 263114 996125 263120 996137
rect 314800 996125 314806 996137
rect 314858 996125 314864 996177
rect 368656 996125 368662 996177
rect 368714 996165 368720 996177
rect 432400 996165 432406 996177
rect 368714 996137 432406 996165
rect 368714 996125 368720 996137
rect 432400 996125 432406 996137
rect 432458 996125 432464 996177
rect 432496 996125 432502 996177
rect 432554 996165 432560 996177
rect 509584 996165 509590 996177
rect 432554 996137 509590 996165
rect 432554 996125 432560 996137
rect 509584 996125 509590 996137
rect 509642 996125 509648 996177
rect 509968 996125 509974 996177
rect 510026 996165 510032 996177
rect 561040 996165 561046 996177
rect 510026 996137 561046 996165
rect 510026 996125 510032 996137
rect 561040 996125 561046 996137
rect 561098 996125 561104 996177
rect 225290 996063 246590 996091
rect 225290 996051 225296 996063
rect 247504 996051 247510 996103
rect 247562 996091 247568 996103
rect 257776 996091 257782 996103
rect 247562 996063 257782 996091
rect 247562 996051 247568 996063
rect 257776 996051 257782 996063
rect 257834 996051 257840 996103
rect 262000 996051 262006 996103
rect 262058 996091 262064 996103
rect 313168 996091 313174 996103
rect 262058 996063 313174 996091
rect 262058 996051 262064 996063
rect 313168 996051 313174 996063
rect 313226 996051 313232 996103
rect 380368 996051 380374 996103
rect 380426 996091 380432 996103
rect 434992 996091 434998 996103
rect 380426 996063 434998 996091
rect 380426 996051 380432 996063
rect 434992 996051 434998 996063
rect 435050 996051 435056 996103
rect 471568 996051 471574 996103
rect 471626 996091 471632 996103
rect 508912 996091 508918 996103
rect 471626 996063 508918 996091
rect 471626 996051 471632 996063
rect 508912 996051 508918 996063
rect 508970 996091 508976 996103
rect 560176 996091 560182 996103
rect 508970 996063 560182 996091
rect 508970 996051 508976 996063
rect 560176 996051 560182 996063
rect 560234 996051 560240 996103
rect 210640 996017 210646 996029
rect 160546 995989 210646 996017
rect 210640 995977 210646 995989
rect 210698 995977 210704 996029
rect 222640 995977 222646 996029
rect 222698 996017 222704 996029
rect 263248 996017 263254 996029
rect 222698 995989 263254 996017
rect 222698 995977 222704 995989
rect 263248 995977 263254 995989
rect 263306 995977 263312 996029
rect 363952 995977 363958 996029
rect 364010 996017 364016 996029
rect 430960 996017 430966 996029
rect 364010 995989 430966 996017
rect 364010 995977 364016 995989
rect 430960 995977 430966 995989
rect 431018 996017 431024 996029
rect 437488 996017 437494 996029
rect 431018 995989 437494 996017
rect 431018 995977 431024 995989
rect 437488 995977 437494 995989
rect 437546 995977 437552 996029
rect 470128 995977 470134 996029
rect 470186 996017 470192 996029
rect 508336 996017 508342 996029
rect 470186 995989 508342 996017
rect 470186 995977 470192 995989
rect 508336 995977 508342 995989
rect 508394 996017 508400 996029
rect 559600 996017 559606 996029
rect 508394 995989 559606 996017
rect 508394 995977 508400 995989
rect 559600 995977 559606 995989
rect 559658 995977 559664 996029
rect 94960 995903 94966 995955
rect 95018 995943 95024 995955
rect 102832 995943 102838 995955
rect 95018 995915 102838 995943
rect 95018 995903 95024 995915
rect 102832 995903 102838 995915
rect 102890 995903 102896 995955
rect 144016 995943 144022 995955
rect 136834 995915 144022 995943
rect 101200 995869 101206 995881
rect 85954 995841 101206 995869
rect 85954 995807 85982 995841
rect 101200 995829 101206 995841
rect 101258 995829 101264 995881
rect 136834 995807 136862 995915
rect 144016 995903 144022 995915
rect 144074 995903 144080 995955
rect 172816 995903 172822 995955
rect 172874 995943 172880 995955
rect 211792 995943 211798 995955
rect 172874 995915 211798 995943
rect 172874 995903 172880 995915
rect 211792 995903 211798 995915
rect 211850 995903 211856 995955
rect 250480 995903 250486 995955
rect 250538 995943 250544 995955
rect 254512 995943 254518 995955
rect 250538 995915 254518 995943
rect 250538 995903 250544 995915
rect 254512 995903 254518 995915
rect 254570 995903 254576 995955
rect 299440 995943 299446 995955
rect 283714 995915 299446 995943
rect 143920 995869 143926 995881
rect 139330 995841 143926 995869
rect 139330 995807 139358 995841
rect 143920 995829 143926 995841
rect 143978 995829 143984 995881
rect 204016 995869 204022 995881
rect 188866 995841 204022 995869
rect 188866 995807 188894 995841
rect 204016 995829 204022 995841
rect 204074 995829 204080 995881
rect 283714 995807 283742 995915
rect 299440 995903 299446 995915
rect 299498 995903 299504 995955
rect 382960 995903 382966 995955
rect 383018 995943 383024 995955
rect 383018 995915 396734 995943
rect 383018 995903 383024 995915
rect 310288 995869 310294 995881
rect 290626 995841 310294 995869
rect 290626 995807 290654 995841
rect 310288 995829 310294 995841
rect 310346 995829 310352 995881
rect 383344 995829 383350 995881
rect 383402 995869 383408 995881
rect 383402 995841 389438 995869
rect 383402 995829 383408 995841
rect 389410 995807 389438 995841
rect 396706 995807 396734 995915
rect 466384 995903 466390 995955
rect 466442 995943 466448 995955
rect 466442 995915 471902 995943
rect 466442 995903 466448 995915
rect 417520 995829 417526 995881
rect 417578 995869 417584 995881
rect 421552 995869 421558 995881
rect 417578 995841 421558 995869
rect 417578 995829 417584 995841
rect 421552 995829 421558 995841
rect 421610 995829 421616 995881
rect 471874 995869 471902 995915
rect 471952 995903 471958 995955
rect 472010 995943 472016 995955
rect 472010 995915 483902 995943
rect 472010 995903 472016 995915
rect 471874 995841 481406 995869
rect 481378 995807 481406 995841
rect 483874 995807 483902 995915
rect 625456 995903 625462 995955
rect 625514 995943 625520 995955
rect 625514 995915 635870 995943
rect 625514 995903 625520 995915
rect 621904 995829 621910 995881
rect 621962 995869 621968 995881
rect 621962 995841 631550 995869
rect 621962 995829 621968 995841
rect 631522 995807 631550 995841
rect 635842 995807 635870 995915
rect 85936 995755 85942 995807
rect 85994 995755 86000 995807
rect 91504 995755 91510 995807
rect 91562 995795 91568 995807
rect 103984 995795 103990 995807
rect 91562 995767 103990 995795
rect 91562 995755 91568 995767
rect 103984 995755 103990 995767
rect 104042 995755 104048 995807
rect 136816 995755 136822 995807
rect 136874 995755 136880 995807
rect 139312 995755 139318 995807
rect 139370 995755 139376 995807
rect 142960 995755 142966 995807
rect 143018 995795 143024 995807
rect 143728 995795 143734 995807
rect 143018 995767 143734 995795
rect 143018 995755 143024 995767
rect 143728 995755 143734 995767
rect 143786 995755 143792 995807
rect 149584 995755 149590 995807
rect 149642 995795 149648 995807
rect 154864 995795 154870 995807
rect 149642 995767 154870 995795
rect 149642 995755 149648 995767
rect 154864 995755 154870 995767
rect 154922 995755 154928 995807
rect 175696 995755 175702 995807
rect 175754 995795 175760 995807
rect 185200 995795 185206 995807
rect 175754 995767 185206 995795
rect 175754 995755 175760 995767
rect 185200 995755 185206 995767
rect 185258 995755 185264 995807
rect 188848 995755 188854 995807
rect 188906 995755 188912 995807
rect 190576 995755 190582 995807
rect 190634 995795 190640 995807
rect 204688 995795 204694 995807
rect 190634 995767 204694 995795
rect 190634 995755 190640 995767
rect 204688 995755 204694 995767
rect 204746 995755 204752 995807
rect 226000 995755 226006 995807
rect 226058 995795 226064 995807
rect 226058 995767 236414 995795
rect 226058 995755 226064 995767
rect 94960 995681 94966 995733
rect 95018 995721 95024 995733
rect 102448 995721 102454 995733
rect 95018 995693 102454 995721
rect 95018 995681 95024 995693
rect 102448 995681 102454 995693
rect 102506 995681 102512 995733
rect 137968 995681 137974 995733
rect 138026 995721 138032 995733
rect 143824 995721 143830 995733
rect 138026 995693 143830 995721
rect 138026 995681 138032 995693
rect 143824 995681 143830 995693
rect 143882 995681 143888 995733
rect 188080 995681 188086 995733
rect 188138 995721 188144 995733
rect 203056 995721 203062 995733
rect 188138 995693 203062 995721
rect 188138 995681 188144 995693
rect 203056 995681 203062 995693
rect 203114 995681 203120 995733
rect 95056 995607 95062 995659
rect 95114 995647 95120 995659
rect 102352 995647 102358 995659
rect 95114 995619 102358 995647
rect 95114 995607 95120 995619
rect 102352 995607 102358 995619
rect 102410 995607 102416 995659
rect 137392 995607 137398 995659
rect 137450 995647 137456 995659
rect 143632 995647 143638 995659
rect 137450 995619 143638 995647
rect 137450 995607 137456 995619
rect 143632 995607 143638 995619
rect 143690 995607 143696 995659
rect 144208 995647 144214 995659
rect 143746 995619 144214 995647
rect 93520 995533 93526 995585
rect 93578 995573 93584 995585
rect 98032 995573 98038 995585
rect 93578 995545 98038 995573
rect 93578 995533 93584 995545
rect 98032 995533 98038 995545
rect 98090 995533 98096 995585
rect 126736 995533 126742 995585
rect 126794 995573 126800 995585
rect 143746 995573 143774 995619
rect 144208 995607 144214 995619
rect 144266 995607 144272 995659
rect 194416 995607 194422 995659
rect 194474 995647 194480 995659
rect 195088 995647 195094 995659
rect 194474 995619 195094 995647
rect 194474 995607 194480 995619
rect 195088 995607 195094 995619
rect 195146 995607 195152 995659
rect 236386 995647 236414 995767
rect 236464 995755 236470 995807
rect 236522 995795 236528 995807
rect 254896 995795 254902 995807
rect 236522 995767 254902 995795
rect 236522 995755 236528 995767
rect 254896 995755 254902 995767
rect 254954 995755 254960 995807
rect 283696 995755 283702 995807
rect 283754 995755 283760 995807
rect 290608 995755 290614 995807
rect 290666 995755 290672 995807
rect 292528 995755 292534 995807
rect 292586 995795 292592 995807
rect 305488 995795 305494 995807
rect 292586 995767 305494 995795
rect 292586 995755 292592 995767
rect 305488 995755 305494 995767
rect 305546 995755 305552 995807
rect 360880 995755 360886 995807
rect 360938 995795 360944 995807
rect 365776 995795 365782 995807
rect 360938 995767 365782 995795
rect 360938 995755 360944 995767
rect 365776 995755 365782 995767
rect 365834 995755 365840 995807
rect 366736 995755 366742 995807
rect 366794 995795 366800 995807
rect 371632 995795 371638 995807
rect 366794 995767 371638 995795
rect 366794 995755 366800 995767
rect 371632 995755 371638 995767
rect 371690 995755 371696 995807
rect 383632 995755 383638 995807
rect 383690 995795 383696 995807
rect 384400 995795 384406 995807
rect 383690 995767 384406 995795
rect 383690 995755 383696 995767
rect 384400 995755 384406 995767
rect 384458 995755 384464 995807
rect 389392 995755 389398 995807
rect 389450 995755 389456 995807
rect 396688 995755 396694 995807
rect 396746 995755 396752 995807
rect 472624 995755 472630 995807
rect 472682 995795 472688 995807
rect 473296 995795 473302 995807
rect 472682 995767 473302 995795
rect 472682 995755 472688 995767
rect 473296 995755 473302 995767
rect 473354 995755 473360 995807
rect 481360 995755 481366 995807
rect 481418 995755 481424 995807
rect 483856 995755 483862 995807
rect 483914 995755 483920 995807
rect 485680 995755 485686 995807
rect 485738 995795 485744 995807
rect 488944 995795 488950 995807
rect 485738 995767 488950 995795
rect 485738 995755 485744 995767
rect 488944 995755 488950 995767
rect 489002 995755 489008 995807
rect 524080 995755 524086 995807
rect 524138 995795 524144 995807
rect 529840 995795 529846 995807
rect 524138 995767 529846 995795
rect 524138 995755 524144 995767
rect 529840 995755 529846 995767
rect 529898 995755 529904 995807
rect 556528 995755 556534 995807
rect 556586 995795 556592 995807
rect 563248 995795 563254 995807
rect 556586 995767 563254 995795
rect 556586 995755 556592 995767
rect 563248 995755 563254 995767
rect 563306 995755 563312 995807
rect 622000 995755 622006 995807
rect 622058 995795 622064 995807
rect 627856 995795 627862 995807
rect 622058 995767 627862 995795
rect 622058 995755 622064 995767
rect 627856 995755 627862 995767
rect 627914 995755 627920 995807
rect 631504 995755 631510 995807
rect 631562 995755 631568 995807
rect 635824 995755 635830 995807
rect 635882 995755 635888 995807
rect 638800 995755 638806 995807
rect 638858 995795 638864 995807
rect 649936 995795 649942 995807
rect 638858 995767 649942 995795
rect 638858 995755 638864 995767
rect 649936 995755 649942 995767
rect 649994 995755 650000 995807
rect 245680 995681 245686 995733
rect 245738 995721 245744 995733
rect 246544 995721 246550 995733
rect 245738 995693 246550 995721
rect 245738 995681 245744 995693
rect 246544 995681 246550 995693
rect 246602 995681 246608 995733
rect 250384 995681 250390 995733
rect 250442 995721 250448 995733
rect 257104 995721 257110 995733
rect 250442 995693 257110 995721
rect 250442 995681 250448 995693
rect 257104 995681 257110 995693
rect 257162 995681 257168 995733
rect 291184 995681 291190 995733
rect 291242 995721 291248 995733
rect 305968 995721 305974 995733
rect 291242 995693 305974 995721
rect 291242 995681 291248 995693
rect 305968 995681 305974 995693
rect 306026 995681 306032 995733
rect 366160 995681 366166 995733
rect 366218 995721 366224 995733
rect 371728 995721 371734 995733
rect 366218 995693 371734 995721
rect 366218 995681 366224 995693
rect 371728 995681 371734 995693
rect 371786 995681 371792 995733
rect 383440 995681 383446 995733
rect 383498 995721 383504 995733
rect 384976 995721 384982 995733
rect 383498 995693 384982 995721
rect 383498 995681 383504 995693
rect 384976 995681 384982 995693
rect 385034 995681 385040 995733
rect 472528 995681 472534 995733
rect 472586 995721 472592 995733
rect 474064 995721 474070 995733
rect 472586 995693 474070 995721
rect 472586 995681 472592 995693
rect 474064 995681 474070 995693
rect 474122 995681 474128 995733
rect 523984 995681 523990 995733
rect 524042 995721 524048 995733
rect 525328 995721 525334 995733
rect 524042 995693 525334 995721
rect 524042 995681 524048 995693
rect 525328 995681 525334 995693
rect 525386 995681 525392 995733
rect 625840 995681 625846 995733
rect 625898 995721 625904 995733
rect 626512 995721 626518 995733
rect 625898 995693 626518 995721
rect 625898 995681 625904 995693
rect 626512 995681 626518 995693
rect 626570 995681 626576 995733
rect 237232 995647 237238 995659
rect 236386 995619 237238 995647
rect 237232 995607 237238 995619
rect 237290 995607 237296 995659
rect 247600 995607 247606 995659
rect 247658 995647 247664 995659
rect 255952 995647 255958 995659
rect 247658 995619 255958 995647
rect 247658 995607 247664 995619
rect 255952 995607 255958 995619
rect 256010 995607 256016 995659
rect 297328 995607 297334 995659
rect 297386 995647 297392 995659
rect 298192 995647 298198 995659
rect 297386 995619 298198 995647
rect 297386 995607 297392 995619
rect 298192 995607 298198 995619
rect 298250 995607 298256 995659
rect 383248 995607 383254 995659
rect 383306 995647 383312 995659
rect 388048 995647 388054 995659
rect 383306 995619 388054 995647
rect 383306 995607 383312 995619
rect 388048 995607 388054 995619
rect 388106 995607 388112 995659
rect 472432 995607 472438 995659
rect 472490 995647 472496 995659
rect 474640 995647 474646 995659
rect 472490 995619 474646 995647
rect 472490 995607 472496 995619
rect 474640 995607 474646 995619
rect 474698 995607 474704 995659
rect 523888 995607 523894 995659
rect 523946 995647 523952 995659
rect 524752 995647 524758 995659
rect 523946 995619 524758 995647
rect 523946 995607 523952 995619
rect 524752 995607 524758 995619
rect 524810 995607 524816 995659
rect 559600 995607 559606 995659
rect 559658 995647 559664 995659
rect 564592 995647 564598 995659
rect 559658 995619 564598 995647
rect 559658 995607 559664 995619
rect 564592 995607 564598 995619
rect 564650 995607 564656 995659
rect 625744 995607 625750 995659
rect 625802 995647 625808 995659
rect 627088 995647 627094 995659
rect 625802 995619 627094 995647
rect 625802 995607 625808 995619
rect 627088 995607 627094 995619
rect 627146 995607 627152 995659
rect 126794 995545 143774 995573
rect 126794 995533 126800 995545
rect 143824 995533 143830 995585
rect 143882 995573 143888 995585
rect 144112 995573 144118 995585
rect 143882 995545 144118 995573
rect 143882 995533 143888 995545
rect 144112 995533 144118 995545
rect 144170 995533 144176 995585
rect 191920 995533 191926 995585
rect 191978 995573 191984 995585
rect 195184 995573 195190 995585
rect 191978 995545 195190 995573
rect 191978 995533 191984 995545
rect 195184 995533 195190 995545
rect 195242 995533 195248 995585
rect 295408 995533 295414 995585
rect 295466 995573 295472 995585
rect 298288 995573 298294 995585
rect 295466 995545 298294 995573
rect 295466 995533 295472 995545
rect 298288 995533 298294 995545
rect 298346 995533 298352 995585
rect 383152 995533 383158 995585
rect 383210 995573 383216 995585
rect 388816 995573 388822 995585
rect 383210 995545 388822 995573
rect 383210 995533 383216 995545
rect 388816 995533 388822 995545
rect 388874 995533 388880 995585
rect 472144 995533 472150 995585
rect 472202 995573 472208 995585
rect 476368 995573 476374 995585
rect 472202 995545 476374 995573
rect 472202 995533 472208 995545
rect 476368 995533 476374 995545
rect 476426 995533 476432 995585
rect 510256 995533 510262 995585
rect 510314 995573 510320 995585
rect 521392 995573 521398 995585
rect 510314 995545 521398 995573
rect 510314 995533 510320 995545
rect 521392 995533 521398 995545
rect 521450 995533 521456 995585
rect 523792 995533 523798 995585
rect 523850 995573 523856 995585
rect 528976 995573 528982 995585
rect 523850 995545 528982 995573
rect 523850 995533 523856 995545
rect 528976 995533 528982 995545
rect 529034 995533 529040 995585
rect 560176 995533 560182 995585
rect 560234 995573 560240 995585
rect 564496 995573 564502 995585
rect 560234 995545 564502 995573
rect 560234 995533 560240 995545
rect 564496 995533 564502 995545
rect 564554 995533 564560 995585
rect 625648 995533 625654 995585
rect 625706 995573 625712 995585
rect 630160 995573 630166 995585
rect 625706 995545 630166 995573
rect 625706 995533 625712 995545
rect 630160 995533 630166 995545
rect 630218 995533 630224 995585
rect 82288 995459 82294 995511
rect 82346 995499 82352 995511
rect 100720 995499 100726 995511
rect 82346 995471 100726 995499
rect 82346 995459 82352 995471
rect 100720 995459 100726 995471
rect 100778 995459 100784 995511
rect 293680 995459 293686 995511
rect 293738 995499 293744 995511
rect 307600 995499 307606 995511
rect 293738 995471 307606 995499
rect 293738 995459 293744 995471
rect 307600 995459 307606 995471
rect 307658 995459 307664 995511
rect 380080 995459 380086 995511
rect 380138 995499 380144 995511
rect 392368 995499 392374 995511
rect 380138 995471 392374 995499
rect 380138 995459 380144 995471
rect 392368 995459 392374 995471
rect 392426 995459 392432 995511
rect 466192 995459 466198 995511
rect 466250 995499 466256 995511
rect 482704 995499 482710 995511
rect 466250 995471 482710 995499
rect 466250 995459 466256 995471
rect 482704 995459 482710 995471
rect 482762 995459 482768 995511
rect 523600 995459 523606 995511
rect 523658 995499 523664 995511
rect 526096 995499 526102 995511
rect 523658 995471 526102 995499
rect 523658 995459 523664 995471
rect 526096 995459 526102 995471
rect 526154 995459 526160 995511
rect 532240 995499 532246 995511
rect 526210 995471 532246 995499
rect 185104 995385 185110 995437
rect 185162 995425 185168 995437
rect 203632 995425 203638 995437
rect 185162 995397 203638 995425
rect 185162 995385 185168 995397
rect 203632 995385 203638 995397
rect 203690 995385 203696 995437
rect 379792 995385 379798 995437
rect 379850 995425 379856 995437
rect 393712 995425 393718 995437
rect 379850 995397 393718 995425
rect 379850 995385 379856 995397
rect 393712 995385 393718 995397
rect 393770 995385 393776 995437
rect 471856 995385 471862 995437
rect 471914 995425 471920 995437
rect 480976 995425 480982 995437
rect 471914 995397 480982 995425
rect 471914 995385 471920 995397
rect 480976 995385 480982 995397
rect 481034 995385 481040 995437
rect 519184 995385 519190 995437
rect 519242 995425 519248 995437
rect 526210 995425 526238 995471
rect 532240 995459 532246 995471
rect 532298 995459 532304 995511
rect 625552 995459 625558 995511
rect 625610 995499 625616 995511
rect 630928 995499 630934 995511
rect 625610 995471 630934 995499
rect 625610 995459 625616 995471
rect 630928 995459 630934 995471
rect 630986 995459 630992 995511
rect 519242 995397 526238 995425
rect 519242 995385 519248 995397
rect 86320 995311 86326 995363
rect 86378 995351 86384 995363
rect 99760 995351 99766 995363
rect 86378 995323 99766 995351
rect 86378 995311 86384 995323
rect 99760 995311 99766 995323
rect 99818 995311 99824 995363
rect 521296 995311 521302 995363
rect 521354 995351 521360 995363
rect 537376 995351 537382 995363
rect 521354 995323 537382 995351
rect 521354 995311 521360 995323
rect 537376 995311 537382 995323
rect 537434 995311 537440 995363
rect 132112 995237 132118 995289
rect 132170 995277 132176 995289
rect 146800 995277 146806 995289
rect 132170 995249 146806 995277
rect 132170 995237 132176 995249
rect 146800 995237 146806 995249
rect 146858 995237 146864 995289
rect 184144 995237 184150 995289
rect 184202 995277 184208 995289
rect 195760 995277 195766 995289
rect 184202 995249 195766 995277
rect 184202 995237 184208 995249
rect 195760 995237 195766 995249
rect 195818 995237 195824 995289
rect 519088 995237 519094 995289
rect 519146 995277 519152 995289
rect 530560 995277 530566 995289
rect 519146 995249 530566 995277
rect 519146 995237 519152 995249
rect 530560 995237 530566 995249
rect 530618 995277 530624 995289
rect 632368 995277 632374 995289
rect 530618 995249 632374 995277
rect 530618 995237 530624 995249
rect 632368 995237 632374 995249
rect 632426 995237 632432 995289
rect 182992 995163 182998 995215
rect 183050 995203 183056 995215
rect 196816 995203 196822 995215
rect 183050 995175 196822 995203
rect 183050 995163 183056 995175
rect 196816 995163 196822 995175
rect 196874 995163 196880 995215
rect 469456 995163 469462 995215
rect 469514 995203 469520 995215
rect 485968 995203 485974 995215
rect 469514 995175 485974 995203
rect 469514 995163 469520 995175
rect 485968 995163 485974 995175
rect 486026 995163 486032 995215
rect 501808 995163 501814 995215
rect 501866 995203 501872 995215
rect 528208 995203 528214 995215
rect 501866 995175 528214 995203
rect 501866 995163 501872 995175
rect 528208 995163 528214 995175
rect 528266 995163 528272 995215
rect 558928 995163 558934 995215
rect 558986 995203 558992 995215
rect 649360 995203 649366 995215
rect 558986 995175 649366 995203
rect 558986 995163 558992 995175
rect 649360 995163 649366 995175
rect 649418 995163 649424 995215
rect 69136 995089 69142 995141
rect 69194 995129 69200 995141
rect 298384 995129 298390 995141
rect 69194 995101 298390 995129
rect 69194 995089 69200 995101
rect 298384 995089 298390 995101
rect 298442 995089 298448 995141
rect 519952 995089 519958 995141
rect 520010 995129 520016 995141
rect 649744 995129 649750 995141
rect 520010 995101 649750 995129
rect 520010 995089 520016 995101
rect 649744 995089 649750 995101
rect 649802 995089 649808 995141
rect 222928 995015 222934 995067
rect 222986 995055 222992 995067
rect 649648 995055 649654 995067
rect 222986 995027 649654 995055
rect 222986 995015 222992 995027
rect 649648 995015 649654 995027
rect 649706 995015 649712 995067
rect 237424 994941 237430 994993
rect 237482 994981 237488 994993
rect 250480 994981 250486 994993
rect 237482 994953 250486 994981
rect 237482 994941 237488 994953
rect 250480 994941 250486 994953
rect 250538 994941 250544 994993
rect 289264 994793 289270 994845
rect 289322 994833 289328 994845
rect 296656 994833 296662 994845
rect 289322 994805 296662 994833
rect 289322 994793 289328 994805
rect 296656 994793 296662 994805
rect 296714 994793 296720 994845
rect 239440 994053 239446 994105
rect 239498 994093 239504 994105
rect 279280 994093 279286 994105
rect 239498 994065 279286 994093
rect 239498 994053 239504 994065
rect 279280 994053 279286 994065
rect 279338 994053 279344 994105
rect 234928 993905 234934 993957
rect 234986 993945 234992 993957
rect 250384 993945 250390 993957
rect 234986 993917 250390 993945
rect 234986 993905 234992 993917
rect 250384 993905 250390 993917
rect 250442 993905 250448 993957
rect 570736 993905 570742 993957
rect 570794 993945 570800 993957
rect 635248 993945 635254 993957
rect 570794 993917 635254 993945
rect 570794 993905 570800 993917
rect 635248 993905 635254 993917
rect 635306 993905 635312 993957
rect 180496 993831 180502 993883
rect 180554 993871 180560 993883
rect 198640 993871 198646 993883
rect 180554 993843 198646 993871
rect 180554 993831 180560 993843
rect 198640 993831 198646 993843
rect 198698 993831 198704 993883
rect 238672 993831 238678 993883
rect 238730 993871 238736 993883
rect 259024 993871 259030 993883
rect 238730 993843 259030 993871
rect 238730 993831 238736 993843
rect 259024 993831 259030 993843
rect 259082 993831 259088 993883
rect 563248 993831 563254 993883
rect 563306 993871 563312 993883
rect 641008 993871 641014 993883
rect 563306 993843 641014 993871
rect 563306 993831 563312 993843
rect 641008 993831 641014 993843
rect 641066 993831 641072 993883
rect 77680 993757 77686 993809
rect 77738 993797 77744 993809
rect 95056 993797 95062 993809
rect 77738 993769 95062 993797
rect 77738 993757 77744 993769
rect 95056 993757 95062 993769
rect 95114 993757 95120 993809
rect 129328 993757 129334 993809
rect 129386 993797 129392 993809
rect 149584 993797 149590 993809
rect 129386 993769 149590 993797
rect 129386 993757 129392 993769
rect 149584 993757 149590 993769
rect 149642 993757 149648 993809
rect 181360 993757 181366 993809
rect 181418 993797 181424 993809
rect 209776 993797 209782 993809
rect 181418 993769 209782 993797
rect 181418 993757 181424 993769
rect 209776 993757 209782 993769
rect 209834 993757 209840 993809
rect 231472 993757 231478 993809
rect 231530 993797 231536 993809
rect 260080 993797 260086 993809
rect 231530 993769 260086 993797
rect 231530 993757 231536 993769
rect 260080 993757 260086 993769
rect 260138 993757 260144 993809
rect 282832 993757 282838 993809
rect 282890 993797 282896 993809
rect 309904 993797 309910 993809
rect 282890 993769 309910 993797
rect 282890 993757 282896 993769
rect 309904 993757 309910 993769
rect 309962 993757 309968 993809
rect 567376 993757 567382 993809
rect 567434 993797 567440 993809
rect 634864 993797 634870 993809
rect 567434 993769 634870 993797
rect 567434 993757 567440 993769
rect 634864 993757 634870 993769
rect 634922 993757 634928 993809
rect 80176 993683 80182 993735
rect 80234 993723 80240 993735
rect 105328 993723 105334 993735
rect 80234 993695 105334 993723
rect 80234 993683 80240 993695
rect 105328 993683 105334 993695
rect 105386 993683 105392 993735
rect 131824 993683 131830 993735
rect 131882 993723 131888 993735
rect 156592 993723 156598 993735
rect 131882 993695 156598 993723
rect 131882 993683 131888 993695
rect 156592 993683 156598 993695
rect 156650 993683 156656 993735
rect 179824 993683 179830 993735
rect 179882 993723 179888 993735
rect 208720 993723 208726 993735
rect 179882 993695 208726 993723
rect 179882 993683 179888 993695
rect 208720 993683 208726 993695
rect 208778 993683 208784 993735
rect 232528 993683 232534 993735
rect 232586 993723 232592 993735
rect 261040 993723 261046 993735
rect 232586 993695 261046 993723
rect 232586 993683 232592 993695
rect 261040 993683 261046 993695
rect 261098 993683 261104 993735
rect 284368 993683 284374 993735
rect 284426 993723 284432 993735
rect 312784 993723 312790 993735
rect 284426 993695 312790 993723
rect 284426 993683 284432 993695
rect 312784 993683 312790 993695
rect 312842 993683 312848 993735
rect 372496 993683 372502 993735
rect 372554 993723 372560 993735
rect 393040 993723 393046 993735
rect 372554 993695 393046 993723
rect 372554 993683 372560 993695
rect 393040 993683 393046 993695
rect 393098 993683 393104 993735
rect 573040 993683 573046 993735
rect 573098 993723 573104 993735
rect 637360 993723 637366 993735
rect 573098 993695 637366 993723
rect 573098 993683 573104 993695
rect 637360 993683 637366 993695
rect 637418 993683 637424 993735
rect 77296 993609 77302 993661
rect 77354 993649 77360 993661
rect 105904 993649 105910 993661
rect 77354 993621 105910 993649
rect 77354 993609 77360 993621
rect 105904 993609 105910 993621
rect 105962 993609 105968 993661
rect 128464 993609 128470 993661
rect 128522 993649 128528 993661
rect 157264 993649 157270 993661
rect 128522 993621 157270 993649
rect 128522 993609 128528 993621
rect 157264 993609 157270 993621
rect 157322 993609 157328 993661
rect 185392 993609 185398 993661
rect 185450 993649 185456 993661
rect 236752 993649 236758 993661
rect 185450 993621 236758 993649
rect 185450 993609 185456 993621
rect 236752 993609 236758 993621
rect 236810 993649 236816 993661
rect 239440 993649 239446 993661
rect 236810 993621 239446 993649
rect 236810 993609 236816 993621
rect 239440 993609 239446 993621
rect 239498 993609 239504 993661
rect 250480 993609 250486 993661
rect 250538 993649 250544 993661
rect 289264 993649 289270 993661
rect 250538 993621 289270 993649
rect 250538 993609 250544 993621
rect 289264 993609 289270 993621
rect 289322 993609 289328 993661
rect 365776 993609 365782 993661
rect 365834 993649 365840 993661
rect 398800 993649 398806 993661
rect 365834 993621 398806 993649
rect 365834 993609 365840 993621
rect 398800 993609 398806 993621
rect 398858 993609 398864 993661
rect 443536 993609 443542 993661
rect 443594 993649 443600 993661
rect 487792 993649 487798 993661
rect 443594 993621 487798 993649
rect 443594 993609 443600 993621
rect 487792 993609 487798 993621
rect 487850 993609 487856 993661
rect 521392 993609 521398 993661
rect 521450 993649 521456 993661
rect 538960 993649 538966 993661
rect 521450 993621 538966 993649
rect 521450 993609 521456 993621
rect 538960 993609 538966 993621
rect 539018 993609 539024 993661
rect 61840 993535 61846 993587
rect 61898 993575 61904 993587
rect 82576 993575 82582 993587
rect 61898 993547 82582 993575
rect 61898 993535 61904 993547
rect 82576 993535 82582 993547
rect 82634 993575 82640 993587
rect 133936 993575 133942 993587
rect 82634 993547 133942 993575
rect 82634 993535 82640 993547
rect 133936 993535 133942 993547
rect 133994 993575 134000 993587
rect 143824 993575 143830 993587
rect 133994 993547 143830 993575
rect 133994 993535 134000 993547
rect 143824 993535 143830 993547
rect 143882 993535 143888 993587
rect 237424 993535 237430 993587
rect 237482 993575 237488 993587
rect 251344 993575 251350 993587
rect 237482 993547 251350 993575
rect 237482 993535 237488 993547
rect 251344 993535 251350 993547
rect 251402 993535 251408 993587
rect 279280 993535 279286 993587
rect 279338 993575 279344 993587
rect 288112 993575 288118 993587
rect 279338 993547 288118 993575
rect 279338 993535 279344 993547
rect 288112 993535 288118 993547
rect 288170 993575 288176 993587
rect 390160 993575 390166 993587
rect 288170 993547 390166 993575
rect 288170 993535 288176 993547
rect 390160 993535 390166 993547
rect 390218 993575 390224 993587
rect 403120 993575 403126 993587
rect 390218 993547 403126 993575
rect 390218 993535 390224 993547
rect 403120 993535 403126 993547
rect 403178 993535 403184 993587
rect 331216 992573 331222 992625
rect 331274 992613 331280 992625
rect 332560 992613 332566 992625
rect 331274 992585 332566 992613
rect 331274 992573 331280 992585
rect 332560 992573 332566 992585
rect 332618 992573 332624 992625
rect 73378 992141 106622 992169
rect 73378 992107 73406 992141
rect 73360 992055 73366 992107
rect 73418 992055 73424 992107
rect 106594 992095 106622 992141
rect 627682 992141 650078 992169
rect 627682 992107 627710 992141
rect 650050 992107 650078 992141
rect 110128 992095 110134 992107
rect 106594 992067 110134 992095
rect 110128 992055 110134 992067
rect 110186 992055 110192 992107
rect 627664 992055 627670 992107
rect 627722 992055 627728 992107
rect 650032 992055 650038 992107
rect 650090 992055 650096 992107
rect 290896 991759 290902 991811
rect 290954 991799 290960 991811
rect 298960 991799 298966 991811
rect 290954 991771 298966 991799
rect 290954 991759 290960 991771
rect 298960 991759 298966 991771
rect 299018 991759 299024 991811
rect 105808 990501 105814 990553
rect 105866 990541 105872 990553
rect 109552 990541 109558 990553
rect 105866 990513 109558 990541
rect 105866 990501 105872 990513
rect 109552 990501 109558 990513
rect 109610 990501 109616 990553
rect 640528 989909 640534 989961
rect 640586 989949 640592 989961
rect 649840 989949 649846 989961
rect 640586 989921 649846 989949
rect 640586 989909 640592 989921
rect 649840 989909 649846 989921
rect 649898 989909 649904 989961
rect 569872 989539 569878 989591
rect 569930 989579 569936 989591
rect 592432 989579 592438 989591
rect 569930 989551 592438 989579
rect 569930 989539 569936 989551
rect 592432 989539 592438 989551
rect 592490 989539 592496 989591
rect 569968 989465 569974 989517
rect 570026 989505 570032 989517
rect 608752 989505 608758 989517
rect 570026 989477 608758 989505
rect 570026 989465 570032 989477
rect 608752 989465 608758 989477
rect 608810 989465 608816 989517
rect 371632 989391 371638 989443
rect 371690 989431 371696 989443
rect 397840 989431 397846 989443
rect 371690 989403 397846 989431
rect 371690 989391 371696 989403
rect 397840 989391 397846 989403
rect 397898 989391 397904 989443
rect 437776 989391 437782 989443
rect 437834 989431 437840 989443
rect 462736 989431 462742 989443
rect 437834 989403 462742 989431
rect 437834 989391 437840 989403
rect 462736 989391 462742 989403
rect 462794 989391 462800 989443
rect 515632 989391 515638 989443
rect 515690 989431 515696 989443
rect 527632 989431 527638 989443
rect 515690 989403 527638 989431
rect 515690 989391 515696 989403
rect 527632 989391 527638 989403
rect 527690 989391 527696 989443
rect 533680 989391 533686 989443
rect 533738 989431 533744 989443
rect 576304 989431 576310 989443
rect 533738 989403 576310 989431
rect 533738 989391 533744 989403
rect 576304 989391 576310 989403
rect 576362 989391 576368 989443
rect 154480 989317 154486 989369
rect 154538 989357 154544 989369
rect 161680 989357 161686 989369
rect 154538 989329 161686 989357
rect 154538 989317 154544 989329
rect 161680 989317 161686 989329
rect 161738 989317 161744 989369
rect 203152 989317 203158 989369
rect 203210 989357 203216 989369
rect 213328 989357 213334 989369
rect 203210 989329 213334 989357
rect 203210 989317 203216 989329
rect 213328 989317 213334 989329
rect 213386 989317 213392 989369
rect 270736 989317 270742 989369
rect 270794 989357 270800 989369
rect 284272 989357 284278 989369
rect 270794 989329 284278 989357
rect 270794 989317 270800 989329
rect 284272 989317 284278 989329
rect 284330 989317 284336 989369
rect 319600 989317 319606 989369
rect 319658 989357 319664 989369
rect 348496 989357 348502 989369
rect 319658 989329 348502 989357
rect 319658 989317 319664 989329
rect 348496 989317 348502 989329
rect 348554 989317 348560 989369
rect 371536 989317 371542 989369
rect 371594 989357 371600 989369
rect 414064 989357 414070 989369
rect 371594 989329 414070 989357
rect 371594 989317 371600 989329
rect 414064 989317 414070 989329
rect 414122 989317 414128 989369
rect 437872 989317 437878 989369
rect 437930 989357 437936 989369
rect 478960 989357 478966 989369
rect 437930 989329 478966 989357
rect 437930 989317 437936 989329
rect 478960 989317 478966 989329
rect 479018 989317 479024 989369
rect 515536 989317 515542 989369
rect 515594 989357 515600 989369
rect 543760 989357 543766 989369
rect 515594 989329 543766 989357
rect 515594 989317 515600 989329
rect 543760 989317 543766 989329
rect 543818 989317 543824 989369
rect 569776 989317 569782 989369
rect 569834 989357 569840 989369
rect 624976 989357 624982 989369
rect 569834 989329 624982 989357
rect 569834 989317 569840 989329
rect 624976 989317 624982 989329
rect 625034 989317 625040 989369
rect 643312 989317 643318 989369
rect 643370 989357 643376 989369
rect 650128 989357 650134 989369
rect 643370 989329 650134 989357
rect 643370 989317 643376 989329
rect 650128 989317 650134 989329
rect 650186 989317 650192 989369
rect 89584 989243 89590 989295
rect 89642 989283 89648 989295
rect 109360 989283 109366 989295
rect 89642 989255 109366 989283
rect 89642 989243 89648 989255
rect 109360 989243 109366 989255
rect 109418 989243 109424 989295
rect 138256 989243 138262 989295
rect 138314 989283 138320 989295
rect 161488 989283 161494 989295
rect 138314 989255 161494 989283
rect 138314 989243 138320 989255
rect 161488 989243 161494 989255
rect 161546 989243 161552 989295
rect 216016 989243 216022 989295
rect 216074 989283 216080 989295
rect 235600 989283 235606 989295
rect 216074 989255 235606 989283
rect 216074 989243 216080 989255
rect 235600 989243 235606 989255
rect 235658 989243 235664 989295
rect 267952 989243 267958 989295
rect 268010 989283 268016 989295
rect 300496 989283 300502 989295
rect 268010 989255 300502 989283
rect 268010 989243 268016 989255
rect 300496 989243 300502 989255
rect 300554 989243 300560 989295
rect 319696 989243 319702 989295
rect 319754 989283 319760 989295
rect 365392 989283 365398 989295
rect 319754 989255 365398 989283
rect 319754 989243 319760 989255
rect 365392 989243 365398 989255
rect 365450 989243 365456 989295
rect 371728 989243 371734 989295
rect 371786 989283 371792 989295
rect 430288 989283 430294 989295
rect 371786 989255 430294 989283
rect 371786 989243 371792 989255
rect 430288 989243 430294 989255
rect 430346 989243 430352 989295
rect 437968 989243 437974 989295
rect 438026 989283 438032 989295
rect 495184 989283 495190 989295
rect 438026 989255 495190 989283
rect 438026 989243 438032 989255
rect 495184 989243 495190 989255
rect 495242 989243 495248 989295
rect 515728 989243 515734 989295
rect 515786 989283 515792 989295
rect 560080 989283 560086 989295
rect 515786 989255 560086 989283
rect 515786 989243 515792 989255
rect 560080 989243 560086 989255
rect 560138 989243 560144 989295
rect 567280 989243 567286 989295
rect 567338 989283 567344 989295
rect 658096 989283 658102 989295
rect 567338 989255 658102 989283
rect 567338 989243 567344 989255
rect 658096 989243 658102 989255
rect 658154 989243 658160 989295
rect 47632 988281 47638 988333
rect 47690 988321 47696 988333
rect 122032 988321 122038 988333
rect 47690 988293 122038 988321
rect 47690 988281 47696 988293
rect 122032 988281 122038 988293
rect 122090 988281 122096 988333
rect 44752 988207 44758 988259
rect 44810 988247 44816 988259
rect 186928 988247 186934 988259
rect 44810 988219 186934 988247
rect 44810 988207 44816 988219
rect 186928 988207 186934 988219
rect 186986 988207 186992 988259
rect 44848 988133 44854 988185
rect 44906 988173 44912 988185
rect 251824 988173 251830 988185
rect 44906 988145 251830 988173
rect 44906 988133 44912 988145
rect 251824 988133 251830 988145
rect 251882 988133 251888 988185
rect 44944 988059 44950 988111
rect 45002 988099 45008 988111
rect 316720 988099 316726 988111
rect 45002 988071 316726 988099
rect 45002 988059 45008 988071
rect 316720 988059 316726 988071
rect 316778 988059 316784 988111
rect 45040 987985 45046 988037
rect 45098 988025 45104 988037
rect 381616 988025 381622 988037
rect 45098 987997 381622 988025
rect 45098 987985 45104 987997
rect 381616 987985 381622 987997
rect 381674 987985 381680 988037
rect 45136 987911 45142 987963
rect 45194 987951 45200 987963
rect 446512 987951 446518 987963
rect 45194 987923 446518 987951
rect 45194 987911 45200 987923
rect 446512 987911 446518 987923
rect 446570 987911 446576 987963
rect 43120 987837 43126 987889
rect 43178 987877 43184 987889
rect 511408 987877 511414 987889
rect 43178 987849 511414 987877
rect 43178 987837 43184 987849
rect 511408 987837 511414 987849
rect 511466 987837 511472 987889
rect 65104 986727 65110 986779
rect 65162 986767 65168 986779
rect 93520 986767 93526 986779
rect 65162 986739 93526 986767
rect 65162 986727 65168 986739
rect 93520 986727 93526 986739
rect 93578 986727 93584 986779
rect 47536 986653 47542 986705
rect 47594 986693 47600 986705
rect 109168 986693 109174 986705
rect 47594 986665 109174 986693
rect 47594 986653 47600 986665
rect 109168 986653 109174 986665
rect 109226 986653 109232 986705
rect 47728 986579 47734 986631
rect 47786 986619 47792 986631
rect 107920 986619 107926 986631
rect 47786 986591 107926 986619
rect 47786 986579 47792 986591
rect 107920 986579 107926 986591
rect 107978 986579 107984 986631
rect 47440 986505 47446 986557
rect 47498 986545 47504 986557
rect 107536 986545 107542 986557
rect 47498 986517 107542 986545
rect 47498 986505 47504 986517
rect 107536 986505 107542 986517
rect 107594 986505 107600 986557
rect 63280 986431 63286 986483
rect 63338 986471 63344 986483
rect 145360 986471 145366 986483
rect 63338 986443 145366 986471
rect 63338 986431 63344 986443
rect 145360 986431 145366 986443
rect 145418 986431 145424 986483
rect 564496 986431 564502 986483
rect 564554 986471 564560 986483
rect 658000 986471 658006 986483
rect 564554 986443 658006 986471
rect 564554 986431 564560 986443
rect 658000 986431 658006 986443
rect 658058 986431 658064 986483
rect 65200 986357 65206 986409
rect 65258 986397 65264 986409
rect 197200 986397 197206 986409
rect 65258 986369 197206 986397
rect 65258 986357 65264 986369
rect 197200 986357 197206 986369
rect 197258 986357 197264 986409
rect 564592 986357 564598 986409
rect 564650 986397 564656 986409
rect 660880 986397 660886 986409
rect 564650 986369 660886 986397
rect 564650 986357 564656 986369
rect 660880 986357 660886 986369
rect 660938 986357 660944 986409
rect 64912 986135 64918 986187
rect 64970 986175 64976 986187
rect 69040 986175 69046 986187
rect 64970 986147 69046 986175
rect 64970 986135 64976 986147
rect 69040 986135 69046 986147
rect 69098 986135 69104 986187
rect 632368 983693 632374 983745
rect 632426 983733 632432 983745
rect 674512 983733 674518 983745
rect 632426 983705 674518 983733
rect 632426 983693 632432 983705
rect 674512 983693 674518 983705
rect 674570 983693 674576 983745
rect 633040 983619 633046 983671
rect 633098 983659 633104 983671
rect 674128 983659 674134 983671
rect 633098 983631 674134 983659
rect 633098 983619 633104 983631
rect 674128 983619 674134 983631
rect 674186 983619 674192 983671
rect 64816 983545 64822 983597
rect 64874 983585 64880 983597
rect 237424 983585 237430 983597
rect 64874 983557 237430 983585
rect 64874 983545 64880 983557
rect 237424 983545 237430 983557
rect 237482 983545 237488 983597
rect 528208 983545 528214 983597
rect 528266 983585 528272 983597
rect 649552 983585 649558 983597
rect 528266 983557 649558 983585
rect 528266 983545 528272 983557
rect 649552 983545 649558 983557
rect 649610 983545 649616 983597
rect 65008 983471 65014 983523
rect 65066 983511 65072 983523
rect 290800 983511 290806 983523
rect 65066 983483 290806 983511
rect 65066 983471 65072 983483
rect 290800 983471 290806 983483
rect 290858 983471 290864 983523
rect 417520 983471 417526 983523
rect 417578 983511 417584 983523
rect 649456 983511 649462 983523
rect 417578 983483 649462 983511
rect 417578 983471 417584 983483
rect 649456 983471 649462 983483
rect 649514 983471 649520 983523
rect 50512 973481 50518 973533
rect 50570 973521 50576 973533
rect 59440 973521 59446 973533
rect 50570 973493 59446 973521
rect 50570 973481 50576 973493
rect 59440 973481 59446 973493
rect 59498 973481 59504 973533
rect 42160 967265 42166 967317
rect 42218 967305 42224 967317
rect 43120 967305 43126 967317
rect 42218 967277 43126 967305
rect 42218 967265 42224 967277
rect 43120 967265 43126 967277
rect 43178 967265 43184 967317
rect 649648 964749 649654 964801
rect 649706 964789 649712 964801
rect 653776 964789 653782 964801
rect 649706 964761 653782 964789
rect 649706 964749 649712 964761
rect 653776 964749 653782 964761
rect 653834 964749 653840 964801
rect 42160 960975 42166 961027
rect 42218 961015 42224 961027
rect 42448 961015 42454 961027
rect 42218 960987 42454 961015
rect 42218 960975 42224 960987
rect 42448 960975 42454 960987
rect 42506 960975 42512 961027
rect 46096 959051 46102 959103
rect 46154 959091 46160 959103
rect 59536 959091 59542 959103
rect 46154 959063 59542 959091
rect 46154 959051 46160 959063
rect 59536 959051 59542 959063
rect 59594 959051 59600 959103
rect 675184 956979 675190 957031
rect 675242 957019 675248 957031
rect 675472 957019 675478 957031
rect 675242 956991 675478 957019
rect 675242 956979 675248 956991
rect 675472 956979 675478 956991
rect 675530 956979 675536 957031
rect 42064 955203 42070 955255
rect 42122 955243 42128 955255
rect 42832 955243 42838 955255
rect 42122 955215 42838 955243
rect 42122 955203 42128 955215
rect 42832 955203 42838 955215
rect 42890 955203 42896 955255
rect 669520 954685 669526 954737
rect 669578 954725 669584 954737
rect 675376 954725 675382 954737
rect 669578 954697 675382 954725
rect 669578 954685 669584 954697
rect 675376 954685 675382 954697
rect 675434 954685 675440 954737
rect 41776 954611 41782 954663
rect 41834 954611 41840 954663
rect 41794 954441 41822 954611
rect 41776 954389 41782 954441
rect 41834 954389 41840 954441
rect 674128 953945 674134 953997
rect 674186 953985 674192 953997
rect 675472 953985 675478 953997
rect 674186 953957 675478 953985
rect 674186 953945 674192 953957
rect 675472 953945 675478 953957
rect 675530 953945 675536 953997
rect 674032 952021 674038 952073
rect 674090 952061 674096 952073
rect 675472 952061 675478 952073
rect 674090 952033 675478 952061
rect 674090 952021 674096 952033
rect 675472 952021 675478 952033
rect 675530 952021 675536 952073
rect 42544 944621 42550 944673
rect 42602 944661 42608 944673
rect 59536 944661 59542 944673
rect 42602 944633 59542 944661
rect 42602 944621 42608 944633
rect 59536 944621 59542 944633
rect 59594 944621 59600 944673
rect 42544 944177 42550 944229
rect 42602 944217 42608 944229
rect 51856 944217 51862 944229
rect 42602 944189 51862 944217
rect 42602 944177 42608 944189
rect 51856 944177 51862 944189
rect 51914 944177 51920 944229
rect 42544 944029 42550 944081
rect 42602 944069 42608 944081
rect 46096 944069 46102 944081
rect 42602 944041 46102 944069
rect 42602 944029 42608 944041
rect 46096 944029 46102 944041
rect 46154 944029 46160 944081
rect 42544 942993 42550 943045
rect 42602 943033 42608 943045
rect 47536 943033 47542 943045
rect 42602 943005 47542 943033
rect 42602 942993 42608 943005
rect 47536 942993 47542 943005
rect 47594 942993 47600 943045
rect 42544 942845 42550 942897
rect 42602 942885 42608 942897
rect 47728 942885 47734 942897
rect 42602 942857 47734 942885
rect 42602 942845 42608 942857
rect 47728 942845 47734 942857
rect 47786 942845 47792 942897
rect 40336 942327 40342 942379
rect 40394 942367 40400 942379
rect 42544 942367 42550 942379
rect 40394 942339 42550 942367
rect 40394 942327 40400 942339
rect 42544 942327 42550 942339
rect 42602 942327 42608 942379
rect 658096 939515 658102 939567
rect 658154 939555 658160 939567
rect 674416 939555 674422 939567
rect 658154 939527 674422 939555
rect 658154 939515 658160 939527
rect 674416 939515 674422 939527
rect 674474 939515 674480 939567
rect 655312 939367 655318 939419
rect 655370 939407 655376 939419
rect 674512 939407 674518 939419
rect 655370 939379 674518 939407
rect 655370 939367 655376 939379
rect 674512 939367 674518 939379
rect 674570 939367 674576 939419
rect 655216 939219 655222 939271
rect 655274 939259 655280 939271
rect 676816 939259 676822 939271
rect 655274 939231 676822 939259
rect 655274 939219 655280 939231
rect 676816 939219 676822 939231
rect 676874 939219 676880 939271
rect 655120 939071 655126 939123
rect 655178 939111 655184 939123
rect 676912 939111 676918 939123
rect 655178 939083 676918 939111
rect 655178 939071 655184 939083
rect 676912 939071 676918 939083
rect 676970 939071 676976 939123
rect 674128 938923 674134 938975
rect 674186 938963 674192 938975
rect 676912 938963 676918 938975
rect 674186 938935 676918 938963
rect 674186 938923 674192 938935
rect 676912 938923 676918 938935
rect 676970 938923 676976 938975
rect 660880 937961 660886 938013
rect 660938 938001 660944 938013
rect 674416 938001 674422 938013
rect 660938 937973 674422 938001
rect 660938 937961 660944 937973
rect 674416 937961 674422 937973
rect 674474 937961 674480 938013
rect 658000 936259 658006 936311
rect 658058 936299 658064 936311
rect 676816 936299 676822 936311
rect 658058 936271 676822 936299
rect 658058 936259 658064 936271
rect 676816 936259 676822 936271
rect 676874 936259 676880 936311
rect 42544 932115 42550 932167
rect 42602 932155 42608 932167
rect 53200 932155 53206 932167
rect 42602 932127 53206 932155
rect 42602 932115 42608 932127
rect 53200 932115 53206 932127
rect 53258 932115 53264 932167
rect 51856 930487 51862 930539
rect 51914 930527 51920 930539
rect 59536 930527 59542 930539
rect 51914 930499 59542 930527
rect 51914 930487 51920 930499
rect 59536 930487 59542 930499
rect 59594 930487 59600 930539
rect 654448 927453 654454 927505
rect 654506 927493 654512 927505
rect 666736 927493 666742 927505
rect 654506 927465 666742 927493
rect 654506 927453 654512 927465
rect 666736 927453 666742 927465
rect 666794 927453 666800 927505
rect 649648 927379 649654 927431
rect 649706 927419 649712 927431
rect 677008 927419 677014 927431
rect 649706 927391 677014 927419
rect 649706 927379 649712 927391
rect 677008 927379 677014 927391
rect 677066 927379 677072 927431
rect 53392 915835 53398 915887
rect 53450 915875 53456 915887
rect 59536 915875 59542 915887
rect 53450 915847 59542 915875
rect 53450 915835 53456 915847
rect 59536 915835 59542 915847
rect 59594 915835 59600 915887
rect 653968 915835 653974 915887
rect 654026 915875 654032 915887
rect 660976 915875 660982 915887
rect 654026 915847 660982 915875
rect 654026 915835 654032 915847
rect 660976 915835 660982 915847
rect 661034 915835 661040 915887
rect 650224 907103 650230 907155
rect 650282 907143 650288 907155
rect 653776 907143 653782 907155
rect 650282 907115 653782 907143
rect 650282 907103 650288 907115
rect 653776 907103 653782 907115
rect 653834 907103 653840 907155
rect 654448 904365 654454 904417
rect 654506 904405 654512 904417
rect 663952 904405 663958 904417
rect 654506 904377 663958 904405
rect 654506 904365 654512 904377
rect 663952 904365 663958 904377
rect 664010 904365 664016 904417
rect 50320 901479 50326 901531
rect 50378 901519 50384 901531
rect 59536 901519 59542 901531
rect 50378 901491 59542 901519
rect 50378 901479 50384 901491
rect 59536 901479 59542 901491
rect 59594 901479 59600 901531
rect 53488 887123 53494 887175
rect 53546 887163 53552 887175
rect 59536 887163 59542 887175
rect 53546 887135 59542 887163
rect 53546 887123 53552 887135
rect 59536 887123 59542 887135
rect 59594 887123 59600 887175
rect 653968 881277 653974 881329
rect 654026 881317 654032 881329
rect 660880 881317 660886 881329
rect 654026 881289 660886 881317
rect 654026 881277 654032 881289
rect 660880 881277 660886 881289
rect 660938 881277 660944 881329
rect 47536 872619 47542 872671
rect 47594 872659 47600 872671
rect 59536 872659 59542 872671
rect 47594 872631 59542 872659
rect 47594 872619 47600 872631
rect 59536 872619 59542 872631
rect 59594 872619 59600 872671
rect 674608 872619 674614 872671
rect 674666 872659 674672 872671
rect 675376 872659 675382 872671
rect 674666 872631 675382 872659
rect 674666 872619 674672 872631
rect 675376 872619 675382 872631
rect 675434 872619 675440 872671
rect 673360 872101 673366 872153
rect 673418 872141 673424 872153
rect 675472 872141 675478 872153
rect 673418 872113 675478 872141
rect 673418 872101 673424 872113
rect 675472 872101 675478 872113
rect 675530 872101 675536 872153
rect 674224 871657 674230 871709
rect 674282 871697 674288 871709
rect 675088 871697 675094 871709
rect 674282 871669 675094 871697
rect 674282 871657 674288 871669
rect 675088 871657 675094 871669
rect 675146 871697 675152 871709
rect 675376 871697 675382 871709
rect 675146 871669 675382 871697
rect 675146 871657 675152 871669
rect 675376 871657 675382 871669
rect 675434 871657 675440 871709
rect 674896 871435 674902 871487
rect 674954 871475 674960 871487
rect 675184 871475 675190 871487
rect 674954 871447 675190 871475
rect 674954 871435 674960 871447
rect 675184 871435 675190 871447
rect 675242 871475 675248 871487
rect 675376 871475 675382 871487
rect 675242 871447 675382 871475
rect 675242 871435 675248 871447
rect 675376 871435 675382 871447
rect 675434 871435 675440 871487
rect 654448 869807 654454 869859
rect 654506 869847 654512 869859
rect 663760 869847 663766 869859
rect 654506 869819 663766 869847
rect 654506 869807 654512 869819
rect 663760 869807 663766 869819
rect 663818 869807 663824 869859
rect 673264 869141 673270 869193
rect 673322 869181 673328 869193
rect 675472 869181 675478 869193
rect 673322 869153 675478 869181
rect 673322 869141 673328 869153
rect 675472 869141 675478 869153
rect 675530 869141 675536 869193
rect 674320 868327 674326 868379
rect 674378 868367 674384 868379
rect 675376 868367 675382 868379
rect 674378 868339 675382 868367
rect 674378 868327 674384 868339
rect 675376 868327 675382 868339
rect 675434 868327 675440 868379
rect 673168 867809 673174 867861
rect 673226 867849 673232 867861
rect 675376 867849 675382 867861
rect 673226 867821 675382 867849
rect 673226 867809 673232 867821
rect 675376 867809 675382 867821
rect 675434 867809 675440 867861
rect 675088 866477 675094 866529
rect 675146 866517 675152 866529
rect 675376 866517 675382 866529
rect 675146 866489 675382 866517
rect 675146 866477 675152 866489
rect 675376 866477 675382 866489
rect 675434 866477 675440 866529
rect 666640 865293 666646 865345
rect 666698 865333 666704 865345
rect 675376 865333 675382 865345
rect 666698 865305 675382 865333
rect 666698 865293 666704 865305
rect 675376 865293 675382 865305
rect 675434 865293 675440 865345
rect 674512 862925 674518 862977
rect 674570 862965 674576 862977
rect 675376 862965 675382 862977
rect 674570 862937 675382 862965
rect 674570 862925 674576 862937
rect 675376 862925 675382 862937
rect 675434 862925 675440 862977
rect 47440 858263 47446 858315
rect 47498 858303 47504 858315
rect 58576 858303 58582 858315
rect 47498 858275 58582 858303
rect 47498 858263 47504 858275
rect 58576 858263 58582 858275
rect 58634 858263 58640 858315
rect 654160 858263 654166 858315
rect 654218 858303 654224 858315
rect 661072 858303 661078 858315
rect 654218 858275 661078 858303
rect 654218 858263 654224 858275
rect 661072 858263 661078 858275
rect 661130 858263 661136 858315
rect 675088 855747 675094 855799
rect 675146 855787 675152 855799
rect 675472 855787 675478 855799
rect 675146 855759 675478 855787
rect 675146 855747 675152 855759
rect 675472 855747 675478 855759
rect 675530 855747 675536 855799
rect 674896 855599 674902 855651
rect 674954 855639 674960 855651
rect 675568 855639 675574 855651
rect 674954 855611 675574 855639
rect 674954 855599 674960 855611
rect 675568 855599 675574 855611
rect 675626 855599 675632 855651
rect 53296 843833 53302 843885
rect 53354 843873 53360 843885
rect 59536 843873 59542 843885
rect 53354 843845 59542 843873
rect 53354 843833 53360 843845
rect 59536 843833 59542 843845
rect 59594 843833 59600 843885
rect 653968 835175 653974 835227
rect 654026 835215 654032 835227
rect 666832 835215 666838 835227
rect 654026 835187 666838 835215
rect 654026 835175 654032 835187
rect 666832 835175 666838 835187
rect 666890 835175 666896 835227
rect 47728 829477 47734 829529
rect 47786 829517 47792 829529
rect 59536 829517 59542 829529
rect 47786 829489 59542 829517
rect 47786 829477 47792 829489
rect 59536 829477 59542 829489
rect 59594 829477 59600 829529
rect 653968 823705 653974 823757
rect 654026 823745 654032 823757
rect 669904 823745 669910 823757
rect 654026 823717 669910 823745
rect 654026 823705 654032 823717
rect 669904 823705 669910 823717
rect 669962 823705 669968 823757
rect 42544 819265 42550 819317
rect 42602 819305 42608 819317
rect 53488 819305 53494 819317
rect 42602 819277 53494 819305
rect 42602 819265 42608 819277
rect 53488 819265 53494 819277
rect 53546 819265 53552 819317
rect 42832 818525 42838 818577
rect 42890 818565 42896 818577
rect 47536 818565 47542 818577
rect 42890 818537 47542 818565
rect 42890 818525 42896 818537
rect 47536 818525 47542 818537
rect 47594 818525 47600 818577
rect 42544 818229 42550 818281
rect 42602 818269 42608 818281
rect 50320 818269 50326 818281
rect 42602 818241 50326 818269
rect 42602 818229 42608 818241
rect 50320 818229 50326 818241
rect 50378 818229 50384 818281
rect 50416 815047 50422 815099
rect 50474 815087 50480 815099
rect 59536 815087 59542 815099
rect 50474 815059 59542 815087
rect 50474 815047 50480 815059
rect 59536 815047 59542 815059
rect 59594 815047 59600 815099
rect 654448 812161 654454 812213
rect 654506 812201 654512 812213
rect 664048 812201 664054 812213
rect 654506 812173 664054 812201
rect 654506 812161 654512 812173
rect 664048 812161 664054 812173
rect 664106 812161 664112 812213
rect 42544 807425 42550 807477
rect 42602 807465 42608 807477
rect 42832 807465 42838 807477
rect 42602 807437 42838 807465
rect 42602 807425 42608 807437
rect 42832 807425 42838 807437
rect 42890 807425 42896 807477
rect 43120 802541 43126 802593
rect 43178 802581 43184 802593
rect 43408 802581 43414 802593
rect 43178 802553 43414 802581
rect 43178 802541 43184 802553
rect 43408 802541 43414 802553
rect 43466 802541 43472 802593
rect 42064 802393 42070 802445
rect 42122 802433 42128 802445
rect 43120 802433 43126 802445
rect 42122 802405 43126 802433
rect 42122 802393 42128 802405
rect 43120 802393 43126 802405
rect 43178 802393 43184 802445
rect 41968 802023 41974 802075
rect 42026 802063 42032 802075
rect 42448 802063 42454 802075
rect 42026 802035 42454 802063
rect 42026 802023 42032 802035
rect 42448 802023 42454 802035
rect 42506 802023 42512 802075
rect 43312 800617 43318 800669
rect 43370 800657 43376 800669
rect 45136 800657 45142 800669
rect 43370 800629 45142 800657
rect 43370 800617 43376 800629
rect 45136 800617 45142 800629
rect 45194 800617 45200 800669
rect 50320 800617 50326 800669
rect 50378 800657 50384 800669
rect 59536 800657 59542 800669
rect 50378 800629 59542 800657
rect 50378 800617 50384 800629
rect 59536 800617 59542 800629
rect 59594 800617 59600 800669
rect 41872 800173 41878 800225
rect 41930 800173 41936 800225
rect 41890 800003 41918 800173
rect 41872 799951 41878 800003
rect 41930 799951 41936 800003
rect 42832 798323 42838 798375
rect 42890 798323 42896 798375
rect 42928 798323 42934 798375
rect 42986 798323 42992 798375
rect 42160 798101 42166 798153
rect 42218 798141 42224 798153
rect 42850 798141 42878 798323
rect 42218 798113 42878 798141
rect 42218 798101 42224 798113
rect 42736 798027 42742 798079
rect 42794 798067 42800 798079
rect 42946 798067 42974 798323
rect 42794 798039 42974 798067
rect 42794 798027 42800 798039
rect 42064 797287 42070 797339
rect 42122 797327 42128 797339
rect 43312 797327 43318 797339
rect 42122 797299 43318 797327
rect 42122 797287 42128 797299
rect 43312 797287 43318 797299
rect 43370 797287 43376 797339
rect 42160 796251 42166 796303
rect 42218 796291 42224 796303
rect 42736 796291 42742 796303
rect 42218 796263 42742 796291
rect 42218 796251 42224 796263
rect 42736 796251 42742 796263
rect 42794 796251 42800 796303
rect 42160 794993 42166 795045
rect 42218 795033 42224 795045
rect 43024 795033 43030 795045
rect 42218 795005 43030 795033
rect 42218 794993 42224 795005
rect 43024 794993 43030 795005
rect 43082 794993 43088 795045
rect 42160 793143 42166 793195
rect 42218 793183 42224 793195
rect 43120 793183 43126 793195
rect 42218 793155 43126 793183
rect 42218 793143 42224 793155
rect 43120 793143 43126 793155
rect 43178 793143 43184 793195
rect 42160 790627 42166 790679
rect 42218 790667 42224 790679
rect 42736 790667 42742 790679
rect 42218 790639 42742 790667
rect 42218 790627 42224 790639
rect 42736 790627 42742 790639
rect 42794 790627 42800 790679
rect 674704 790553 674710 790605
rect 674762 790593 674768 790605
rect 675472 790593 675478 790605
rect 674762 790565 675478 790593
rect 674762 790553 674768 790565
rect 675472 790553 675478 790565
rect 675530 790553 675536 790605
rect 42160 789887 42166 789939
rect 42218 789927 42224 789939
rect 42832 789927 42838 789939
rect 42218 789899 42838 789927
rect 42218 789887 42224 789899
rect 42832 789887 42838 789899
rect 42890 789887 42896 789939
rect 42160 789443 42166 789495
rect 42218 789483 42224 789495
rect 43408 789483 43414 789495
rect 42218 789455 43414 789483
rect 42218 789443 42224 789455
rect 43408 789443 43414 789455
rect 43466 789443 43472 789495
rect 674992 789221 674998 789273
rect 675050 789261 675056 789273
rect 675568 789261 675574 789273
rect 675050 789233 675574 789261
rect 675050 789221 675056 789233
rect 675568 789221 675574 789233
rect 675626 789221 675632 789273
rect 674224 789147 674230 789199
rect 674282 789187 674288 789199
rect 675088 789187 675094 789199
rect 674282 789159 675094 789187
rect 674282 789147 674288 789159
rect 675088 789147 675094 789159
rect 675146 789147 675152 789199
rect 42160 788777 42166 788829
rect 42218 788817 42224 788829
rect 42448 788817 42454 788829
rect 42218 788789 42454 788817
rect 42218 788777 42224 788789
rect 42448 788777 42454 788789
rect 42506 788777 42512 788829
rect 42160 787001 42166 787053
rect 42218 787041 42224 787053
rect 42928 787041 42934 787053
rect 42218 787013 42934 787041
rect 42218 787001 42224 787013
rect 42928 787001 42934 787013
rect 42986 787001 42992 787053
rect 42160 786409 42166 786461
rect 42218 786449 42224 786461
rect 42736 786449 42742 786461
rect 42218 786421 42742 786449
rect 42218 786409 42224 786421
rect 42736 786409 42742 786421
rect 42794 786409 42800 786461
rect 47536 786261 47542 786313
rect 47594 786301 47600 786313
rect 59536 786301 59542 786313
rect 47594 786273 59542 786301
rect 47594 786261 47600 786273
rect 59536 786261 59542 786273
rect 59594 786261 59600 786313
rect 654064 786261 654070 786313
rect 654122 786301 654128 786313
rect 669712 786301 669718 786313
rect 654122 786273 669718 786301
rect 654122 786261 654128 786273
rect 669712 786261 669718 786273
rect 669770 786261 669776 786313
rect 42064 785595 42070 785647
rect 42122 785635 42128 785647
rect 42832 785635 42838 785647
rect 42122 785607 42838 785635
rect 42122 785595 42128 785607
rect 42832 785595 42838 785607
rect 42890 785595 42896 785647
rect 672304 783449 672310 783501
rect 672362 783489 672368 783501
rect 675376 783489 675382 783501
rect 672362 783461 675382 783489
rect 672362 783449 672368 783461
rect 675376 783449 675382 783461
rect 675434 783449 675440 783501
rect 672880 783079 672886 783131
rect 672938 783119 672944 783131
rect 675088 783119 675094 783131
rect 672938 783091 675094 783119
rect 672938 783079 672944 783091
rect 675088 783079 675094 783091
rect 675146 783119 675152 783131
rect 675472 783119 675478 783131
rect 675146 783091 675478 783119
rect 675146 783079 675152 783091
rect 675472 783079 675478 783091
rect 675530 783079 675536 783131
rect 673456 782931 673462 782983
rect 673514 782971 673520 782983
rect 675376 782971 675382 782983
rect 673514 782943 675382 782971
rect 673514 782931 673520 782943
rect 675376 782931 675382 782943
rect 675434 782931 675440 782983
rect 672496 782487 672502 782539
rect 672554 782527 672560 782539
rect 674992 782527 674998 782539
rect 672554 782499 674998 782527
rect 672554 782487 672560 782499
rect 674992 782487 674998 782499
rect 675050 782527 675056 782539
rect 675472 782527 675478 782539
rect 675050 782499 675478 782527
rect 675050 782487 675056 782499
rect 675472 782487 675478 782499
rect 675530 782487 675536 782539
rect 663856 780489 663862 780541
rect 663914 780529 663920 780541
rect 675088 780529 675094 780541
rect 663914 780501 675094 780529
rect 663914 780489 663920 780501
rect 675088 780489 675094 780501
rect 675146 780489 675152 780541
rect 673072 779749 673078 779801
rect 673130 779789 673136 779801
rect 675376 779789 675382 779801
rect 673130 779761 675382 779789
rect 673130 779749 673136 779761
rect 675376 779749 675382 779761
rect 675434 779749 675440 779801
rect 672208 779305 672214 779357
rect 672266 779345 672272 779357
rect 675472 779345 675478 779357
rect 672266 779317 675478 779345
rect 672266 779305 672272 779317
rect 675472 779305 675478 779317
rect 675530 779305 675536 779357
rect 672976 778565 672982 778617
rect 673034 778605 673040 778617
rect 675376 778605 675382 778617
rect 673034 778577 675382 778605
rect 673034 778565 673040 778577
rect 675376 778565 675382 778577
rect 675434 778565 675440 778617
rect 672688 777603 672694 777655
rect 672746 777643 672752 777655
rect 675472 777643 675478 777655
rect 672746 777615 675478 777643
rect 672746 777603 672752 777615
rect 675472 777603 675478 777615
rect 675530 777603 675536 777655
rect 675088 777011 675094 777063
rect 675146 777051 675152 777063
rect 675376 777051 675382 777063
rect 675146 777023 675382 777051
rect 675146 777011 675152 777023
rect 675376 777011 675382 777023
rect 675434 777011 675440 777063
rect 42736 775901 42742 775953
rect 42794 775941 42800 775953
rect 47728 775941 47734 775953
rect 42794 775913 47734 775941
rect 42794 775901 42800 775913
rect 47728 775901 47734 775913
rect 47786 775901 47792 775953
rect 42736 775309 42742 775361
rect 42794 775349 42800 775361
rect 50416 775349 50422 775361
rect 42794 775321 50422 775349
rect 42794 775309 42800 775321
rect 50416 775309 50422 775321
rect 50474 775309 50480 775361
rect 42736 774791 42742 774843
rect 42794 774831 42800 774843
rect 53296 774831 53302 774843
rect 42794 774803 53302 774831
rect 42794 774791 42800 774803
rect 53296 774791 53302 774803
rect 53354 774791 53360 774843
rect 654064 774717 654070 774769
rect 654122 774757 654128 774769
rect 672400 774757 672406 774769
rect 654122 774729 672406 774757
rect 654122 774717 654128 774729
rect 672400 774717 672406 774729
rect 672458 774717 672464 774769
rect 53488 771831 53494 771883
rect 53546 771871 53552 771883
rect 59536 771871 59542 771883
rect 53546 771843 59542 771871
rect 53546 771831 53552 771843
rect 59536 771831 59542 771843
rect 59594 771831 59600 771883
rect 653968 763247 653974 763299
rect 654026 763287 654032 763299
rect 661168 763287 661174 763299
rect 654026 763259 661174 763287
rect 654026 763247 654032 763259
rect 661168 763247 661174 763259
rect 661226 763247 661232 763299
rect 660976 762877 660982 762929
rect 661034 762917 661040 762929
rect 674416 762917 674422 762929
rect 661034 762889 674422 762917
rect 661034 762877 661040 762889
rect 674416 762877 674422 762889
rect 674474 762877 674480 762929
rect 666736 762285 666742 762337
rect 666794 762325 666800 762337
rect 674416 762325 674422 762337
rect 666794 762297 674422 762325
rect 666794 762285 666800 762297
rect 674416 762285 674422 762297
rect 674474 762285 674480 762337
rect 663952 761989 663958 762041
rect 664010 762029 664016 762041
rect 674608 762029 674614 762041
rect 664010 762001 674614 762029
rect 664010 761989 664016 762001
rect 674608 761989 674614 762001
rect 674666 761989 674672 762041
rect 42832 758585 42838 758637
rect 42890 758625 42896 758637
rect 43024 758625 43030 758637
rect 42890 758597 43030 758625
rect 42890 758585 42896 758597
rect 43024 758585 43030 758597
rect 43082 758585 43088 758637
rect 43024 757623 43030 757675
rect 43082 757663 43088 757675
rect 45040 757663 45046 757675
rect 43082 757635 45046 757663
rect 43082 757623 43088 757635
rect 45040 757623 45046 757635
rect 45098 757623 45104 757675
rect 53680 757475 53686 757527
rect 53738 757515 53744 757527
rect 59536 757515 59542 757527
rect 53738 757487 59542 757515
rect 53738 757475 53744 757487
rect 59536 757475 59542 757487
rect 59594 757475 59600 757527
rect 41584 757327 41590 757379
rect 41642 757367 41648 757379
rect 43504 757367 43510 757379
rect 41642 757339 43510 757367
rect 41642 757327 41648 757339
rect 43504 757327 43510 757339
rect 43562 757327 43568 757379
rect 41680 757253 41686 757305
rect 41738 757293 41744 757305
rect 43408 757293 43414 757305
rect 41738 757265 43414 757293
rect 41738 757253 41744 757265
rect 43408 757253 43414 757265
rect 43466 757253 43472 757305
rect 41872 756957 41878 757009
rect 41930 756957 41936 757009
rect 42064 756957 42070 757009
rect 42122 756997 42128 757009
rect 43312 756997 43318 757009
rect 42122 756969 43318 756997
rect 42122 756957 42128 756969
rect 43312 756957 43318 756969
rect 43370 756957 43376 757009
rect 41890 756787 41918 756957
rect 41872 756735 41878 756787
rect 41930 756735 41936 756787
rect 42832 756661 42838 756713
rect 42890 756701 42896 756713
rect 43216 756701 43222 756713
rect 42890 756673 43222 756701
rect 42890 756661 42896 756673
rect 43216 756661 43222 756673
rect 43274 756661 43280 756713
rect 43024 754219 43030 754271
rect 43082 754219 43088 754271
rect 43042 754185 43070 754219
rect 42178 754157 43070 754185
rect 42178 754123 42206 754157
rect 42160 754071 42166 754123
rect 42218 754071 42224 754123
rect 43024 754071 43030 754123
rect 43082 754111 43088 754123
rect 43216 754111 43222 754123
rect 43082 754083 43222 754111
rect 43082 754071 43088 754083
rect 43216 754071 43222 754083
rect 43274 754071 43280 754123
rect 42064 753035 42070 753087
rect 42122 753075 42128 753087
rect 43120 753075 43126 753087
rect 42122 753047 43126 753075
rect 42122 753035 42128 753047
rect 43120 753035 43126 753047
rect 43178 753035 43184 753087
rect 43120 751817 43126 751829
rect 42946 751789 43126 751817
rect 42946 751755 42974 751789
rect 43120 751777 43126 751789
rect 43178 751777 43184 751829
rect 42928 751703 42934 751755
rect 42986 751703 42992 751755
rect 43408 751629 43414 751681
rect 43466 751669 43472 751681
rect 43696 751669 43702 751681
rect 43466 751641 43702 751669
rect 43466 751629 43472 751641
rect 43696 751629 43702 751641
rect 43754 751629 43760 751681
rect 42064 751111 42070 751163
rect 42122 751151 42128 751163
rect 42928 751151 42934 751163
rect 42122 751123 42934 751151
rect 42122 751111 42128 751123
rect 42928 751111 42934 751123
rect 42986 751111 42992 751163
rect 42160 750371 42166 750423
rect 42218 750411 42224 750423
rect 43024 750411 43030 750423
rect 42218 750383 43030 750411
rect 42218 750371 42224 750383
rect 43024 750371 43030 750383
rect 43082 750371 43088 750423
rect 43024 750223 43030 750275
rect 43082 750263 43088 750275
rect 43504 750263 43510 750275
rect 43082 750235 43510 750263
rect 43082 750223 43088 750235
rect 43504 750223 43510 750235
rect 43562 750223 43568 750275
rect 649744 748817 649750 748869
rect 649802 748857 649808 748869
rect 677008 748857 677014 748869
rect 649802 748829 677014 748857
rect 649802 748817 649808 748829
rect 677008 748817 677014 748829
rect 677066 748817 677072 748869
rect 42160 747263 42166 747315
rect 42218 747303 42224 747315
rect 43120 747303 43126 747315
rect 42218 747275 43126 747303
rect 42218 747263 42224 747275
rect 43120 747263 43126 747275
rect 43178 747263 43184 747315
rect 43024 747007 43030 747019
rect 42178 746979 43030 747007
rect 42178 746945 42206 746979
rect 43024 746967 43030 746979
rect 43082 746967 43088 747019
rect 42160 746893 42166 746945
rect 42218 746893 42224 746945
rect 672880 745931 672886 745983
rect 672938 745971 672944 745983
rect 675088 745971 675094 745983
rect 672938 745943 675094 745971
rect 672938 745931 672944 745943
rect 675088 745931 675094 745943
rect 675146 745931 675152 745983
rect 42160 745635 42166 745687
rect 42218 745675 42224 745687
rect 42928 745675 42934 745687
rect 42218 745647 42934 745675
rect 42218 745635 42224 745647
rect 42928 745635 42934 745647
rect 42986 745635 42992 745687
rect 42448 745487 42454 745539
rect 42506 745527 42512 745539
rect 42928 745527 42934 745539
rect 42506 745499 42934 745527
rect 42506 745487 42512 745499
rect 42928 745487 42934 745499
rect 42986 745487 42992 745539
rect 42160 743785 42166 743837
rect 42218 743825 42224 743837
rect 42928 743825 42934 743837
rect 42218 743797 42934 743825
rect 42218 743785 42224 743797
rect 42928 743785 42934 743797
rect 42986 743785 42992 743837
rect 42064 743193 42070 743245
rect 42122 743233 42128 743245
rect 43120 743233 43126 743245
rect 42122 743205 43126 743233
rect 42122 743193 42128 743205
rect 43120 743193 43126 743205
rect 43178 743193 43184 743245
rect 53584 743045 53590 743097
rect 53642 743085 53648 743097
rect 59536 743085 59542 743097
rect 53642 743057 59542 743085
rect 53642 743045 53648 743057
rect 59536 743045 59542 743057
rect 59594 743045 59600 743097
rect 42160 742601 42166 742653
rect 42218 742641 42224 742653
rect 43024 742641 43030 742653
rect 42218 742613 43030 742641
rect 42218 742601 42224 742613
rect 43024 742601 43030 742613
rect 43082 742601 43088 742653
rect 653968 740159 653974 740211
rect 654026 740199 654032 740211
rect 663952 740199 663958 740211
rect 654026 740171 663958 740199
rect 654026 740159 654032 740171
rect 663952 740159 663958 740171
rect 664010 740159 664016 740211
rect 672496 740159 672502 740211
rect 672554 740199 672560 740211
rect 674704 740199 674710 740211
rect 672554 740171 674710 740199
rect 672554 740159 672560 740171
rect 674704 740159 674710 740171
rect 674762 740159 674768 740211
rect 673168 738087 673174 738139
rect 673226 738127 673232 738139
rect 675088 738127 675094 738139
rect 673226 738099 675094 738127
rect 673226 738087 673232 738099
rect 675088 738087 675094 738099
rect 675146 738127 675152 738139
rect 675472 738127 675478 738139
rect 675146 738099 675478 738127
rect 675146 738087 675152 738099
rect 675472 738087 675478 738099
rect 675530 738087 675536 738139
rect 673360 737865 673366 737917
rect 673418 737905 673424 737917
rect 675376 737905 675382 737917
rect 673418 737877 675382 737905
rect 673418 737865 673424 737877
rect 675376 737865 675382 737877
rect 675434 737865 675440 737917
rect 674704 737643 674710 737695
rect 674762 737683 674768 737695
rect 675376 737683 675382 737695
rect 674762 737655 675382 737683
rect 674762 737643 674768 737655
rect 675376 737643 675382 737655
rect 675434 737643 675440 737695
rect 660976 737273 660982 737325
rect 661034 737313 661040 737325
rect 675088 737313 675094 737325
rect 661034 737285 675094 737313
rect 661034 737273 661040 737285
rect 675088 737273 675094 737285
rect 675146 737273 675152 737325
rect 674608 735423 674614 735475
rect 674666 735463 674672 735475
rect 675472 735463 675478 735475
rect 674666 735435 675478 735463
rect 674666 735423 674672 735435
rect 675472 735423 675478 735435
rect 675530 735423 675536 735475
rect 673264 734757 673270 734809
rect 673322 734797 673328 734809
rect 675376 734797 675382 734809
rect 673322 734769 675382 734797
rect 673322 734757 673328 734769
rect 675376 734757 675382 734769
rect 675434 734757 675440 734809
rect 672784 734387 672790 734439
rect 672842 734427 672848 734439
rect 675376 734427 675382 734439
rect 672842 734399 675382 734427
rect 672842 734387 672848 734399
rect 675376 734387 675382 734399
rect 675434 734387 675440 734439
rect 672880 733573 672886 733625
rect 672938 733613 672944 733625
rect 675472 733613 675478 733625
rect 672938 733585 675478 733613
rect 672938 733573 672944 733585
rect 675472 733573 675478 733585
rect 675530 733573 675536 733625
rect 42832 732685 42838 732737
rect 42890 732725 42896 732737
rect 53488 732725 53494 732737
rect 42890 732697 53494 732725
rect 42890 732685 42896 732697
rect 53488 732685 53494 732697
rect 53546 732685 53552 732737
rect 672592 732315 672598 732367
rect 672650 732355 672656 732367
rect 675472 732355 675478 732367
rect 672650 732327 675478 732355
rect 672650 732315 672656 732327
rect 675472 732315 675478 732327
rect 675530 732315 675536 732367
rect 42832 732093 42838 732145
rect 42890 732133 42896 732145
rect 53680 732133 53686 732145
rect 42890 732105 53686 732133
rect 42890 732093 42896 732105
rect 53680 732093 53686 732105
rect 53738 732093 53744 732145
rect 675088 732019 675094 732071
rect 675146 732059 675152 732071
rect 675376 732059 675382 732071
rect 675146 732031 675382 732059
rect 675146 732019 675152 732031
rect 675376 732019 675382 732031
rect 675434 732019 675440 732071
rect 42832 731797 42838 731849
rect 42890 731837 42896 731849
rect 47536 731837 47542 731849
rect 42890 731809 47542 731837
rect 42890 731797 42896 731809
rect 47536 731797 47542 731809
rect 47594 731797 47600 731849
rect 674608 731501 674614 731553
rect 674666 731541 674672 731553
rect 674800 731541 674806 731553
rect 674666 731513 674806 731541
rect 674666 731501 674672 731513
rect 674800 731501 674806 731513
rect 674858 731501 674864 731553
rect 674512 730465 674518 730517
rect 674570 730505 674576 730517
rect 675472 730505 675478 730517
rect 674570 730477 675478 730505
rect 674570 730465 674576 730477
rect 675472 730465 675478 730477
rect 675530 730465 675536 730517
rect 47536 728615 47542 728667
rect 47594 728655 47600 728667
rect 59536 728655 59542 728667
rect 47594 728627 59542 728655
rect 47594 728615 47600 728627
rect 59536 728615 59542 728627
rect 59594 728615 59600 728667
rect 674032 728615 674038 728667
rect 674090 728655 674096 728667
rect 675472 728655 675478 728667
rect 674090 728627 675478 728655
rect 674090 728615 674096 728627
rect 675472 728615 675478 728627
rect 675530 728615 675536 728667
rect 663760 718033 663766 718085
rect 663818 718073 663824 718085
rect 674608 718073 674614 718085
rect 663818 718045 674614 718073
rect 663818 718033 663824 718045
rect 674608 718033 674614 718045
rect 674666 718033 674672 718085
rect 660880 717589 660886 717641
rect 660938 717629 660944 717641
rect 674608 717629 674614 717641
rect 660938 717601 674614 717629
rect 660938 717589 660944 717601
rect 674608 717589 674614 717601
rect 674666 717589 674672 717641
rect 43120 717219 43126 717271
rect 43178 717259 43184 717271
rect 43792 717259 43798 717271
rect 43178 717231 43798 717259
rect 43178 717219 43184 717231
rect 43792 717219 43798 717231
rect 43850 717219 43856 717271
rect 654256 717145 654262 717197
rect 654314 717185 654320 717197
rect 666928 717185 666934 717197
rect 654314 717157 666934 717185
rect 654314 717145 654320 717157
rect 666928 717145 666934 717157
rect 666986 717145 666992 717197
rect 43120 717071 43126 717123
rect 43178 717111 43184 717123
rect 44944 717111 44950 717123
rect 43178 717083 44950 717111
rect 43178 717071 43184 717083
rect 44944 717071 44950 717083
rect 45002 717071 45008 717123
rect 661072 716997 661078 717049
rect 661130 717037 661136 717049
rect 674608 717037 674614 717049
rect 661130 717009 674614 717037
rect 661130 716997 661136 717009
rect 674608 716997 674614 717009
rect 674666 716997 674672 717049
rect 674608 715665 674614 715717
rect 674666 715705 674672 715717
rect 674800 715705 674806 715717
rect 674666 715677 674806 715705
rect 674666 715665 674672 715677
rect 674800 715665 674806 715677
rect 674858 715665 674864 715717
rect 50416 714259 50422 714311
rect 50474 714299 50480 714311
rect 59536 714299 59542 714311
rect 50474 714271 59542 714299
rect 50474 714259 50480 714271
rect 59536 714259 59542 714271
rect 59594 714259 59600 714311
rect 41488 714185 41494 714237
rect 41546 714225 41552 714237
rect 43504 714225 43510 714237
rect 41546 714197 43510 714225
rect 41546 714185 41552 714197
rect 43504 714185 43510 714197
rect 43562 714185 43568 714237
rect 41584 714111 41590 714163
rect 41642 714151 41648 714163
rect 43600 714151 43606 714163
rect 41642 714123 43606 714151
rect 41642 714111 41648 714123
rect 43600 714111 43606 714123
rect 43658 714111 43664 714163
rect 41680 714037 41686 714089
rect 41738 714077 41744 714089
rect 43408 714077 43414 714089
rect 41738 714049 43414 714077
rect 41738 714037 41744 714049
rect 43408 714037 43414 714049
rect 43466 714037 43472 714089
rect 41872 713815 41878 713867
rect 41930 713815 41936 713867
rect 41968 713815 41974 713867
rect 42026 713855 42032 713867
rect 43216 713855 43222 713867
rect 42026 713827 43222 713855
rect 42026 713815 42032 713827
rect 43216 713815 43222 713827
rect 43274 713815 43280 713867
rect 41890 713571 41918 713815
rect 41872 713519 41878 713571
rect 41930 713519 41936 713571
rect 42064 711669 42070 711721
rect 42122 711709 42128 711721
rect 43312 711709 43318 711721
rect 42122 711681 43318 711709
rect 42122 711669 42128 711681
rect 43312 711669 43318 711681
rect 43370 711669 43376 711721
rect 43216 711595 43222 711647
rect 43274 711595 43280 711647
rect 43408 711635 43414 711647
rect 43330 711607 43414 711635
rect 43120 711373 43126 711425
rect 43178 711413 43184 711425
rect 43234 711413 43262 711595
rect 43330 711425 43358 711607
rect 43408 711595 43414 711607
rect 43466 711595 43472 711647
rect 43178 711385 43262 711413
rect 43178 711373 43184 711385
rect 43312 711373 43318 711425
rect 43370 711373 43376 711425
rect 674320 711299 674326 711351
rect 674378 711339 674384 711351
rect 674512 711339 674518 711351
rect 674378 711311 674518 711339
rect 674378 711299 674384 711311
rect 674512 711299 674518 711311
rect 674570 711299 674576 711351
rect 42160 710855 42166 710907
rect 42218 710895 42224 710907
rect 43408 710895 43414 710907
rect 42218 710867 43414 710895
rect 42218 710855 42224 710867
rect 43408 710855 43414 710867
rect 43466 710855 43472 710907
rect 42160 709893 42166 709945
rect 42218 709933 42224 709945
rect 43120 709933 43126 709945
rect 42218 709905 43126 709933
rect 42218 709893 42224 709905
rect 43120 709893 43126 709905
rect 43178 709893 43184 709945
rect 672304 709893 672310 709945
rect 672362 709933 672368 709945
rect 674608 709933 674614 709945
rect 672362 709905 674614 709933
rect 672362 709893 672368 709905
rect 674608 709893 674614 709905
rect 674666 709893 674672 709945
rect 674416 709301 674422 709353
rect 674474 709341 674480 709353
rect 674608 709341 674614 709353
rect 674474 709313 674614 709341
rect 674474 709301 674480 709313
rect 674608 709301 674614 709313
rect 674666 709301 674672 709353
rect 672688 709153 672694 709205
rect 672746 709193 672752 709205
rect 674416 709193 674422 709205
rect 672746 709165 674422 709193
rect 672746 709153 672752 709165
rect 674416 709153 674422 709165
rect 674474 709153 674480 709205
rect 672208 708635 672214 708687
rect 672266 708675 672272 708687
rect 674416 708675 674422 708687
rect 672266 708647 674422 708675
rect 672266 708635 672272 708647
rect 674416 708635 674422 708647
rect 674474 708635 674480 708687
rect 672976 707007 672982 707059
rect 673034 707047 673040 707059
rect 674416 707047 674422 707059
rect 673034 707019 674422 707047
rect 673034 707007 673040 707019
rect 674416 707007 674422 707019
rect 674474 707007 674480 707059
rect 42160 706711 42166 706763
rect 42218 706751 42224 706763
rect 43792 706751 43798 706763
rect 42218 706723 43798 706751
rect 42218 706711 42224 706723
rect 43792 706711 43798 706723
rect 43850 706711 43856 706763
rect 43216 706563 43222 706615
rect 43274 706563 43280 706615
rect 43234 706393 43262 706563
rect 43216 706341 43222 706393
rect 43274 706341 43280 706393
rect 674704 705601 674710 705653
rect 674762 705641 674768 705653
rect 674992 705641 674998 705653
rect 674762 705613 674998 705641
rect 674762 705601 674768 705613
rect 674992 705601 674998 705613
rect 675050 705601 675056 705653
rect 42160 704269 42166 704321
rect 42218 704309 42224 704321
rect 42736 704309 42742 704321
rect 42218 704281 42742 704309
rect 42218 704269 42224 704281
rect 42736 704269 42742 704281
rect 42794 704269 42800 704321
rect 42736 704121 42742 704173
rect 42794 704161 42800 704173
rect 43600 704161 43606 704173
rect 42794 704133 43606 704161
rect 42794 704121 42800 704133
rect 43600 704121 43606 704133
rect 43658 704121 43664 704173
rect 42064 703677 42070 703729
rect 42122 703717 42128 703729
rect 43024 703717 43030 703729
rect 42122 703689 43030 703717
rect 42122 703677 42128 703689
rect 43024 703677 43030 703689
rect 43082 703677 43088 703729
rect 42160 702863 42166 702915
rect 42218 702903 42224 702915
rect 43120 702903 43126 702915
rect 42218 702875 43126 702903
rect 42218 702863 42224 702875
rect 43120 702863 43126 702875
rect 43178 702863 43184 702915
rect 43120 702715 43126 702767
rect 43178 702755 43184 702767
rect 43504 702755 43510 702767
rect 43178 702727 43510 702755
rect 43178 702715 43184 702727
rect 43504 702715 43510 702727
rect 43562 702715 43568 702767
rect 649840 702715 649846 702767
rect 649898 702755 649904 702767
rect 677008 702755 677014 702767
rect 649898 702727 677014 702755
rect 649898 702715 649904 702727
rect 677008 702715 677014 702727
rect 677066 702715 677072 702767
rect 42160 702271 42166 702323
rect 42218 702311 42224 702323
rect 42736 702311 42742 702323
rect 42218 702283 42742 702311
rect 42218 702271 42224 702283
rect 42736 702271 42742 702283
rect 42794 702271 42800 702323
rect 42064 700421 42070 700473
rect 42122 700461 42128 700473
rect 43120 700461 43126 700473
rect 42122 700433 43126 700461
rect 42122 700421 42128 700433
rect 43120 700421 43126 700433
rect 43178 700421 43184 700473
rect 42160 700051 42166 700103
rect 42218 700091 42224 700103
rect 42448 700091 42454 700103
rect 42218 700063 42454 700091
rect 42218 700051 42224 700063
rect 42448 700051 42454 700063
rect 42506 700051 42512 700103
rect 42448 699829 42454 699881
rect 42506 699869 42512 699881
rect 59536 699869 59542 699881
rect 42506 699841 59542 699869
rect 42506 699829 42512 699841
rect 59536 699829 59542 699841
rect 59594 699829 59600 699881
rect 672688 699829 672694 699881
rect 672746 699869 672752 699881
rect 673168 699869 673174 699881
rect 672746 699841 673174 699869
rect 672746 699829 672752 699841
rect 673168 699829 673174 699841
rect 673226 699829 673232 699881
rect 42160 699163 42166 699215
rect 42218 699203 42224 699215
rect 43024 699203 43030 699215
rect 42218 699175 43030 699203
rect 42218 699163 42224 699175
rect 43024 699163 43030 699175
rect 43082 699163 43088 699215
rect 654448 694057 654454 694109
rect 654506 694097 654512 694109
rect 669808 694097 669814 694109
rect 654506 694069 669814 694097
rect 654506 694057 654512 694069
rect 669808 694057 669814 694069
rect 669866 694057 669872 694109
rect 672688 692947 672694 692999
rect 672746 692987 672752 692999
rect 675472 692987 675478 692999
rect 672746 692959 675478 692987
rect 672746 692947 672752 692959
rect 675472 692947 675478 692959
rect 675530 692947 675536 692999
rect 672304 692873 672310 692925
rect 672362 692913 672368 692925
rect 675376 692913 675382 692925
rect 672362 692885 675382 692913
rect 672362 692873 672368 692885
rect 675376 692873 675382 692885
rect 675434 692873 675440 692925
rect 674608 692651 674614 692703
rect 674666 692691 674672 692703
rect 675376 692691 675382 692703
rect 674666 692663 675382 692691
rect 674666 692651 674672 692663
rect 675376 692651 675382 692663
rect 675434 692651 675440 692703
rect 674800 690653 674806 690705
rect 674858 690693 674864 690705
rect 675472 690693 675478 690705
rect 674858 690665 675478 690693
rect 674858 690653 674864 690665
rect 675472 690653 675478 690665
rect 675530 690653 675536 690705
rect 673072 689765 673078 689817
rect 673130 689805 673136 689817
rect 675376 689805 675382 689817
rect 673130 689777 675382 689805
rect 673130 689765 673136 689777
rect 675376 689765 675382 689777
rect 675434 689765 675440 689817
rect 42832 689469 42838 689521
rect 42890 689509 42896 689521
rect 50416 689509 50422 689521
rect 42890 689481 50422 689509
rect 42890 689469 42896 689481
rect 50416 689469 50422 689481
rect 50474 689469 50480 689521
rect 672976 689321 672982 689373
rect 673034 689361 673040 689373
rect 675376 689361 675382 689373
rect 673034 689333 675382 689361
rect 673034 689321 673040 689333
rect 675376 689321 675382 689333
rect 675434 689321 675440 689373
rect 42448 688581 42454 688633
rect 42506 688621 42512 688633
rect 47536 688621 47542 688633
rect 42506 688593 47542 688621
rect 42506 688581 42512 688593
rect 47536 688581 47542 688593
rect 47594 688581 47600 688633
rect 673168 688581 673174 688633
rect 673226 688621 673232 688633
rect 675472 688621 675478 688633
rect 673226 688593 675478 688621
rect 673226 688581 673232 688593
rect 675472 688581 675478 688593
rect 675530 688581 675536 688633
rect 674704 687323 674710 687375
rect 674762 687363 674768 687375
rect 675472 687363 675478 687375
rect 674762 687335 675478 687363
rect 674762 687323 674768 687335
rect 675472 687323 675478 687335
rect 675530 687323 675536 687375
rect 669616 686213 669622 686265
rect 669674 686253 669680 686265
rect 675376 686253 675382 686265
rect 669674 686225 675382 686253
rect 669674 686213 669680 686225
rect 675376 686213 675382 686225
rect 675434 686213 675440 686265
rect 47536 685473 47542 685525
rect 47594 685513 47600 685525
rect 59536 685513 59542 685525
rect 47594 685485 59542 685513
rect 47594 685473 47600 685485
rect 59536 685473 59542 685485
rect 59594 685473 59600 685525
rect 673936 685473 673942 685525
rect 673994 685513 674000 685525
rect 675472 685513 675478 685525
rect 673994 685485 675478 685513
rect 673994 685473 674000 685485
rect 675472 685473 675478 685485
rect 675530 685473 675536 685525
rect 675472 683623 675478 683675
rect 675530 683623 675536 683675
rect 675490 683379 675518 683623
rect 675472 683327 675478 683379
rect 675530 683327 675536 683379
rect 43408 673855 43414 673907
rect 43466 673895 43472 673907
rect 44848 673895 44854 673907
rect 43466 673867 44854 673895
rect 43466 673855 43472 673867
rect 44848 673855 44854 673867
rect 44906 673855 44912 673907
rect 674704 673041 674710 673093
rect 674762 673081 674768 673093
rect 674992 673081 674998 673093
rect 674762 673053 674998 673081
rect 674762 673041 674768 673053
rect 674992 673041 674998 673053
rect 675050 673041 675056 673093
rect 669904 672893 669910 672945
rect 669962 672933 669968 672945
rect 674704 672933 674710 672945
rect 669962 672905 674710 672933
rect 669962 672893 669968 672905
rect 674704 672893 674710 672905
rect 674762 672893 674768 672945
rect 666832 672301 666838 672353
rect 666890 672341 666896 672353
rect 674704 672341 674710 672353
rect 666890 672313 674710 672341
rect 666890 672301 666896 672313
rect 674704 672301 674710 672313
rect 674762 672301 674768 672353
rect 664048 671857 664054 671909
rect 664106 671897 664112 671909
rect 674704 671897 674710 671909
rect 664106 671869 674710 671897
rect 664106 671857 664112 671869
rect 674704 671857 674710 671869
rect 674762 671857 674768 671909
rect 50416 671043 50422 671095
rect 50474 671083 50480 671095
rect 59536 671083 59542 671095
rect 50474 671055 59542 671083
rect 50474 671043 50480 671055
rect 59536 671043 59542 671055
rect 59594 671043 59600 671095
rect 654448 671043 654454 671095
rect 654506 671083 654512 671095
rect 661072 671083 661078 671095
rect 654506 671055 661078 671083
rect 654506 671043 654512 671055
rect 661072 671043 661078 671055
rect 661130 671043 661136 671095
rect 41680 670969 41686 671021
rect 41738 670969 41744 671021
rect 42160 670969 42166 671021
rect 42218 671009 42224 671021
rect 43696 671009 43702 671021
rect 42218 670981 43702 671009
rect 42218 670969 42224 670981
rect 43696 670969 43702 670981
rect 43754 670969 43760 671021
rect 674320 670969 674326 671021
rect 674378 671009 674384 671021
rect 674704 671009 674710 671021
rect 674378 670981 674710 671009
rect 674378 670969 674384 670981
rect 674704 670969 674710 670981
rect 674762 670969 674768 671021
rect 41698 670935 41726 670969
rect 41698 670907 43550 670935
rect 41488 670821 41494 670873
rect 41546 670861 41552 670873
rect 43408 670861 43414 670873
rect 41546 670833 43414 670861
rect 41546 670821 41552 670833
rect 43408 670821 43414 670833
rect 43466 670821 43472 670873
rect 43522 670799 43550 670907
rect 43504 670747 43510 670799
rect 43562 670747 43568 670799
rect 41968 670599 41974 670651
rect 42026 670599 42032 670651
rect 42064 670599 42070 670651
rect 42122 670639 42128 670651
rect 43120 670639 43126 670651
rect 42122 670611 43126 670639
rect 42122 670599 42128 670611
rect 43120 670599 43126 670611
rect 43178 670599 43184 670651
rect 41986 670355 42014 670599
rect 41968 670303 41974 670355
rect 42026 670303 42032 670355
rect 43024 670229 43030 670281
rect 43082 670269 43088 670281
rect 43312 670269 43318 670281
rect 43082 670241 43318 670269
rect 43082 670229 43088 670241
rect 43312 670229 43318 670241
rect 43370 670229 43376 670281
rect 42448 670081 42454 670133
rect 42506 670121 42512 670133
rect 43024 670121 43030 670133
rect 42506 670093 43030 670121
rect 42506 670081 42512 670093
rect 43024 670081 43030 670093
rect 43082 670081 43088 670133
rect 43024 668897 43030 668949
rect 43082 668897 43088 668949
rect 42160 668527 42166 668579
rect 42218 668567 42224 668579
rect 43042 668567 43070 668897
rect 42218 668539 43070 668567
rect 42218 668527 42224 668539
rect 42832 668453 42838 668505
rect 42890 668493 42896 668505
rect 43312 668493 43318 668505
rect 42890 668465 43318 668493
rect 42890 668453 42896 668465
rect 43312 668453 43318 668465
rect 43370 668453 43376 668505
rect 42160 667861 42166 667913
rect 42218 667901 42224 667913
rect 43600 667901 43606 667913
rect 42218 667873 43606 667901
rect 42218 667861 42224 667873
rect 43600 667861 43606 667873
rect 43658 667861 43664 667913
rect 42160 666677 42166 666729
rect 42218 666717 42224 666729
rect 42832 666717 42838 666729
rect 42218 666689 42838 666717
rect 42218 666677 42224 666689
rect 42832 666677 42838 666689
rect 42890 666677 42896 666729
rect 42832 666529 42838 666581
rect 42890 666569 42896 666581
rect 43408 666569 43414 666581
rect 42890 666541 43414 666569
rect 42890 666529 42896 666541
rect 43408 666529 43414 666541
rect 43466 666529 43472 666581
rect 42160 665345 42166 665397
rect 42218 665385 42224 665397
rect 43120 665385 43126 665397
rect 42218 665357 43126 665385
rect 42218 665345 42224 665357
rect 43120 665345 43126 665357
rect 43178 665345 43184 665397
rect 43120 665197 43126 665249
rect 43178 665237 43184 665249
rect 43504 665237 43510 665249
rect 43178 665209 43510 665237
rect 43178 665197 43184 665209
rect 43504 665197 43510 665209
rect 43562 665197 43568 665249
rect 672784 665197 672790 665249
rect 672842 665237 672848 665249
rect 673840 665237 673846 665249
rect 672842 665209 673846 665237
rect 672842 665197 672848 665209
rect 673840 665197 673846 665209
rect 673898 665197 673904 665249
rect 672592 664161 672598 664213
rect 672650 664201 672656 664213
rect 674704 664201 674710 664213
rect 672650 664173 674710 664201
rect 672650 664161 672656 664173
rect 674704 664161 674710 664173
rect 674762 664161 674768 664213
rect 42736 663495 42742 663547
rect 42794 663495 42800 663547
rect 42754 663461 42782 663495
rect 42562 663433 42782 663461
rect 42160 663347 42166 663399
rect 42218 663387 42224 663399
rect 42562 663387 42590 663433
rect 42218 663359 42590 663387
rect 42218 663347 42224 663359
rect 42736 663347 42742 663399
rect 42794 663387 42800 663399
rect 43696 663387 43702 663399
rect 42794 663359 43702 663387
rect 42794 663347 42800 663359
rect 43696 663347 43702 663359
rect 43754 663347 43760 663399
rect 672880 662311 672886 662363
rect 672938 662351 672944 662363
rect 673840 662351 673846 662363
rect 672938 662323 673846 662351
rect 672938 662311 672944 662323
rect 673840 662311 673846 662323
rect 673898 662311 673904 662363
rect 42064 661053 42070 661105
rect 42122 661093 42128 661105
rect 42832 661093 42838 661105
rect 42122 661065 42838 661093
rect 42122 661053 42128 661065
rect 42832 661053 42838 661065
rect 42890 661053 42896 661105
rect 42160 659869 42166 659921
rect 42218 659909 42224 659921
rect 42736 659909 42742 659921
rect 42218 659881 42742 659909
rect 42218 659869 42224 659881
rect 42736 659869 42742 659881
rect 42794 659869 42800 659921
rect 650032 659499 650038 659551
rect 650090 659539 650096 659551
rect 674704 659539 674710 659551
rect 650090 659511 674710 659539
rect 650090 659499 650096 659511
rect 674704 659499 674710 659511
rect 674762 659499 674768 659551
rect 42160 659203 42166 659255
rect 42218 659243 42224 659255
rect 43120 659243 43126 659255
rect 42218 659215 43126 659243
rect 42218 659203 42224 659215
rect 43120 659203 43126 659215
rect 43178 659203 43184 659255
rect 674416 658463 674422 658515
rect 674474 658503 674480 658515
rect 675472 658503 675478 658515
rect 674474 658475 675478 658503
rect 674474 658463 674480 658475
rect 675472 658463 675478 658475
rect 675530 658463 675536 658515
rect 42064 657353 42070 657405
rect 42122 657393 42128 657405
rect 42448 657393 42454 657405
rect 42122 657365 42454 657393
rect 42122 657353 42128 657365
rect 42448 657353 42454 657365
rect 42506 657353 42512 657405
rect 42928 656687 42934 656739
rect 42986 656727 42992 656739
rect 59536 656727 59542 656739
rect 42986 656699 59542 656727
rect 42986 656687 42992 656699
rect 59536 656687 59542 656699
rect 59594 656687 59600 656739
rect 42160 656613 42166 656665
rect 42218 656653 42224 656665
rect 43120 656653 43126 656665
rect 42218 656625 43126 656653
rect 42218 656613 42224 656625
rect 43120 656613 43126 656625
rect 43178 656613 43184 656665
rect 672688 653727 672694 653779
rect 672746 653767 672752 653779
rect 674512 653767 674518 653779
rect 672746 653739 674518 653767
rect 672746 653727 672752 653739
rect 674512 653727 674518 653739
rect 674570 653727 674576 653779
rect 673264 648251 673270 648303
rect 673322 648291 673328 648303
rect 675376 648291 675382 648303
rect 673322 648263 675382 648291
rect 673322 648251 673328 648263
rect 675376 648251 675382 648263
rect 675434 648251 675440 648303
rect 654256 648029 654262 648081
rect 654314 648069 654320 648081
rect 664048 648069 664054 648081
rect 654314 648041 664054 648069
rect 654314 648029 654320 648041
rect 664048 648029 664054 648041
rect 664106 648029 664112 648081
rect 673744 648029 673750 648081
rect 673802 648069 673808 648081
rect 675376 648069 675382 648081
rect 673802 648041 675382 648069
rect 673802 648029 673808 648041
rect 675376 648029 675382 648041
rect 675434 648029 675440 648081
rect 673360 647067 673366 647119
rect 673418 647107 673424 647119
rect 674512 647107 674518 647119
rect 673418 647079 674518 647107
rect 673418 647067 673424 647079
rect 674512 647067 674518 647079
rect 674570 647107 674576 647119
rect 675376 647107 675382 647119
rect 674570 647079 675382 647107
rect 674570 647067 674576 647079
rect 675376 647067 675382 647079
rect 675434 647067 675440 647119
rect 675376 646401 675382 646453
rect 675434 646401 675440 646453
rect 674800 646327 674806 646379
rect 674858 646367 674864 646379
rect 675394 646367 675422 646401
rect 674858 646339 675422 646367
rect 674858 646327 674864 646339
rect 674512 645883 674518 645935
rect 674570 645923 674576 645935
rect 674992 645923 674998 645935
rect 674570 645895 674998 645923
rect 674570 645883 674576 645895
rect 674992 645883 674998 645895
rect 675050 645883 675056 645935
rect 42928 645217 42934 645269
rect 42986 645257 42992 645269
rect 50416 645257 50422 645269
rect 42986 645229 50422 645257
rect 42986 645217 42992 645229
rect 50416 645217 50422 645229
rect 50474 645217 50480 645269
rect 42448 645069 42454 645121
rect 42506 645109 42512 645121
rect 59536 645109 59542 645121
rect 42506 645081 59542 645109
rect 42506 645069 42512 645081
rect 59536 645069 59542 645081
rect 59594 645069 59600 645121
rect 672784 644551 672790 644603
rect 672842 644591 672848 644603
rect 675472 644591 675478 644603
rect 672842 644563 675478 644591
rect 672842 644551 672848 644563
rect 675472 644551 675478 644563
rect 675530 644551 675536 644603
rect 672496 644033 672502 644085
rect 672554 644073 672560 644085
rect 675472 644073 675478 644085
rect 672554 644045 675478 644073
rect 672554 644033 672560 644045
rect 675472 644033 675478 644045
rect 675530 644033 675536 644085
rect 672880 643367 672886 643419
rect 672938 643407 672944 643419
rect 675376 643407 675382 643419
rect 672938 643379 675382 643407
rect 672938 643367 672944 643379
rect 675376 643367 675382 643379
rect 675434 643367 675440 643419
rect 672688 642257 672694 642309
rect 672746 642297 672752 642309
rect 675472 642297 675478 642309
rect 672746 642269 675478 642297
rect 672746 642257 672752 642269
rect 675472 642257 675478 642269
rect 675530 642257 675536 642309
rect 673936 642109 673942 642161
rect 673994 642149 674000 642161
rect 674128 642149 674134 642161
rect 673994 642121 674134 642149
rect 673994 642109 674000 642121
rect 674128 642109 674134 642121
rect 674186 642109 674192 642161
rect 666736 641073 666742 641125
rect 666794 641113 666800 641125
rect 675472 641113 675478 641125
rect 666794 641085 675478 641113
rect 666794 641073 666800 641085
rect 675472 641073 675478 641085
rect 675530 641073 675536 641125
rect 674800 638187 674806 638239
rect 674858 638227 674864 638239
rect 675472 638227 675478 638239
rect 674858 638199 675478 638227
rect 674858 638187 674864 638199
rect 675472 638187 675478 638199
rect 675530 638187 675536 638239
rect 43120 627975 43126 628027
rect 43178 628015 43184 628027
rect 43696 628015 43702 628027
rect 43178 627987 43702 628015
rect 43178 627975 43184 627987
rect 43696 627975 43702 627987
rect 43754 627975 43760 628027
rect 43504 627901 43510 627953
rect 43562 627941 43568 627953
rect 44752 627941 44758 627953
rect 43562 627913 44758 627941
rect 43562 627901 43568 627913
rect 44752 627901 44758 627913
rect 44810 627901 44816 627953
rect 43024 627827 43030 627879
rect 43082 627867 43088 627879
rect 43408 627867 43414 627879
rect 43082 627839 43414 627867
rect 43082 627827 43088 627839
rect 43408 627827 43414 627839
rect 43466 627827 43472 627879
rect 50416 627827 50422 627879
rect 50474 627867 50480 627879
rect 59536 627867 59542 627879
rect 50474 627839 59542 627867
rect 50474 627827 50480 627839
rect 59536 627827 59542 627839
rect 59594 627827 59600 627879
rect 674416 627827 674422 627879
rect 674474 627867 674480 627879
rect 675088 627867 675094 627879
rect 674474 627839 675094 627867
rect 674474 627827 674480 627839
rect 675088 627827 675094 627839
rect 675146 627827 675152 627879
rect 41680 627679 41686 627731
rect 41738 627719 41744 627731
rect 43024 627719 43030 627731
rect 41738 627691 43030 627719
rect 41738 627679 41744 627691
rect 43024 627679 43030 627691
rect 43082 627679 43088 627731
rect 672400 627679 672406 627731
rect 672458 627719 672464 627731
rect 674416 627719 674422 627731
rect 672458 627691 674422 627719
rect 672458 627679 672464 627691
rect 674416 627679 674422 627691
rect 674474 627679 674480 627731
rect 42160 627605 42166 627657
rect 42218 627645 42224 627657
rect 43120 627645 43126 627657
rect 42218 627617 43126 627645
rect 42218 627605 42224 627617
rect 43120 627605 43126 627617
rect 43178 627605 43184 627657
rect 41872 627383 41878 627435
rect 41930 627383 41936 627435
rect 42064 627383 42070 627435
rect 42122 627423 42128 627435
rect 43120 627423 43126 627435
rect 42122 627395 43126 627423
rect 42122 627383 42128 627395
rect 43120 627383 43126 627395
rect 43178 627383 43184 627435
rect 41890 627213 41918 627383
rect 669712 627309 669718 627361
rect 669770 627349 669776 627361
rect 674896 627349 674902 627361
rect 669770 627321 674902 627349
rect 669770 627309 669776 627321
rect 674896 627309 674902 627321
rect 674954 627309 674960 627361
rect 41872 627161 41878 627213
rect 41930 627161 41936 627213
rect 661168 626569 661174 626621
rect 661226 626609 661232 626621
rect 674416 626609 674422 626621
rect 661226 626581 674422 626609
rect 661226 626569 661232 626581
rect 674416 626569 674422 626581
rect 674474 626569 674480 626621
rect 670960 625459 670966 625511
rect 671018 625499 671024 625511
rect 674416 625499 674422 625511
rect 671018 625471 674422 625499
rect 671018 625459 671024 625471
rect 674416 625459 674422 625471
rect 674474 625459 674480 625511
rect 42160 625311 42166 625363
rect 42218 625351 42224 625363
rect 42928 625351 42934 625363
rect 42218 625323 42934 625351
rect 42218 625311 42224 625323
rect 42928 625311 42934 625323
rect 42986 625311 42992 625363
rect 42928 625163 42934 625215
rect 42986 625203 42992 625215
rect 43216 625203 43222 625215
rect 42986 625175 43222 625203
rect 42986 625163 42992 625175
rect 43216 625163 43222 625175
rect 43274 625163 43280 625215
rect 42160 624645 42166 624697
rect 42218 624685 42224 624697
rect 43504 624685 43510 624697
rect 42218 624657 43510 624685
rect 42218 624645 42224 624657
rect 43504 624645 43510 624657
rect 43562 624645 43568 624697
rect 42160 622203 42166 622255
rect 42218 622243 42224 622255
rect 43408 622243 43414 622255
rect 42218 622215 43414 622243
rect 42218 622203 42224 622215
rect 43408 622203 43414 622215
rect 43466 622203 43472 622255
rect 654352 622203 654358 622255
rect 654410 622243 654416 622255
rect 672592 622243 672598 622255
rect 654410 622215 672598 622243
rect 654410 622203 654416 622215
rect 672592 622203 672598 622215
rect 672650 622203 672656 622255
rect 671920 622129 671926 622181
rect 671978 622169 671984 622181
rect 676912 622169 676918 622181
rect 671978 622141 676918 622169
rect 671978 622129 671984 622141
rect 676912 622129 676918 622141
rect 676970 622129 676976 622181
rect 672016 622055 672022 622107
rect 672074 622095 672080 622107
rect 676816 622095 676822 622107
rect 672074 622067 676822 622095
rect 672074 622055 672080 622067
rect 676816 622055 676822 622067
rect 676874 622055 676880 622107
rect 42160 621611 42166 621663
rect 42218 621651 42224 621663
rect 43120 621651 43126 621663
rect 42218 621623 43126 621651
rect 42218 621611 42224 621623
rect 43120 621611 43126 621623
rect 43178 621611 43184 621663
rect 42064 620871 42070 620923
rect 42122 620911 42128 620923
rect 42928 620911 42934 620923
rect 42122 620883 42934 620911
rect 42122 620871 42128 620883
rect 42928 620871 42934 620883
rect 42986 620871 42992 620923
rect 42160 620353 42166 620405
rect 42218 620393 42224 620405
rect 43024 620393 43030 620405
rect 42218 620365 43030 620393
rect 42218 620353 42224 620365
rect 43024 620353 43030 620365
rect 43082 620353 43088 620405
rect 672976 618429 672982 618481
rect 673034 618469 673040 618481
rect 674416 618469 674422 618481
rect 673034 618441 674422 618469
rect 673034 618429 673040 618441
rect 674416 618429 674422 618441
rect 674474 618429 674480 618481
rect 672304 617837 672310 617889
rect 672362 617877 672368 617889
rect 674416 617877 674422 617889
rect 672362 617849 674422 617877
rect 672362 617837 672368 617849
rect 674416 617837 674422 617849
rect 674474 617837 674480 617889
rect 673072 617541 673078 617593
rect 673130 617581 673136 617593
rect 674704 617581 674710 617593
rect 673130 617553 674710 617581
rect 673130 617541 673136 617553
rect 674704 617541 674710 617553
rect 674762 617541 674768 617593
rect 42160 617171 42166 617223
rect 42218 617211 42224 617223
rect 43696 617211 43702 617223
rect 42218 617183 43702 617211
rect 42218 617171 42224 617183
rect 43696 617171 43702 617183
rect 43754 617171 43760 617223
rect 42160 615987 42166 616039
rect 42218 616027 42224 616039
rect 42448 616027 42454 616039
rect 42218 615999 42454 616027
rect 42218 615987 42224 615999
rect 42448 615987 42454 615999
rect 42506 615987 42512 616039
rect 42160 614137 42166 614189
rect 42218 614177 42224 614189
rect 43120 614177 43126 614189
rect 42218 614149 43126 614177
rect 42218 614137 42224 614149
rect 43120 614137 43126 614149
rect 43178 614137 43184 614189
rect 42832 613471 42838 613523
rect 42890 613511 42896 613523
rect 59536 613511 59542 613523
rect 42890 613483 59542 613511
rect 42890 613471 42896 613483
rect 59536 613471 59542 613483
rect 59594 613471 59600 613523
rect 649936 613471 649942 613523
rect 649994 613511 650000 613523
rect 677104 613511 677110 613523
rect 649994 613483 677110 613511
rect 649994 613471 650000 613483
rect 677104 613471 677110 613483
rect 677162 613471 677168 613523
rect 654352 613397 654358 613449
rect 654410 613437 654416 613449
rect 669520 613437 669526 613449
rect 654410 613409 669526 613437
rect 654410 613397 654416 613409
rect 669520 613397 669526 613409
rect 669578 613397 669584 613449
rect 673360 613397 673366 613449
rect 673418 613437 673424 613449
rect 674992 613437 674998 613449
rect 673418 613409 674998 613437
rect 673418 613397 673424 613409
rect 674992 613397 674998 613409
rect 675050 613397 675056 613449
rect 675088 612139 675094 612191
rect 675146 612179 675152 612191
rect 675472 612179 675478 612191
rect 675146 612151 675478 612179
rect 675146 612139 675152 612151
rect 675472 612139 675478 612151
rect 675530 612139 675536 612191
rect 671824 604073 671830 604125
rect 671882 604113 671888 604125
rect 675472 604113 675478 604125
rect 671882 604085 675478 604113
rect 671882 604073 671888 604085
rect 675472 604073 675478 604085
rect 675530 604073 675536 604125
rect 673552 603259 673558 603311
rect 673610 603299 673616 603311
rect 675376 603299 675382 603311
rect 673610 603271 675382 603299
rect 673610 603259 673616 603271
rect 675376 603259 675382 603271
rect 675434 603259 675440 603311
rect 42160 603111 42166 603163
rect 42218 603151 42224 603163
rect 42832 603151 42838 603163
rect 42218 603123 42838 603151
rect 42218 603111 42224 603123
rect 42832 603111 42838 603123
rect 42890 603111 42896 603163
rect 672112 602815 672118 602867
rect 672170 602855 672176 602867
rect 674992 602855 674998 602867
rect 672170 602827 674998 602855
rect 672170 602815 672176 602827
rect 674992 602815 674998 602827
rect 675050 602855 675056 602867
rect 675472 602855 675478 602867
rect 675050 602827 675478 602855
rect 675050 602815 675056 602827
rect 675472 602815 675478 602827
rect 675530 602815 675536 602867
rect 673360 602667 673366 602719
rect 673418 602707 673424 602719
rect 675376 602707 675382 602719
rect 673418 602679 675382 602707
rect 673418 602667 673424 602679
rect 675376 602667 675382 602679
rect 675434 602667 675440 602719
rect 672304 602445 672310 602497
rect 672362 602485 672368 602497
rect 675088 602485 675094 602497
rect 672362 602457 675094 602485
rect 672362 602445 672368 602457
rect 675088 602445 675094 602457
rect 675146 602485 675152 602497
rect 675376 602485 675382 602497
rect 675146 602457 675382 602485
rect 675146 602445 675152 602457
rect 675376 602445 675382 602457
rect 675434 602445 675440 602497
rect 42736 602223 42742 602275
rect 42794 602263 42800 602275
rect 51856 602263 51862 602275
rect 42794 602235 51862 602263
rect 42794 602223 42800 602235
rect 51856 602223 51862 602235
rect 51914 602223 51920 602275
rect 663760 601927 663766 601979
rect 663818 601967 663824 601979
rect 674416 601967 674422 601979
rect 663818 601939 674422 601967
rect 663818 601927 663824 601939
rect 674416 601927 674422 601939
rect 674474 601927 674480 601979
rect 42832 601853 42838 601905
rect 42890 601893 42896 601905
rect 59536 601893 59542 601905
rect 42890 601865 59542 601893
rect 42890 601853 42896 601865
rect 59536 601853 59542 601865
rect 59594 601853 59600 601905
rect 673072 599781 673078 599833
rect 673130 599821 673136 599833
rect 675376 599821 675382 599833
rect 673130 599793 675382 599821
rect 673130 599781 673136 599793
rect 675376 599781 675382 599793
rect 675434 599781 675440 599833
rect 672976 599263 672982 599315
rect 673034 599303 673040 599315
rect 675376 599303 675382 599315
rect 673034 599275 675382 599303
rect 673034 599263 673040 599275
rect 675376 599263 675382 599275
rect 675434 599263 675440 599315
rect 654448 599041 654454 599093
rect 654506 599081 654512 599093
rect 672400 599081 672406 599093
rect 654506 599053 672406 599081
rect 654506 599041 654512 599053
rect 672400 599041 672406 599053
rect 672458 599041 672464 599093
rect 673168 598375 673174 598427
rect 673226 598415 673232 598427
rect 675472 598415 675478 598427
rect 673226 598387 675478 598415
rect 673226 598375 673232 598387
rect 675472 598375 675478 598387
rect 675530 598375 675536 598427
rect 672208 597117 672214 597169
rect 672266 597157 672272 597169
rect 675472 597157 675478 597169
rect 672266 597129 675478 597157
rect 672266 597117 672272 597129
rect 675472 597117 675478 597129
rect 675530 597117 675536 597169
rect 674416 596821 674422 596873
rect 674474 596861 674480 596873
rect 675376 596861 675382 596873
rect 674474 596833 675382 596861
rect 674474 596821 674480 596833
rect 675376 596821 675382 596833
rect 675434 596821 675440 596873
rect 654448 587497 654454 587549
rect 654506 587537 654512 587549
rect 666832 587537 666838 587549
rect 654506 587509 666838 587537
rect 654506 587497 654512 587509
rect 666832 587497 666838 587509
rect 666890 587497 666896 587549
rect 671920 587497 671926 587549
rect 671978 587537 671984 587549
rect 676816 587537 676822 587549
rect 671978 587509 676822 587537
rect 671978 587497 671984 587509
rect 676816 587497 676822 587509
rect 676874 587497 676880 587549
rect 51856 585943 51862 585995
rect 51914 585983 51920 585995
rect 59536 585983 59542 585995
rect 51914 585955 59542 585983
rect 51914 585943 51920 585955
rect 59536 585943 59542 585955
rect 59594 585943 59600 585995
rect 43120 584685 43126 584737
rect 43178 584725 43184 584737
rect 47632 584725 47638 584737
rect 43178 584697 47638 584725
rect 43178 584685 43184 584697
rect 47632 584685 47638 584697
rect 47690 584685 47696 584737
rect 41488 584463 41494 584515
rect 41546 584503 41552 584515
rect 43216 584503 43222 584515
rect 41546 584475 43222 584503
rect 41546 584463 41552 584475
rect 43216 584463 43222 584475
rect 43274 584463 43280 584515
rect 41776 584241 41782 584293
rect 41834 584281 41840 584293
rect 43408 584281 43414 584293
rect 41834 584253 43414 584281
rect 41834 584241 41840 584253
rect 43408 584241 43414 584253
rect 43466 584241 43472 584293
rect 41872 584167 41878 584219
rect 41930 584167 41936 584219
rect 41890 583997 41918 584167
rect 41872 583945 41878 583997
rect 41930 583945 41936 583997
rect 42832 583797 42838 583849
rect 42890 583837 42896 583849
rect 43312 583837 43318 583849
rect 42890 583809 43318 583837
rect 42890 583797 42896 583809
rect 43312 583797 43318 583809
rect 43370 583797 43376 583849
rect 663952 582021 663958 582073
rect 664010 582061 664016 582073
rect 674416 582061 674422 582073
rect 664010 582033 674422 582061
rect 664010 582021 664016 582033
rect 674416 582021 674422 582033
rect 674474 582021 674480 582073
rect 655216 581947 655222 581999
rect 655274 581987 655280 581999
rect 674608 581987 674614 581999
rect 655274 581959 674614 581987
rect 655274 581947 655280 581959
rect 674608 581947 674614 581959
rect 674666 581947 674672 581999
rect 666928 581577 666934 581629
rect 666986 581617 666992 581629
rect 674608 581617 674614 581629
rect 666986 581589 674614 581617
rect 666986 581577 666992 581589
rect 674608 581577 674614 581589
rect 674666 581577 674672 581629
rect 43024 581503 43030 581555
rect 43082 581543 43088 581555
rect 43312 581543 43318 581555
rect 43082 581515 43318 581543
rect 43082 581503 43088 581515
rect 43312 581503 43318 581515
rect 43370 581503 43376 581555
rect 42064 581429 42070 581481
rect 42122 581469 42128 581481
rect 43120 581469 43126 581481
rect 42122 581441 43126 581469
rect 42122 581429 42128 581441
rect 43120 581429 43126 581441
rect 43178 581429 43184 581481
rect 670960 580837 670966 580889
rect 671018 580877 671024 580889
rect 674416 580877 674422 580889
rect 671018 580849 674422 580877
rect 671018 580837 671024 580849
rect 674416 580837 674422 580849
rect 674474 580837 674480 580889
rect 671920 579135 671926 579187
rect 671978 579175 671984 579187
rect 673840 579175 673846 579187
rect 671978 579147 673846 579175
rect 671978 579135 671984 579147
rect 673840 579135 673846 579147
rect 673898 579135 673904 579187
rect 42160 578987 42166 579039
rect 42218 579027 42224 579039
rect 43024 579027 43030 579039
rect 42218 578999 43030 579027
rect 42218 578987 42224 578999
rect 43024 578987 43030 578999
rect 43082 578987 43088 579039
rect 43024 578839 43030 578891
rect 43082 578879 43088 578891
rect 43408 578879 43414 578891
rect 43082 578851 43414 578879
rect 43082 578839 43088 578851
rect 43408 578839 43414 578851
rect 43466 578839 43472 578891
rect 42160 577137 42166 577189
rect 42218 577177 42224 577189
rect 43120 577177 43126 577189
rect 42218 577149 43126 577177
rect 42218 577137 42224 577149
rect 43120 577137 43126 577149
rect 43178 577137 43184 577189
rect 654448 576027 654454 576079
rect 654506 576067 654512 576079
rect 669904 576067 669910 576079
rect 654506 576039 669910 576067
rect 654506 576027 654512 576039
rect 669904 576027 669910 576039
rect 669962 576027 669968 576079
rect 672688 575953 672694 576005
rect 672746 575993 672752 576005
rect 673840 575993 673846 576005
rect 672746 575965 673846 575993
rect 672746 575953 672752 575965
rect 673840 575953 673846 575965
rect 673898 575953 673904 576005
rect 672496 573585 672502 573637
rect 672554 573625 672560 573637
rect 673840 573625 673846 573637
rect 672554 573597 673846 573625
rect 672554 573585 672560 573597
rect 673840 573585 673846 573597
rect 673898 573585 673904 573637
rect 42160 573437 42166 573489
rect 42218 573477 42224 573489
rect 43024 573477 43030 573489
rect 42218 573449 43030 573477
rect 42218 573437 42224 573449
rect 43024 573437 43030 573449
rect 43082 573437 43088 573489
rect 672784 573067 672790 573119
rect 672842 573107 672848 573119
rect 673840 573107 673846 573119
rect 672842 573079 673846 573107
rect 672842 573067 672848 573079
rect 673840 573067 673846 573079
rect 673898 573067 673904 573119
rect 42160 572623 42166 572675
rect 42218 572663 42224 572675
rect 42928 572663 42934 572675
rect 42218 572635 42934 572663
rect 42218 572623 42224 572635
rect 42928 572623 42934 572635
rect 42986 572623 42992 572675
rect 672880 571587 672886 571639
rect 672938 571627 672944 571639
rect 674416 571627 674422 571639
rect 672938 571599 674422 571627
rect 672938 571587 672944 571599
rect 674416 571587 674422 571599
rect 674474 571587 674480 571639
rect 42160 570995 42166 571047
rect 42218 571035 42224 571047
rect 43120 571035 43126 571047
rect 42218 571007 43126 571035
rect 42218 570995 42224 571007
rect 43120 570995 43126 571007
rect 43178 570995 43184 571047
rect 42928 570255 42934 570307
rect 42986 570295 42992 570307
rect 59536 570295 59542 570307
rect 42986 570267 59542 570295
rect 42986 570255 42992 570267
rect 59536 570255 59542 570267
rect 59594 570255 59600 570307
rect 42064 569663 42070 569715
rect 42122 569703 42128 569715
rect 43120 569703 43126 569715
rect 42122 569675 43126 569703
rect 42122 569663 42128 569675
rect 43120 569663 43126 569675
rect 43178 569663 43184 569715
rect 650128 567369 650134 567421
rect 650186 567409 650192 567421
rect 677008 567409 677014 567421
rect 650186 567381 677014 567409
rect 650186 567369 650192 567381
rect 677008 567369 677014 567381
rect 677066 567369 677072 567421
rect 654448 567295 654454 567347
rect 654506 567335 654512 567347
rect 666640 567335 666646 567347
rect 654506 567307 666646 567335
rect 654506 567295 654512 567307
rect 666640 567295 666646 567307
rect 666698 567295 666704 567347
rect 672304 564409 672310 564461
rect 672362 564449 672368 564461
rect 675088 564449 675094 564461
rect 672362 564421 675094 564449
rect 672362 564409 672368 564421
rect 675088 564409 675094 564421
rect 675146 564409 675152 564461
rect 672112 564335 672118 564387
rect 672170 564375 672176 564387
rect 674992 564375 674998 564387
rect 672170 564347 674998 564375
rect 672170 564335 672176 564347
rect 674992 564335 674998 564347
rect 675050 564335 675056 564387
rect 674224 559525 674230 559577
rect 674282 559565 674288 559577
rect 675376 559565 675382 559577
rect 674282 559537 675382 559565
rect 674282 559525 674288 559537
rect 675376 559525 675382 559537
rect 675434 559525 675440 559577
rect 43024 559303 43030 559355
rect 43082 559343 43088 559355
rect 48880 559343 48886 559355
rect 43082 559315 48886 559343
rect 43082 559303 43088 559315
rect 48880 559303 48886 559315
rect 48938 559303 48944 559355
rect 42832 558859 42838 558911
rect 42890 558899 42896 558911
rect 59536 558899 59542 558911
rect 42890 558871 59542 558899
rect 42890 558859 42896 558871
rect 59536 558859 59542 558871
rect 59594 558859 59600 558911
rect 674704 558045 674710 558097
rect 674762 558085 674768 558097
rect 675376 558085 675382 558097
rect 674762 558057 675382 558085
rect 674762 558045 674768 558057
rect 675376 558045 675382 558057
rect 675434 558045 675440 558097
rect 674992 557823 674998 557875
rect 675050 557863 675056 557875
rect 675376 557863 675382 557875
rect 675050 557835 675382 557863
rect 675050 557823 675056 557835
rect 675376 557823 675382 557835
rect 675434 557823 675440 557875
rect 673744 557601 673750 557653
rect 673802 557641 673808 557653
rect 675472 557641 675478 557653
rect 673802 557613 675478 557641
rect 673802 557601 673808 557613
rect 675472 557601 675478 557613
rect 675530 557601 675536 557653
rect 675088 557083 675094 557135
rect 675146 557123 675152 557135
rect 675472 557123 675478 557135
rect 675146 557095 675478 557123
rect 675146 557083 675152 557095
rect 675472 557083 675478 557095
rect 675530 557083 675536 557135
rect 660880 555825 660886 555877
rect 660938 555865 660944 555877
rect 674992 555865 674998 555877
rect 660938 555837 674998 555865
rect 660938 555825 660944 555837
rect 674992 555825 674998 555837
rect 675050 555825 675056 555877
rect 674416 555233 674422 555285
rect 674474 555273 674480 555285
rect 675472 555273 675478 555285
rect 674474 555245 675478 555273
rect 674474 555233 674480 555245
rect 675472 555233 675478 555245
rect 675530 555233 675536 555285
rect 673264 553753 673270 553805
rect 673322 553793 673328 553805
rect 675472 553793 675478 553805
rect 673322 553765 675478 553793
rect 673322 553753 673328 553765
rect 675472 553753 675478 553765
rect 675530 553753 675536 553805
rect 672880 553161 672886 553213
rect 672938 553201 672944 553213
rect 675376 553201 675382 553213
rect 672938 553173 675382 553201
rect 672938 553161 672944 553173
rect 675376 553161 675382 553173
rect 675434 553161 675440 553213
rect 654448 552939 654454 552991
rect 654506 552979 654512 552991
rect 666640 552979 666646 552991
rect 654506 552951 666646 552979
rect 654506 552939 654512 552951
rect 666640 552939 666646 552951
rect 666698 552939 666704 552991
rect 674320 551903 674326 551955
rect 674378 551943 674384 551955
rect 675472 551943 675478 551955
rect 674378 551915 675478 551943
rect 674378 551903 674384 551915
rect 675472 551903 675478 551915
rect 675530 551903 675536 551955
rect 674992 551607 674998 551659
rect 675050 551647 675056 551659
rect 675376 551647 675382 551659
rect 675050 551619 675382 551647
rect 675050 551607 675056 551619
rect 675376 551607 675382 551619
rect 675434 551607 675440 551659
rect 674512 550053 674518 550105
rect 674570 550093 674576 550105
rect 675472 550093 675478 550105
rect 674570 550065 675478 550093
rect 674570 550053 674576 550065
rect 675472 550053 675478 550065
rect 675530 550053 675536 550105
rect 674608 548203 674614 548255
rect 674666 548243 674672 548255
rect 675472 548243 675478 548255
rect 674666 548215 675478 548243
rect 674666 548203 674672 548215
rect 675472 548203 675478 548215
rect 675530 548203 675536 548255
rect 48880 544651 48886 544703
rect 48938 544691 48944 544703
rect 59536 544691 59542 544703
rect 48938 544663 59542 544691
rect 48938 544651 48944 544663
rect 59536 544651 59542 544663
rect 59594 544651 59600 544703
rect 41872 544207 41878 544259
rect 41930 544247 41936 544259
rect 42928 544247 42934 544259
rect 41930 544219 42934 544247
rect 41930 544207 41936 544219
rect 42928 544207 42934 544219
rect 42986 544207 42992 544259
rect 43024 541469 43030 541521
rect 43082 541509 43088 541521
rect 50512 541509 50518 541521
rect 43082 541481 50518 541509
rect 43082 541469 43088 541481
rect 50512 541469 50518 541481
rect 50570 541469 50576 541521
rect 654448 541469 654454 541521
rect 654506 541509 654512 541521
rect 669712 541509 669718 541521
rect 654506 541481 669718 541509
rect 654506 541469 654512 541481
rect 669712 541469 669718 541481
rect 669770 541469 669776 541521
rect 41584 541247 41590 541299
rect 41642 541287 41648 541299
rect 43600 541287 43606 541299
rect 41642 541259 43606 541287
rect 41642 541247 41648 541259
rect 43600 541247 43606 541259
rect 43658 541247 43664 541299
rect 42064 541173 42070 541225
rect 42122 541213 42128 541225
rect 43216 541213 43222 541225
rect 42122 541185 43222 541213
rect 42122 541173 42128 541185
rect 43216 541173 43222 541185
rect 43274 541173 43280 541225
rect 42448 541099 42454 541151
rect 42506 541139 42512 541151
rect 42506 541111 42590 541139
rect 42506 541099 42512 541111
rect 41968 540951 41974 541003
rect 42026 540991 42032 541003
rect 42448 540991 42454 541003
rect 42026 540963 42454 540991
rect 42026 540951 42032 540963
rect 42448 540951 42454 540963
rect 42506 540951 42512 541003
rect 42160 540729 42166 540781
rect 42218 540769 42224 540781
rect 42562 540769 42590 541111
rect 42218 540741 42590 540769
rect 42218 540729 42224 540741
rect 42064 538879 42070 538931
rect 42122 538919 42128 538931
rect 42928 538919 42934 538931
rect 42122 538891 42934 538919
rect 42122 538879 42128 538891
rect 42928 538879 42934 538891
rect 42986 538879 42992 538931
rect 42928 538731 42934 538783
rect 42986 538771 42992 538783
rect 43216 538771 43222 538783
rect 42986 538743 43222 538771
rect 42986 538731 42992 538743
rect 43216 538731 43222 538743
rect 43274 538731 43280 538783
rect 42160 538139 42166 538191
rect 42218 538179 42224 538191
rect 43024 538179 43030 538191
rect 42218 538151 43030 538179
rect 42218 538139 42224 538151
rect 43024 538139 43030 538151
rect 43082 538139 43088 538191
rect 669808 537177 669814 537229
rect 669866 537217 669872 537229
rect 674800 537217 674806 537229
rect 669866 537189 674806 537217
rect 669866 537177 669872 537189
rect 674800 537177 674806 537189
rect 674858 537177 674864 537229
rect 661072 536585 661078 536637
rect 661130 536625 661136 536637
rect 674800 536625 674806 536637
rect 661130 536597 674806 536625
rect 661130 536585 661136 536597
rect 674800 536585 674806 536597
rect 674858 536585 674864 536637
rect 671920 536141 671926 536193
rect 671978 536181 671984 536193
rect 674800 536181 674806 536193
rect 671978 536153 674806 536181
rect 671978 536141 671984 536153
rect 674800 536141 674806 536153
rect 674858 536141 674864 536193
rect 42064 535771 42070 535823
rect 42122 535811 42128 535823
rect 43120 535811 43126 535823
rect 42122 535783 43126 535811
rect 42122 535771 42128 535783
rect 43120 535771 43126 535783
rect 43178 535771 43184 535823
rect 655120 535771 655126 535823
rect 655178 535811 655184 535823
rect 676816 535811 676822 535823
rect 655178 535783 676822 535811
rect 655178 535771 655184 535783
rect 676816 535771 676822 535783
rect 676874 535771 676880 535823
rect 43120 535623 43126 535675
rect 43178 535663 43184 535675
rect 43600 535663 43606 535675
rect 43178 535635 43606 535663
rect 43178 535623 43184 535635
rect 43600 535623 43606 535635
rect 43658 535623 43664 535675
rect 42160 535031 42166 535083
rect 42218 535071 42224 535083
rect 42928 535071 42934 535083
rect 42218 535043 42934 535071
rect 42218 535031 42224 535043
rect 42928 535031 42934 535043
rect 42986 535031 42992 535083
rect 42160 530887 42166 530939
rect 42218 530927 42224 530939
rect 43024 530927 43030 530939
rect 42218 530899 43030 530927
rect 42218 530887 42224 530899
rect 43024 530887 43030 530899
rect 43082 530887 43088 530939
rect 42064 530221 42070 530273
rect 42122 530261 42128 530273
rect 42448 530261 42454 530273
rect 42122 530233 42454 530261
rect 42122 530221 42128 530233
rect 42448 530221 42454 530233
rect 42506 530221 42512 530273
rect 43120 530147 43126 530199
rect 43178 530147 43184 530199
rect 42448 530073 42454 530125
rect 42506 530113 42512 530125
rect 43138 530113 43166 530147
rect 42506 530085 43166 530113
rect 42506 530073 42512 530085
rect 43312 529999 43318 530051
rect 43370 530039 43376 530051
rect 43696 530039 43702 530051
rect 43370 530011 43702 530039
rect 43370 529999 43376 530011
rect 43696 529999 43702 530011
rect 43754 529999 43760 530051
rect 43024 529925 43030 529977
rect 43082 529965 43088 529977
rect 59536 529965 59542 529977
rect 43082 529937 59542 529965
rect 43082 529925 43088 529937
rect 59536 529925 59542 529937
rect 59594 529925 59600 529977
rect 654064 529925 654070 529977
rect 654122 529965 654128 529977
rect 672496 529965 672502 529977
rect 654122 529937 672502 529965
rect 654122 529925 654128 529937
rect 672496 529925 672502 529937
rect 672554 529925 672560 529977
rect 671824 529851 671830 529903
rect 671882 529891 671888 529903
rect 673648 529891 673654 529903
rect 671882 529863 673654 529891
rect 671882 529851 671888 529863
rect 673648 529851 673654 529863
rect 673706 529851 673712 529903
rect 43120 529481 43126 529533
rect 43178 529481 43184 529533
rect 43138 529447 43166 529481
rect 43138 529419 43262 529447
rect 42928 529333 42934 529385
rect 42986 529373 42992 529385
rect 43120 529373 43126 529385
rect 42986 529345 43126 529373
rect 42986 529333 42992 529345
rect 43120 529333 43126 529345
rect 43178 529333 43184 529385
rect 42448 529185 42454 529237
rect 42506 529225 42512 529237
rect 42928 529225 42934 529237
rect 42506 529197 42934 529225
rect 42506 529185 42512 529197
rect 42928 529185 42934 529197
rect 42986 529185 42992 529237
rect 42832 528889 42838 528941
rect 42890 528929 42896 528941
rect 43234 528929 43262 529419
rect 672208 529037 672214 529089
rect 672266 529077 672272 529089
rect 674800 529077 674806 529089
rect 672266 529049 674806 529077
rect 672266 529037 672272 529049
rect 674800 529037 674806 529049
rect 674858 529037 674864 529089
rect 42890 528901 43262 528929
rect 42890 528889 42896 528901
rect 672976 528445 672982 528497
rect 673034 528485 673040 528497
rect 674800 528485 674806 528497
rect 673034 528457 674806 528485
rect 673034 528445 673040 528457
rect 674800 528445 674806 528457
rect 674858 528445 674864 528497
rect 42160 527631 42166 527683
rect 42218 527671 42224 527683
rect 42928 527671 42934 527683
rect 42218 527643 42934 527671
rect 42218 527631 42224 527643
rect 42928 527631 42934 527643
rect 42986 527631 42992 527683
rect 42064 527039 42070 527091
rect 42122 527079 42128 527091
rect 43120 527079 43126 527091
rect 42122 527051 43126 527079
rect 42122 527039 42128 527051
rect 43120 527039 43126 527051
rect 43178 527039 43184 527091
rect 42160 526447 42166 526499
rect 42218 526487 42224 526499
rect 42832 526487 42838 526499
rect 42218 526459 42838 526487
rect 42218 526447 42224 526459
rect 42832 526447 42838 526459
rect 42890 526447 42896 526499
rect 677200 525929 677206 525981
rect 677258 525969 677264 525981
rect 677392 525969 677398 525981
rect 677258 525941 677398 525969
rect 677258 525929 677264 525941
rect 677392 525929 677398 525941
rect 677450 525929 677456 525981
rect 650224 524301 650230 524353
rect 650282 524341 650288 524353
rect 677008 524341 677014 524353
rect 650282 524313 677014 524341
rect 650282 524301 650288 524313
rect 677008 524301 677014 524313
rect 677066 524301 677072 524353
rect 41872 519787 41878 519839
rect 41930 519827 41936 519839
rect 43024 519827 43030 519839
rect 41930 519799 43030 519827
rect 41930 519787 41936 519799
rect 43024 519787 43030 519799
rect 43082 519787 43088 519839
rect 654448 519269 654454 519321
rect 654506 519309 654512 519321
rect 663856 519309 663862 519321
rect 654506 519281 663862 519309
rect 654506 519269 654512 519281
rect 663856 519269 663862 519281
rect 663914 519269 663920 519321
rect 53968 515495 53974 515547
rect 54026 515535 54032 515547
rect 59536 515535 59542 515547
rect 54026 515507 59542 515535
rect 54026 515495 54032 515507
rect 59536 515495 59542 515507
rect 59594 515495 59600 515547
rect 43120 509723 43126 509775
rect 43178 509763 43184 509775
rect 43312 509763 43318 509775
rect 43178 509735 43318 509763
rect 43178 509723 43184 509735
rect 43312 509723 43318 509735
rect 43370 509723 43376 509775
rect 654448 506911 654454 506963
rect 654506 506951 654512 506963
rect 663856 506951 663862 506963
rect 654506 506923 663862 506951
rect 654506 506911 654512 506923
rect 663856 506911 663862 506923
rect 663914 506911 663920 506963
rect 47728 501139 47734 501191
rect 47786 501179 47792 501191
rect 59536 501179 59542 501191
rect 47786 501151 59542 501179
rect 47786 501139 47792 501151
rect 59536 501139 59542 501151
rect 59594 501139 59600 501191
rect 654352 495367 654358 495419
rect 654410 495407 654416 495419
rect 661168 495407 661174 495419
rect 654410 495379 661174 495407
rect 654410 495367 654416 495379
rect 661168 495367 661174 495379
rect 661226 495367 661232 495419
rect 664048 493221 664054 493273
rect 664106 493261 664112 493273
rect 675088 493261 675094 493273
rect 664106 493233 675094 493261
rect 664106 493221 664112 493233
rect 675088 493221 675094 493233
rect 675146 493221 675152 493273
rect 655312 492481 655318 492533
rect 655370 492521 655376 492533
rect 674896 492521 674902 492533
rect 655370 492493 674902 492521
rect 655370 492481 655376 492493
rect 674896 492481 674902 492493
rect 674954 492481 674960 492533
rect 672592 492407 672598 492459
rect 672650 492447 672656 492459
rect 673840 492447 673846 492459
rect 672650 492419 673846 492447
rect 672650 492407 672656 492419
rect 673840 492407 673846 492419
rect 673898 492407 673904 492459
rect 44752 486709 44758 486761
rect 44810 486749 44816 486761
rect 58576 486749 58582 486761
rect 44810 486721 58582 486749
rect 44810 486709 44816 486721
rect 58576 486709 58582 486721
rect 58634 486709 58640 486761
rect 654256 483823 654262 483875
rect 654314 483863 654320 483875
rect 666928 483863 666934 483875
rect 654314 483835 666934 483863
rect 654314 483823 654320 483835
rect 666928 483823 666934 483835
rect 666986 483823 666992 483875
rect 672880 483749 672886 483801
rect 672938 483789 672944 483801
rect 673840 483789 673846 483801
rect 672938 483761 673846 483789
rect 672938 483749 672944 483761
rect 673840 483749 673846 483761
rect 673898 483749 673904 483801
rect 650320 479457 650326 479509
rect 650378 479497 650384 479509
rect 677008 479497 677014 479509
rect 650378 479469 677014 479497
rect 650378 479457 650384 479469
rect 677008 479457 677014 479469
rect 677066 479457 677072 479509
rect 44848 472353 44854 472405
rect 44906 472393 44912 472405
rect 59536 472393 59542 472405
rect 44906 472365 59542 472393
rect 44906 472353 44912 472365
rect 59536 472353 59542 472365
rect 59594 472353 59600 472405
rect 654448 472205 654454 472257
rect 654506 472245 654512 472257
rect 660976 472245 660982 472257
rect 654506 472217 660982 472245
rect 654506 472205 654512 472217
rect 660976 472205 660982 472217
rect 661034 472205 661040 472257
rect 43312 469393 43318 469445
rect 43370 469433 43376 469445
rect 43600 469433 43606 469445
rect 43370 469405 43606 469433
rect 43370 469393 43376 469405
rect 43600 469393 43606 469405
rect 43658 469393 43664 469445
rect 50512 457923 50518 457975
rect 50570 457963 50576 457975
rect 59536 457963 59542 457975
rect 50570 457935 59542 457963
rect 50570 457923 50576 457935
rect 59536 457923 59542 457935
rect 59594 457923 59600 457975
rect 654448 457923 654454 457975
rect 654506 457963 654512 457975
rect 660976 457963 660982 457975
rect 654506 457935 660982 457963
rect 654506 457923 654512 457935
rect 660976 457923 660982 457935
rect 661034 457923 661040 457975
rect 43216 449265 43222 449317
rect 43274 449305 43280 449317
rect 43600 449305 43606 449317
rect 43274 449277 43606 449305
rect 43274 449265 43280 449277
rect 43600 449265 43606 449277
rect 43658 449265 43664 449317
rect 654352 446379 654358 446431
rect 654410 446419 654416 446431
rect 669808 446419 669814 446431
rect 654410 446391 669814 446419
rect 654410 446379 654416 446391
rect 669808 446379 669814 446391
rect 669866 446379 669872 446431
rect 53872 443567 53878 443619
rect 53930 443607 53936 443619
rect 59536 443607 59542 443619
rect 53930 443579 59542 443607
rect 53930 443567 53936 443579
rect 59536 443567 59542 443579
rect 59594 443567 59600 443619
rect 654448 434909 654454 434961
rect 654506 434949 654512 434961
rect 663952 434949 663958 434961
rect 654506 434921 663958 434949
rect 654506 434909 654512 434921
rect 663952 434909 663958 434921
rect 664010 434909 664016 434961
rect 42832 432245 42838 432297
rect 42890 432285 42896 432297
rect 53968 432285 53974 432297
rect 42890 432257 53974 432285
rect 42890 432245 42896 432257
rect 53968 432245 53974 432257
rect 54026 432245 54032 432297
rect 42544 431949 42550 432001
rect 42602 431989 42608 432001
rect 47728 431989 47734 432001
rect 42602 431961 47734 431989
rect 42602 431949 42608 431961
rect 47728 431949 47734 431961
rect 47786 431949 47792 432001
rect 47632 429137 47638 429189
rect 47690 429177 47696 429189
rect 59536 429177 59542 429189
rect 47690 429149 59542 429177
rect 47690 429137 47696 429149
rect 59536 429137 59542 429149
rect 59594 429137 59600 429189
rect 654448 426177 654454 426229
rect 654506 426217 654512 426229
rect 669616 426217 669622 426229
rect 654506 426189 669622 426217
rect 654506 426177 654512 426189
rect 669616 426177 669622 426189
rect 669674 426177 669680 426229
rect 42928 423365 42934 423417
rect 42986 423405 42992 423417
rect 43696 423405 43702 423417
rect 42986 423377 43702 423405
rect 42986 423365 42992 423377
rect 43696 423365 43702 423377
rect 43754 423365 43760 423417
rect 40240 420479 40246 420531
rect 40298 420519 40304 420531
rect 41776 420519 41782 420531
rect 40298 420491 41782 420519
rect 40298 420479 40304 420491
rect 41776 420479 41782 420491
rect 41834 420479 41840 420531
rect 42448 417593 42454 417645
rect 42506 417633 42512 417645
rect 56176 417633 56182 417645
rect 42506 417605 56182 417633
rect 42506 417593 42512 417605
rect 56176 417593 56182 417605
rect 56234 417593 56240 417645
rect 39952 415891 39958 415943
rect 40010 415931 40016 415943
rect 42448 415931 42454 415943
rect 40010 415903 42454 415931
rect 40010 415891 40016 415903
rect 42448 415891 42454 415903
rect 42506 415891 42512 415943
rect 40048 415373 40054 415425
rect 40106 415413 40112 415425
rect 43120 415413 43126 415425
rect 40106 415385 43126 415413
rect 40106 415373 40112 415385
rect 43120 415373 43126 415385
rect 43178 415373 43184 415425
rect 40144 414707 40150 414759
rect 40202 414747 40208 414759
rect 43024 414747 43030 414759
rect 40202 414719 43030 414747
rect 40202 414707 40208 414719
rect 43024 414707 43030 414719
rect 43082 414707 43088 414759
rect 45040 414707 45046 414759
rect 45098 414747 45104 414759
rect 58384 414747 58390 414759
rect 45098 414719 58390 414747
rect 45098 414707 45104 414719
rect 58384 414707 58390 414719
rect 58442 414707 58448 414759
rect 41776 413375 41782 413427
rect 41834 413375 41840 413427
rect 41794 413205 41822 413375
rect 41776 413153 41782 413205
rect 41834 413153 41840 413205
rect 653872 411821 653878 411873
rect 653930 411861 653936 411873
rect 669520 411861 669526 411873
rect 653930 411833 669526 411861
rect 653930 411821 653936 411833
rect 669520 411821 669526 411833
rect 669578 411821 669584 411873
rect 42448 411377 42454 411429
rect 42506 411417 42512 411429
rect 43216 411417 43222 411429
rect 42506 411389 43222 411417
rect 42506 411377 42512 411389
rect 43216 411377 43222 411389
rect 43274 411377 43280 411429
rect 42160 410933 42166 410985
rect 42218 410973 42224 410985
rect 42544 410973 42550 410985
rect 42218 410945 42550 410973
rect 42218 410933 42224 410945
rect 42544 410933 42550 410945
rect 42602 410933 42608 410985
rect 42160 409675 42166 409727
rect 42218 409715 42224 409727
rect 42544 409715 42550 409727
rect 42218 409687 42550 409715
rect 42218 409675 42224 409687
rect 42544 409675 42550 409687
rect 42602 409675 42608 409727
rect 42160 409453 42166 409505
rect 42218 409493 42224 409505
rect 42352 409493 42358 409505
rect 42218 409465 42358 409493
rect 42218 409453 42224 409465
rect 42352 409453 42358 409465
rect 42410 409453 42416 409505
rect 42352 409305 42358 409357
rect 42410 409345 42416 409357
rect 42928 409345 42934 409357
rect 42410 409317 42934 409345
rect 42410 409305 42416 409317
rect 42928 409305 42934 409317
rect 42986 409305 42992 409357
rect 43312 409123 43318 409135
rect 43042 409095 43318 409123
rect 43042 409061 43070 409095
rect 43312 409083 43318 409095
rect 43370 409083 43376 409135
rect 43024 409009 43030 409061
rect 43082 409009 43088 409061
rect 42160 408195 42166 408247
rect 42218 408235 42224 408247
rect 42352 408235 42358 408247
rect 42218 408207 42358 408235
rect 42218 408195 42224 408207
rect 42352 408195 42358 408207
rect 42410 408195 42416 408247
rect 42064 407455 42070 407507
rect 42122 407495 42128 407507
rect 43120 407495 43126 407507
rect 42122 407467 43126 407495
rect 42122 407455 42128 407467
rect 43120 407455 43126 407467
rect 43178 407455 43184 407507
rect 42160 407011 42166 407063
rect 42218 407051 42224 407063
rect 42928 407051 42934 407063
rect 42218 407023 42934 407051
rect 42218 407011 42224 407023
rect 42928 407011 42934 407023
rect 42986 407011 42992 407063
rect 42544 406049 42550 406101
rect 42602 406089 42608 406101
rect 53392 406089 53398 406101
rect 42602 406061 53398 406089
rect 42602 406049 42608 406061
rect 53392 406049 53398 406061
rect 53450 406049 53456 406101
rect 672400 406049 672406 406101
rect 672458 406089 672464 406101
rect 673840 406089 673846 406101
rect 672458 406061 673846 406089
rect 672458 406049 672464 406061
rect 673840 406049 673846 406061
rect 673898 406049 673904 406101
rect 666832 405457 666838 405509
rect 666890 405497 666896 405509
rect 674704 405497 674710 405509
rect 666890 405469 674710 405497
rect 666890 405457 666896 405469
rect 674704 405457 674710 405469
rect 674762 405457 674768 405509
rect 669904 404421 669910 404473
rect 669962 404461 669968 404473
rect 674704 404461 674710 404473
rect 669962 404433 674710 404461
rect 669962 404421 669968 404433
rect 674704 404421 674710 404433
rect 674762 404421 674768 404473
rect 42160 403163 42166 403215
rect 42218 403203 42224 403215
rect 43024 403203 43030 403215
rect 42218 403175 43030 403203
rect 42218 403163 42224 403175
rect 43024 403163 43030 403175
rect 43082 403163 43088 403215
rect 43312 403163 43318 403215
rect 43370 403163 43376 403215
rect 42928 403089 42934 403141
rect 42986 403129 42992 403141
rect 43330 403129 43358 403163
rect 42986 403101 43358 403129
rect 42986 403089 42992 403101
rect 673360 400425 673366 400477
rect 673418 400465 673424 400477
rect 676912 400465 676918 400477
rect 673418 400437 676918 400465
rect 673418 400425 673424 400437
rect 676912 400425 676918 400437
rect 676970 400425 676976 400477
rect 56272 400351 56278 400403
rect 56330 400391 56336 400403
rect 57616 400391 57622 400403
rect 56330 400363 57622 400391
rect 56330 400351 56336 400363
rect 57616 400351 57622 400363
rect 57674 400351 57680 400403
rect 654448 400351 654454 400403
rect 654506 400391 654512 400403
rect 666832 400391 666838 400403
rect 654506 400363 666838 400391
rect 654506 400351 654512 400363
rect 666832 400351 666838 400363
rect 666890 400351 666896 400403
rect 673744 400351 673750 400403
rect 673802 400391 673808 400403
rect 677200 400391 677206 400403
rect 673802 400363 677206 400391
rect 673802 400351 673808 400363
rect 677200 400351 677206 400363
rect 677258 400351 677264 400403
rect 650416 391767 650422 391819
rect 650474 391807 650480 391819
rect 677104 391807 677110 391819
rect 650474 391779 677110 391807
rect 650474 391767 650480 391779
rect 677104 391767 677110 391779
rect 677162 391767 677168 391819
rect 42352 389325 42358 389377
rect 42410 389365 42416 389377
rect 44848 389365 44854 389377
rect 42410 389337 44854 389365
rect 42410 389325 42416 389337
rect 44848 389325 44854 389337
rect 44906 389325 44912 389377
rect 654448 388807 654454 388859
rect 654506 388847 654512 388859
rect 669616 388847 669622 388859
rect 654506 388819 669622 388847
rect 654506 388807 654512 388819
rect 669616 388807 669622 388819
rect 669674 388807 669680 388859
rect 42640 388733 42646 388785
rect 42698 388773 42704 388785
rect 50512 388773 50518 388785
rect 42698 388745 50518 388773
rect 42698 388733 42704 388745
rect 50512 388733 50518 388745
rect 50570 388733 50576 388785
rect 42640 387993 42646 388045
rect 42698 388033 42704 388045
rect 44752 388033 44758 388045
rect 42698 388005 44758 388033
rect 42698 387993 42704 388005
rect 44752 387993 44758 388005
rect 44810 387993 44816 388045
rect 675376 386365 675382 386417
rect 675434 386365 675440 386417
rect 675394 386195 675422 386365
rect 675376 386143 675382 386195
rect 675434 386143 675440 386195
rect 44944 385921 44950 385973
rect 45002 385961 45008 385973
rect 59248 385961 59254 385973
rect 45002 385933 59254 385961
rect 45002 385921 45008 385933
rect 59248 385921 59254 385933
rect 59306 385921 59312 385973
rect 675184 385403 675190 385455
rect 675242 385443 675248 385455
rect 675472 385443 675478 385455
rect 675242 385415 675478 385443
rect 675242 385403 675248 385415
rect 675472 385403 675478 385415
rect 675530 385403 675536 385455
rect 675088 384811 675094 384863
rect 675146 384851 675152 384863
rect 675376 384851 675382 384863
rect 675146 384823 675382 384851
rect 675146 384811 675152 384823
rect 675376 384811 675382 384823
rect 675434 384811 675440 384863
rect 674896 384663 674902 384715
rect 674954 384703 674960 384715
rect 675088 384703 675094 384715
rect 674954 384675 675094 384703
rect 674954 384663 674960 384675
rect 675088 384663 675094 384675
rect 675146 384663 675152 384715
rect 674128 383109 674134 383161
rect 674186 383149 674192 383161
rect 675280 383149 675286 383161
rect 674186 383121 675286 383149
rect 674186 383109 674192 383121
rect 675280 383109 675286 383121
rect 675338 383109 675344 383161
rect 674224 382443 674230 382495
rect 674282 382483 674288 382495
rect 675472 382483 675478 382495
rect 674282 382455 675478 382483
rect 674282 382443 674288 382455
rect 675472 382443 675478 382455
rect 675530 382443 675536 382495
rect 654448 380075 654454 380127
rect 654506 380115 654512 380127
rect 666736 380115 666742 380127
rect 654506 380087 666742 380115
rect 654506 380075 654512 380087
rect 666736 380075 666742 380087
rect 666794 380075 666800 380127
rect 674800 378151 674806 378203
rect 674858 378191 674864 378203
rect 675376 378191 675382 378203
rect 674858 378163 675382 378191
rect 674858 378151 674864 378163
rect 675376 378151 675382 378163
rect 675434 378151 675440 378203
rect 674512 377559 674518 377611
rect 674570 377599 674576 377611
rect 675376 377599 675382 377611
rect 674570 377571 675382 377599
rect 674570 377559 674576 377571
rect 675376 377559 675382 377571
rect 675434 377559 675440 377611
rect 674608 376893 674614 376945
rect 674666 376933 674672 376945
rect 675472 376933 675478 376945
rect 674666 376905 675478 376933
rect 674666 376893 674672 376905
rect 675472 376893 675478 376905
rect 675530 376893 675536 376945
rect 42640 376523 42646 376575
rect 42698 376563 42704 376575
rect 44752 376563 44758 376575
rect 42698 376535 44758 376563
rect 42698 376523 42704 376535
rect 44752 376523 44758 376535
rect 44810 376523 44816 376575
rect 673936 375709 673942 375761
rect 673994 375749 674000 375761
rect 675472 375749 675478 375761
rect 673994 375721 675478 375749
rect 673994 375709 674000 375721
rect 675472 375709 675478 375721
rect 675530 375709 675536 375761
rect 40048 374303 40054 374355
rect 40106 374343 40112 374355
rect 43120 374343 43126 374355
rect 40106 374315 43126 374343
rect 40106 374303 40112 374315
rect 43120 374303 43126 374315
rect 43178 374303 43184 374355
rect 40240 373637 40246 373689
rect 40298 373677 40304 373689
rect 42832 373677 42838 373689
rect 40298 373649 42838 373677
rect 40298 373637 40304 373649
rect 42832 373637 42838 373649
rect 42890 373637 42896 373689
rect 39952 371565 39958 371617
rect 40010 371605 40016 371617
rect 43312 371605 43318 371617
rect 40010 371577 43318 371605
rect 40010 371565 40016 371577
rect 43312 371565 43318 371577
rect 43370 371565 43376 371617
rect 47728 371565 47734 371617
rect 47786 371605 47792 371617
rect 59536 371605 59542 371617
rect 47786 371577 59542 371605
rect 47786 371565 47792 371577
rect 59536 371565 59542 371577
rect 59594 371565 59600 371617
rect 42736 370455 42742 370507
rect 42794 370495 42800 370507
rect 43216 370495 43222 370507
rect 42794 370467 43222 370495
rect 42794 370455 42800 370467
rect 43216 370455 43222 370467
rect 43274 370455 43280 370507
rect 42160 369937 42166 369989
rect 42218 369977 42224 369989
rect 42352 369977 42358 369989
rect 42218 369949 42358 369977
rect 42218 369937 42224 369949
rect 42352 369937 42358 369949
rect 42410 369937 42416 369989
rect 42352 369789 42358 369841
rect 42410 369829 42416 369841
rect 42832 369829 42838 369841
rect 42410 369801 42838 369829
rect 42410 369789 42416 369801
rect 42832 369789 42838 369801
rect 42890 369789 42896 369841
rect 42928 369493 42934 369545
rect 42986 369533 42992 369545
rect 43120 369533 43126 369545
rect 42986 369505 43126 369533
rect 42986 369493 42992 369505
rect 43120 369493 43126 369505
rect 43178 369493 43184 369545
rect 43216 369197 43222 369249
rect 43274 369237 43280 369249
rect 43408 369237 43414 369249
rect 43274 369209 43414 369237
rect 43274 369197 43280 369209
rect 43408 369197 43414 369209
rect 43466 369197 43472 369249
rect 42064 368087 42070 368139
rect 42122 368127 42128 368139
rect 43120 368127 43126 368139
rect 42122 368099 43126 368127
rect 42122 368087 42128 368099
rect 43120 368087 43126 368099
rect 43178 368087 43184 368139
rect 43216 368087 43222 368139
rect 43274 368087 43280 368139
rect 43234 367917 43262 368087
rect 43216 367865 43222 367917
rect 43274 367865 43280 367917
rect 42064 367347 42070 367399
rect 42122 367387 42128 367399
rect 47440 367387 47446 367399
rect 42122 367359 47446 367387
rect 42122 367347 42128 367359
rect 47440 367347 47446 367359
rect 47498 367347 47504 367399
rect 42064 366237 42070 366289
rect 42122 366277 42128 366289
rect 42928 366277 42934 366289
rect 42122 366249 42934 366277
rect 42122 366237 42128 366249
rect 42928 366237 42934 366249
rect 42986 366237 42992 366289
rect 654448 365793 654454 365845
rect 654506 365833 654512 365845
rect 661072 365833 661078 365845
rect 654506 365805 661078 365833
rect 654506 365793 654512 365805
rect 661072 365793 661078 365805
rect 661130 365793 661136 365845
rect 42160 364979 42166 365031
rect 42218 365019 42224 365031
rect 42832 365019 42838 365031
rect 42218 364991 42838 365019
rect 42218 364979 42224 364991
rect 42832 364979 42838 364991
rect 42890 364979 42896 365031
rect 42064 364239 42070 364291
rect 42122 364279 42128 364291
rect 43024 364279 43030 364291
rect 42122 364251 43030 364279
rect 42122 364239 42128 364251
rect 43024 364239 43030 364251
rect 43082 364239 43088 364291
rect 42160 363795 42166 363847
rect 42218 363835 42224 363847
rect 42352 363835 42358 363847
rect 42218 363807 42358 363835
rect 42218 363795 42224 363807
rect 42352 363795 42358 363807
rect 42410 363795 42416 363847
rect 42160 360095 42166 360147
rect 42218 360135 42224 360147
rect 43120 360135 43126 360147
rect 42218 360107 43126 360135
rect 42218 360095 42224 360107
rect 43120 360095 43126 360107
rect 43178 360095 43184 360147
rect 669712 360021 669718 360073
rect 669770 360061 669776 360073
rect 674416 360061 674422 360073
rect 669770 360033 674422 360061
rect 669770 360021 669776 360033
rect 674416 360021 674422 360033
rect 674474 360021 674480 360073
rect 666640 359725 666646 359777
rect 666698 359765 666704 359777
rect 674704 359765 674710 359777
rect 666698 359737 674710 359765
rect 666698 359725 666704 359737
rect 674704 359725 674710 359737
rect 674762 359725 674768 359777
rect 672496 358985 672502 359037
rect 672554 359025 672560 359037
rect 674416 359025 674422 359037
rect 672554 358997 674422 359025
rect 672554 358985 672560 358997
rect 674416 358985 674422 358997
rect 674474 358985 674480 359037
rect 47440 357135 47446 357187
rect 47498 357175 47504 357187
rect 59536 357175 59542 357187
rect 47498 357147 59542 357175
rect 47498 357135 47504 357147
rect 59536 357135 59542 357147
rect 59594 357135 59600 357187
rect 42832 345887 42838 345939
rect 42890 345927 42896 345939
rect 47632 345927 47638 345939
rect 42890 345899 47638 345927
rect 42890 345887 42896 345899
rect 47632 345887 47638 345899
rect 47690 345887 47696 345939
rect 650512 345591 650518 345643
rect 650570 345631 650576 345643
rect 677008 345631 677014 345643
rect 650570 345603 677014 345631
rect 650570 345591 650576 345603
rect 677008 345591 677014 345603
rect 677066 345591 677072 345643
rect 42832 345369 42838 345421
rect 42890 345409 42896 345421
rect 45040 345409 45046 345421
rect 42890 345381 45046 345409
rect 42890 345369 42896 345381
rect 45040 345369 45046 345381
rect 45098 345369 45104 345421
rect 42832 344777 42838 344829
rect 42890 344817 42896 344829
rect 53872 344817 53878 344829
rect 42890 344789 53878 344817
rect 42890 344777 42896 344789
rect 53872 344777 53878 344789
rect 53930 344777 53936 344829
rect 50512 342779 50518 342831
rect 50570 342819 50576 342831
rect 58384 342819 58390 342831
rect 50570 342791 58390 342819
rect 50570 342779 50576 342791
rect 58384 342779 58390 342791
rect 58442 342779 58448 342831
rect 654448 342705 654454 342757
rect 654506 342745 654512 342757
rect 666640 342745 666646 342757
rect 654506 342717 666646 342745
rect 654506 342705 654512 342717
rect 666640 342705 666646 342717
rect 666698 342705 666704 342757
rect 675184 340929 675190 340981
rect 675242 340969 675248 340981
rect 675472 340969 675478 340981
rect 675242 340941 675478 340969
rect 675242 340929 675248 340941
rect 675472 340929 675478 340941
rect 675530 340929 675536 340981
rect 674992 340781 674998 340833
rect 675050 340821 675056 340833
rect 675184 340821 675190 340833
rect 675050 340793 675190 340821
rect 675050 340781 675056 340793
rect 675184 340781 675190 340793
rect 675242 340781 675248 340833
rect 674896 339523 674902 339575
rect 674954 339563 674960 339575
rect 675376 339563 675382 339575
rect 674954 339535 675382 339563
rect 674954 339523 674960 339535
rect 675376 339523 675382 339535
rect 675434 339523 675440 339575
rect 674320 336563 674326 336615
rect 674378 336603 674384 336615
rect 675376 336603 675382 336615
rect 674378 336575 675382 336603
rect 674378 336563 674384 336575
rect 675376 336563 675382 336575
rect 675434 336563 675440 336615
rect 673936 333529 673942 333581
rect 673994 333569 674000 333581
rect 675376 333569 675382 333581
rect 673994 333541 675382 333569
rect 673994 333529 674000 333541
rect 675376 333529 675382 333541
rect 675434 333529 675440 333581
rect 674032 332715 674038 332767
rect 674090 332755 674096 332767
rect 675376 332755 675382 332767
rect 674090 332727 675382 332755
rect 674090 332715 674096 332727
rect 675376 332715 675382 332727
rect 675434 332715 675440 332767
rect 654448 332271 654454 332323
rect 654506 332311 654512 332323
rect 663760 332311 663766 332323
rect 654506 332283 663766 332311
rect 654506 332271 654512 332283
rect 663760 332271 663766 332283
rect 663818 332271 663824 332323
rect 43216 332197 43222 332249
rect 43274 332237 43280 332249
rect 45040 332237 45046 332249
rect 43274 332209 45046 332237
rect 43274 332197 43280 332209
rect 45040 332197 45046 332209
rect 45098 332197 45104 332249
rect 674128 332197 674134 332249
rect 674186 332237 674192 332249
rect 675472 332237 675478 332249
rect 674186 332209 675478 332237
rect 674186 332197 674192 332209
rect 675472 332197 675478 332209
rect 675530 332197 675536 332249
rect 674512 331753 674518 331805
rect 674570 331793 674576 331805
rect 675376 331793 675382 331805
rect 674570 331765 675382 331793
rect 674570 331753 674576 331765
rect 675376 331753 675382 331765
rect 675434 331753 675440 331805
rect 40144 329533 40150 329585
rect 40202 329573 40208 329585
rect 43024 329573 43030 329585
rect 40202 329545 43030 329573
rect 40202 329533 40208 329545
rect 43024 329533 43030 329545
rect 43082 329533 43088 329585
rect 40048 329311 40054 329363
rect 40106 329351 40112 329363
rect 43120 329351 43126 329363
rect 40106 329323 43126 329351
rect 40106 329311 40112 329323
rect 43120 329311 43126 329323
rect 43178 329311 43184 329363
rect 53392 328349 53398 328401
rect 53450 328389 53456 328401
rect 57808 328389 57814 328401
rect 53450 328361 57814 328389
rect 53450 328349 53456 328361
rect 57808 328349 57814 328361
rect 57866 328349 57872 328401
rect 41776 327017 41782 327069
rect 41834 327017 41840 327069
rect 41794 326773 41822 327017
rect 42256 326943 42262 326995
rect 42314 326983 42320 326995
rect 42928 326983 42934 326995
rect 42314 326955 42934 326983
rect 42314 326943 42320 326955
rect 42928 326943 42934 326955
rect 42986 326943 42992 326995
rect 41776 326721 41782 326773
rect 41834 326721 41840 326773
rect 42064 324871 42070 324923
rect 42122 324911 42128 324923
rect 42832 324911 42838 324923
rect 42122 324883 42838 324911
rect 42122 324871 42128 324883
rect 42832 324871 42838 324883
rect 42890 324871 42896 324923
rect 42160 324131 42166 324183
rect 42218 324171 42224 324183
rect 50320 324171 50326 324183
rect 42218 324143 50326 324171
rect 42218 324131 42224 324143
rect 50320 324131 50326 324143
rect 50378 324131 50384 324183
rect 42160 323095 42166 323147
rect 42218 323135 42224 323147
rect 43120 323135 43126 323147
rect 42218 323107 43126 323135
rect 42218 323095 42224 323107
rect 43120 323095 43126 323107
rect 43178 323095 43184 323147
rect 42064 321763 42070 321815
rect 42122 321803 42128 321815
rect 42544 321803 42550 321815
rect 42122 321775 42550 321803
rect 42122 321763 42128 321775
rect 42544 321763 42550 321775
rect 42602 321763 42608 321815
rect 42160 321023 42166 321075
rect 42218 321063 42224 321075
rect 43024 321063 43030 321075
rect 42218 321035 43030 321063
rect 42218 321023 42224 321035
rect 43024 321023 43030 321035
rect 43082 321023 43088 321075
rect 42256 318729 42262 318781
rect 42314 318769 42320 318781
rect 42832 318769 42838 318781
rect 42314 318741 42838 318769
rect 42314 318729 42320 318741
rect 42832 318729 42838 318741
rect 42890 318729 42896 318781
rect 42064 316879 42070 316931
rect 42122 316919 42128 316931
rect 42928 316919 42934 316931
rect 42122 316891 42934 316919
rect 42122 316879 42128 316891
rect 42928 316879 42934 316891
rect 42986 316879 42992 316931
rect 661168 315029 661174 315081
rect 661226 315069 661232 315081
rect 674416 315069 674422 315081
rect 661226 315041 674422 315069
rect 661226 315029 661232 315041
rect 674416 315029 674422 315041
rect 674474 315029 674480 315081
rect 663856 314733 663862 314785
rect 663914 314773 663920 314785
rect 674704 314773 674710 314785
rect 663914 314745 674710 314773
rect 663914 314733 663920 314745
rect 674704 314733 674710 314745
rect 674762 314733 674768 314785
rect 666928 313993 666934 314045
rect 666986 314033 666992 314045
rect 674416 314033 674422 314045
rect 666986 314005 674422 314033
rect 666986 313993 666992 314005
rect 674416 313993 674422 314005
rect 674474 313993 674480 314045
rect 44848 313919 44854 313971
rect 44906 313959 44912 313971
rect 58000 313959 58006 313971
rect 44906 313931 58006 313959
rect 44906 313919 44912 313931
rect 58000 313919 58006 313931
rect 58058 313919 58064 313971
rect 42832 302671 42838 302723
rect 42890 302711 42896 302723
rect 44944 302711 44950 302723
rect 42890 302683 44950 302711
rect 42890 302671 42896 302683
rect 44944 302671 44950 302683
rect 45002 302671 45008 302723
rect 650608 302597 650614 302649
rect 650666 302637 650672 302649
rect 674416 302637 674422 302649
rect 650666 302609 674422 302637
rect 650666 302597 650672 302609
rect 674416 302597 674422 302609
rect 674474 302597 674480 302649
rect 42448 302301 42454 302353
rect 42506 302341 42512 302353
rect 47728 302341 47734 302353
rect 42506 302313 47734 302341
rect 42506 302301 42512 302313
rect 47728 302301 47734 302313
rect 47786 302301 47792 302353
rect 42832 301635 42838 301687
rect 42890 301675 42896 301687
rect 56272 301675 56278 301687
rect 42890 301647 56278 301675
rect 42890 301635 42896 301647
rect 56272 301635 56278 301647
rect 56330 301635 56336 301687
rect 44944 299563 44950 299615
rect 45002 299603 45008 299615
rect 59440 299603 59446 299615
rect 45002 299575 59446 299603
rect 45002 299563 45008 299575
rect 59440 299563 59446 299575
rect 59498 299563 59504 299615
rect 674896 295419 674902 295471
rect 674954 295459 674960 295471
rect 675088 295459 675094 295471
rect 674954 295431 675094 295459
rect 674954 295419 674960 295431
rect 675088 295419 675094 295431
rect 675146 295419 675152 295471
rect 674032 294753 674038 294805
rect 674090 294793 674096 294805
rect 675088 294793 675094 294805
rect 674090 294765 675094 294793
rect 674090 294753 674096 294765
rect 675088 294753 675094 294765
rect 675146 294753 675152 294805
rect 654544 293791 654550 293843
rect 654602 293831 654608 293843
rect 663760 293831 663766 293843
rect 654602 293803 663766 293831
rect 654602 293791 654608 293803
rect 663760 293791 663766 293803
rect 663818 293791 663824 293843
rect 674800 293495 674806 293547
rect 674858 293535 674864 293547
rect 675088 293535 675094 293547
rect 674858 293507 675094 293535
rect 674858 293495 674864 293507
rect 675088 293495 675094 293507
rect 675146 293495 675152 293547
rect 674320 292903 674326 292955
rect 674378 292943 674384 292955
rect 675376 292943 675382 292955
rect 674378 292915 675382 292943
rect 674378 292903 674384 292915
rect 675376 292903 675382 292915
rect 675434 292903 675440 292955
rect 674704 291719 674710 291771
rect 674762 291759 674768 291771
rect 675088 291759 675094 291771
rect 674762 291731 675094 291759
rect 674762 291719 674768 291731
rect 675088 291719 675094 291731
rect 675146 291719 675152 291771
rect 674512 291645 674518 291697
rect 674570 291685 674576 291697
rect 675184 291685 675190 291697
rect 674570 291657 675190 291685
rect 674570 291645 674576 291657
rect 675184 291645 675190 291657
rect 675242 291645 675248 291697
rect 42832 290091 42838 290143
rect 42890 290131 42896 290143
rect 47632 290131 47638 290143
rect 42890 290103 47638 290131
rect 42890 290091 42896 290103
rect 47632 290091 47638 290103
rect 47690 290091 47696 290143
rect 673936 289425 673942 289477
rect 673994 289465 674000 289477
rect 675376 289465 675382 289477
rect 673994 289437 675382 289465
rect 673994 289425 674000 289437
rect 675376 289425 675382 289437
rect 675434 289425 675440 289477
rect 674992 288537 674998 288589
rect 675050 288577 675056 288589
rect 675472 288577 675478 288589
rect 675050 288549 675478 288577
rect 675050 288537 675056 288549
rect 675472 288537 675478 288549
rect 675530 288537 675536 288589
rect 674416 287723 674422 287775
rect 674474 287763 674480 287775
rect 675376 287763 675382 287775
rect 674474 287735 675382 287763
rect 674474 287723 674480 287735
rect 675376 287723 675382 287735
rect 675434 287723 675440 287775
rect 674128 287205 674134 287257
rect 674186 287245 674192 287257
rect 675472 287245 675478 287257
rect 674186 287217 675478 287245
rect 674186 287205 674192 287217
rect 675472 287205 675478 287217
rect 675530 287205 675536 287257
rect 674224 286761 674230 286813
rect 674282 286801 674288 286813
rect 675376 286801 675382 286813
rect 674282 286773 675382 286801
rect 674282 286761 674288 286773
rect 675376 286761 675382 286773
rect 675434 286761 675440 286813
rect 39952 285355 39958 285407
rect 40010 285395 40016 285407
rect 43312 285395 43318 285407
rect 40010 285367 43318 285395
rect 40010 285355 40016 285367
rect 43312 285355 43318 285367
rect 43370 285355 43376 285407
rect 40048 285281 40054 285333
rect 40106 285321 40112 285333
rect 43120 285321 43126 285333
rect 40106 285293 43126 285321
rect 40106 285281 40112 285293
rect 43120 285281 43126 285293
rect 43178 285281 43184 285333
rect 40144 285207 40150 285259
rect 40202 285247 40208 285259
rect 43024 285247 43030 285259
rect 40202 285219 43030 285247
rect 40202 285207 40208 285219
rect 43024 285207 43030 285219
rect 43082 285207 43088 285259
rect 40240 285133 40246 285185
rect 40298 285173 40304 285185
rect 42928 285173 42934 285185
rect 40298 285145 42934 285173
rect 40298 285133 40304 285145
rect 42928 285133 42934 285145
rect 42986 285133 42992 285185
rect 45136 285133 45142 285185
rect 45194 285173 45200 285185
rect 58096 285173 58102 285185
rect 45194 285145 58102 285173
rect 45194 285133 45200 285145
rect 58096 285133 58102 285145
rect 58154 285133 58160 285185
rect 654064 284763 654070 284815
rect 654122 284803 654128 284815
rect 660880 284803 660886 284815
rect 654122 284775 660886 284803
rect 654122 284763 654128 284775
rect 660880 284763 660886 284775
rect 660938 284763 660944 284815
rect 42160 282913 42166 282965
rect 42218 282953 42224 282965
rect 42448 282953 42454 282965
rect 42218 282925 42454 282953
rect 42218 282913 42224 282925
rect 42448 282913 42454 282925
rect 42506 282913 42512 282965
rect 42160 281729 42166 281781
rect 42218 281769 42224 281781
rect 42352 281769 42358 281781
rect 42218 281741 42358 281769
rect 42218 281729 42224 281741
rect 42352 281729 42358 281741
rect 42410 281729 42416 281781
rect 42160 281063 42166 281115
rect 42218 281103 42224 281115
rect 53584 281103 53590 281115
rect 42218 281075 53590 281103
rect 42218 281063 42224 281075
rect 53584 281063 53590 281075
rect 53642 281063 53648 281115
rect 42160 279879 42166 279931
rect 42218 279919 42224 279931
rect 42928 279919 42934 279931
rect 42218 279891 42934 279919
rect 42218 279879 42224 279891
rect 42928 279879 42934 279891
rect 42986 279879 42992 279931
rect 42928 279731 42934 279783
rect 42986 279771 42992 279783
rect 43312 279771 43318 279783
rect 42986 279743 43318 279771
rect 42986 279731 42992 279743
rect 43312 279731 43318 279743
rect 43370 279731 43376 279783
rect 255202 278633 332798 278661
rect 64816 278547 64822 278599
rect 64874 278587 64880 278599
rect 67216 278587 67222 278599
rect 64874 278559 67222 278587
rect 64874 278547 64880 278559
rect 67216 278547 67222 278559
rect 67274 278547 67280 278599
rect 255202 278525 255230 278633
rect 332770 278599 332798 278633
rect 348802 278633 380798 278661
rect 348802 278599 348830 278633
rect 268144 278547 268150 278599
rect 268202 278587 268208 278599
rect 293776 278587 293782 278599
rect 268202 278559 293782 278587
rect 268202 278547 268208 278559
rect 293776 278547 293782 278559
rect 293834 278547 293840 278599
rect 299536 278547 299542 278599
rect 299594 278587 299600 278599
rect 330160 278587 330166 278599
rect 299594 278559 330166 278587
rect 299594 278547 299600 278559
rect 330160 278547 330166 278559
rect 330218 278547 330224 278599
rect 332752 278547 332758 278599
rect 332810 278547 332816 278599
rect 348784 278547 348790 278599
rect 348842 278547 348848 278599
rect 350320 278547 350326 278599
rect 350378 278587 350384 278599
rect 380656 278587 380662 278599
rect 350378 278559 380662 278587
rect 350378 278547 350384 278559
rect 380656 278547 380662 278559
rect 380714 278547 380720 278599
rect 255184 278473 255190 278525
rect 255242 278473 255248 278525
rect 287248 278473 287254 278525
rect 287306 278513 287312 278525
rect 335536 278513 335542 278525
rect 287306 278485 299870 278513
rect 287306 278473 287312 278485
rect 233776 278399 233782 278451
rect 233834 278439 233840 278451
rect 267760 278439 267766 278451
rect 233834 278411 267766 278439
rect 233834 278399 233840 278411
rect 267760 278399 267766 278411
rect 267818 278399 267824 278451
rect 267856 278399 267862 278451
rect 267914 278439 267920 278451
rect 268144 278439 268150 278451
rect 267914 278411 268150 278439
rect 267914 278399 267920 278411
rect 268144 278399 268150 278411
rect 268202 278399 268208 278451
rect 293776 278399 293782 278451
rect 293834 278439 293840 278451
rect 299728 278439 299734 278451
rect 293834 278411 299734 278439
rect 293834 278399 293840 278411
rect 299728 278399 299734 278411
rect 299786 278399 299792 278451
rect 293200 278325 293206 278377
rect 293258 278365 293264 278377
rect 299536 278365 299542 278377
rect 293258 278337 299542 278365
rect 293258 278325 293264 278337
rect 299536 278325 299542 278337
rect 299594 278325 299600 278377
rect 299842 278365 299870 278485
rect 300226 278485 335542 278513
rect 300226 278365 300254 278485
rect 335536 278473 335542 278485
rect 335594 278473 335600 278525
rect 380770 278513 380798 278633
rect 380866 278633 393854 278661
rect 380866 278599 380894 278633
rect 393826 278599 393854 278633
rect 380848 278547 380854 278599
rect 380906 278547 380912 278599
rect 381232 278547 381238 278599
rect 381290 278587 381296 278599
rect 390256 278587 390262 278599
rect 381290 278559 390262 278587
rect 381290 278547 381296 278559
rect 390256 278547 390262 278559
rect 390314 278547 390320 278599
rect 393808 278547 393814 278599
rect 393866 278547 393872 278599
rect 383056 278513 383062 278525
rect 380290 278485 380702 278513
rect 380770 278485 383062 278513
rect 300400 278399 300406 278451
rect 300458 278439 300464 278451
rect 380290 278439 380318 278485
rect 300458 278411 380318 278439
rect 380674 278439 380702 278485
rect 383056 278473 383062 278485
rect 383114 278473 383120 278525
rect 440656 278473 440662 278525
rect 440714 278513 440720 278525
rect 489616 278513 489622 278525
rect 440714 278485 489622 278513
rect 440714 278473 440720 278485
rect 489616 278473 489622 278485
rect 489674 278473 489680 278525
rect 495376 278473 495382 278525
rect 495434 278513 495440 278525
rect 501328 278513 501334 278525
rect 495434 278485 501334 278513
rect 495434 278473 495440 278485
rect 501328 278473 501334 278485
rect 501386 278473 501392 278525
rect 625072 278473 625078 278525
rect 625130 278513 625136 278525
rect 631024 278513 631030 278525
rect 625130 278485 631030 278513
rect 625130 278473 625136 278485
rect 631024 278473 631030 278485
rect 631082 278473 631088 278525
rect 380674 278411 382046 278439
rect 300458 278399 300464 278411
rect 299842 278337 300254 278365
rect 300304 278325 300310 278377
rect 300362 278365 300368 278377
rect 380272 278365 380278 278377
rect 300362 278337 380278 278365
rect 300362 278325 300368 278337
rect 380272 278325 380278 278337
rect 380330 278325 380336 278377
rect 380656 278325 380662 278377
rect 380714 278365 380720 278377
rect 381904 278365 381910 278377
rect 380714 278337 381910 278365
rect 380714 278325 380720 278337
rect 381904 278325 381910 278337
rect 381962 278325 381968 278377
rect 382018 278365 382046 278411
rect 397456 278399 397462 278451
rect 397514 278439 397520 278451
rect 417424 278439 417430 278451
rect 397514 278411 417430 278439
rect 397514 278399 397520 278411
rect 417424 278399 417430 278411
rect 417482 278399 417488 278451
rect 525520 278399 525526 278451
rect 525578 278439 525584 278451
rect 551248 278439 551254 278451
rect 525578 278411 551254 278439
rect 525578 278399 525584 278411
rect 551248 278399 551254 278411
rect 551306 278399 551312 278451
rect 610480 278399 610486 278451
rect 610538 278439 610544 278451
rect 610768 278439 610774 278451
rect 610538 278411 610774 278439
rect 610538 278399 610544 278411
rect 610768 278399 610774 278411
rect 610826 278399 610832 278451
rect 389008 278365 389014 278377
rect 382018 278337 389014 278365
rect 389008 278325 389014 278337
rect 389066 278325 389072 278377
rect 290800 278251 290806 278303
rect 290858 278291 290864 278303
rect 364144 278291 364150 278303
rect 290858 278263 364150 278291
rect 290858 278251 290864 278263
rect 364144 278251 364150 278263
rect 364202 278251 364208 278303
rect 365776 278251 365782 278303
rect 365834 278291 365840 278303
rect 368848 278291 368854 278303
rect 365834 278263 368854 278291
rect 365834 278251 365840 278263
rect 368848 278251 368854 278263
rect 368906 278251 368912 278303
rect 378256 278251 378262 278303
rect 378314 278291 378320 278303
rect 387760 278291 387766 278303
rect 378314 278263 387766 278291
rect 378314 278251 378320 278263
rect 387760 278251 387766 278263
rect 387818 278251 387824 278303
rect 396688 278251 396694 278303
rect 396746 278291 396752 278303
rect 440656 278291 440662 278303
rect 396746 278263 440662 278291
rect 396746 278251 396752 278263
rect 440656 278251 440662 278263
rect 440714 278251 440720 278303
rect 440752 278251 440758 278303
rect 440810 278291 440816 278303
rect 490192 278291 490198 278303
rect 440810 278263 490198 278291
rect 440810 278251 440816 278263
rect 490192 278251 490198 278263
rect 490250 278251 490256 278303
rect 294736 278177 294742 278229
rect 294794 278217 294800 278229
rect 299536 278217 299542 278229
rect 294794 278189 299542 278217
rect 294794 278177 294800 278189
rect 299536 278177 299542 278189
rect 299594 278177 299600 278229
rect 299824 278177 299830 278229
rect 299882 278217 299888 278229
rect 396208 278217 396214 278229
rect 299882 278189 396214 278217
rect 299882 278177 299888 278189
rect 396208 278177 396214 278189
rect 396266 278177 396272 278229
rect 240976 278103 240982 278155
rect 241034 278143 241040 278155
rect 241034 278115 299774 278143
rect 241034 278103 241040 278115
rect 266032 278029 266038 278081
rect 266090 278069 266096 278081
rect 299746 278069 299774 278115
rect 299920 278103 299926 278155
rect 299978 278143 299984 278155
rect 331312 278143 331318 278155
rect 299978 278115 331318 278143
rect 299978 278103 299984 278115
rect 331312 278103 331318 278115
rect 331370 278103 331376 278155
rect 352912 278103 352918 278155
rect 352970 278143 352976 278155
rect 352970 278115 357374 278143
rect 352970 278103 352976 278115
rect 299824 278069 299830 278081
rect 266090 278041 299678 278069
rect 299746 278041 299830 278069
rect 266090 278029 266096 278041
rect 299650 278007 299678 278041
rect 299824 278029 299830 278041
rect 299882 278029 299888 278081
rect 300400 278029 300406 278081
rect 300458 278069 300464 278081
rect 334384 278069 334390 278081
rect 300458 278041 334390 278069
rect 300458 278029 300464 278041
rect 334384 278029 334390 278041
rect 334442 278029 334448 278081
rect 353488 278029 353494 278081
rect 353546 278069 353552 278081
rect 357346 278069 357374 278115
rect 369616 278103 369622 278155
rect 369674 278143 369680 278155
rect 380176 278143 380182 278155
rect 369674 278115 380182 278143
rect 369674 278103 369680 278115
rect 380176 278103 380182 278115
rect 380234 278103 380240 278155
rect 380656 278103 380662 278155
rect 380714 278143 380720 278155
rect 390160 278143 390166 278155
rect 380714 278115 390166 278143
rect 380714 278103 380720 278115
rect 390160 278103 390166 278115
rect 390218 278103 390224 278155
rect 390256 278103 390262 278155
rect 390314 278143 390320 278155
rect 636496 278143 636502 278155
rect 390314 278115 636502 278143
rect 390314 278103 390320 278115
rect 636496 278103 636502 278115
rect 636554 278103 636560 278155
rect 415312 278069 415318 278081
rect 353546 278041 357182 278069
rect 357346 278041 415318 278069
rect 353546 278029 353552 278041
rect 223120 277955 223126 278007
rect 223178 277995 223184 278007
rect 299488 277995 299494 278007
rect 223178 277967 299494 277995
rect 223178 277955 223184 277967
rect 299488 277955 299494 277967
rect 299546 277955 299552 278007
rect 299632 277955 299638 278007
rect 299690 277955 299696 278007
rect 300304 277955 300310 278007
rect 300362 277995 300368 278007
rect 329104 277995 329110 278007
rect 300362 277967 329110 277995
rect 300362 277955 300368 277967
rect 329104 277955 329110 277967
rect 329162 277955 329168 278007
rect 355504 277955 355510 278007
rect 355562 277995 355568 278007
rect 357154 277995 357182 278041
rect 415312 278029 415318 278041
rect 415370 278029 415376 278081
rect 422320 277995 422326 278007
rect 355562 277967 357086 277995
rect 357154 277967 422326 277995
rect 355562 277955 355568 277967
rect 64912 277881 64918 277933
rect 64970 277921 64976 277933
rect 184336 277921 184342 277933
rect 64970 277893 184342 277921
rect 64970 277881 64976 277893
rect 184336 277881 184342 277893
rect 184394 277881 184400 277933
rect 291472 277881 291478 277933
rect 291530 277921 291536 277933
rect 356944 277921 356950 277933
rect 291530 277893 356950 277921
rect 291530 277881 291536 277893
rect 356944 277881 356950 277893
rect 357002 277881 357008 277933
rect 357058 277921 357086 277967
rect 422320 277955 422326 277967
rect 422378 277955 422384 278007
rect 436624 277921 436630 277933
rect 357058 277893 436630 277921
rect 436624 277881 436630 277893
rect 436682 277881 436688 277933
rect 42160 277807 42166 277859
rect 42218 277847 42224 277859
rect 43120 277847 43126 277859
rect 42218 277819 43126 277847
rect 42218 277807 42224 277819
rect 43120 277807 43126 277819
rect 43178 277807 43184 277859
rect 288400 277807 288406 277859
rect 288458 277847 288464 277859
rect 342736 277847 342742 277859
rect 288458 277819 342742 277847
rect 288458 277807 288464 277819
rect 342736 277807 342742 277819
rect 342794 277807 342800 277859
rect 356848 277807 356854 277859
rect 356906 277847 356912 277859
rect 450832 277847 450838 277859
rect 356906 277819 450838 277847
rect 356906 277807 356912 277819
rect 450832 277807 450838 277819
rect 450890 277807 450896 277859
rect 289936 277733 289942 277785
rect 289994 277773 290000 277785
rect 357040 277773 357046 277785
rect 289994 277745 357046 277773
rect 289994 277733 290000 277745
rect 357040 277733 357046 277745
rect 357098 277733 357104 277785
rect 358768 277733 358774 277785
rect 358826 277773 358832 277785
rect 465232 277773 465238 277785
rect 358826 277745 465238 277773
rect 358826 277733 358832 277745
rect 465232 277733 465238 277745
rect 465290 277733 465296 277785
rect 295792 277659 295798 277711
rect 295850 277699 295856 277711
rect 403600 277699 403606 277711
rect 295850 277671 403606 277699
rect 295850 277659 295856 277671
rect 403600 277659 403606 277671
rect 403658 277659 403664 277711
rect 296464 277585 296470 277637
rect 296522 277625 296528 277637
rect 410800 277625 410806 277637
rect 296522 277597 410806 277625
rect 296522 277585 296528 277597
rect 410800 277585 410806 277597
rect 410858 277585 410864 277637
rect 297520 277511 297526 277563
rect 297578 277551 297584 277563
rect 417904 277551 417910 277563
rect 297578 277523 417910 277551
rect 297578 277511 297584 277523
rect 417904 277511 417910 277523
rect 417962 277511 417968 277563
rect 292048 277437 292054 277489
rect 292106 277477 292112 277489
rect 375088 277477 375094 277489
rect 292106 277449 375094 277477
rect 292106 277437 292112 277449
rect 375088 277437 375094 277449
rect 375146 277437 375152 277489
rect 375184 277437 375190 277489
rect 375242 277477 375248 277489
rect 385168 277477 385174 277489
rect 375242 277449 385174 277477
rect 375242 277437 375248 277449
rect 385168 277437 385174 277449
rect 385226 277437 385232 277489
rect 42064 277363 42070 277415
rect 42122 277403 42128 277415
rect 43024 277403 43030 277415
rect 42122 277375 43030 277403
rect 42122 277363 42128 277375
rect 43024 277363 43030 277375
rect 43082 277363 43088 277415
rect 247888 277363 247894 277415
rect 247946 277403 247952 277415
rect 332176 277403 332182 277415
rect 247946 277375 332182 277403
rect 247946 277363 247952 277375
rect 332176 277363 332182 277375
rect 332234 277363 332240 277415
rect 363760 277363 363766 277415
rect 363818 277403 363824 277415
rect 378736 277403 378742 277415
rect 363818 277375 378742 277403
rect 363818 277363 363824 277375
rect 378736 277363 378742 277375
rect 378794 277363 378800 277415
rect 378832 277363 378838 277415
rect 378890 277403 378896 277415
rect 486832 277403 486838 277415
rect 378890 277375 486838 277403
rect 378890 277363 378896 277375
rect 486832 277363 486838 277375
rect 486890 277363 486896 277415
rect 298192 277289 298198 277341
rect 298250 277329 298256 277341
rect 425008 277329 425014 277341
rect 298250 277301 425014 277329
rect 298250 277289 298256 277301
rect 425008 277289 425014 277301
rect 425066 277289 425072 277341
rect 299056 277215 299062 277267
rect 299114 277255 299120 277267
rect 432208 277255 432214 277267
rect 299114 277227 432214 277255
rect 299114 277215 299120 277227
rect 432208 277215 432214 277227
rect 432266 277215 432272 277267
rect 314704 277141 314710 277193
rect 314762 277181 314768 277193
rect 328048 277181 328054 277193
rect 314762 277153 328054 277181
rect 314762 277141 314768 277153
rect 328048 277141 328054 277153
rect 328106 277141 328112 277193
rect 328144 277141 328150 277193
rect 328202 277181 328208 277193
rect 460720 277181 460726 277193
rect 328202 277153 460726 277181
rect 328202 277141 328208 277153
rect 460720 277141 460726 277153
rect 460778 277141 460784 277193
rect 225232 277067 225238 277119
rect 225290 277107 225296 277119
rect 273616 277107 273622 277119
rect 225290 277079 273622 277107
rect 225290 277067 225296 277079
rect 273616 277067 273622 277079
rect 273674 277067 273680 277119
rect 300208 277067 300214 277119
rect 300266 277107 300272 277119
rect 439312 277107 439318 277119
rect 300266 277079 439318 277107
rect 300266 277067 300272 277079
rect 439312 277067 439318 277079
rect 439370 277067 439376 277119
rect 301264 276993 301270 277045
rect 301322 277033 301328 277045
rect 338800 277033 338806 277045
rect 301322 277005 338806 277033
rect 301322 276993 301328 277005
rect 338800 276993 338806 277005
rect 338858 276993 338864 277045
rect 364816 276993 364822 277045
rect 364874 277033 364880 277045
rect 378640 277033 378646 277045
rect 364874 277005 378646 277033
rect 364874 276993 364880 277005
rect 378640 276993 378646 277005
rect 378698 276993 378704 277045
rect 378736 276993 378742 277045
rect 378794 277033 378800 277045
rect 504688 277033 504694 277045
rect 378794 277005 504694 277033
rect 378794 276993 378800 277005
rect 504688 276993 504694 277005
rect 504746 276993 504752 277045
rect 300784 276919 300790 276971
rect 300842 276959 300848 276971
rect 446512 276959 446518 276971
rect 300842 276931 446518 276959
rect 300842 276919 300848 276931
rect 446512 276919 446518 276931
rect 446570 276919 446576 276971
rect 289264 276845 289270 276897
rect 289322 276885 289328 276897
rect 350032 276885 350038 276897
rect 289322 276857 350038 276885
rect 289322 276845 289328 276857
rect 350032 276845 350038 276857
rect 350090 276845 350096 276897
rect 376624 276845 376630 276897
rect 376682 276885 376688 276897
rect 378544 276885 378550 276897
rect 376682 276857 378550 276885
rect 376682 276845 376688 276857
rect 378544 276845 378550 276857
rect 378602 276845 378608 276897
rect 378640 276845 378646 276897
rect 378698 276885 378704 276897
rect 515440 276885 515446 276897
rect 378698 276857 515446 276885
rect 378698 276845 378704 276857
rect 515440 276845 515446 276857
rect 515498 276845 515504 276897
rect 301840 276771 301846 276823
rect 301898 276811 301904 276823
rect 453520 276811 453526 276823
rect 301898 276783 453526 276811
rect 301898 276771 301904 276783
rect 453520 276771 453526 276783
rect 453578 276771 453584 276823
rect 215728 276697 215734 276749
rect 215786 276737 215792 276749
rect 314704 276737 314710 276749
rect 215786 276709 314710 276737
rect 215786 276697 215792 276709
rect 314704 276697 314710 276709
rect 314762 276697 314768 276749
rect 327376 276737 327382 276749
rect 317794 276709 327382 276737
rect 208528 276623 208534 276675
rect 208586 276663 208592 276675
rect 317794 276663 317822 276709
rect 327376 276697 327382 276709
rect 327434 276697 327440 276749
rect 349168 276697 349174 276749
rect 349226 276737 349232 276749
rect 366928 276737 366934 276749
rect 349226 276709 366934 276737
rect 349226 276697 349232 276709
rect 366928 276697 366934 276709
rect 366986 276697 366992 276749
rect 367024 276697 367030 276749
rect 367082 276737 367088 276749
rect 518992 276737 518998 276749
rect 367082 276709 518998 276737
rect 367082 276697 367088 276709
rect 518992 276697 518998 276709
rect 519050 276697 519056 276749
rect 208586 276635 317822 276663
rect 208586 276623 208592 276635
rect 324976 276623 324982 276675
rect 325034 276663 325040 276675
rect 365776 276663 365782 276675
rect 325034 276635 365782 276663
rect 325034 276623 325040 276635
rect 365776 276623 365782 276635
rect 365834 276623 365840 276675
rect 378832 276663 378838 276675
rect 365890 276635 378838 276663
rect 197872 276549 197878 276601
rect 197930 276589 197936 276601
rect 325840 276589 325846 276601
rect 197930 276561 325846 276589
rect 197930 276549 197936 276561
rect 325840 276549 325846 276561
rect 325898 276549 325904 276601
rect 325936 276549 325942 276601
rect 325994 276589 326000 276601
rect 328144 276589 328150 276601
rect 325994 276561 328150 276589
rect 325994 276549 326000 276561
rect 328144 276549 328150 276561
rect 328202 276549 328208 276601
rect 361552 276549 361558 276601
rect 361610 276589 361616 276601
rect 365890 276589 365918 276635
rect 378832 276623 378838 276635
rect 378890 276623 378896 276675
rect 378928 276623 378934 276675
rect 378986 276663 378992 276675
rect 378986 276635 387134 276663
rect 378986 276623 378992 276635
rect 361610 276561 365918 276589
rect 366850 276561 378686 276589
rect 361610 276549 361616 276561
rect 114640 276475 114646 276527
rect 114698 276515 114704 276527
rect 322096 276515 322102 276527
rect 114698 276487 322102 276515
rect 114698 276475 114704 276487
rect 322096 276475 322102 276487
rect 322154 276475 322160 276527
rect 327184 276515 327190 276527
rect 325378 276487 327190 276515
rect 230608 276401 230614 276453
rect 230666 276441 230672 276453
rect 325378 276441 325406 276487
rect 327184 276475 327190 276487
rect 327242 276475 327248 276527
rect 351088 276475 351094 276527
rect 351146 276515 351152 276527
rect 366850 276515 366878 276561
rect 351146 276487 366878 276515
rect 351146 276475 351152 276487
rect 366928 276475 366934 276527
rect 366986 276515 366992 276527
rect 378658 276515 378686 276561
rect 379024 276549 379030 276601
rect 379082 276589 379088 276601
rect 386992 276589 386998 276601
rect 379082 276561 386998 276589
rect 379082 276549 379088 276561
rect 386992 276549 386998 276561
rect 387050 276549 387056 276601
rect 387106 276589 387134 276635
rect 390160 276623 390166 276675
rect 390218 276663 390224 276675
rect 554704 276663 554710 276675
rect 390218 276635 554710 276663
rect 390218 276623 390224 276635
rect 554704 276623 554710 276635
rect 554762 276623 554768 276675
rect 611824 276589 611830 276601
rect 387106 276561 611830 276589
rect 611824 276549 611830 276561
rect 611882 276549 611888 276601
rect 401200 276515 401206 276527
rect 366986 276487 378590 276515
rect 378658 276487 401206 276515
rect 366986 276475 366992 276487
rect 230666 276413 325406 276441
rect 230666 276401 230672 276413
rect 325456 276401 325462 276453
rect 325514 276441 325520 276453
rect 372016 276441 372022 276453
rect 325514 276413 372022 276441
rect 325514 276401 325520 276413
rect 372016 276401 372022 276413
rect 372074 276401 372080 276453
rect 372112 276401 372118 276453
rect 372170 276441 372176 276453
rect 378448 276441 378454 276453
rect 372170 276413 378454 276441
rect 372170 276401 372176 276413
rect 378448 276401 378454 276413
rect 378506 276401 378512 276453
rect 378562 276441 378590 276487
rect 401200 276475 401206 276487
rect 401258 276475 401264 276527
rect 642256 276475 642262 276527
rect 642314 276515 642320 276527
rect 649552 276515 649558 276527
rect 642314 276487 649558 276515
rect 642314 276475 642320 276487
rect 649552 276475 649558 276487
rect 649610 276475 649616 276527
rect 379024 276441 379030 276453
rect 378562 276413 379030 276441
rect 379024 276401 379030 276413
rect 379082 276401 379088 276453
rect 379600 276401 379606 276453
rect 379658 276441 379664 276453
rect 398896 276441 398902 276453
rect 379658 276413 398902 276441
rect 379658 276401 379664 276413
rect 398896 276401 398902 276413
rect 398954 276401 398960 276453
rect 243760 276327 243766 276379
rect 243818 276367 243824 276379
rect 434512 276367 434518 276379
rect 243818 276339 434518 276367
rect 243818 276327 243824 276339
rect 434512 276327 434518 276339
rect 434570 276327 434576 276379
rect 231952 276253 231958 276305
rect 232010 276293 232016 276305
rect 338224 276293 338230 276305
rect 232010 276265 338230 276293
rect 232010 276253 232016 276265
rect 338224 276253 338230 276265
rect 338282 276253 338288 276305
rect 346480 276253 346486 276305
rect 346538 276293 346544 276305
rect 365584 276293 365590 276305
rect 346538 276265 365590 276293
rect 346538 276253 346544 276265
rect 365584 276253 365590 276265
rect 365642 276253 365648 276305
rect 372208 276253 372214 276305
rect 372266 276293 372272 276305
rect 382960 276293 382966 276305
rect 372266 276265 382966 276293
rect 372266 276253 372272 276265
rect 382960 276253 382966 276265
rect 383018 276253 383024 276305
rect 383056 276253 383062 276305
rect 383114 276293 383120 276305
rect 383114 276265 385118 276293
rect 383114 276253 383120 276265
rect 232336 276179 232342 276231
rect 232394 276219 232400 276231
rect 341776 276219 341782 276231
rect 232394 276191 341782 276219
rect 232394 276179 232400 276191
rect 341776 276179 341782 276191
rect 341834 276179 341840 276231
rect 348400 276179 348406 276231
rect 348458 276219 348464 276231
rect 379888 276219 379894 276231
rect 348458 276191 379894 276219
rect 348458 276179 348464 276191
rect 379888 276179 379894 276191
rect 379946 276179 379952 276231
rect 379984 276179 379990 276231
rect 380042 276219 380048 276231
rect 384976 276219 384982 276231
rect 380042 276191 384982 276219
rect 380042 276179 380048 276191
rect 384976 276179 384982 276191
rect 385034 276179 385040 276231
rect 385090 276219 385118 276265
rect 385168 276253 385174 276305
rect 385226 276293 385232 276305
rect 565456 276293 565462 276305
rect 385226 276265 565462 276293
rect 385226 276253 385232 276265
rect 565456 276253 565462 276265
rect 565514 276253 565520 276305
rect 572464 276219 572470 276231
rect 385090 276191 572470 276219
rect 572464 276179 572470 276191
rect 572522 276179 572528 276231
rect 244720 276105 244726 276157
rect 244778 276145 244784 276157
rect 441712 276145 441718 276157
rect 244778 276117 441718 276145
rect 244778 276105 244784 276117
rect 441712 276105 441718 276117
rect 441770 276105 441776 276157
rect 245392 276031 245398 276083
rect 245450 276071 245456 276083
rect 448816 276071 448822 276083
rect 245450 276043 448822 276071
rect 245450 276031 245456 276043
rect 448816 276031 448822 276043
rect 448874 276031 448880 276083
rect 246352 275957 246358 276009
rect 246410 275997 246416 276009
rect 455920 275997 455926 276009
rect 246410 275969 455926 275997
rect 246410 275957 246416 275969
rect 455920 275957 455926 275969
rect 455978 275957 455984 276009
rect 233488 275883 233494 275935
rect 233546 275923 233552 275935
rect 348976 275923 348982 275935
rect 233546 275895 348982 275923
rect 233546 275883 233552 275895
rect 348976 275883 348982 275895
rect 349034 275883 349040 275935
rect 369520 275883 369526 275935
rect 369578 275923 369584 275935
rect 384880 275923 384886 275935
rect 369578 275895 384886 275923
rect 369578 275883 369584 275895
rect 384880 275883 384886 275895
rect 384938 275883 384944 275935
rect 384976 275883 384982 275935
rect 385034 275923 385040 275935
rect 579664 275923 579670 275935
rect 385034 275895 579670 275923
rect 385034 275883 385040 275895
rect 579664 275883 579670 275895
rect 579722 275883 579728 275935
rect 247408 275809 247414 275861
rect 247466 275849 247472 275861
rect 463120 275849 463126 275861
rect 247466 275821 463126 275849
rect 247466 275809 247472 275821
rect 463120 275809 463126 275821
rect 463178 275809 463184 275861
rect 227440 275735 227446 275787
rect 227498 275775 227504 275787
rect 298960 275775 298966 275787
rect 227498 275747 298966 275775
rect 227498 275735 227504 275747
rect 298960 275735 298966 275747
rect 299018 275735 299024 275787
rect 311536 275735 311542 275787
rect 311594 275775 311600 275787
rect 532144 275775 532150 275787
rect 311594 275747 532150 275775
rect 311594 275735 311600 275747
rect 532144 275735 532150 275747
rect 532202 275735 532208 275787
rect 248080 275661 248086 275713
rect 248138 275701 248144 275713
rect 470224 275701 470230 275713
rect 248138 275673 470230 275701
rect 248138 275661 248144 275673
rect 470224 275661 470230 275673
rect 470282 275661 470288 275713
rect 234064 275587 234070 275639
rect 234122 275627 234128 275639
rect 356080 275627 356086 275639
rect 234122 275599 356086 275627
rect 234122 275587 234128 275599
rect 356080 275587 356086 275599
rect 356138 275587 356144 275639
rect 364240 275587 364246 275639
rect 364298 275627 364304 275639
rect 378736 275627 378742 275639
rect 364298 275599 378742 275627
rect 364298 275587 364304 275599
rect 378736 275587 378742 275599
rect 378794 275587 378800 275639
rect 378832 275587 378838 275639
rect 378890 275627 378896 275639
rect 601072 275627 601078 275639
rect 378890 275599 601078 275627
rect 378890 275587 378896 275599
rect 601072 275587 601078 275599
rect 601130 275587 601136 275639
rect 249136 275513 249142 275565
rect 249194 275553 249200 275565
rect 477424 275553 477430 275565
rect 249194 275525 477430 275553
rect 249194 275513 249200 275525
rect 477424 275513 477430 275525
rect 477482 275513 477488 275565
rect 42256 275439 42262 275491
rect 42314 275479 42320 275491
rect 42928 275479 42934 275491
rect 42314 275451 42934 275479
rect 42314 275439 42320 275451
rect 42928 275439 42934 275451
rect 42986 275439 42992 275491
rect 196720 275439 196726 275491
rect 196778 275479 196784 275491
rect 270256 275479 270262 275491
rect 196778 275451 270262 275479
rect 196778 275439 196784 275451
rect 270256 275439 270262 275451
rect 270314 275439 270320 275491
rect 322576 275439 322582 275491
rect 322634 275479 322640 275491
rect 564208 275479 564214 275491
rect 322634 275451 564214 275479
rect 322634 275439 322640 275451
rect 564208 275439 564214 275451
rect 564266 275439 564272 275491
rect 235024 275365 235030 275417
rect 235082 275405 235088 275417
rect 363184 275405 363190 275417
rect 235082 275377 363190 275405
rect 235082 275365 235088 275377
rect 363184 275365 363190 275377
rect 363242 275365 363248 275417
rect 368560 275365 368566 275417
rect 368618 275405 368624 275417
rect 372976 275405 372982 275417
rect 368618 275377 372982 275405
rect 368618 275365 368624 275377
rect 372976 275365 372982 275377
rect 373034 275365 373040 275417
rect 375568 275365 375574 275417
rect 375626 275405 375632 275417
rect 378832 275405 378838 275417
rect 375626 275377 378838 275405
rect 375626 275365 375632 275377
rect 378832 275365 378838 275377
rect 378890 275365 378896 275417
rect 378928 275365 378934 275417
rect 378986 275405 378992 275417
rect 379984 275405 379990 275417
rect 378986 275377 379990 275405
rect 378986 275365 378992 275377
rect 379984 275365 379990 275377
rect 380042 275365 380048 275417
rect 380944 275365 380950 275417
rect 381002 275405 381008 275417
rect 381002 275377 384734 275405
rect 381002 275365 381008 275377
rect 235984 275291 235990 275343
rect 236042 275331 236048 275343
rect 370288 275331 370294 275343
rect 236042 275303 370294 275331
rect 236042 275291 236048 275303
rect 370288 275291 370294 275303
rect 370346 275291 370352 275343
rect 372592 275291 372598 275343
rect 372650 275331 372656 275343
rect 384592 275331 384598 275343
rect 372650 275303 384598 275331
rect 372650 275291 372656 275303
rect 384592 275291 384598 275303
rect 384650 275291 384656 275343
rect 384706 275331 384734 275377
rect 384784 275365 384790 275417
rect 384842 275405 384848 275417
rect 622480 275405 622486 275417
rect 384842 275377 622486 275405
rect 384842 275365 384848 275377
rect 622480 275365 622486 275377
rect 622538 275365 622544 275417
rect 398800 275331 398806 275343
rect 384706 275303 398806 275331
rect 398800 275291 398806 275303
rect 398858 275291 398864 275343
rect 398896 275291 398902 275343
rect 398954 275331 398960 275343
rect 633136 275331 633142 275343
rect 398954 275303 633142 275331
rect 398954 275291 398960 275303
rect 633136 275291 633142 275303
rect 633194 275291 633200 275343
rect 200176 275217 200182 275269
rect 200234 275257 200240 275269
rect 270832 275257 270838 275269
rect 200234 275229 270838 275257
rect 200234 275217 200240 275229
rect 270832 275217 270838 275229
rect 270890 275217 270896 275269
rect 284944 275217 284950 275269
rect 285002 275257 285008 275269
rect 314416 275257 314422 275269
rect 285002 275229 314422 275257
rect 285002 275217 285008 275229
rect 314416 275217 314422 275229
rect 314474 275217 314480 275269
rect 316624 275217 316630 275269
rect 316682 275257 316688 275269
rect 571312 275257 571318 275269
rect 316682 275229 571318 275257
rect 316682 275217 316688 275229
rect 571312 275217 571318 275229
rect 571370 275217 571376 275269
rect 228016 275143 228022 275195
rect 228074 275183 228080 275195
rect 306064 275183 306070 275195
rect 228074 275155 306070 275183
rect 228074 275143 228080 275155
rect 306064 275143 306070 275155
rect 306122 275143 306128 275195
rect 316912 275143 316918 275195
rect 316970 275183 316976 275195
rect 578512 275183 578518 275195
rect 316970 275155 578518 275183
rect 316970 275143 316976 275155
rect 578512 275143 578518 275155
rect 578570 275143 578576 275195
rect 236752 275069 236758 275121
rect 236810 275109 236816 275121
rect 377488 275109 377494 275121
rect 236810 275081 377494 275109
rect 236810 275069 236816 275081
rect 377488 275069 377494 275081
rect 377546 275069 377552 275121
rect 377680 275069 377686 275121
rect 377738 275109 377744 275121
rect 397456 275109 397462 275121
rect 377738 275081 397462 275109
rect 377738 275069 377744 275081
rect 397456 275069 397462 275081
rect 397514 275069 397520 275121
rect 398800 275069 398806 275121
rect 398858 275109 398864 275121
rect 647536 275109 647542 275121
rect 398858 275081 647542 275109
rect 398858 275069 398864 275081
rect 647536 275069 647542 275081
rect 647594 275069 647600 275121
rect 229072 274995 229078 275047
rect 229130 275035 229136 275047
rect 313264 275035 313270 275047
rect 229130 275007 313270 275035
rect 229130 274995 229136 275007
rect 313264 274995 313270 275007
rect 313322 274995 313328 275047
rect 317968 274995 317974 275047
rect 318026 275035 318032 275047
rect 585616 275035 585622 275047
rect 318026 275007 585622 275035
rect 318026 274995 318032 275007
rect 585616 274995 585622 275007
rect 585674 274995 585680 275047
rect 242992 274921 242998 274973
rect 243050 274961 243056 274973
rect 427408 274961 427414 274973
rect 243050 274933 427414 274961
rect 243050 274921 243056 274933
rect 427408 274921 427414 274933
rect 427466 274921 427472 274973
rect 258544 274847 258550 274899
rect 258602 274887 258608 274899
rect 333136 274887 333142 274899
rect 258602 274859 333142 274887
rect 258602 274847 258608 274859
rect 333136 274847 333142 274859
rect 333194 274847 333200 274899
rect 368080 274847 368086 274899
rect 368138 274887 368144 274899
rect 378640 274887 378646 274899
rect 368138 274859 378646 274887
rect 368138 274847 368144 274859
rect 378640 274847 378646 274859
rect 378698 274847 378704 274899
rect 378736 274847 378742 274899
rect 378794 274887 378800 274899
rect 384784 274887 384790 274899
rect 378794 274859 384790 274887
rect 378794 274847 378800 274859
rect 384784 274847 384790 274859
rect 384842 274847 384848 274899
rect 384880 274847 384886 274899
rect 384938 274887 384944 274899
rect 551056 274887 551062 274899
rect 384938 274859 551062 274887
rect 384938 274847 384944 274859
rect 551056 274847 551062 274859
rect 551114 274847 551120 274899
rect 242224 274773 242230 274825
rect 242282 274813 242288 274825
rect 420208 274813 420214 274825
rect 242282 274785 420214 274813
rect 242282 274773 242288 274785
rect 420208 274773 420214 274785
rect 420266 274773 420272 274825
rect 241072 274699 241078 274751
rect 241130 274739 241136 274751
rect 413200 274739 413206 274751
rect 241130 274711 413206 274739
rect 241130 274699 241136 274711
rect 413200 274699 413206 274711
rect 413258 274699 413264 274751
rect 223024 274625 223030 274677
rect 223082 274665 223088 274677
rect 263344 274665 263350 274677
rect 223082 274637 263350 274665
rect 223082 274625 223088 274637
rect 263344 274625 263350 274637
rect 263402 274625 263408 274677
rect 269200 274625 269206 274677
rect 269258 274665 269264 274677
rect 334480 274665 334486 274677
rect 269258 274637 334486 274665
rect 269258 274625 269264 274637
rect 334480 274625 334486 274637
rect 334538 274625 334544 274677
rect 370960 274625 370966 274677
rect 371018 274665 371024 274677
rect 375184 274665 375190 274677
rect 371018 274637 375190 274665
rect 371018 274625 371024 274637
rect 375184 274625 375190 274637
rect 375242 274625 375248 274677
rect 375952 274625 375958 274677
rect 376010 274665 376016 274677
rect 378352 274665 378358 274677
rect 376010 274637 378358 274665
rect 376010 274625 376016 274637
rect 378352 274625 378358 274637
rect 378410 274625 378416 274677
rect 378640 274625 378646 274677
rect 378698 274665 378704 274677
rect 540400 274665 540406 274677
rect 378698 274637 540406 274665
rect 378698 274625 378704 274637
rect 540400 274625 540406 274637
rect 540458 274625 540464 274677
rect 240496 274551 240502 274603
rect 240554 274591 240560 274603
rect 406000 274591 406006 274603
rect 240554 274563 406006 274591
rect 240554 274551 240560 274563
rect 406000 274551 406006 274563
rect 406058 274551 406064 274603
rect 239344 274477 239350 274529
rect 239402 274517 239408 274529
rect 398608 274517 398614 274529
rect 239402 274489 398614 274517
rect 239402 274477 239408 274489
rect 398608 274477 398614 274489
rect 398666 274477 398672 274529
rect 238480 274403 238486 274455
rect 238538 274443 238544 274455
rect 372784 274443 372790 274455
rect 238538 274415 372790 274443
rect 238538 274403 238544 274415
rect 372784 274403 372790 274415
rect 372842 274403 372848 274455
rect 372880 274403 372886 274455
rect 372938 274443 372944 274455
rect 378640 274443 378646 274455
rect 372938 274415 378646 274443
rect 372938 274403 372944 274415
rect 378640 274403 378646 274415
rect 378698 274403 378704 274455
rect 379024 274403 379030 274455
rect 379082 274443 379088 274455
rect 398896 274443 398902 274455
rect 379082 274415 398902 274443
rect 379082 274403 379088 274415
rect 398896 274403 398902 274415
rect 398954 274403 398960 274455
rect 237808 274329 237814 274381
rect 237866 274369 237872 274381
rect 372592 274369 372598 274381
rect 237866 274341 372598 274369
rect 237866 274329 237872 274341
rect 372592 274329 372598 274341
rect 372650 274329 372656 274381
rect 372976 274329 372982 274381
rect 373034 274369 373040 274381
rect 381616 274369 381622 274381
rect 373034 274341 381622 274369
rect 373034 274329 373040 274341
rect 381616 274329 381622 274341
rect 381674 274329 381680 274381
rect 382768 274329 382774 274381
rect 382826 274369 382832 274381
rect 400048 274369 400054 274381
rect 382826 274341 400054 274369
rect 382826 274329 382832 274341
rect 400048 274329 400054 274341
rect 400106 274329 400112 274381
rect 408976 274329 408982 274381
rect 409034 274369 409040 274381
rect 449296 274369 449302 274381
rect 409034 274341 449302 274369
rect 409034 274329 409040 274341
rect 449296 274329 449302 274341
rect 449354 274329 449360 274381
rect 226288 274255 226294 274307
rect 226346 274295 226352 274307
rect 291856 274295 291862 274307
rect 226346 274267 291862 274295
rect 226346 274255 226352 274267
rect 291856 274255 291862 274267
rect 291914 274255 291920 274307
rect 297808 274255 297814 274307
rect 297866 274295 297872 274307
rect 337936 274295 337942 274307
rect 297866 274267 337942 274295
rect 297866 274255 297872 274267
rect 337936 274255 337942 274267
rect 337994 274255 338000 274307
rect 358288 274255 358294 274307
rect 358346 274295 358352 274307
rect 378640 274295 378646 274307
rect 358346 274267 378646 274295
rect 358346 274255 358352 274267
rect 378640 274255 378646 274267
rect 378698 274255 378704 274307
rect 378736 274255 378742 274307
rect 378794 274295 378800 274307
rect 383536 274295 383542 274307
rect 378794 274267 383542 274295
rect 378794 274255 378800 274267
rect 383536 274255 383542 274267
rect 383594 274255 383600 274307
rect 385072 274255 385078 274307
rect 385130 274295 385136 274307
rect 390544 274295 390550 274307
rect 385130 274267 390550 274295
rect 385130 274255 385136 274267
rect 390544 274255 390550 274267
rect 390602 274255 390608 274307
rect 511888 274295 511894 274307
rect 391810 274267 511894 274295
rect 184336 274181 184342 274233
rect 184394 274221 184400 274233
rect 200080 274221 200086 274233
rect 184394 274193 200086 274221
rect 184394 274181 184400 274193
rect 200080 274181 200086 274193
rect 200138 274181 200144 274233
rect 207376 274181 207382 274233
rect 207434 274221 207440 274233
rect 271312 274221 271318 274233
rect 207434 274193 271318 274221
rect 207434 274181 207440 274193
rect 271312 274181 271318 274193
rect 271370 274181 271376 274233
rect 271408 274181 271414 274233
rect 271466 274221 271472 274233
rect 271466 274193 272606 274221
rect 271466 274181 271472 274193
rect 214576 274107 214582 274159
rect 214634 274147 214640 274159
rect 272464 274147 272470 274159
rect 214634 274119 272470 274147
rect 214634 274107 214640 274119
rect 272464 274107 272470 274119
rect 272522 274107 272528 274159
rect 272578 274147 272606 274193
rect 276400 274181 276406 274233
rect 276458 274221 276464 274233
rect 335632 274221 335638 274233
rect 276458 274193 335638 274221
rect 276458 274181 276464 274193
rect 335632 274181 335638 274193
rect 335690 274181 335696 274233
rect 364336 274181 364342 274233
rect 364394 274221 364400 274233
rect 391810 274221 391838 274267
rect 511888 274255 511894 274267
rect 511946 274255 511952 274307
rect 645712 274255 645718 274307
rect 645770 274295 645776 274307
rect 649456 274295 649462 274307
rect 645770 274267 649462 274295
rect 645770 274255 645776 274267
rect 649456 274255 649462 274267
rect 649514 274255 649520 274307
rect 364394 274193 391838 274221
rect 364394 274181 364400 274193
rect 398896 274181 398902 274233
rect 398954 274221 398960 274233
rect 408976 274221 408982 274233
rect 398954 274193 408982 274221
rect 398954 274181 398960 274193
rect 408976 274181 408982 274193
rect 409034 274181 409040 274233
rect 449296 274181 449302 274233
rect 449354 274221 449360 274233
rect 469456 274221 469462 274233
rect 449354 274193 469462 274221
rect 449354 274181 449360 274193
rect 469456 274181 469462 274193
rect 469514 274181 469520 274233
rect 272578 274119 284990 274147
rect 225424 274033 225430 274085
rect 225482 274073 225488 274085
rect 284656 274073 284662 274085
rect 225482 274045 284662 274073
rect 225482 274033 225488 274045
rect 284656 274033 284662 274045
rect 284714 274033 284720 274085
rect 225232 273959 225238 274011
rect 225290 273999 225296 274011
rect 281104 273999 281110 274011
rect 225290 273971 281110 273999
rect 225290 273959 225296 273971
rect 281104 273959 281110 273971
rect 281162 273959 281168 274011
rect 284962 273999 284990 274119
rect 287056 274107 287062 274159
rect 287114 274147 287120 274159
rect 337072 274147 337078 274159
rect 287114 274119 337078 274147
rect 287114 274107 287120 274119
rect 337072 274107 337078 274119
rect 337130 274107 337136 274159
rect 360496 274107 360502 274159
rect 360554 274147 360560 274159
rect 479728 274147 479734 274159
rect 360554 274119 479734 274147
rect 360554 274107 360560 274119
rect 479728 274107 479734 274119
rect 479786 274107 479792 274159
rect 286672 274033 286678 274085
rect 286730 274073 286736 274085
rect 328720 274073 328726 274085
rect 286730 274045 328726 274073
rect 286730 274033 286736 274045
rect 328720 274033 328726 274045
rect 328778 274033 328784 274085
rect 360016 274033 360022 274085
rect 360074 274073 360080 274085
rect 476176 274073 476182 274085
rect 360074 274045 476182 274073
rect 360074 274033 360080 274045
rect 476176 274033 476182 274045
rect 476234 274033 476240 274085
rect 284962 273971 287966 273999
rect 239440 273885 239446 273937
rect 239498 273925 239504 273937
rect 275248 273925 275254 273937
rect 239498 273897 275254 273925
rect 239498 273885 239504 273897
rect 275248 273885 275254 273897
rect 275306 273885 275312 273937
rect 287938 273925 287966 273971
rect 304912 273959 304918 274011
rect 304970 273999 304976 274011
rect 338896 273999 338902 274011
rect 304970 273971 338902 273999
rect 304970 273959 304976 273971
rect 338896 273959 338902 273971
rect 338954 273959 338960 274011
rect 374320 273999 374326 274011
rect 349186 273971 374326 273999
rect 349186 273925 349214 273971
rect 374320 273959 374326 273971
rect 374378 273959 374384 274011
rect 378544 273999 378550 274011
rect 374434 273971 378550 273999
rect 287938 273897 349214 273925
rect 352240 273885 352246 273937
rect 352298 273925 352304 273937
rect 365872 273925 365878 273937
rect 352298 273897 365878 273925
rect 352298 273885 352304 273897
rect 365872 273885 365878 273897
rect 365930 273885 365936 273937
rect 370288 273885 370294 273937
rect 370346 273925 370352 273937
rect 374434 273925 374462 273971
rect 378544 273959 378550 273971
rect 378602 273959 378608 274011
rect 378640 273959 378646 274011
rect 378698 273999 378704 274011
rect 461968 273999 461974 274011
rect 378698 273971 461974 273999
rect 378698 273959 378704 273971
rect 461968 273959 461974 273971
rect 462026 273959 462032 274011
rect 469456 273959 469462 274011
rect 469514 273999 469520 274011
rect 508336 273999 508342 274011
rect 469514 273971 508342 273999
rect 469514 273959 469520 273971
rect 508336 273959 508342 273971
rect 508394 273959 508400 274011
rect 370346 273897 374462 273925
rect 370346 273885 370352 273897
rect 375664 273885 375670 273937
rect 375722 273925 375728 273937
rect 383440 273925 383446 273937
rect 375722 273897 383446 273925
rect 375722 273885 375728 273897
rect 383440 273885 383446 273897
rect 383498 273885 383504 273937
rect 383536 273885 383542 273937
rect 383594 273925 383600 273937
rect 558256 273925 558262 273937
rect 383594 273897 558262 273925
rect 383594 273885 383600 273897
rect 558256 273885 558262 273897
rect 558314 273885 558320 273937
rect 232432 273811 232438 273863
rect 232490 273851 232496 273863
rect 274672 273851 274678 273863
rect 232490 273823 274678 273851
rect 232490 273811 232496 273823
rect 274672 273811 274678 273823
rect 274730 273811 274736 273863
rect 308848 273811 308854 273863
rect 308906 273851 308912 273863
rect 308906 273823 329726 273851
rect 308906 273811 308912 273823
rect 229744 273737 229750 273789
rect 229802 273777 229808 273789
rect 320080 273777 320086 273789
rect 229802 273749 320086 273777
rect 229802 273737 229808 273749
rect 320080 273737 320086 273749
rect 320138 273737 320144 273789
rect 329698 273777 329726 273823
rect 356176 273811 356182 273863
rect 356234 273851 356240 273863
rect 444112 273851 444118 273863
rect 356234 273823 444118 273851
rect 356234 273811 356240 273823
rect 444112 273811 444118 273823
rect 444170 273811 444176 273863
rect 365104 273777 365110 273789
rect 329698 273749 365110 273777
rect 365104 273737 365110 273749
rect 365162 273737 365168 273789
rect 365200 273737 365206 273789
rect 365258 273777 365264 273789
rect 382384 273777 382390 273789
rect 365258 273749 382390 273777
rect 365258 273737 365264 273749
rect 382384 273737 382390 273749
rect 382442 273737 382448 273789
rect 382480 273737 382486 273789
rect 382538 273777 382544 273789
rect 383152 273777 383158 273789
rect 382538 273749 383158 273777
rect 382538 273737 382544 273749
rect 383152 273737 383158 273749
rect 383210 273737 383216 273789
rect 383248 273737 383254 273789
rect 383306 273777 383312 273789
rect 391696 273777 391702 273789
rect 383306 273749 391702 273777
rect 383306 273737 383312 273749
rect 391696 273737 391702 273749
rect 391754 273737 391760 273789
rect 403120 273737 403126 273789
rect 403178 273777 403184 273789
rect 417328 273777 417334 273789
rect 403178 273749 417334 273777
rect 403178 273737 403184 273749
rect 417328 273737 417334 273749
rect 417386 273737 417392 273789
rect 231760 273663 231766 273715
rect 231818 273703 231824 273715
rect 325456 273703 325462 273715
rect 231818 273675 325462 273703
rect 231818 273663 231824 273675
rect 325456 273663 325462 273675
rect 325514 273663 325520 273715
rect 354448 273663 354454 273715
rect 354506 273703 354512 273715
rect 429808 273703 429814 273715
rect 354506 273675 429814 273703
rect 354506 273663 354512 273675
rect 429808 273663 429814 273675
rect 429866 273663 429872 273715
rect 262672 273589 262678 273641
rect 262730 273629 262736 273641
rect 365776 273629 365782 273641
rect 262730 273601 365782 273629
rect 262730 273589 262736 273601
rect 365776 273589 365782 273601
rect 365834 273589 365840 273641
rect 365872 273589 365878 273641
rect 365930 273629 365936 273641
rect 411952 273629 411958 273641
rect 365930 273601 411958 273629
rect 365930 273589 365936 273601
rect 411952 273589 411958 273601
rect 412010 273589 412016 273641
rect 67216 273515 67222 273567
rect 67274 273555 67280 273567
rect 79024 273555 79030 273567
rect 67274 273527 79030 273555
rect 67274 273515 67280 273527
rect 79024 273515 79030 273527
rect 79082 273515 79088 273567
rect 153808 273515 153814 273567
rect 153866 273555 153872 273567
rect 163120 273555 163126 273567
rect 153866 273527 163126 273555
rect 153866 273515 153872 273527
rect 163120 273515 163126 273527
rect 163178 273515 163184 273567
rect 165808 273515 165814 273567
rect 165866 273555 165872 273567
rect 166960 273555 166966 273567
rect 165866 273527 166966 273555
rect 165866 273515 165872 273527
rect 166960 273515 166966 273527
rect 167018 273515 167024 273567
rect 170512 273515 170518 273567
rect 170570 273555 170576 273567
rect 172720 273555 172726 273567
rect 170570 273527 172726 273555
rect 170570 273515 170576 273527
rect 172720 273515 172726 273527
rect 172778 273515 172784 273567
rect 174064 273515 174070 273567
rect 174122 273555 174128 273567
rect 175504 273555 175510 273567
rect 174122 273527 175510 273555
rect 174122 273515 174128 273527
rect 175504 273515 175510 273527
rect 175562 273515 175568 273567
rect 177616 273515 177622 273567
rect 177674 273555 177680 273567
rect 178384 273555 178390 273567
rect 177674 273527 178390 273555
rect 177674 273515 177680 273527
rect 178384 273515 178390 273527
rect 178442 273515 178448 273567
rect 180016 273515 180022 273567
rect 180074 273555 180080 273567
rect 181360 273555 181366 273567
rect 180074 273527 181366 273555
rect 180074 273515 180080 273527
rect 181360 273515 181366 273527
rect 181418 273515 181424 273567
rect 184720 273515 184726 273567
rect 184778 273555 184784 273567
rect 187024 273555 187030 273567
rect 184778 273527 187030 273555
rect 184778 273515 184784 273527
rect 187024 273515 187030 273527
rect 187082 273515 187088 273567
rect 198640 273515 198646 273567
rect 198698 273555 198704 273567
rect 212368 273555 212374 273567
rect 198698 273527 212374 273555
rect 198698 273515 198704 273527
rect 212368 273515 212374 273527
rect 212426 273515 212432 273567
rect 257872 273515 257878 273567
rect 257930 273555 257936 273567
rect 282448 273555 282454 273567
rect 257930 273527 282454 273555
rect 257930 273515 257936 273527
rect 282448 273515 282454 273527
rect 282506 273515 282512 273567
rect 315376 273515 315382 273567
rect 315434 273555 315440 273567
rect 322576 273555 322582 273567
rect 315434 273527 322582 273555
rect 315434 273515 315440 273527
rect 322576 273515 322582 273527
rect 322634 273515 322640 273567
rect 322672 273515 322678 273567
rect 322730 273555 322736 273567
rect 325264 273555 325270 273567
rect 322730 273527 325270 273555
rect 322730 273515 322736 273527
rect 325264 273515 325270 273527
rect 325322 273515 325328 273567
rect 325456 273515 325462 273567
rect 325514 273555 325520 273567
rect 334576 273555 334582 273567
rect 325514 273527 334582 273555
rect 325514 273515 325520 273527
rect 334576 273515 334582 273527
rect 334634 273515 334640 273567
rect 340624 273515 340630 273567
rect 340682 273555 340688 273567
rect 343504 273555 343510 273567
rect 340682 273527 343510 273555
rect 340682 273515 340688 273527
rect 343504 273515 343510 273527
rect 343562 273515 343568 273567
rect 344656 273515 344662 273567
rect 344714 273555 344720 273567
rect 347728 273555 347734 273567
rect 344714 273527 347734 273555
rect 344714 273515 344720 273527
rect 347728 273515 347734 273527
rect 347786 273515 347792 273567
rect 356944 273515 356950 273567
rect 357002 273555 357008 273567
rect 367888 273555 367894 273567
rect 357002 273527 367894 273555
rect 357002 273515 357008 273527
rect 367888 273515 367894 273527
rect 367946 273515 367952 273567
rect 374128 273515 374134 273567
rect 374186 273555 374192 273567
rect 378064 273555 378070 273567
rect 374186 273527 378070 273555
rect 374186 273515 374192 273527
rect 378064 273515 378070 273527
rect 378122 273515 378128 273567
rect 378352 273515 378358 273567
rect 378410 273555 378416 273567
rect 396208 273555 396214 273567
rect 378410 273527 396214 273555
rect 378410 273515 378416 273527
rect 396208 273515 396214 273527
rect 396266 273515 396272 273567
rect 397360 273515 397366 273567
rect 397418 273555 397424 273567
rect 595120 273555 595126 273567
rect 397418 273527 595126 273555
rect 397418 273515 397424 273527
rect 595120 273515 595126 273527
rect 595178 273515 595184 273567
rect 91984 273441 91990 273493
rect 92042 273481 92048 273493
rect 206032 273481 206038 273493
rect 92042 273453 206038 273481
rect 92042 273441 92048 273453
rect 206032 273441 206038 273453
rect 206090 273441 206096 273493
rect 224560 273441 224566 273493
rect 224618 273481 224624 273493
rect 271504 273481 271510 273493
rect 224618 273453 271510 273481
rect 224618 273441 224624 273453
rect 271504 273441 271510 273453
rect 271562 273441 271568 273493
rect 271600 273441 271606 273493
rect 271658 273481 271664 273493
rect 279472 273481 279478 273493
rect 271658 273453 279478 273481
rect 271658 273441 271664 273453
rect 279472 273441 279478 273453
rect 279530 273441 279536 273493
rect 281200 273441 281206 273493
rect 281258 273481 281264 273493
rect 285808 273481 285814 273493
rect 281258 273453 285814 273481
rect 281258 273441 281264 273453
rect 285808 273441 285814 273453
rect 285866 273441 285872 273493
rect 285904 273441 285910 273493
rect 285962 273481 285968 273493
rect 310864 273481 310870 273493
rect 285962 273453 310870 273481
rect 285962 273441 285968 273453
rect 310864 273441 310870 273453
rect 310922 273441 310928 273493
rect 314512 273441 314518 273493
rect 314570 273481 314576 273493
rect 557008 273481 557014 273493
rect 314570 273453 557014 273481
rect 314570 273441 314576 273453
rect 557008 273441 557014 273453
rect 557066 273441 557072 273493
rect 146512 273367 146518 273419
rect 146570 273407 146576 273419
rect 151120 273407 151126 273419
rect 146570 273379 151126 273407
rect 146570 273367 146576 273379
rect 151120 273367 151126 273379
rect 151178 273367 151184 273419
rect 161008 273367 161014 273419
rect 161066 273407 161072 273419
rect 394576 273407 394582 273419
rect 161066 273379 394582 273407
rect 161066 273367 161072 273379
rect 394576 273367 394582 273379
rect 394634 273367 394640 273419
rect 404080 273407 404086 273419
rect 394690 273379 404086 273407
rect 144400 273293 144406 273345
rect 144458 273333 144464 273345
rect 146800 273333 146806 273345
rect 144458 273305 146806 273333
rect 144458 273293 144464 273305
rect 146800 273293 146806 273305
rect 146858 273293 146864 273345
rect 157456 273293 157462 273345
rect 157514 273333 157520 273345
rect 394690 273333 394718 273379
rect 404080 273367 404086 273379
rect 404138 273367 404144 273419
rect 403984 273333 403990 273345
rect 157514 273305 394718 273333
rect 394786 273305 403990 273333
rect 157514 273293 157520 273305
rect 158608 273219 158614 273271
rect 158666 273259 158672 273271
rect 161200 273259 161206 273271
rect 158666 273231 161206 273259
rect 158666 273219 158672 273231
rect 161200 273219 161206 273231
rect 161258 273219 161264 273271
rect 163120 273219 163126 273271
rect 163178 273259 163184 273271
rect 394786 273259 394814 273305
rect 403984 273293 403990 273305
rect 404042 273293 404048 273345
rect 163178 273231 394814 273259
rect 163178 273219 163184 273231
rect 394864 273219 394870 273271
rect 394922 273259 394928 273271
rect 408208 273259 408214 273271
rect 394922 273231 408214 273259
rect 394922 273219 394928 273231
rect 408208 273219 408214 273231
rect 408266 273219 408272 273271
rect 128944 273145 128950 273197
rect 129002 273185 129008 273197
rect 146512 273185 146518 273197
rect 129002 273157 146518 273185
rect 129002 273145 129008 273157
rect 146512 273145 146518 273157
rect 146570 273145 146576 273197
rect 147856 273185 147862 273197
rect 146626 273157 147862 273185
rect 95632 273071 95638 273123
rect 95690 273111 95696 273123
rect 100720 273111 100726 273123
rect 95690 273083 100726 273111
rect 95690 273071 95696 273083
rect 100720 273071 100726 273083
rect 100778 273071 100784 273123
rect 132496 273071 132502 273123
rect 132554 273111 132560 273123
rect 146626 273111 146654 273157
rect 147856 273145 147862 273157
rect 147914 273145 147920 273197
rect 147952 273145 147958 273197
rect 148010 273185 148016 273197
rect 149680 273185 149686 273197
rect 148010 273157 149686 273185
rect 148010 273145 148016 273157
rect 149680 273145 149686 273157
rect 149738 273145 149744 273197
rect 151408 273145 151414 273197
rect 151466 273185 151472 273197
rect 152560 273185 152566 273197
rect 151466 273157 152566 273185
rect 151466 273145 151472 273157
rect 152560 273145 152566 273157
rect 152618 273145 152624 273197
rect 152656 273145 152662 273197
rect 152714 273185 152720 273197
rect 155344 273185 155350 273197
rect 152714 273157 155350 273185
rect 152714 273145 152720 273157
rect 155344 273145 155350 273157
rect 155402 273145 155408 273197
rect 156208 273145 156214 273197
rect 156266 273185 156272 273197
rect 158320 273185 158326 273197
rect 156266 273157 158326 273185
rect 156266 273145 156272 273157
rect 158320 273145 158326 273157
rect 158378 273145 158384 273197
rect 159856 273145 159862 273197
rect 159914 273185 159920 273197
rect 161104 273185 161110 273197
rect 159914 273157 161110 273185
rect 159914 273145 159920 273157
rect 161104 273145 161110 273157
rect 161162 273145 161168 273197
rect 162160 273145 162166 273197
rect 162218 273185 162224 273197
rect 164080 273185 164086 273197
rect 162218 273157 164086 273185
rect 162218 273145 162224 273157
rect 164080 273145 164086 273157
rect 164138 273145 164144 273197
rect 164176 273145 164182 273197
rect 164234 273185 164240 273197
rect 378448 273185 378454 273197
rect 164234 273157 378454 273185
rect 164234 273145 164240 273157
rect 378448 273145 378454 273157
rect 378506 273145 378512 273197
rect 400624 273185 400630 273197
rect 378562 273157 400630 273185
rect 132554 273083 146654 273111
rect 132554 273071 132560 273083
rect 146704 273071 146710 273123
rect 146762 273111 146768 273123
rect 377968 273111 377974 273123
rect 146762 273083 377974 273111
rect 146762 273071 146768 273083
rect 377968 273071 377974 273083
rect 378026 273071 378032 273123
rect 143152 272997 143158 273049
rect 143210 273037 143216 273049
rect 378562 273037 378590 273157
rect 400624 273145 400630 273157
rect 400682 273145 400688 273197
rect 399664 273111 399670 273123
rect 143210 273009 378590 273037
rect 378658 273083 399670 273111
rect 143210 272997 143216 273009
rect 130096 272923 130102 272975
rect 130154 272963 130160 272975
rect 132400 272963 132406 272975
rect 130154 272935 132406 272963
rect 130154 272923 130160 272935
rect 132400 272923 132406 272935
rect 132458 272923 132464 272975
rect 133552 272923 133558 272975
rect 133610 272963 133616 272975
rect 135280 272963 135286 272975
rect 133610 272935 135286 272963
rect 133610 272923 133616 272935
rect 135280 272923 135286 272935
rect 135338 272923 135344 272975
rect 139600 272923 139606 272975
rect 139658 272963 139664 272975
rect 378658 272963 378686 273083
rect 399664 273071 399670 273083
rect 399722 273071 399728 273123
rect 378736 272997 378742 273049
rect 378794 273037 378800 273049
rect 398608 273037 398614 273049
rect 378794 273009 398614 273037
rect 378794 272997 378800 273009
rect 398608 272997 398614 273009
rect 398666 272997 398672 273049
rect 398032 272963 398038 272975
rect 139658 272935 378686 272963
rect 378754 272935 398038 272963
rect 139658 272923 139664 272935
rect 65872 272849 65878 272901
rect 65930 272889 65936 272901
rect 198640 272889 198646 272901
rect 65930 272861 198646 272889
rect 65930 272849 65936 272861
rect 198640 272849 198646 272861
rect 198698 272849 198704 272901
rect 198736 272849 198742 272901
rect 198794 272889 198800 272901
rect 211600 272889 211606 272901
rect 198794 272861 211606 272889
rect 198794 272849 198800 272861
rect 211600 272849 211606 272861
rect 211658 272849 211664 272901
rect 220816 272849 220822 272901
rect 220874 272889 220880 272901
rect 245488 272889 245494 272901
rect 220874 272861 245494 272889
rect 220874 272849 220880 272861
rect 245488 272849 245494 272861
rect 245546 272849 245552 272901
rect 267856 272849 267862 272901
rect 267914 272889 267920 272901
rect 270352 272889 270358 272901
rect 267914 272861 270358 272889
rect 267914 272849 267920 272861
rect 270352 272849 270358 272861
rect 270410 272849 270416 272901
rect 270448 272849 270454 272901
rect 270506 272889 270512 272901
rect 271408 272889 271414 272901
rect 270506 272861 271414 272889
rect 270506 272849 270512 272861
rect 271408 272849 271414 272861
rect 271466 272849 271472 272901
rect 271504 272849 271510 272901
rect 271562 272889 271568 272901
rect 277552 272889 277558 272901
rect 271562 272861 277558 272889
rect 271562 272849 271568 272861
rect 277552 272849 277558 272861
rect 277610 272849 277616 272901
rect 278800 272849 278806 272901
rect 278858 272889 278864 272901
rect 280048 272889 280054 272901
rect 278858 272861 280054 272889
rect 278858 272849 278864 272861
rect 280048 272849 280054 272861
rect 280106 272849 280112 272901
rect 280720 272849 280726 272901
rect 280778 272889 280784 272901
rect 282352 272889 282358 272901
rect 280778 272861 282358 272889
rect 280778 272849 280784 272861
rect 282352 272849 282358 272861
rect 282410 272849 282416 272901
rect 282448 272849 282454 272901
rect 282506 272889 282512 272901
rect 378256 272889 378262 272901
rect 282506 272861 378262 272889
rect 282506 272849 282512 272861
rect 378256 272849 378262 272861
rect 378314 272849 378320 272901
rect 378640 272889 378646 272901
rect 378466 272861 378646 272889
rect 101488 272775 101494 272827
rect 101546 272815 101552 272827
rect 103600 272815 103606 272827
rect 101546 272787 103606 272815
rect 101546 272775 101552 272787
rect 103600 272775 103606 272787
rect 103658 272775 103664 272827
rect 105040 272775 105046 272827
rect 105098 272815 105104 272827
rect 106480 272815 106486 272827
rect 105098 272787 106486 272815
rect 105098 272775 105104 272787
rect 106480 272775 106486 272787
rect 106538 272775 106544 272827
rect 115792 272775 115798 272827
rect 115850 272815 115856 272827
rect 118000 272815 118006 272827
rect 115850 272787 118006 272815
rect 115850 272775 115856 272787
rect 118000 272775 118006 272787
rect 118058 272775 118064 272827
rect 119344 272775 119350 272827
rect 119402 272815 119408 272827
rect 120880 272815 120886 272827
rect 119402 272787 120886 272815
rect 119402 272775 119408 272787
rect 120880 272775 120886 272787
rect 120938 272775 120944 272827
rect 122896 272775 122902 272827
rect 122954 272815 122960 272827
rect 123760 272815 123766 272827
rect 122954 272787 123766 272815
rect 122954 272775 122960 272787
rect 123760 272775 123766 272787
rect 123818 272775 123824 272827
rect 124144 272775 124150 272827
rect 124202 272815 124208 272827
rect 126544 272815 126550 272827
rect 124202 272787 126550 272815
rect 124202 272775 124208 272787
rect 126544 272775 126550 272787
rect 126602 272775 126608 272827
rect 127696 272775 127702 272827
rect 127754 272815 127760 272827
rect 129520 272815 129526 272827
rect 127754 272787 129526 272815
rect 127754 272775 127760 272787
rect 129520 272775 129526 272787
rect 129578 272775 129584 272827
rect 131248 272775 131254 272827
rect 131306 272815 131312 272827
rect 132304 272815 132310 272827
rect 131306 272787 132310 272815
rect 131306 272775 131312 272787
rect 132304 272775 132310 272787
rect 132362 272775 132368 272827
rect 137200 272775 137206 272827
rect 137258 272815 137264 272827
rect 138160 272815 138166 272827
rect 137258 272787 138166 272815
rect 137258 272775 137264 272787
rect 138160 272775 138166 272787
rect 138218 272775 138224 272827
rect 142000 272775 142006 272827
rect 142058 272815 142064 272827
rect 143920 272815 143926 272827
rect 142058 272787 143926 272815
rect 142058 272775 142064 272787
rect 143920 272775 143926 272787
rect 143978 272775 143984 272827
rect 146704 272775 146710 272827
rect 146762 272815 146768 272827
rect 378466 272815 378494 272861
rect 378640 272849 378646 272861
rect 378698 272849 378704 272901
rect 378754 272815 378782 272935
rect 398032 272923 398038 272935
rect 398090 272923 398096 272975
rect 378928 272849 378934 272901
rect 378986 272889 378992 272901
rect 380752 272889 380758 272901
rect 378986 272861 380758 272889
rect 378986 272849 378992 272861
rect 380752 272849 380758 272861
rect 380810 272849 380816 272901
rect 380848 272849 380854 272901
rect 380906 272889 380912 272901
rect 643888 272889 643894 272901
rect 380906 272861 643894 272889
rect 380906 272849 380912 272861
rect 643888 272849 643894 272861
rect 643946 272849 643952 272901
rect 146762 272787 378494 272815
rect 378562 272787 378782 272815
rect 146762 272775 146768 272787
rect 135952 272701 135958 272753
rect 136010 272741 136016 272753
rect 146608 272741 146614 272753
rect 136010 272713 146614 272741
rect 136010 272701 136016 272713
rect 146608 272701 146614 272713
rect 146666 272701 146672 272753
rect 147856 272701 147862 272753
rect 147914 272741 147920 272753
rect 378562 272741 378590 272787
rect 378832 272775 378838 272827
rect 378890 272815 378896 272827
rect 378890 272787 387806 272815
rect 378890 272775 378896 272787
rect 387568 272741 387574 272753
rect 147914 272713 378590 272741
rect 378658 272713 387574 272741
rect 147914 272701 147920 272713
rect 151120 272627 151126 272679
rect 151178 272667 151184 272679
rect 378658 272667 378686 272713
rect 387568 272701 387574 272713
rect 387626 272701 387632 272753
rect 387778 272741 387806 272787
rect 391408 272775 391414 272827
rect 391466 272815 391472 272827
rect 412240 272815 412246 272827
rect 391466 272787 412246 272815
rect 391466 272775 391472 272787
rect 412240 272775 412246 272787
rect 412298 272775 412304 272827
rect 596176 272775 596182 272827
rect 596234 272815 596240 272827
rect 598480 272815 598486 272827
rect 596234 272787 598486 272815
rect 596234 272775 596240 272787
rect 598480 272775 598486 272787
rect 598538 272775 598544 272827
rect 387778 272713 387998 272741
rect 151178 272639 378686 272667
rect 151178 272627 151184 272639
rect 378736 272627 378742 272679
rect 378794 272667 378800 272679
rect 380368 272667 380374 272679
rect 378794 272639 380374 272667
rect 378794 272627 378800 272639
rect 380368 272627 380374 272639
rect 380426 272627 380432 272679
rect 380752 272627 380758 272679
rect 380810 272667 380816 272679
rect 381328 272667 381334 272679
rect 380810 272639 381334 272667
rect 380810 272627 380816 272639
rect 381328 272627 381334 272639
rect 381386 272627 381392 272679
rect 381616 272627 381622 272679
rect 381674 272667 381680 272679
rect 386416 272667 386422 272679
rect 381674 272639 386422 272667
rect 381674 272627 381680 272639
rect 386416 272627 386422 272639
rect 386474 272627 386480 272679
rect 386512 272627 386518 272679
rect 386570 272667 386576 272679
rect 387856 272667 387862 272679
rect 386570 272639 387862 272667
rect 386570 272627 386576 272639
rect 387856 272627 387862 272639
rect 387914 272627 387920 272679
rect 387970 272667 387998 272713
rect 397264 272701 397270 272753
rect 397322 272741 397328 272753
rect 397322 272713 398942 272741
rect 397322 272701 397328 272713
rect 398800 272667 398806 272679
rect 387970 272639 398806 272667
rect 398800 272627 398806 272639
rect 398858 272627 398864 272679
rect 398914 272667 398942 272713
rect 612976 272667 612982 272679
rect 398914 272639 612982 272667
rect 612976 272627 612982 272639
rect 613034 272627 613040 272679
rect 125296 272553 125302 272605
rect 125354 272593 125360 272605
rect 378352 272593 378358 272605
rect 125354 272565 378358 272593
rect 125354 272553 125360 272565
rect 378352 272553 378358 272565
rect 378410 272553 378416 272605
rect 378544 272553 378550 272605
rect 378602 272593 378608 272605
rect 391888 272593 391894 272605
rect 378602 272565 391894 272593
rect 378602 272553 378608 272565
rect 391888 272553 391894 272565
rect 391946 272553 391952 272605
rect 394576 272553 394582 272605
rect 394634 272593 394640 272605
rect 396880 272593 396886 272605
rect 394634 272565 396886 272593
rect 394634 272553 394640 272565
rect 396880 272553 396886 272565
rect 396938 272553 396944 272605
rect 397360 272553 397366 272605
rect 397418 272593 397424 272605
rect 591568 272593 591574 272605
rect 397418 272565 591574 272593
rect 397418 272553 397424 272565
rect 591568 272553 591574 272565
rect 591626 272553 591632 272605
rect 121744 272479 121750 272531
rect 121802 272519 121808 272531
rect 380272 272519 380278 272531
rect 121802 272491 380278 272519
rect 121802 272479 121808 272491
rect 380272 272479 380278 272491
rect 380330 272479 380336 272531
rect 380368 272479 380374 272531
rect 380426 272519 380432 272531
rect 402352 272519 402358 272531
rect 380426 272491 402358 272519
rect 380426 272479 380432 272491
rect 402352 272479 402358 272491
rect 402410 272479 402416 272531
rect 118096 272405 118102 272457
rect 118154 272445 118160 272457
rect 394192 272445 394198 272457
rect 118154 272417 394198 272445
rect 118154 272405 118160 272417
rect 394192 272405 394198 272417
rect 394250 272405 394256 272457
rect 394288 272405 394294 272457
rect 394346 272445 394352 272457
rect 584368 272445 584374 272457
rect 394346 272417 584374 272445
rect 394346 272405 394352 272417
rect 584368 272405 584374 272417
rect 584426 272405 584432 272457
rect 84880 272331 84886 272383
rect 84938 272371 84944 272383
rect 86320 272371 86326 272383
rect 84938 272343 86326 272371
rect 84938 272331 84944 272343
rect 86320 272331 86326 272343
rect 86378 272331 86384 272383
rect 111088 272331 111094 272383
rect 111146 272371 111152 272383
rect 111146 272343 392414 272371
rect 111146 272331 111152 272343
rect 107440 272257 107446 272309
rect 107498 272297 107504 272309
rect 378544 272297 378550 272309
rect 107498 272269 378550 272297
rect 107498 272257 107504 272269
rect 378544 272257 378550 272269
rect 378602 272257 378608 272309
rect 390928 272297 390934 272309
rect 378658 272269 390934 272297
rect 103888 272183 103894 272235
rect 103946 272223 103952 272235
rect 378658 272223 378686 272269
rect 390928 272257 390934 272269
rect 390986 272257 390992 272309
rect 392386 272297 392414 272343
rect 392464 272331 392470 272383
rect 392522 272371 392528 272383
rect 587920 272371 587926 272383
rect 392522 272343 587926 272371
rect 392522 272331 392528 272343
rect 587920 272331 587926 272343
rect 587978 272331 587984 272383
rect 392560 272297 392566 272309
rect 392386 272269 392566 272297
rect 392560 272257 392566 272269
rect 392618 272257 392624 272309
rect 393808 272257 393814 272309
rect 393866 272297 393872 272309
rect 573712 272297 573718 272309
rect 393866 272269 573718 272297
rect 393866 272257 393872 272269
rect 573712 272257 573718 272269
rect 573770 272257 573776 272309
rect 103946 272195 378686 272223
rect 103946 272183 103952 272195
rect 378736 272183 378742 272235
rect 378794 272223 378800 272235
rect 378928 272223 378934 272235
rect 378794 272195 378934 272223
rect 378794 272183 378800 272195
rect 378928 272183 378934 272195
rect 378986 272183 378992 272235
rect 379984 272183 379990 272235
rect 380042 272223 380048 272235
rect 381424 272223 381430 272235
rect 380042 272195 381430 272223
rect 380042 272183 380048 272195
rect 381424 272183 381430 272195
rect 381482 272183 381488 272235
rect 381520 272183 381526 272235
rect 381578 272223 381584 272235
rect 382480 272223 382486 272235
rect 381578 272195 382486 272223
rect 381578 272183 381584 272195
rect 382480 272183 382486 272195
rect 382538 272183 382544 272235
rect 382672 272183 382678 272235
rect 382730 272223 382736 272235
rect 541552 272223 541558 272235
rect 382730 272195 541558 272223
rect 382730 272183 382736 272195
rect 541552 272183 541558 272195
rect 541610 272183 541616 272235
rect 67024 272109 67030 272161
rect 67082 272149 67088 272161
rect 213232 272149 213238 272161
rect 67082 272121 213238 272149
rect 67082 272109 67088 272121
rect 213232 272109 213238 272121
rect 213290 272109 213296 272161
rect 221008 272109 221014 272161
rect 221066 272149 221072 272161
rect 249040 272149 249046 272161
rect 221066 272121 249046 272149
rect 221066 272109 221072 272121
rect 249040 272109 249046 272121
rect 249098 272109 249104 272161
rect 258352 272109 258358 272161
rect 258410 272149 258416 272161
rect 552304 272149 552310 272161
rect 258410 272121 552310 272149
rect 258410 272109 258416 272121
rect 552304 272109 552310 272121
rect 552362 272109 552368 272161
rect 89584 272035 89590 272087
rect 89642 272075 89648 272087
rect 92080 272075 92086 272087
rect 89642 272047 92086 272075
rect 89642 272035 89648 272047
rect 92080 272035 92086 272047
rect 92138 272035 92144 272087
rect 145552 272035 145558 272087
rect 145610 272075 145616 272087
rect 146704 272075 146710 272087
rect 145610 272047 146710 272075
rect 145610 272035 145616 272047
rect 146704 272035 146710 272047
rect 146762 272035 146768 272087
rect 150256 272035 150262 272087
rect 150314 272075 150320 272087
rect 164176 272075 164182 272087
rect 150314 272047 164182 272075
rect 150314 272035 150320 272047
rect 164176 272035 164182 272047
rect 164234 272035 164240 272087
rect 164560 272035 164566 272087
rect 164618 272075 164624 272087
rect 405904 272075 405910 272087
rect 164618 272047 405910 272075
rect 164618 272035 164624 272047
rect 405904 272035 405910 272047
rect 405962 272035 405968 272087
rect 99184 271961 99190 272013
rect 99242 272001 99248 272013
rect 198736 272001 198742 272013
rect 99242 271973 198742 272001
rect 99242 271961 99248 271973
rect 198736 271961 198742 271973
rect 198794 271961 198800 272013
rect 198832 271961 198838 272013
rect 198890 272001 198896 272013
rect 212176 272001 212182 272013
rect 198890 271973 212182 272001
rect 198890 271961 198896 271973
rect 212176 271961 212182 271973
rect 212234 271961 212240 272013
rect 224080 271961 224086 272013
rect 224138 272001 224144 272013
rect 267952 272001 267958 272013
rect 224138 271973 267958 272001
rect 224138 271961 224144 271973
rect 267952 271961 267958 271973
rect 268010 271961 268016 272013
rect 268048 271961 268054 272013
rect 268106 272001 268112 272013
rect 278992 272001 278998 272013
rect 268106 271973 278998 272001
rect 268106 271961 268112 271973
rect 278992 271961 278998 271973
rect 279050 271961 279056 272013
rect 285520 271961 285526 272013
rect 285578 272001 285584 272013
rect 321520 272001 321526 272013
rect 285578 271973 321526 272001
rect 285578 271961 285584 271973
rect 321520 271961 321526 271973
rect 321578 271961 321584 272013
rect 321616 271961 321622 272013
rect 321674 272001 321680 272013
rect 329776 272001 329782 272013
rect 321674 271973 329782 272001
rect 321674 271961 321680 271973
rect 329776 271961 329782 271973
rect 329834 271961 329840 272013
rect 336976 271961 336982 272013
rect 337034 272001 337040 272013
rect 343024 272001 343030 272013
rect 337034 271973 343030 272001
rect 337034 271961 337040 271973
rect 343024 271961 343030 271973
rect 343082 271961 343088 272013
rect 347920 271961 347926 272013
rect 347978 272001 347984 272013
rect 358480 272001 358486 272013
rect 347978 271973 358486 272001
rect 347978 271961 347984 271973
rect 358480 271961 358486 271973
rect 358538 271961 358544 272013
rect 365776 271961 365782 272013
rect 365834 272001 365840 272013
rect 380176 272001 380182 272013
rect 365834 271973 380182 272001
rect 365834 271961 365840 271973
rect 380176 271961 380182 271973
rect 380234 271961 380240 272013
rect 380272 271961 380278 272013
rect 380330 272001 380336 272013
rect 395248 272001 395254 272013
rect 380330 271973 395254 272001
rect 380330 271961 380336 271973
rect 395248 271961 395254 271973
rect 395306 271961 395312 272013
rect 396880 271961 396886 272013
rect 396938 272001 396944 272013
rect 398704 272001 398710 272013
rect 396938 271973 398710 272001
rect 396938 271961 396944 271973
rect 398704 271961 398710 271973
rect 398762 271961 398768 272013
rect 398800 271961 398806 272013
rect 398858 272001 398864 272013
rect 618832 272001 618838 272013
rect 398858 271973 618838 272001
rect 398858 271961 398864 271973
rect 618832 271961 618838 271973
rect 618890 271961 618896 272013
rect 172912 271887 172918 271939
rect 172970 271927 172976 271939
rect 175600 271927 175606 271939
rect 172970 271899 175606 271927
rect 172970 271887 172976 271899
rect 175600 271887 175606 271899
rect 175658 271887 175664 271939
rect 176464 271887 176470 271939
rect 176522 271927 176528 271939
rect 178480 271927 178486 271939
rect 176522 271899 178486 271927
rect 176522 271887 176528 271899
rect 178480 271887 178486 271899
rect 178538 271887 178544 271939
rect 407536 271927 407542 271939
rect 178786 271899 407542 271927
rect 171664 271739 171670 271791
rect 171722 271779 171728 271791
rect 178786 271779 178814 271899
rect 407536 271887 407542 271899
rect 407594 271887 407600 271939
rect 409648 271887 409654 271939
rect 409706 271927 409712 271939
rect 433456 271927 433462 271939
rect 409706 271899 433462 271927
rect 409706 271887 409712 271899
rect 433456 271887 433462 271899
rect 433514 271887 433520 271939
rect 633616 271887 633622 271939
rect 633674 271927 633680 271939
rect 642256 271927 642262 271939
rect 633674 271899 642262 271927
rect 633674 271887 633680 271899
rect 642256 271887 642262 271899
rect 642314 271887 642320 271939
rect 394864 271853 394870 271865
rect 171722 271751 178814 271779
rect 181186 271825 394870 271853
rect 171722 271739 171728 271751
rect 100834 271677 106622 271705
rect 100720 271591 100726 271643
rect 100778 271631 100784 271643
rect 100834 271631 100862 271677
rect 100778 271603 100862 271631
rect 100778 271591 100784 271603
rect 106594 271483 106622 271677
rect 175312 271665 175318 271717
rect 175370 271705 175376 271717
rect 181186 271705 181214 271825
rect 394864 271813 394870 271825
rect 394922 271813 394928 271865
rect 394960 271813 394966 271865
rect 395018 271853 395024 271865
rect 406672 271853 406678 271865
rect 395018 271825 406678 271853
rect 395018 271813 395024 271825
rect 406672 271813 406678 271825
rect 406730 271813 406736 271865
rect 409264 271779 409270 271791
rect 175370 271677 181214 271705
rect 182338 271751 409270 271779
rect 175370 271665 175376 271677
rect 121168 271591 121174 271643
rect 121226 271631 121232 271643
rect 121226 271603 126878 271631
rect 121226 271591 121232 271603
rect 126850 271557 126878 271603
rect 156880 271591 156886 271643
rect 156938 271631 156944 271643
rect 156938 271603 177182 271631
rect 156938 271591 156944 271603
rect 126850 271529 146942 271557
rect 120976 271483 120982 271495
rect 106594 271455 120982 271483
rect 120976 271443 120982 271455
rect 121034 271443 121040 271495
rect 146914 271483 146942 271529
rect 177040 271483 177046 271495
rect 146914 271455 177046 271483
rect 177040 271443 177046 271455
rect 177098 271443 177104 271495
rect 102640 271369 102646 271421
rect 102698 271409 102704 271421
rect 156880 271409 156886 271421
rect 102698 271381 156886 271409
rect 102698 271369 102704 271381
rect 156880 271369 156886 271381
rect 156938 271369 156944 271421
rect 177154 271409 177182 271603
rect 178864 271591 178870 271643
rect 178922 271631 178928 271643
rect 182338 271631 182366 271751
rect 409264 271739 409270 271751
rect 409322 271739 409328 271791
rect 182416 271665 182422 271717
rect 182474 271705 182480 271717
rect 403168 271705 403174 271717
rect 182474 271677 403174 271705
rect 182474 271665 182480 271677
rect 403168 271665 403174 271677
rect 403226 271665 403232 271717
rect 178922 271603 182366 271631
rect 178922 271591 178928 271603
rect 185968 271591 185974 271643
rect 186026 271631 186032 271643
rect 403024 271631 403030 271643
rect 186026 271603 403030 271631
rect 186026 271591 186032 271603
rect 403024 271591 403030 271603
rect 403082 271591 403088 271643
rect 189520 271517 189526 271569
rect 189578 271557 189584 271569
rect 403120 271557 403126 271569
rect 189578 271529 403126 271557
rect 189578 271517 189584 271529
rect 403120 271517 403126 271529
rect 403178 271517 403184 271569
rect 403312 271517 403318 271569
rect 403370 271557 403376 271569
rect 403370 271529 403550 271557
rect 403370 271517 403376 271529
rect 195760 271443 195766 271495
rect 195818 271483 195824 271495
rect 206608 271483 206614 271495
rect 195818 271455 206614 271483
rect 195818 271443 195824 271455
rect 206608 271443 206614 271455
rect 206666 271443 206672 271495
rect 209776 271443 209782 271495
rect 209834 271483 209840 271495
rect 209834 271455 212222 271483
rect 209834 271443 209840 271455
rect 198832 271409 198838 271421
rect 177154 271381 198838 271409
rect 198832 271369 198838 271381
rect 198890 271369 198896 271421
rect 212080 271409 212086 271421
rect 198946 271381 212086 271409
rect 113488 271295 113494 271347
rect 113546 271335 113552 271347
rect 198946 271335 198974 271381
rect 212080 271369 212086 271381
rect 212138 271369 212144 271421
rect 212194 271409 212222 271455
rect 223696 271443 223702 271495
rect 223754 271483 223760 271495
rect 267856 271483 267862 271495
rect 223754 271455 267862 271483
rect 223754 271443 223760 271455
rect 267856 271443 267862 271455
rect 267914 271443 267920 271495
rect 267952 271443 267958 271495
rect 268010 271483 268016 271495
rect 274000 271483 274006 271495
rect 268010 271455 274006 271483
rect 268010 271443 268016 271455
rect 274000 271443 274006 271455
rect 274058 271443 274064 271495
rect 275152 271443 275158 271495
rect 275210 271483 275216 271495
rect 279664 271483 279670 271495
rect 275210 271455 279670 271483
rect 275210 271443 275216 271455
rect 279664 271443 279670 271455
rect 279722 271443 279728 271495
rect 283792 271443 283798 271495
rect 283850 271483 283856 271495
rect 307312 271483 307318 271495
rect 283850 271455 307318 271483
rect 283850 271443 283856 271455
rect 307312 271443 307318 271455
rect 307370 271443 307376 271495
rect 313648 271443 313654 271495
rect 313706 271483 313712 271495
rect 321616 271483 321622 271495
rect 313706 271455 321622 271483
rect 313706 271443 313712 271455
rect 321616 271443 321622 271455
rect 321674 271443 321680 271495
rect 333328 271483 333334 271495
rect 321730 271455 333334 271483
rect 216112 271409 216118 271421
rect 212194 271381 216118 271409
rect 216112 271369 216118 271381
rect 216170 271369 216176 271421
rect 220336 271369 220342 271421
rect 220394 271409 220400 271421
rect 241840 271409 241846 271421
rect 220394 271381 241846 271409
rect 220394 271369 220400 271381
rect 241840 271369 241846 271381
rect 241898 271369 241904 271421
rect 246640 271369 246646 271421
rect 246698 271409 246704 271421
rect 246698 271381 247742 271409
rect 246698 271369 246704 271381
rect 211888 271335 211894 271347
rect 113546 271307 198974 271335
rect 199042 271307 211894 271335
rect 113546 271295 113552 271307
rect 116944 271221 116950 271273
rect 117002 271261 117008 271273
rect 199042 271261 199070 271307
rect 211888 271295 211894 271307
rect 211946 271295 211952 271347
rect 213328 271295 213334 271347
rect 213386 271335 213392 271347
rect 216688 271335 216694 271347
rect 213386 271307 216694 271335
rect 213386 271295 213392 271307
rect 216688 271295 216694 271307
rect 216746 271295 216752 271347
rect 219760 271295 219766 271347
rect 219818 271335 219824 271347
rect 238288 271335 238294 271347
rect 219818 271307 238294 271335
rect 219818 271295 219824 271307
rect 238288 271295 238294 271307
rect 238346 271295 238352 271347
rect 117002 271233 199070 271261
rect 117002 271221 117008 271233
rect 199120 271221 199126 271273
rect 199178 271261 199184 271273
rect 214960 271261 214966 271273
rect 199178 271233 214966 271261
rect 199178 271221 199184 271233
rect 214960 271221 214966 271233
rect 215018 271221 215024 271273
rect 247714 271261 247742 271381
rect 253744 271369 253750 271421
rect 253802 271409 253808 271421
rect 277264 271409 277270 271421
rect 253802 271381 277270 271409
rect 253802 271369 253808 271381
rect 277264 271369 277270 271381
rect 277322 271369 277328 271421
rect 282736 271369 282742 271421
rect 282794 271409 282800 271421
rect 296656 271409 296662 271421
rect 282794 271381 296662 271409
rect 282794 271369 282800 271381
rect 296656 271369 296662 271381
rect 296714 271369 296720 271421
rect 312112 271369 312118 271421
rect 312170 271409 312176 271421
rect 321730 271409 321758 271455
rect 333328 271443 333334 271455
rect 333386 271443 333392 271495
rect 333424 271443 333430 271495
rect 333482 271483 333488 271495
rect 342640 271483 342646 271495
rect 333482 271455 342646 271483
rect 333482 271443 333488 271455
rect 342640 271443 342646 271455
rect 342698 271443 342704 271495
rect 345712 271443 345718 271495
rect 345770 271483 345776 271495
rect 358384 271483 358390 271495
rect 345770 271455 358390 271483
rect 345770 271443 345776 271455
rect 358384 271443 358390 271455
rect 358442 271443 358448 271495
rect 358480 271443 358486 271495
rect 358538 271483 358544 271495
rect 374416 271483 374422 271495
rect 358538 271455 374422 271483
rect 358538 271443 358544 271455
rect 374416 271443 374422 271455
rect 374474 271443 374480 271495
rect 374704 271443 374710 271495
rect 374762 271483 374768 271495
rect 403216 271483 403222 271495
rect 374762 271455 403222 271483
rect 374762 271443 374768 271455
rect 403216 271443 403222 271455
rect 403274 271443 403280 271495
rect 403522 271483 403550 271529
rect 459280 271517 459286 271569
rect 459338 271557 459344 271569
rect 479440 271557 479446 271569
rect 459338 271529 479446 271557
rect 459338 271517 459344 271529
rect 479440 271517 479446 271529
rect 479498 271517 479504 271569
rect 499600 271517 499606 271569
rect 499658 271557 499664 271569
rect 518320 271557 518326 271569
rect 499658 271529 518326 271557
rect 499658 271517 499664 271529
rect 518320 271517 518326 271529
rect 518378 271517 518384 271569
rect 593968 271483 593974 271495
rect 403522 271455 593974 271483
rect 593968 271443 593974 271455
rect 594026 271443 594032 271495
rect 312170 271381 321758 271409
rect 312170 271369 312176 271381
rect 324112 271369 324118 271421
rect 324170 271409 324176 271421
rect 325552 271409 325558 271421
rect 324170 271381 325558 271409
rect 324170 271369 324176 271381
rect 325552 271369 325558 271381
rect 325610 271369 325616 271421
rect 329968 271369 329974 271421
rect 330026 271409 330032 271421
rect 341968 271409 341974 271421
rect 330026 271381 341974 271409
rect 330026 271369 330032 271381
rect 341968 271369 341974 271381
rect 342026 271369 342032 271421
rect 347440 271369 347446 271421
rect 347498 271409 347504 271421
rect 372688 271409 372694 271421
rect 347498 271381 372694 271409
rect 347498 271369 347504 271381
rect 372688 271369 372694 271381
rect 372746 271369 372752 271421
rect 374032 271369 374038 271421
rect 374090 271409 374096 271421
rect 590320 271409 590326 271421
rect 374090 271381 590326 271409
rect 374090 271369 374096 271381
rect 590320 271369 590326 271381
rect 590378 271369 590384 271421
rect 264496 271295 264502 271347
rect 264554 271335 264560 271347
rect 278512 271335 278518 271347
rect 264554 271307 278518 271335
rect 264554 271295 264560 271307
rect 278512 271295 278518 271307
rect 278570 271295 278576 271347
rect 282928 271295 282934 271347
rect 282986 271335 282992 271347
rect 300112 271335 300118 271347
rect 282986 271307 300118 271335
rect 282986 271295 282992 271307
rect 300112 271295 300118 271307
rect 300170 271295 300176 271347
rect 308176 271295 308182 271347
rect 308234 271335 308240 271347
rect 319408 271335 319414 271347
rect 308234 271307 319414 271335
rect 308234 271295 308240 271307
rect 319408 271295 319414 271307
rect 319466 271295 319472 271347
rect 320368 271295 320374 271347
rect 320426 271335 320432 271347
rect 325648 271335 325654 271347
rect 320426 271307 325654 271335
rect 320426 271295 320432 271307
rect 325648 271295 325654 271307
rect 325706 271295 325712 271347
rect 339376 271335 339382 271347
rect 328210 271307 339382 271335
rect 247714 271233 267710 271261
rect 120496 271147 120502 271199
rect 120554 271187 120560 271199
rect 211792 271187 211798 271199
rect 120554 271159 211798 271187
rect 120554 271147 120560 271159
rect 211792 271147 211798 271159
rect 211850 271147 211856 271199
rect 219280 271147 219286 271199
rect 219338 271187 219344 271199
rect 234640 271187 234646 271199
rect 219338 271159 234646 271187
rect 219338 271147 219344 271159
rect 234640 271147 234646 271159
rect 234698 271147 234704 271199
rect 109840 271073 109846 271125
rect 109898 271113 109904 271125
rect 201520 271113 201526 271125
rect 109898 271085 201526 271113
rect 109898 271073 109904 271085
rect 201520 271073 201526 271085
rect 201578 271073 201584 271125
rect 202576 271073 202582 271125
rect 202634 271113 202640 271125
rect 215440 271113 215446 271125
rect 202634 271085 215446 271113
rect 202634 271073 202640 271085
rect 215440 271073 215446 271085
rect 215498 271073 215504 271125
rect 218896 271073 218902 271125
rect 218954 271113 218960 271125
rect 231184 271113 231190 271125
rect 218954 271085 231190 271113
rect 218954 271073 218960 271085
rect 231184 271073 231190 271085
rect 231242 271073 231248 271125
rect 267682 271113 267710 271233
rect 283408 271221 283414 271273
rect 283466 271261 283472 271273
rect 303664 271261 303670 271273
rect 283466 271233 303670 271261
rect 283466 271221 283472 271233
rect 303664 271221 303670 271233
rect 303722 271221 303728 271273
rect 308464 271221 308470 271273
rect 308522 271261 308528 271273
rect 328210 271261 328238 271307
rect 339376 271295 339382 271307
rect 339434 271295 339440 271347
rect 345328 271335 345334 271347
rect 341026 271307 345334 271335
rect 340912 271261 340918 271273
rect 308522 271233 328238 271261
rect 329794 271233 340918 271261
rect 308522 271221 308528 271233
rect 276400 271187 276406 271199
rect 268642 271159 276406 271187
rect 268642 271113 268670 271159
rect 276400 271147 276406 271159
rect 276458 271147 276464 271199
rect 284464 271147 284470 271199
rect 284522 271187 284528 271199
rect 285904 271187 285910 271199
rect 284522 271159 285910 271187
rect 284522 271147 284528 271159
rect 285904 271147 285910 271159
rect 285962 271147 285968 271199
rect 319120 271147 319126 271199
rect 319178 271187 319184 271199
rect 329794 271187 329822 271233
rect 340912 271221 340918 271233
rect 340970 271221 340976 271273
rect 341026 271187 341054 271307
rect 345328 271295 345334 271307
rect 345386 271295 345392 271347
rect 347248 271295 347254 271347
rect 347306 271335 347312 271347
rect 347306 271307 362174 271335
rect 347306 271295 347312 271307
rect 346384 271221 346390 271273
rect 346442 271261 346448 271273
rect 362032 271261 362038 271273
rect 346442 271233 362038 271261
rect 346442 271221 346448 271233
rect 362032 271221 362038 271233
rect 362090 271221 362096 271273
rect 319178 271159 329822 271187
rect 329986 271159 341054 271187
rect 319178 271147 319184 271159
rect 267682 271085 268670 271113
rect 268720 271073 268726 271125
rect 268778 271113 268784 271125
rect 270448 271113 270454 271125
rect 268778 271085 270454 271113
rect 268778 271073 268784 271085
rect 270448 271073 270454 271085
rect 270506 271073 270512 271125
rect 292528 271073 292534 271125
rect 292586 271113 292592 271125
rect 292586 271085 312446 271113
rect 292586 271073 292592 271085
rect 106288 270999 106294 271051
rect 106346 271039 106352 271051
rect 191440 271039 191446 271051
rect 106346 271011 191446 271039
rect 106346 270999 106352 271011
rect 191440 270999 191446 271011
rect 191498 270999 191504 271051
rect 193072 270999 193078 271051
rect 193130 271039 193136 271051
rect 269872 271039 269878 271051
rect 193130 271011 269878 271039
rect 193130 270999 193136 271011
rect 269872 270999 269878 271011
rect 269930 270999 269936 271051
rect 282160 270999 282166 271051
rect 282218 271039 282224 271051
rect 293008 271039 293014 271051
rect 282218 271011 293014 271039
rect 282218 270999 282224 271011
rect 293008 270999 293014 271011
rect 293066 270999 293072 271051
rect 302512 270999 302518 271051
rect 302570 271039 302576 271051
rect 312418 271039 312446 271085
rect 315952 271073 315958 271125
rect 316010 271113 316016 271125
rect 322000 271113 322006 271125
rect 316010 271085 322006 271113
rect 316010 271073 316016 271085
rect 322000 271073 322006 271085
rect 322058 271073 322064 271125
rect 322768 271073 322774 271125
rect 322826 271113 322832 271125
rect 329488 271113 329494 271125
rect 322826 271085 329494 271113
rect 322826 271073 322832 271085
rect 329488 271073 329494 271085
rect 329546 271073 329552 271125
rect 329680 271073 329686 271125
rect 329738 271113 329744 271125
rect 329986 271113 330014 271159
rect 345232 271147 345238 271199
rect 345290 271187 345296 271199
rect 354832 271187 354838 271199
rect 345290 271159 354838 271187
rect 345290 271147 345296 271159
rect 354832 271147 354838 271159
rect 354890 271147 354896 271199
rect 362146 271187 362174 271307
rect 366160 271295 366166 271347
rect 366218 271335 366224 271347
rect 370384 271335 370390 271347
rect 366218 271307 370390 271335
rect 366218 271295 366224 271307
rect 370384 271295 370390 271307
rect 370442 271295 370448 271347
rect 370480 271295 370486 271347
rect 370538 271335 370544 271347
rect 403408 271335 403414 271347
rect 370538 271307 403414 271335
rect 370538 271295 370544 271307
rect 403408 271295 403414 271307
rect 403466 271295 403472 271347
rect 413200 271295 413206 271347
rect 413258 271335 413264 271347
rect 559408 271335 559414 271347
rect 413258 271307 559414 271335
rect 413258 271295 413264 271307
rect 559408 271295 559414 271307
rect 559466 271295 559472 271347
rect 365104 271221 365110 271273
rect 365162 271261 365168 271273
rect 381520 271261 381526 271273
rect 365162 271233 381526 271261
rect 365162 271221 365168 271233
rect 381520 271221 381526 271233
rect 381578 271221 381584 271273
rect 381904 271221 381910 271273
rect 381962 271261 381968 271273
rect 409648 271261 409654 271273
rect 381962 271233 409654 271261
rect 381962 271221 381968 271233
rect 409648 271221 409654 271233
rect 409706 271221 409712 271273
rect 433456 271221 433462 271273
rect 433514 271261 433520 271273
rect 459280 271261 459286 271273
rect 433514 271233 459286 271261
rect 433514 271221 433520 271233
rect 459280 271221 459286 271233
rect 459338 271221 459344 271273
rect 479440 271221 479446 271273
rect 479498 271261 479504 271273
rect 499600 271261 499606 271273
rect 479498 271233 499606 271261
rect 479498 271221 479504 271233
rect 499600 271221 499606 271233
rect 499658 271221 499664 271273
rect 518320 271221 518326 271273
rect 518378 271261 518384 271273
rect 543952 271261 543958 271273
rect 518378 271233 543958 271261
rect 518378 271221 518384 271233
rect 543952 271221 543958 271233
rect 544010 271221 544016 271273
rect 369136 271187 369142 271199
rect 362146 271159 369142 271187
rect 369136 271147 369142 271159
rect 369194 271147 369200 271199
rect 369232 271147 369238 271199
rect 369290 271187 369296 271199
rect 373648 271187 373654 271199
rect 369290 271159 373654 271187
rect 369290 271147 369296 271159
rect 373648 271147 373654 271159
rect 373706 271147 373712 271199
rect 374416 271147 374422 271199
rect 374474 271187 374480 271199
rect 376240 271187 376246 271199
rect 374474 271159 376246 271187
rect 374474 271147 374480 271159
rect 376240 271147 376246 271159
rect 376298 271147 376304 271199
rect 376336 271147 376342 271199
rect 376394 271187 376400 271199
rect 378064 271187 378070 271199
rect 376394 271159 378070 271187
rect 376394 271147 376400 271159
rect 378064 271147 378070 271159
rect 378122 271147 378128 271199
rect 378160 271147 378166 271199
rect 378218 271187 378224 271199
rect 395056 271187 395062 271199
rect 378218 271159 395062 271187
rect 378218 271147 378224 271159
rect 395056 271147 395062 271159
rect 395114 271147 395120 271199
rect 395440 271147 395446 271199
rect 395498 271187 395504 271199
rect 534448 271187 534454 271199
rect 395498 271159 534454 271187
rect 395498 271147 395504 271159
rect 534448 271147 534454 271159
rect 534506 271147 534512 271199
rect 329738 271085 330014 271113
rect 329738 271073 329744 271085
rect 333328 271073 333334 271125
rect 333386 271113 333392 271125
rect 336688 271113 336694 271125
rect 333386 271085 336694 271113
rect 333386 271073 333392 271085
rect 336688 271073 336694 271085
rect 336746 271073 336752 271125
rect 393616 271113 393622 271125
rect 336802 271085 393622 271113
rect 320272 271039 320278 271051
rect 302570 271011 308318 271039
rect 312418 271011 320278 271039
rect 302570 270999 302576 271011
rect 191920 270925 191926 270977
rect 191978 270965 191984 270977
rect 213808 270965 213814 270977
rect 191978 270937 213814 270965
rect 191978 270925 191984 270937
rect 213808 270925 213814 270937
rect 213866 270925 213872 270977
rect 218704 270925 218710 270977
rect 218762 270965 218768 270977
rect 227632 270965 227638 270977
rect 218762 270937 227638 270965
rect 218762 270925 218768 270937
rect 227632 270925 227638 270937
rect 227690 270925 227696 270977
rect 257296 270925 257302 270977
rect 257354 270965 257360 270977
rect 277456 270965 277462 270977
rect 257354 270937 277462 270965
rect 257354 270925 257360 270937
rect 277456 270925 277462 270937
rect 277514 270925 277520 270977
rect 281680 270925 281686 270977
rect 281738 270965 281744 270977
rect 289456 270965 289462 270977
rect 281738 270937 289462 270965
rect 281738 270925 281744 270937
rect 289456 270925 289462 270937
rect 289514 270925 289520 270977
rect 294256 270925 294262 270977
rect 294314 270965 294320 270977
rect 308176 270965 308182 270977
rect 294314 270937 308182 270965
rect 294314 270925 294320 270937
rect 308176 270925 308182 270937
rect 308234 270925 308240 270977
rect 308290 270965 308318 271011
rect 320272 270999 320278 271011
rect 320330 270999 320336 271051
rect 322096 270999 322102 271051
rect 322154 271039 322160 271051
rect 336802 271039 336830 271085
rect 393616 271073 393622 271085
rect 393674 271073 393680 271125
rect 394480 271073 394486 271125
rect 394538 271113 394544 271125
rect 580912 271113 580918 271125
rect 394538 271085 580918 271113
rect 394538 271073 394544 271085
rect 580912 271073 580918 271085
rect 580970 271073 580976 271125
rect 322154 271011 336830 271039
rect 322154 270999 322160 271011
rect 336880 270999 336886 271051
rect 336938 271039 336944 271051
rect 383056 271039 383062 271051
rect 336938 271011 383062 271039
rect 336938 270999 336944 271011
rect 383056 270999 383062 271011
rect 383114 270999 383120 271051
rect 383152 270999 383158 271051
rect 383210 271039 383216 271051
rect 510640 271039 510646 271051
rect 383210 271011 510646 271039
rect 383210 270999 383216 271011
rect 510640 270999 510646 271011
rect 510698 270999 510704 271051
rect 322672 270965 322678 270977
rect 308290 270937 322678 270965
rect 322672 270925 322678 270937
rect 322730 270925 322736 270977
rect 322960 270925 322966 270977
rect 323018 270965 323024 270977
rect 324880 270965 324886 270977
rect 323018 270937 324886 270965
rect 323018 270925 323024 270937
rect 324880 270925 324886 270937
rect 324938 270925 324944 270977
rect 326320 270925 326326 270977
rect 326378 270965 326384 270977
rect 341488 270965 341494 270977
rect 326378 270937 341494 270965
rect 326378 270925 326384 270937
rect 341488 270925 341494 270937
rect 341546 270925 341552 270977
rect 344752 270925 344758 270977
rect 344810 270965 344816 270977
rect 351280 270965 351286 270977
rect 344810 270937 351286 270965
rect 344810 270925 344816 270937
rect 351280 270925 351286 270937
rect 351338 270925 351344 270977
rect 363856 270925 363862 270977
rect 363914 270965 363920 270977
rect 371536 270965 371542 270977
rect 363914 270937 371542 270965
rect 363914 270925 363920 270937
rect 371536 270925 371542 270937
rect 371594 270925 371600 270977
rect 373456 270925 373462 270977
rect 373514 270965 373520 270977
rect 388624 270965 388630 270977
rect 373514 270937 388630 270965
rect 373514 270925 373520 270937
rect 388624 270925 388630 270937
rect 388682 270925 388688 270977
rect 388720 270925 388726 270977
rect 388778 270965 388784 270977
rect 545200 270965 545206 270977
rect 388778 270937 545206 270965
rect 388778 270925 388784 270937
rect 545200 270925 545206 270937
rect 545258 270925 545264 270977
rect 168112 270851 168118 270903
rect 168170 270891 168176 270903
rect 394960 270891 394966 270903
rect 168170 270863 394966 270891
rect 168170 270851 168176 270863
rect 394960 270851 394966 270863
rect 395018 270851 395024 270903
rect 395056 270851 395062 270903
rect 395114 270891 395120 270903
rect 401296 270891 401302 270903
rect 395114 270863 401302 270891
rect 395114 270851 395120 270863
rect 401296 270851 401302 270863
rect 401354 270851 401360 270903
rect 403408 270851 403414 270903
rect 403466 270891 403472 270903
rect 413200 270891 413206 270903
rect 403466 270863 413206 270891
rect 403466 270851 403472 270863
rect 413200 270851 413206 270863
rect 413258 270851 413264 270903
rect 177040 270777 177046 270829
rect 177098 270817 177104 270829
rect 177098 270789 193022 270817
rect 177098 270777 177104 270789
rect 68176 270703 68182 270755
rect 68234 270743 68240 270755
rect 69040 270743 69046 270755
rect 68234 270715 69046 270743
rect 68234 270703 68240 270715
rect 69040 270703 69046 270715
rect 69098 270703 69104 270755
rect 75376 270703 75382 270755
rect 75434 270743 75440 270755
rect 77680 270743 77686 270755
rect 75434 270715 77686 270743
rect 75434 270703 75440 270715
rect 77680 270703 77686 270715
rect 77738 270703 77744 270755
rect 188368 270703 188374 270755
rect 188426 270743 188432 270755
rect 190000 270743 190006 270755
rect 188426 270715 190006 270743
rect 188426 270703 188432 270715
rect 190000 270703 190006 270715
rect 190058 270703 190064 270755
rect 190768 270703 190774 270755
rect 190826 270743 190832 270755
rect 192880 270743 192886 270755
rect 190826 270715 192886 270743
rect 190826 270703 190832 270715
rect 192880 270703 192886 270715
rect 192938 270703 192944 270755
rect 192994 270743 193022 270789
rect 195472 270777 195478 270829
rect 195530 270817 195536 270829
rect 214480 270817 214486 270829
rect 195530 270789 214486 270817
rect 195530 270777 195536 270789
rect 214480 270777 214486 270789
rect 214538 270777 214544 270829
rect 218224 270777 218230 270829
rect 218282 270817 218288 270829
rect 223984 270817 223990 270829
rect 218282 270789 223990 270817
rect 218282 270777 218288 270789
rect 223984 270777 223990 270789
rect 224042 270777 224048 270829
rect 260944 270777 260950 270829
rect 261002 270817 261008 270829
rect 277936 270817 277942 270829
rect 261002 270789 277942 270817
rect 261002 270777 261008 270789
rect 277936 270777 277942 270789
rect 277994 270777 278000 270829
rect 314800 270777 314806 270829
rect 314858 270817 314864 270829
rect 319696 270817 319702 270829
rect 314858 270789 319702 270817
rect 314858 270777 314864 270789
rect 319696 270777 319702 270789
rect 319754 270777 319760 270829
rect 322000 270777 322006 270829
rect 322058 270817 322064 270829
rect 340432 270817 340438 270829
rect 322058 270789 340438 270817
rect 322058 270777 322064 270789
rect 340432 270777 340438 270789
rect 340490 270777 340496 270829
rect 342736 270777 342742 270829
rect 342794 270817 342800 270829
rect 359632 270817 359638 270829
rect 342794 270789 359638 270817
rect 342794 270777 342800 270789
rect 359632 270777 359638 270789
rect 359690 270777 359696 270829
rect 362032 270777 362038 270829
rect 362090 270817 362096 270829
rect 365200 270817 365206 270829
rect 362090 270789 365206 270817
rect 362090 270777 362096 270789
rect 365200 270777 365206 270789
rect 365258 270777 365264 270829
rect 365296 270777 365302 270829
rect 365354 270817 365360 270829
rect 367024 270817 367030 270829
rect 365354 270789 367030 270817
rect 365354 270777 365360 270789
rect 367024 270777 367030 270789
rect 367082 270777 367088 270829
rect 367120 270777 367126 270829
rect 367178 270817 367184 270829
rect 369232 270817 369238 270829
rect 367178 270789 369238 270817
rect 367178 270777 367184 270789
rect 369232 270777 369238 270789
rect 369290 270777 369296 270829
rect 370672 270777 370678 270829
rect 370730 270817 370736 270829
rect 373552 270817 373558 270829
rect 370730 270789 373558 270817
rect 370730 270777 370736 270789
rect 373552 270777 373558 270789
rect 373610 270777 373616 270829
rect 373648 270777 373654 270829
rect 373706 270817 373712 270829
rect 376144 270817 376150 270829
rect 373706 270789 376150 270817
rect 373706 270777 373712 270789
rect 376144 270777 376150 270789
rect 376202 270777 376208 270829
rect 377584 270777 377590 270829
rect 377642 270817 377648 270829
rect 378832 270817 378838 270829
rect 377642 270789 378838 270817
rect 377642 270777 377648 270789
rect 378832 270777 378838 270789
rect 378890 270777 378896 270829
rect 378928 270777 378934 270829
rect 378986 270817 378992 270829
rect 386896 270817 386902 270829
rect 378986 270789 386902 270817
rect 378986 270777 378992 270789
rect 386896 270777 386902 270789
rect 386954 270777 386960 270829
rect 388048 270777 388054 270829
rect 388106 270817 388112 270829
rect 395440 270817 395446 270829
rect 388106 270789 395446 270817
rect 388106 270777 388112 270789
rect 395440 270777 395446 270789
rect 395498 270777 395504 270829
rect 398896 270777 398902 270829
rect 398954 270817 398960 270829
rect 404944 270817 404950 270829
rect 398954 270789 404950 270817
rect 398954 270777 398960 270789
rect 404944 270777 404950 270789
rect 405002 270777 405008 270829
rect 195760 270743 195766 270755
rect 192994 270715 195766 270743
rect 195760 270703 195766 270715
rect 195818 270703 195824 270755
rect 206224 270703 206230 270755
rect 206282 270743 206288 270755
rect 215536 270743 215542 270755
rect 206282 270715 215542 270743
rect 206282 270703 206288 270715
rect 215536 270703 215542 270715
rect 215594 270703 215600 270755
rect 217552 270703 217558 270755
rect 217610 270743 217616 270755
rect 220432 270743 220438 270755
rect 217610 270715 220438 270743
rect 217610 270703 217616 270715
rect 220432 270703 220438 270715
rect 220490 270703 220496 270755
rect 250192 270703 250198 270755
rect 250250 270743 250256 270755
rect 276784 270743 276790 270755
rect 250250 270715 276790 270743
rect 250250 270703 250256 270715
rect 276784 270703 276790 270715
rect 276842 270703 276848 270755
rect 317488 270703 317494 270755
rect 317546 270743 317552 270755
rect 392080 270743 392086 270755
rect 317546 270715 392086 270743
rect 317546 270703 317552 270715
rect 392080 270703 392086 270715
rect 392138 270703 392144 270755
rect 394480 270703 394486 270755
rect 394538 270743 394544 270755
rect 570160 270743 570166 270755
rect 394538 270715 570166 270743
rect 394538 270703 394544 270715
rect 570160 270703 570166 270715
rect 570218 270703 570224 270755
rect 230224 270629 230230 270681
rect 230282 270669 230288 270681
rect 310288 270669 310294 270681
rect 230282 270641 310294 270669
rect 230282 270629 230288 270641
rect 310288 270629 310294 270641
rect 310346 270629 310352 270681
rect 310384 270629 310390 270681
rect 310442 270669 310448 270681
rect 325648 270669 325654 270681
rect 310442 270641 325654 270669
rect 310442 270629 310448 270641
rect 325648 270629 325654 270641
rect 325706 270629 325712 270681
rect 328336 270629 328342 270681
rect 328394 270669 328400 270681
rect 329680 270669 329686 270681
rect 328394 270641 329686 270669
rect 328394 270629 328400 270641
rect 329680 270629 329686 270641
rect 329738 270629 329744 270681
rect 329776 270629 329782 270681
rect 329834 270669 329840 270681
rect 549904 270669 549910 270681
rect 329834 270641 549910 270669
rect 329834 270629 329840 270641
rect 549904 270629 549910 270641
rect 549962 270629 549968 270681
rect 231280 270555 231286 270607
rect 231338 270595 231344 270607
rect 328528 270595 328534 270607
rect 231338 270567 328534 270595
rect 231338 270555 231344 270567
rect 328528 270555 328534 270567
rect 328586 270555 328592 270607
rect 328624 270555 328630 270607
rect 328682 270595 328688 270607
rect 332272 270595 332278 270607
rect 328682 270567 332278 270595
rect 328682 270555 328688 270567
rect 332272 270555 332278 270567
rect 332330 270555 332336 270607
rect 336688 270555 336694 270607
rect 336746 270595 336752 270607
rect 339856 270595 339862 270607
rect 336746 270567 339862 270595
rect 336746 270555 336752 270567
rect 339856 270555 339862 270567
rect 339914 270555 339920 270607
rect 348304 270555 348310 270607
rect 348362 270595 348368 270607
rect 352720 270595 352726 270607
rect 348362 270567 352726 270595
rect 348362 270555 348368 270567
rect 352720 270555 352726 270567
rect 352778 270555 352784 270607
rect 358480 270555 358486 270607
rect 358538 270595 358544 270607
rect 370672 270595 370678 270607
rect 358538 270567 370678 270595
rect 358538 270555 358544 270567
rect 370672 270555 370678 270567
rect 370730 270555 370736 270607
rect 370768 270555 370774 270607
rect 370826 270595 370832 270607
rect 373456 270595 373462 270607
rect 370826 270567 373462 270595
rect 370826 270555 370832 270567
rect 373456 270555 373462 270567
rect 373514 270555 373520 270607
rect 373552 270555 373558 270607
rect 373610 270595 373616 270607
rect 379120 270595 379126 270607
rect 373610 270567 379126 270595
rect 373610 270555 373616 270567
rect 379120 270555 379126 270567
rect 379178 270555 379184 270607
rect 379792 270555 379798 270607
rect 379850 270595 379856 270607
rect 388720 270595 388726 270607
rect 379850 270567 388726 270595
rect 379850 270555 379856 270567
rect 388720 270555 388726 270567
rect 388778 270555 388784 270607
rect 388816 270555 388822 270607
rect 388874 270595 388880 270607
rect 561808 270595 561814 270607
rect 388874 270567 561814 270595
rect 388874 270555 388880 270567
rect 561808 270555 561814 270567
rect 561866 270555 561872 270607
rect 623056 270555 623062 270607
rect 623114 270595 623120 270607
rect 641488 270595 641494 270607
rect 623114 270567 641494 270595
rect 623114 270555 623120 270567
rect 641488 270555 641494 270567
rect 641546 270555 641552 270607
rect 203824 270481 203830 270533
rect 203882 270521 203888 270533
rect 270928 270521 270934 270533
rect 203882 270493 270934 270521
rect 203882 270481 203888 270493
rect 270928 270481 270934 270493
rect 270986 270481 270992 270533
rect 307792 270481 307798 270533
rect 307850 270521 307856 270533
rect 503536 270521 503542 270533
rect 307850 270493 503542 270521
rect 307850 270481 307856 270493
rect 503536 270481 503542 270493
rect 503594 270481 503600 270533
rect 544432 270481 544438 270533
rect 544490 270521 544496 270533
rect 564400 270521 564406 270533
rect 544490 270493 564406 270521
rect 544490 270481 544496 270493
rect 564400 270481 564406 270493
rect 564458 270481 564464 270533
rect 244144 270407 244150 270459
rect 244202 270447 244208 270459
rect 438064 270447 438070 270459
rect 244202 270419 438070 270447
rect 244202 270407 244208 270419
rect 438064 270407 438070 270419
rect 438122 270407 438128 270459
rect 440656 270407 440662 270459
rect 440714 270447 440720 270459
rect 460720 270447 460726 270459
rect 440714 270419 460726 270447
rect 440714 270407 440720 270419
rect 460720 270407 460726 270419
rect 460778 270407 460784 270459
rect 469168 270407 469174 270459
rect 469226 270447 469232 270459
rect 469648 270447 469654 270459
rect 469226 270419 469654 270447
rect 469226 270407 469232 270419
rect 469648 270407 469654 270419
rect 469706 270407 469712 270459
rect 232816 270333 232822 270385
rect 232874 270373 232880 270385
rect 328336 270373 328342 270385
rect 232874 270345 328342 270373
rect 232874 270333 232880 270345
rect 328336 270333 328342 270345
rect 328394 270333 328400 270385
rect 328528 270333 328534 270385
rect 328586 270373 328592 270385
rect 331120 270373 331126 270385
rect 328586 270345 331126 270373
rect 328586 270333 328592 270345
rect 331120 270333 331126 270345
rect 331178 270333 331184 270385
rect 338992 270333 338998 270385
rect 339050 270373 339056 270385
rect 352432 270373 352438 270385
rect 339050 270345 352438 270373
rect 339050 270333 339056 270345
rect 352432 270333 352438 270345
rect 352490 270333 352496 270385
rect 355600 270333 355606 270385
rect 355658 270373 355664 270385
rect 373840 270373 373846 270385
rect 355658 270345 373846 270373
rect 355658 270333 355664 270345
rect 373840 270333 373846 270345
rect 373898 270333 373904 270385
rect 375088 270333 375094 270385
rect 375146 270373 375152 270385
rect 379024 270373 379030 270385
rect 375146 270345 379030 270373
rect 375146 270333 375152 270345
rect 379024 270333 379030 270345
rect 379082 270333 379088 270385
rect 379216 270333 379222 270385
rect 379274 270373 379280 270385
rect 568912 270373 568918 270385
rect 379274 270345 568918 270373
rect 379274 270333 379280 270345
rect 568912 270333 568918 270345
rect 568970 270333 568976 270385
rect 245296 270259 245302 270311
rect 245354 270299 245360 270311
rect 332560 270299 332566 270311
rect 245354 270271 332566 270299
rect 245354 270259 245360 270271
rect 332560 270259 332566 270271
rect 332618 270259 332624 270311
rect 339184 270259 339190 270311
rect 339242 270299 339248 270311
rect 445264 270299 445270 270311
rect 339242 270271 379070 270299
rect 339242 270259 339248 270271
rect 233968 270185 233974 270237
rect 234026 270225 234032 270237
rect 338992 270225 338998 270237
rect 234026 270197 338998 270225
rect 234026 270185 234032 270197
rect 338992 270185 338998 270197
rect 339050 270185 339056 270237
rect 357616 270185 357622 270237
rect 357674 270225 357680 270237
rect 366160 270225 366166 270237
rect 357674 270197 366166 270225
rect 357674 270185 357680 270197
rect 366160 270185 366166 270197
rect 366218 270185 366224 270237
rect 367504 270185 367510 270237
rect 367562 270225 367568 270237
rect 378832 270225 378838 270237
rect 367562 270197 378838 270225
rect 367562 270185 367568 270197
rect 378832 270185 378838 270197
rect 378890 270185 378896 270237
rect 379042 270225 379070 270271
rect 379234 270271 445270 270299
rect 379234 270225 379262 270271
rect 445264 270259 445270 270271
rect 445322 270259 445328 270311
rect 469072 270259 469078 270311
rect 469130 270299 469136 270311
rect 469552 270299 469558 270311
rect 469130 270271 469558 270299
rect 469130 270259 469136 270271
rect 469552 270259 469558 270271
rect 469610 270259 469616 270311
rect 379042 270197 379262 270225
rect 379312 270185 379318 270237
rect 379370 270225 379376 270237
rect 576112 270225 576118 270237
rect 379370 270197 576118 270225
rect 379370 270185 379376 270197
rect 576112 270185 576118 270197
rect 576170 270185 576176 270237
rect 245872 270111 245878 270163
rect 245930 270151 245936 270163
rect 348304 270151 348310 270163
rect 245930 270123 348310 270151
rect 245930 270111 245936 270123
rect 348304 270111 348310 270123
rect 348362 270111 348368 270163
rect 352720 270111 352726 270163
rect 352778 270151 352784 270163
rect 452368 270151 452374 270163
rect 352778 270123 452374 270151
rect 352778 270111 352784 270123
rect 452368 270111 452374 270123
rect 452426 270111 452432 270163
rect 469360 270111 469366 270163
rect 469418 270151 469424 270163
rect 469552 270151 469558 270163
rect 469418 270123 469558 270151
rect 469418 270111 469424 270123
rect 469552 270111 469558 270123
rect 469610 270111 469616 270163
rect 234544 270037 234550 270089
rect 234602 270077 234608 270089
rect 342736 270077 342742 270089
rect 234602 270049 342742 270077
rect 234602 270037 234608 270049
rect 342736 270037 342742 270049
rect 342794 270037 342800 270089
rect 363088 270037 363094 270089
rect 363146 270077 363152 270089
rect 378928 270077 378934 270089
rect 363146 270049 378934 270077
rect 363146 270037 363152 270049
rect 378928 270037 378934 270049
rect 378986 270037 378992 270089
rect 379120 270037 379126 270089
rect 379178 270077 379184 270089
rect 379178 270049 387518 270077
rect 379178 270037 379184 270049
rect 98032 269963 98038 270015
rect 98090 270003 98096 270015
rect 100720 270003 100726 270015
rect 98090 269975 100726 270003
rect 98090 269963 98096 269975
rect 100720 269963 100726 269975
rect 100778 269963 100784 270015
rect 140752 269963 140758 270015
rect 140810 270003 140816 270015
rect 141040 270003 141046 270015
rect 140810 269975 141046 270003
rect 140810 269963 140816 269975
rect 141040 269963 141046 269975
rect 141098 269963 141104 270015
rect 194320 269963 194326 270015
rect 194378 270003 194384 270015
rect 314032 270003 314038 270015
rect 194378 269975 314038 270003
rect 194378 269963 194384 269975
rect 314032 269963 314038 269975
rect 314090 269963 314096 270015
rect 314416 269963 314422 270015
rect 314474 270003 314480 270015
rect 325456 270003 325462 270015
rect 314474 269975 325462 270003
rect 314474 269963 314480 269975
rect 325456 269963 325462 269975
rect 325514 269963 325520 270015
rect 325552 269963 325558 270015
rect 325610 270003 325616 270015
rect 371440 270003 371446 270015
rect 325610 269975 371446 270003
rect 325610 269963 325616 269975
rect 371440 269963 371446 269975
rect 371498 269963 371504 270015
rect 375760 269963 375766 270015
rect 375818 270003 375824 270015
rect 387376 270003 387382 270015
rect 375818 269975 387382 270003
rect 375818 269963 375824 269975
rect 387376 269963 387382 269975
rect 387434 269963 387440 270015
rect 387490 270003 387518 270049
rect 387568 270037 387574 270089
rect 387626 270077 387632 270089
rect 583216 270077 583222 270089
rect 387626 270049 583222 270077
rect 387626 270037 387632 270049
rect 583216 270037 583222 270049
rect 583274 270037 583280 270089
rect 669808 270037 669814 270089
rect 669866 270077 669872 270089
rect 674416 270077 674422 270089
rect 669866 270049 674422 270077
rect 669866 270037 669872 270049
rect 674416 270037 674422 270049
rect 674474 270037 674480 270089
rect 586768 270003 586774 270015
rect 387490 269975 586774 270003
rect 586768 269963 586774 269975
rect 586826 269963 586832 270015
rect 79024 269889 79030 269941
rect 79082 269929 79088 269941
rect 83440 269929 83446 269941
rect 79082 269901 83446 269929
rect 79082 269889 79088 269901
rect 83440 269889 83446 269901
rect 83498 269889 83504 269941
rect 247024 269889 247030 269941
rect 247082 269929 247088 269941
rect 459568 269929 459574 269941
rect 247082 269901 459574 269929
rect 247082 269889 247088 269901
rect 459568 269889 459574 269901
rect 459626 269889 459632 269941
rect 469456 269889 469462 269941
rect 469514 269929 469520 269941
rect 488272 269929 488278 269941
rect 469514 269901 488278 269929
rect 469514 269889 469520 269901
rect 488272 269889 488278 269901
rect 488330 269889 488336 269941
rect 226960 269815 226966 269867
rect 227018 269855 227024 269867
rect 295408 269855 295414 269867
rect 227018 269827 295414 269855
rect 227018 269815 227024 269827
rect 295408 269815 295414 269827
rect 295466 269815 295472 269867
rect 310288 269815 310294 269867
rect 310346 269855 310352 269867
rect 323344 269855 323350 269867
rect 310346 269827 323350 269855
rect 310346 269815 310352 269827
rect 323344 269815 323350 269827
rect 323402 269815 323408 269867
rect 323440 269815 323446 269867
rect 323498 269855 323504 269867
rect 325552 269855 325558 269867
rect 323498 269827 325558 269855
rect 323498 269815 323504 269827
rect 325552 269815 325558 269827
rect 325610 269815 325616 269867
rect 325648 269815 325654 269867
rect 325706 269855 325712 269867
rect 524944 269855 524950 269867
rect 325706 269827 524950 269855
rect 325706 269815 325712 269827
rect 524944 269815 524950 269827
rect 525002 269815 525008 269867
rect 235696 269741 235702 269793
rect 235754 269781 235760 269793
rect 366448 269781 366454 269793
rect 235754 269753 366454 269781
rect 235754 269741 235760 269753
rect 366448 269741 366454 269753
rect 366506 269741 366512 269793
rect 366544 269741 366550 269793
rect 366602 269781 366608 269793
rect 379024 269781 379030 269793
rect 366602 269753 379030 269781
rect 366602 269741 366608 269753
rect 379024 269741 379030 269753
rect 379082 269741 379088 269793
rect 379120 269741 379126 269793
rect 379178 269781 379184 269793
rect 597520 269781 597526 269793
rect 379178 269753 597526 269781
rect 379178 269741 379184 269753
rect 597520 269741 597526 269753
rect 597578 269741 597584 269793
rect 660976 269741 660982 269793
rect 661034 269781 661040 269793
rect 674704 269781 674710 269793
rect 661034 269753 674710 269781
rect 661034 269741 661040 269753
rect 674704 269741 674710 269753
rect 674762 269741 674768 269793
rect 247600 269667 247606 269719
rect 247658 269707 247664 269719
rect 466576 269707 466582 269719
rect 247658 269679 466582 269707
rect 247658 269667 247664 269679
rect 466576 269667 466582 269679
rect 466634 269667 466640 269719
rect 248560 269593 248566 269645
rect 248618 269633 248624 269645
rect 473776 269633 473782 269645
rect 248618 269605 473782 269633
rect 248618 269593 248624 269605
rect 473776 269593 473782 269605
rect 473834 269593 473840 269645
rect 236272 269519 236278 269571
rect 236330 269559 236336 269571
rect 358480 269559 358486 269571
rect 236330 269531 358486 269559
rect 236330 269519 236336 269531
rect 358480 269519 358486 269531
rect 358538 269519 358544 269571
rect 358576 269519 358582 269571
rect 358634 269559 358640 269571
rect 387280 269559 387286 269571
rect 358634 269531 387286 269559
rect 358634 269519 358640 269531
rect 387280 269519 387286 269531
rect 387338 269519 387344 269571
rect 387376 269519 387382 269571
rect 387434 269559 387440 269571
rect 604624 269559 604630 269571
rect 387434 269531 604630 269559
rect 387434 269519 387440 269531
rect 604624 269519 604630 269531
rect 604682 269519 604688 269571
rect 227536 269445 227542 269497
rect 227594 269485 227600 269497
rect 302608 269485 302614 269497
rect 227594 269457 302614 269485
rect 227594 269445 227600 269457
rect 302608 269445 302614 269457
rect 302666 269445 302672 269497
rect 312592 269445 312598 269497
rect 312650 269485 312656 269497
rect 542800 269485 542806 269497
rect 312650 269457 542806 269485
rect 312650 269445 312656 269457
rect 542800 269445 542806 269457
rect 542858 269445 542864 269497
rect 249616 269371 249622 269423
rect 249674 269411 249680 269423
rect 480976 269411 480982 269423
rect 249674 269383 480982 269411
rect 249674 269371 249680 269383
rect 480976 269371 480982 269383
rect 481034 269371 481040 269423
rect 228496 269297 228502 269349
rect 228554 269337 228560 269349
rect 309712 269337 309718 269349
rect 228554 269309 309718 269337
rect 228554 269297 228560 269309
rect 309712 269297 309718 269309
rect 309770 269297 309776 269349
rect 313840 269297 313846 269349
rect 313898 269337 313904 269349
rect 553456 269337 553462 269349
rect 313898 269309 553462 269337
rect 313898 269297 313904 269309
rect 553456 269297 553462 269309
rect 553514 269297 553520 269349
rect 221488 269223 221494 269275
rect 221546 269263 221552 269275
rect 251248 269263 251254 269275
rect 221546 269235 251254 269263
rect 221546 269223 221552 269235
rect 251248 269223 251254 269235
rect 251306 269223 251312 269275
rect 251344 269223 251350 269275
rect 251402 269263 251408 269275
rect 495184 269263 495190 269275
rect 251402 269235 495190 269263
rect 251402 269223 251408 269235
rect 495184 269223 495190 269235
rect 495242 269223 495248 269275
rect 243280 269149 243286 269201
rect 243338 269189 243344 269201
rect 431056 269189 431062 269201
rect 243338 269161 431062 269189
rect 243338 269149 243344 269161
rect 431056 269149 431062 269161
rect 431114 269149 431120 269201
rect 663952 269149 663958 269201
rect 664010 269189 664016 269201
rect 674704 269189 674710 269201
rect 664010 269161 674710 269189
rect 664010 269149 664016 269161
rect 674704 269149 674710 269161
rect 674762 269149 674768 269201
rect 242608 269075 242614 269127
rect 242666 269115 242672 269127
rect 423856 269115 423862 269127
rect 242666 269087 423862 269115
rect 242666 269075 242672 269087
rect 423856 269075 423862 269087
rect 423914 269075 423920 269127
rect 241552 269001 241558 269053
rect 241610 269041 241616 269053
rect 416656 269041 416662 269053
rect 241610 269013 416662 269041
rect 241610 269001 241616 269013
rect 416656 269001 416662 269013
rect 416714 269001 416720 269053
rect 428944 269001 428950 269053
rect 429002 269041 429008 269053
rect 429232 269041 429238 269053
rect 429002 269013 429238 269041
rect 429002 269001 429008 269013
rect 429232 269001 429238 269013
rect 429290 269001 429296 269053
rect 229552 268927 229558 268979
rect 229610 268967 229616 268979
rect 313936 268967 313942 268979
rect 229610 268939 313942 268967
rect 229610 268927 229616 268939
rect 313936 268927 313942 268939
rect 313994 268927 314000 268979
rect 314032 268927 314038 268979
rect 314090 268967 314096 268979
rect 325168 268967 325174 268979
rect 314090 268939 325174 268967
rect 314090 268927 314096 268939
rect 325168 268927 325174 268939
rect 325226 268927 325232 268979
rect 325264 268927 325270 268979
rect 325322 268967 325328 268979
rect 327088 268967 327094 268979
rect 325322 268939 327094 268967
rect 325322 268927 325328 268939
rect 327088 268927 327094 268939
rect 327146 268927 327152 268979
rect 327184 268927 327190 268979
rect 327242 268967 327248 268979
rect 336400 268967 336406 268979
rect 327242 268939 336406 268967
rect 327242 268927 327248 268939
rect 336400 268927 336406 268939
rect 336458 268927 336464 268979
rect 351760 268927 351766 268979
rect 351818 268967 351824 268979
rect 378352 268967 378358 268979
rect 351818 268939 378358 268967
rect 351818 268927 351824 268939
rect 378352 268927 378358 268939
rect 378410 268927 378416 268979
rect 378466 268939 378686 268967
rect 240880 268853 240886 268905
rect 240938 268893 240944 268905
rect 378466 268893 378494 268939
rect 240938 268865 378494 268893
rect 378658 268893 378686 268939
rect 378736 268927 378742 268979
rect 378794 268967 378800 268979
rect 387568 268967 387574 268979
rect 378794 268939 387574 268967
rect 378794 268927 378800 268939
rect 387568 268927 387574 268939
rect 387626 268927 387632 268979
rect 388624 268927 388630 268979
rect 388682 268967 388688 268979
rect 388912 268967 388918 268979
rect 388682 268939 388918 268967
rect 388682 268927 388688 268939
rect 388912 268927 388918 268939
rect 388970 268927 388976 268979
rect 390160 268927 390166 268979
rect 390218 268967 390224 268979
rect 395440 268967 395446 268979
rect 390218 268939 395446 268967
rect 390218 268927 390224 268939
rect 395440 268927 395446 268939
rect 395498 268927 395504 268979
rect 398800 268927 398806 268979
rect 398858 268967 398864 268979
rect 536848 268967 536854 268979
rect 398858 268939 536854 268967
rect 398858 268927 398864 268939
rect 536848 268927 536854 268939
rect 536906 268927 536912 268979
rect 409552 268893 409558 268905
rect 378658 268865 409558 268893
rect 240938 268853 240944 268865
rect 409552 268853 409558 268865
rect 409610 268853 409616 268905
rect 225808 268779 225814 268831
rect 225866 268819 225872 268831
rect 288208 268819 288214 268831
rect 225866 268791 288214 268819
rect 225866 268779 225872 268791
rect 288208 268779 288214 268791
rect 288266 268779 288272 268831
rect 313936 268779 313942 268831
rect 313994 268819 314000 268831
rect 316432 268819 316438 268831
rect 313994 268791 316438 268819
rect 313994 268779 314000 268791
rect 316432 268779 316438 268791
rect 316490 268779 316496 268831
rect 317680 268779 317686 268831
rect 317738 268819 317744 268831
rect 371440 268819 371446 268831
rect 317738 268791 371446 268819
rect 317738 268779 317744 268791
rect 371440 268779 371446 268791
rect 371498 268779 371504 268831
rect 371536 268779 371542 268831
rect 371594 268819 371600 268831
rect 372976 268819 372982 268831
rect 371594 268791 372982 268819
rect 371594 268779 371600 268791
rect 372976 268779 372982 268791
rect 373034 268779 373040 268831
rect 373360 268779 373366 268831
rect 373418 268819 373424 268831
rect 378736 268819 378742 268831
rect 373418 268791 378742 268819
rect 373418 268779 373424 268791
rect 378736 268779 378742 268791
rect 378794 268779 378800 268831
rect 379024 268779 379030 268831
rect 379082 268819 379088 268831
rect 529744 268819 529750 268831
rect 379082 268791 529750 268819
rect 379082 268779 379088 268791
rect 529744 268779 529750 268791
rect 529802 268779 529808 268831
rect 240016 268705 240022 268757
rect 240074 268745 240080 268757
rect 378640 268745 378646 268757
rect 240074 268717 378646 268745
rect 240074 268705 240080 268717
rect 378640 268705 378646 268717
rect 378698 268705 378704 268757
rect 378832 268705 378838 268757
rect 378890 268745 378896 268757
rect 398800 268745 398806 268757
rect 378890 268717 398806 268745
rect 378890 268705 378896 268717
rect 398800 268705 398806 268717
rect 398858 268705 398864 268757
rect 403216 268705 403222 268757
rect 403274 268745 403280 268757
rect 403984 268745 403990 268757
rect 403274 268717 403990 268745
rect 403274 268705 403280 268717
rect 403984 268705 403990 268717
rect 404042 268705 404048 268757
rect 210928 268631 210934 268683
rect 210986 268671 210992 268683
rect 271984 268671 271990 268683
rect 210986 268643 271990 268671
rect 210986 268631 210992 268643
rect 271984 268631 271990 268643
rect 272042 268631 272048 268683
rect 272752 268631 272758 268683
rect 272810 268671 272816 268683
rect 334960 268671 334966 268683
rect 272810 268643 334966 268671
rect 272810 268631 272816 268643
rect 334960 268631 334966 268643
rect 335018 268631 335024 268683
rect 348592 268631 348598 268683
rect 348650 268671 348656 268683
rect 373072 268671 373078 268683
rect 348650 268643 373078 268671
rect 348650 268631 348656 268643
rect 373072 268631 373078 268643
rect 373130 268631 373136 268683
rect 373168 268631 373174 268683
rect 373226 268671 373232 268683
rect 377008 268671 377014 268683
rect 373226 268643 377014 268671
rect 373226 268631 373232 268643
rect 377008 268631 377014 268643
rect 377066 268631 377072 268683
rect 377104 268631 377110 268683
rect 377162 268671 377168 268683
rect 526096 268671 526102 268683
rect 377162 268643 526102 268671
rect 377162 268631 377168 268643
rect 526096 268631 526102 268643
rect 526154 268631 526160 268683
rect 238864 268557 238870 268609
rect 238922 268597 238928 268609
rect 372976 268597 372982 268609
rect 238922 268569 372982 268597
rect 238922 268557 238928 268569
rect 372976 268557 372982 268569
rect 373034 268557 373040 268609
rect 378544 268597 378550 268609
rect 373090 268569 378550 268597
rect 238288 268483 238294 268535
rect 238346 268523 238352 268535
rect 371056 268523 371062 268535
rect 238346 268495 371062 268523
rect 238346 268483 238352 268495
rect 371056 268483 371062 268495
rect 371114 268483 371120 268535
rect 371344 268483 371350 268535
rect 371402 268523 371408 268535
rect 373090 268523 373118 268569
rect 378544 268557 378550 268569
rect 378602 268557 378608 268609
rect 378640 268557 378646 268609
rect 378698 268597 378704 268609
rect 402448 268597 402454 268609
rect 378698 268569 402454 268597
rect 378698 268557 378704 268569
rect 402448 268557 402454 268569
rect 402506 268557 402512 268609
rect 403696 268557 403702 268609
rect 403754 268597 403760 268609
rect 409936 268597 409942 268609
rect 403754 268569 409942 268597
rect 403754 268557 403760 268569
rect 409936 268557 409942 268569
rect 409994 268557 410000 268609
rect 371402 268495 373118 268523
rect 371402 268483 371408 268495
rect 373168 268483 373174 268535
rect 373226 268523 373232 268535
rect 382384 268523 382390 268535
rect 373226 268495 382390 268523
rect 373226 268483 373232 268495
rect 382384 268483 382390 268495
rect 382442 268483 382448 268535
rect 382480 268483 382486 268535
rect 382538 268523 382544 268535
rect 395344 268523 395350 268535
rect 382538 268495 395350 268523
rect 382538 268483 382544 268495
rect 395344 268483 395350 268495
rect 395402 268483 395408 268535
rect 395440 268483 395446 268535
rect 395498 268523 395504 268535
rect 408112 268523 408118 268535
rect 395498 268495 408118 268523
rect 395498 268483 395504 268495
rect 408112 268483 408118 268495
rect 408170 268483 408176 268535
rect 237136 268409 237142 268461
rect 237194 268449 237200 268461
rect 357616 268449 357622 268461
rect 237194 268421 357622 268449
rect 237194 268409 237200 268421
rect 357616 268409 357622 268421
rect 357674 268409 357680 268461
rect 357712 268409 357718 268461
rect 357770 268449 357776 268461
rect 358576 268449 358582 268461
rect 357770 268421 358582 268449
rect 357770 268409 357776 268421
rect 358576 268409 358582 268421
rect 358634 268409 358640 268461
rect 366352 268409 366358 268461
rect 366410 268449 366416 268461
rect 377104 268449 377110 268461
rect 366410 268421 377110 268449
rect 366410 268409 366416 268421
rect 377104 268409 377110 268421
rect 377162 268409 377168 268461
rect 377200 268409 377206 268461
rect 377258 268449 377264 268461
rect 390448 268449 390454 268461
rect 377258 268421 390454 268449
rect 377258 268409 377264 268421
rect 390448 268409 390454 268421
rect 390506 268409 390512 268461
rect 403696 268409 403702 268461
rect 403754 268449 403760 268461
rect 406096 268449 406102 268461
rect 403754 268421 406102 268449
rect 403754 268409 403760 268421
rect 406096 268409 406102 268421
rect 406154 268409 406160 268461
rect 499408 268409 499414 268461
rect 499466 268449 499472 268461
rect 502000 268449 502006 268461
rect 499466 268421 502006 268449
rect 499466 268409 499472 268421
rect 502000 268409 502006 268421
rect 502058 268409 502064 268461
rect 218032 268335 218038 268387
rect 218090 268375 218096 268387
rect 272656 268375 272662 268387
rect 218090 268347 272662 268375
rect 218090 268335 218096 268347
rect 272656 268335 272662 268347
rect 272714 268335 272720 268387
rect 283504 268335 283510 268387
rect 283562 268375 283568 268387
rect 336496 268375 336502 268387
rect 283562 268347 336502 268375
rect 283562 268335 283568 268347
rect 336496 268335 336502 268347
rect 336554 268335 336560 268387
rect 357232 268335 357238 268387
rect 357290 268375 357296 268387
rect 358864 268375 358870 268387
rect 357290 268347 358870 268375
rect 357290 268335 357296 268347
rect 358864 268335 358870 268347
rect 358922 268335 358928 268387
rect 359440 268335 359446 268387
rect 359498 268375 359504 268387
rect 378640 268375 378646 268387
rect 359498 268347 378646 268375
rect 359498 268335 359504 268347
rect 378640 268335 378646 268347
rect 378698 268335 378704 268387
rect 378928 268335 378934 268387
rect 378986 268375 378992 268387
rect 501136 268375 501142 268387
rect 378986 268347 501142 268375
rect 378986 268335 378992 268347
rect 501136 268335 501142 268347
rect 501194 268335 501200 268387
rect 228784 268261 228790 268313
rect 228842 268301 228848 268313
rect 274192 268301 274198 268313
rect 228842 268273 274198 268301
rect 228842 268261 228848 268273
rect 274192 268261 274198 268273
rect 274250 268261 274256 268313
rect 290608 268261 290614 268313
rect 290666 268301 290672 268313
rect 337456 268301 337462 268313
rect 290666 268273 337462 268301
rect 290666 268261 290672 268273
rect 337456 268261 337462 268273
rect 337514 268261 337520 268313
rect 353968 268261 353974 268313
rect 354026 268301 354032 268313
rect 354026 268273 359102 268301
rect 354026 268261 354032 268273
rect 222544 268187 222550 268239
rect 222602 268227 222608 268239
rect 259696 268227 259702 268239
rect 222602 268199 259702 268227
rect 222602 268187 222608 268199
rect 259696 268187 259702 268199
rect 259754 268187 259760 268239
rect 260080 268187 260086 268239
rect 260138 268227 260144 268239
rect 355600 268227 355606 268239
rect 260138 268199 355606 268227
rect 260138 268187 260144 268199
rect 355600 268187 355606 268199
rect 355658 268187 355664 268239
rect 358384 268187 358390 268239
rect 358442 268227 358448 268239
rect 359074 268227 359102 268273
rect 360976 268261 360982 268313
rect 361034 268301 361040 268313
rect 483280 268301 483286 268313
rect 361034 268273 483286 268301
rect 361034 268261 361040 268273
rect 483280 268261 483286 268273
rect 483338 268261 483344 268313
rect 426256 268227 426262 268239
rect 358442 268199 358910 268227
rect 359074 268199 426262 268227
rect 358442 268187 358448 268199
rect 223216 268113 223222 268165
rect 223274 268153 223280 268165
rect 266800 268153 266806 268165
rect 223274 268125 266806 268153
rect 223274 268113 223280 268125
rect 266800 268113 266806 268125
rect 266858 268113 266864 268165
rect 287056 268113 287062 268165
rect 287114 268153 287120 268165
rect 287114 268125 316286 268153
rect 287114 268113 287120 268125
rect 235888 268039 235894 268091
rect 235946 268079 235952 268091
rect 274864 268079 274870 268091
rect 235946 268051 274870 268079
rect 235946 268039 235952 268051
rect 274864 268039 274870 268051
rect 274922 268039 274928 268091
rect 294544 268039 294550 268091
rect 294602 268079 294608 268091
rect 315952 268079 315958 268091
rect 294602 268051 315958 268079
rect 294602 268039 294608 268051
rect 315952 268039 315958 268051
rect 316010 268039 316016 268091
rect 221968 267965 221974 268017
rect 222026 268005 222032 268017
rect 256144 268005 256150 268017
rect 222026 267977 256150 268005
rect 222026 267965 222032 267977
rect 256144 267965 256150 267977
rect 256202 267965 256208 268017
rect 286000 267965 286006 268017
rect 286058 268005 286064 268017
rect 316144 268005 316150 268017
rect 286058 267977 316150 268005
rect 286058 267965 286064 267977
rect 316144 267965 316150 267977
rect 316202 267965 316208 268017
rect 316258 268005 316286 268125
rect 316528 268113 316534 268165
rect 316586 268153 316592 268165
rect 337840 268153 337846 268165
rect 316586 268125 337846 268153
rect 316586 268113 316592 268125
rect 337840 268113 337846 268125
rect 337898 268113 337904 268165
rect 358882 268153 358910 268199
rect 426256 268187 426262 268199
rect 426314 268187 426320 268239
rect 499312 268187 499318 268239
rect 499370 268227 499376 268239
rect 499792 268227 499798 268239
rect 499370 268199 499798 268227
rect 499370 268187 499376 268199
rect 499792 268187 499798 268199
rect 499850 268187 499856 268239
rect 370864 268153 370870 268165
rect 358882 268125 370870 268153
rect 370864 268113 370870 268125
rect 370922 268113 370928 268165
rect 372496 268113 372502 268165
rect 372554 268153 372560 268165
rect 378544 268153 378550 268165
rect 372554 268125 378550 268153
rect 372554 268113 372560 268125
rect 378544 268113 378550 268125
rect 378602 268113 378608 268165
rect 378640 268113 378646 268165
rect 378698 268153 378704 268165
rect 468976 268153 468982 268165
rect 378698 268125 468982 268153
rect 378698 268113 378704 268125
rect 468976 268113 468982 268125
rect 469034 268113 469040 268165
rect 316432 268039 316438 268091
rect 316490 268079 316496 268091
rect 322960 268079 322966 268091
rect 316490 268051 322966 268079
rect 316490 268039 316496 268051
rect 322960 268039 322966 268051
rect 323018 268039 323024 268091
rect 323056 268039 323062 268091
rect 323114 268079 323120 268091
rect 326896 268079 326902 268091
rect 323114 268051 326902 268079
rect 323114 268039 323120 268051
rect 326896 268039 326902 268051
rect 326954 268039 326960 268091
rect 326992 268039 326998 268091
rect 327050 268079 327056 268091
rect 327050 268051 328958 268079
rect 327050 268039 327056 268051
rect 324496 268005 324502 268017
rect 316258 267977 324502 268005
rect 324496 267965 324502 267977
rect 324554 267965 324560 268017
rect 324592 267965 324598 268017
rect 324650 268005 324656 268017
rect 328624 268005 328630 268017
rect 324650 267977 328630 268005
rect 324650 267965 324656 267977
rect 328624 267965 328630 267977
rect 328682 267965 328688 268017
rect 328930 268005 328958 268051
rect 329008 268039 329014 268091
rect 329066 268079 329072 268091
rect 348592 268079 348598 268091
rect 329066 268051 348598 268079
rect 329066 268039 329072 268051
rect 348592 268039 348598 268051
rect 348650 268039 348656 268091
rect 371536 268079 371542 268091
rect 348802 268051 371542 268079
rect 336112 268005 336118 268017
rect 328930 267977 336118 268005
rect 336112 267965 336118 267977
rect 336170 267965 336176 268017
rect 336208 267965 336214 268017
rect 336266 268005 336272 268017
rect 348802 268005 348830 268051
rect 371536 268039 371542 268051
rect 371594 268039 371600 268091
rect 371632 268039 371638 268091
rect 371690 268079 371696 268091
rect 387184 268079 387190 268091
rect 371690 268051 387190 268079
rect 371690 268039 371696 268051
rect 387184 268039 387190 268051
rect 387242 268039 387248 268091
rect 387280 268039 387286 268091
rect 387338 268079 387344 268091
rect 454768 268079 454774 268091
rect 387338 268051 454774 268079
rect 387338 268039 387344 268051
rect 454768 268039 454774 268051
rect 454826 268039 454832 268091
rect 336266 267977 348830 268005
rect 336266 267965 336272 267977
rect 355696 267965 355702 268017
rect 355754 268005 355760 268017
rect 440464 268005 440470 268017
rect 355754 267977 440470 268005
rect 355754 267965 355760 267977
rect 440464 267965 440470 267977
rect 440522 267965 440528 268017
rect 243088 267891 243094 267943
rect 243146 267931 243152 267943
rect 275728 267931 275734 267943
rect 243146 267903 275734 267931
rect 243146 267891 243152 267903
rect 275728 267891 275734 267903
rect 275786 267891 275792 267943
rect 285040 267891 285046 267943
rect 285098 267931 285104 267943
rect 317776 267931 317782 267943
rect 285098 267903 317782 267931
rect 285098 267891 285104 267903
rect 317776 267891 317782 267903
rect 317834 267891 317840 267943
rect 322384 267891 322390 267943
rect 322442 267931 322448 267943
rect 326800 267931 326806 267943
rect 322442 267903 326806 267931
rect 322442 267891 322448 267903
rect 326800 267891 326806 267903
rect 326858 267891 326864 267943
rect 326896 267891 326902 267943
rect 326954 267931 326960 267943
rect 377776 267931 377782 267943
rect 326954 267903 358526 267931
rect 326954 267891 326960 267903
rect 65008 267817 65014 267869
rect 65066 267857 65072 267869
rect 67600 267857 67606 267869
rect 65066 267829 67606 267857
rect 65066 267817 65072 267829
rect 67600 267817 67606 267829
rect 67658 267817 67664 267869
rect 258544 267817 258550 267869
rect 258602 267857 258608 267869
rect 358384 267857 358390 267869
rect 258602 267829 358390 267857
rect 258602 267817 258608 267829
rect 358384 267817 358390 267829
rect 358442 267817 358448 267869
rect 358498 267857 358526 267903
rect 358786 267903 377782 267931
rect 358786 267857 358814 267903
rect 377776 267891 377782 267903
rect 377834 267891 377840 267943
rect 378352 267891 378358 267943
rect 378410 267931 378416 267943
rect 378410 267903 378590 267931
rect 378410 267891 378416 267903
rect 358498 267829 358814 267857
rect 358864 267817 358870 267869
rect 358922 267857 358928 267869
rect 371632 267857 371638 267869
rect 358922 267829 371638 267857
rect 358922 267817 358928 267829
rect 371632 267817 371638 267829
rect 371690 267817 371696 267869
rect 372976 267817 372982 267869
rect 373034 267857 373040 267869
rect 377296 267857 377302 267869
rect 373034 267829 377302 267857
rect 373034 267817 373040 267829
rect 377296 267817 377302 267829
rect 377354 267817 377360 267869
rect 377488 267817 377494 267869
rect 377546 267857 377552 267869
rect 378448 267857 378454 267869
rect 377546 267829 378454 267857
rect 377546 267817 377552 267829
rect 378448 267817 378454 267829
rect 378506 267817 378512 267869
rect 378562 267857 378590 267903
rect 379312 267891 379318 267943
rect 379370 267931 379376 267943
rect 386512 267931 386518 267943
rect 379370 267903 386518 267931
rect 379370 267891 379376 267903
rect 386512 267891 386518 267903
rect 386570 267891 386576 267943
rect 388720 267891 388726 267943
rect 388778 267931 388784 267943
rect 390352 267931 390358 267943
rect 388778 267903 390358 267931
rect 388778 267891 388784 267903
rect 390352 267891 390358 267903
rect 390410 267891 390416 267943
rect 390448 267891 390454 267943
rect 390506 267931 390512 267943
rect 413392 267931 413398 267943
rect 390506 267903 413398 267931
rect 390506 267891 390512 267903
rect 413392 267891 413398 267903
rect 413450 267891 413456 267943
rect 390160 267857 390166 267869
rect 378562 267829 390166 267857
rect 390160 267817 390166 267829
rect 390218 267817 390224 267869
rect 390256 267817 390262 267869
rect 390314 267857 390320 267869
rect 413296 267857 413302 267869
rect 390314 267829 413302 267857
rect 390314 267817 390320 267829
rect 413296 267817 413302 267829
rect 413354 267817 413360 267869
rect 204976 267743 204982 267795
rect 205034 267783 205040 267795
rect 312688 267783 312694 267795
rect 205034 267755 312694 267783
rect 205034 267743 205040 267755
rect 312688 267743 312694 267755
rect 312746 267743 312752 267795
rect 319408 267743 319414 267795
rect 319466 267783 319472 267795
rect 322384 267783 322390 267795
rect 319466 267755 322390 267783
rect 319466 267743 319472 267755
rect 322384 267743 322390 267755
rect 322442 267743 322448 267795
rect 322480 267743 322486 267795
rect 322538 267783 322544 267795
rect 621232 267783 621238 267795
rect 322538 267755 621238 267783
rect 322538 267743 322544 267755
rect 621232 267743 621238 267755
rect 621290 267743 621296 267795
rect 276208 267669 276214 267721
rect 276266 267709 276272 267721
rect 298000 267709 298006 267721
rect 276266 267681 298006 267709
rect 276266 267669 276272 267681
rect 298000 267669 298006 267681
rect 298058 267669 298064 267721
rect 326704 267709 326710 267721
rect 298114 267681 326710 267709
rect 287728 267595 287734 267647
rect 287786 267635 287792 267647
rect 297808 267635 297814 267647
rect 287786 267607 297814 267635
rect 287786 267595 287792 267607
rect 297808 267595 297814 267607
rect 297866 267595 297872 267647
rect 279952 267521 279958 267573
rect 280010 267561 280016 267573
rect 298114 267561 298142 267681
rect 326704 267669 326710 267681
rect 326762 267669 326768 267721
rect 326800 267669 326806 267721
rect 326858 267709 326864 267721
rect 376048 267709 376054 267721
rect 326858 267681 376054 267709
rect 326858 267669 326864 267681
rect 376048 267669 376054 267681
rect 376106 267669 376112 267721
rect 378448 267669 378454 267721
rect 378506 267709 378512 267721
rect 379312 267709 379318 267721
rect 378506 267681 379318 267709
rect 378506 267669 378512 267681
rect 379312 267669 379318 267681
rect 379370 267669 379376 267721
rect 379408 267669 379414 267721
rect 379466 267709 379472 267721
rect 389104 267709 389110 267721
rect 379466 267681 389110 267709
rect 379466 267669 379472 267681
rect 389104 267669 389110 267681
rect 389162 267669 389168 267721
rect 389200 267669 389206 267721
rect 389258 267709 389264 267721
rect 414352 267709 414358 267721
rect 389258 267681 414358 267709
rect 389258 267669 389264 267681
rect 414352 267669 414358 267681
rect 414410 267669 414416 267721
rect 298384 267595 298390 267647
rect 298442 267635 298448 267647
rect 327952 267635 327958 267647
rect 298442 267607 327958 267635
rect 298442 267595 298448 267607
rect 327952 267595 327958 267607
rect 328010 267595 328016 267647
rect 377200 267635 377206 267647
rect 328546 267607 377206 267635
rect 280010 267533 298142 267561
rect 280010 267521 280016 267533
rect 311920 267521 311926 267573
rect 311978 267561 311984 267573
rect 320560 267561 320566 267573
rect 311978 267533 320566 267561
rect 311978 267521 311984 267533
rect 320560 267521 320566 267533
rect 320618 267521 320624 267573
rect 321520 267521 321526 267573
rect 321578 267561 321584 267573
rect 328546 267561 328574 267607
rect 377200 267595 377206 267607
rect 377258 267595 377264 267647
rect 377296 267595 377302 267647
rect 377354 267635 377360 267647
rect 382480 267635 382486 267647
rect 377354 267607 382486 267635
rect 377354 267595 377360 267607
rect 382480 267595 382486 267607
rect 382538 267595 382544 267647
rect 383056 267595 383062 267647
rect 383114 267635 383120 267647
rect 385456 267635 385462 267647
rect 383114 267607 385462 267635
rect 383114 267595 383120 267607
rect 385456 267595 385462 267607
rect 385514 267595 385520 267647
rect 387184 267595 387190 267647
rect 387242 267635 387248 267647
rect 389008 267635 389014 267647
rect 387242 267607 389014 267635
rect 387242 267595 387248 267607
rect 389008 267595 389014 267607
rect 389066 267595 389072 267647
rect 390352 267595 390358 267647
rect 390410 267635 390416 267647
rect 399856 267635 399862 267647
rect 390410 267607 399862 267635
rect 390410 267595 390416 267607
rect 399856 267595 399862 267607
rect 399914 267595 399920 267647
rect 403024 267595 403030 267647
rect 403082 267635 403088 267647
rect 410992 267635 410998 267647
rect 403082 267607 410998 267635
rect 403082 267595 403088 267607
rect 410992 267595 410998 267607
rect 411050 267595 411056 267647
rect 321578 267533 328574 267561
rect 321578 267521 321584 267533
rect 328624 267521 328630 267573
rect 328682 267561 328688 267573
rect 328682 267533 338462 267561
rect 328682 267521 328688 267533
rect 138352 267447 138358 267499
rect 138410 267487 138416 267499
rect 140944 267487 140950 267499
rect 138410 267459 140950 267487
rect 138410 267447 138416 267459
rect 140944 267447 140950 267459
rect 141002 267447 141008 267499
rect 290320 267447 290326 267499
rect 290378 267487 290384 267499
rect 338320 267487 338326 267499
rect 290378 267459 338326 267487
rect 290378 267447 290384 267459
rect 338320 267447 338326 267459
rect 338378 267447 338384 267499
rect 338434 267487 338462 267533
rect 353296 267521 353302 267573
rect 353354 267561 353360 267573
rect 419056 267561 419062 267573
rect 353354 267533 419062 267561
rect 353354 267521 353360 267533
rect 419056 267521 419062 267533
rect 419114 267521 419120 267573
rect 357232 267487 357238 267499
rect 338434 267459 357238 267487
rect 357232 267447 357238 267459
rect 357290 267447 357296 267499
rect 357328 267447 357334 267499
rect 357386 267487 357392 267499
rect 368272 267487 368278 267499
rect 357386 267459 368278 267487
rect 357386 267447 357392 267459
rect 368272 267447 368278 267459
rect 368330 267447 368336 267499
rect 368368 267447 368374 267499
rect 368426 267487 368432 267499
rect 377680 267487 377686 267499
rect 368426 267459 377686 267487
rect 368426 267447 368432 267459
rect 377680 267447 377686 267459
rect 377738 267447 377744 267499
rect 377776 267447 377782 267499
rect 377834 267487 377840 267499
rect 378928 267487 378934 267499
rect 377834 267459 378934 267487
rect 377834 267447 377840 267459
rect 378928 267447 378934 267459
rect 378986 267447 378992 267499
rect 379024 267447 379030 267499
rect 379082 267487 379088 267499
rect 382768 267487 382774 267499
rect 379082 267459 382774 267487
rect 379082 267447 379088 267459
rect 382768 267447 382774 267459
rect 382826 267447 382832 267499
rect 389008 267447 389014 267499
rect 389066 267487 389072 267499
rect 390256 267487 390262 267499
rect 389066 267459 390262 267487
rect 389066 267447 389072 267459
rect 390256 267447 390262 267459
rect 390314 267447 390320 267499
rect 395632 267447 395638 267499
rect 395690 267487 395696 267499
rect 398704 267487 398710 267499
rect 395690 267459 398710 267487
rect 395690 267447 395696 267459
rect 398704 267447 398710 267459
rect 398762 267447 398768 267499
rect 398800 267447 398806 267499
rect 398858 267487 398864 267499
rect 421456 267487 421462 267499
rect 398858 267459 421462 267487
rect 398858 267447 398864 267459
rect 421456 267447 421462 267459
rect 421514 267447 421520 267499
rect 288784 267373 288790 267425
rect 288842 267413 288848 267425
rect 346576 267413 346582 267425
rect 288842 267385 346582 267413
rect 288842 267373 288848 267385
rect 346576 267373 346582 267385
rect 346634 267373 346640 267425
rect 355024 267373 355030 267425
rect 355082 267413 355088 267425
rect 433360 267413 433366 267425
rect 355082 267385 433366 267413
rect 355082 267373 355088 267385
rect 433360 267373 433366 267385
rect 433418 267373 433424 267425
rect 291664 267299 291670 267351
rect 291722 267339 291728 267351
rect 363856 267339 363862 267351
rect 291722 267311 363862 267339
rect 291722 267299 291728 267311
rect 363856 267299 363862 267311
rect 363914 267299 363920 267351
rect 368272 267299 368278 267351
rect 368330 267339 368336 267351
rect 378640 267339 378646 267351
rect 368330 267311 378646 267339
rect 368330 267299 368336 267311
rect 378640 267299 378646 267311
rect 378698 267299 378704 267351
rect 379504 267299 379510 267351
rect 379562 267339 379568 267351
rect 383056 267339 383062 267351
rect 379562 267311 383062 267339
rect 379562 267299 379568 267311
rect 383056 267299 383062 267311
rect 383114 267299 383120 267351
rect 387856 267299 387862 267351
rect 387914 267339 387920 267351
rect 629680 267339 629686 267351
rect 387914 267311 629686 267339
rect 387914 267299 387920 267311
rect 629680 267299 629686 267311
rect 629738 267299 629744 267351
rect 289456 267225 289462 267277
rect 289514 267265 289520 267277
rect 353680 267265 353686 267277
rect 289514 267237 353686 267265
rect 289514 267225 289520 267237
rect 353680 267225 353686 267237
rect 353738 267225 353744 267277
rect 356560 267225 356566 267277
rect 356618 267265 356624 267277
rect 447664 267265 447670 267277
rect 356618 267237 447670 267265
rect 356618 267225 356624 267237
rect 447664 267225 447670 267237
rect 447722 267225 447728 267277
rect 293584 267151 293590 267203
rect 293642 267191 293648 267203
rect 379024 267191 379030 267203
rect 293642 267163 379030 267191
rect 293642 267151 293648 267163
rect 379024 267151 379030 267163
rect 379082 267151 379088 267203
rect 379120 267151 379126 267203
rect 379178 267191 379184 267203
rect 387856 267191 387862 267203
rect 379178 267163 387862 267191
rect 379178 267151 379184 267163
rect 387856 267151 387862 267163
rect 387914 267151 387920 267203
rect 388528 267151 388534 267203
rect 388586 267191 388592 267203
rect 419344 267191 419350 267203
rect 388586 267163 419350 267191
rect 388586 267151 388592 267163
rect 419344 267151 419350 267163
rect 419402 267151 419408 267203
rect 262384 267077 262390 267129
rect 262442 267117 262448 267129
rect 333904 267117 333910 267129
rect 262442 267089 333910 267117
rect 262442 267077 262448 267089
rect 333904 267077 333910 267089
rect 333962 267077 333968 267129
rect 351280 267077 351286 267129
rect 351338 267117 351344 267129
rect 357328 267117 357334 267129
rect 351338 267089 357334 267117
rect 351338 267077 351344 267089
rect 357328 267077 357334 267089
rect 357386 267077 357392 267129
rect 357808 267077 357814 267129
rect 357866 267117 357872 267129
rect 458320 267117 458326 267129
rect 357866 267089 458326 267117
rect 357866 267077 357872 267089
rect 458320 267077 458326 267089
rect 458378 267077 458384 267129
rect 295312 267003 295318 267055
rect 295370 267043 295376 267055
rect 378736 267043 378742 267055
rect 295370 267015 378742 267043
rect 295370 267003 295376 267015
rect 378736 267003 378742 267015
rect 378794 267003 378800 267055
rect 378832 267003 378838 267055
rect 378890 267043 378896 267055
rect 398896 267043 398902 267055
rect 378890 267015 398902 267043
rect 378890 267003 378896 267015
rect 398896 267003 398902 267015
rect 398954 267003 398960 267055
rect 403120 267003 403126 267055
rect 403178 267043 403184 267055
rect 411952 267043 411958 267055
rect 403178 267015 411958 267043
rect 403178 267003 403184 267015
rect 411952 267003 411958 267015
rect 412010 267003 412016 267055
rect 295984 266929 295990 266981
rect 296042 266969 296048 266981
rect 389008 266969 389014 266981
rect 296042 266941 389014 266969
rect 296042 266929 296048 266941
rect 389008 266929 389014 266941
rect 389066 266929 389072 266981
rect 389104 266929 389110 266981
rect 389162 266969 389168 266981
rect 404752 266969 404758 266981
rect 389162 266941 404758 266969
rect 389162 266929 389168 266941
rect 404752 266929 404758 266941
rect 404810 266929 404816 266981
rect 408208 266929 408214 266981
rect 408266 266969 408272 266981
rect 408688 266969 408694 266981
rect 408266 266941 408694 266969
rect 408266 266929 408272 266941
rect 408688 266929 408694 266941
rect 408746 266929 408752 266981
rect 251152 266855 251158 266907
rect 251210 266895 251216 266907
rect 332368 266895 332374 266907
rect 251210 266867 332374 266895
rect 251210 266855 251216 266867
rect 332368 266855 332374 266867
rect 332426 266855 332432 266907
rect 359824 266855 359830 266907
rect 359882 266895 359888 266907
rect 472624 266895 472630 266907
rect 359882 266867 472630 266895
rect 359882 266855 359888 266867
rect 472624 266855 472630 266867
rect 472682 266855 472688 266907
rect 296848 266781 296854 266833
rect 296906 266821 296912 266833
rect 389200 266821 389206 266833
rect 296906 266793 389206 266821
rect 296906 266781 296912 266793
rect 389200 266781 389206 266793
rect 389258 266781 389264 266833
rect 389296 266781 389302 266833
rect 389354 266821 389360 266833
rect 412912 266821 412918 266833
rect 389354 266793 412918 266821
rect 389354 266781 389360 266793
rect 412912 266781 412918 266793
rect 412970 266781 412976 266833
rect 298000 266707 298006 266759
rect 298058 266747 298064 266759
rect 398800 266747 398806 266759
rect 298058 266719 398806 266747
rect 298058 266707 298064 266719
rect 398800 266707 398806 266719
rect 398858 266707 398864 266759
rect 398992 266707 398998 266759
rect 399050 266747 399056 266759
rect 408208 266747 408214 266759
rect 399050 266719 408214 266747
rect 399050 266707 399056 266719
rect 408208 266707 408214 266719
rect 408266 266707 408272 266759
rect 408400 266707 408406 266759
rect 408458 266747 408464 266759
rect 413296 266747 413302 266759
rect 408458 266719 413302 266747
rect 408458 266707 408464 266719
rect 413296 266707 413302 266719
rect 413354 266707 413360 266759
rect 298576 266633 298582 266685
rect 298634 266673 298640 266685
rect 428656 266673 428662 266685
rect 298634 266645 428662 266673
rect 298634 266633 298640 266645
rect 428656 266633 428662 266645
rect 428714 266633 428720 266685
rect 244240 266559 244246 266611
rect 244298 266599 244304 266611
rect 331696 266599 331702 266611
rect 244298 266571 331702 266599
rect 244298 266559 244304 266571
rect 331696 266559 331702 266571
rect 331754 266559 331760 266611
rect 338320 266559 338326 266611
rect 338378 266599 338384 266611
rect 360784 266599 360790 266611
rect 338378 266571 360790 266599
rect 338378 266559 338384 266571
rect 360784 266559 360790 266571
rect 360842 266559 360848 266611
rect 362224 266559 362230 266611
rect 362282 266599 362288 266611
rect 494032 266599 494038 266611
rect 362282 266571 494038 266599
rect 362282 266559 362288 266571
rect 494032 266559 494038 266571
rect 494090 266559 494096 266611
rect 237424 266485 237430 266537
rect 237482 266525 237488 266537
rect 330640 266525 330646 266537
rect 237482 266497 330646 266525
rect 237482 266485 237488 266497
rect 330640 266485 330646 266497
rect 330698 266485 330704 266537
rect 362704 266485 362710 266537
rect 362762 266525 362768 266537
rect 497584 266525 497590 266537
rect 362762 266497 497590 266525
rect 362762 266485 362768 266497
rect 497584 266485 497590 266497
rect 497642 266485 497648 266537
rect 299728 266411 299734 266463
rect 299786 266451 299792 266463
rect 435664 266451 435670 266463
rect 299786 266423 435670 266451
rect 299786 266411 299792 266423
rect 435664 266411 435670 266423
rect 435722 266411 435728 266463
rect 300304 266337 300310 266389
rect 300362 266377 300368 266389
rect 442864 266377 442870 266389
rect 300362 266349 442870 266377
rect 300362 266337 300368 266349
rect 442864 266337 442870 266349
rect 442922 266337 442928 266389
rect 521584 266337 521590 266389
rect 521642 266377 521648 266389
rect 523504 266377 523510 266389
rect 521642 266349 523510 266377
rect 521642 266337 521648 266349
rect 523504 266337 523510 266349
rect 523562 266337 523568 266389
rect 301264 266263 301270 266315
rect 301322 266303 301328 266315
rect 449968 266303 449974 266315
rect 301322 266275 449974 266303
rect 301322 266263 301328 266275
rect 449968 266263 449974 266275
rect 450026 266263 450032 266315
rect 230032 266189 230038 266241
rect 230090 266229 230096 266241
rect 329968 266229 329974 266241
rect 230090 266201 329974 266229
rect 230090 266189 230096 266201
rect 329968 266189 329974 266201
rect 330026 266189 330032 266241
rect 365968 266189 365974 266241
rect 366026 266229 366032 266241
rect 522544 266229 522550 266241
rect 366026 266201 522550 266229
rect 366026 266189 366032 266201
rect 522544 266189 522550 266201
rect 522602 266189 522608 266241
rect 302320 266115 302326 266167
rect 302378 266155 302384 266167
rect 457168 266155 457174 266167
rect 302378 266127 457174 266155
rect 302378 266115 302384 266127
rect 457168 266115 457174 266127
rect 457226 266115 457232 266167
rect 302992 266041 302998 266093
rect 303050 266081 303056 266093
rect 464272 266081 464278 266093
rect 303050 266053 464278 266081
rect 303050 266041 303056 266053
rect 464272 266041 464278 266053
rect 464330 266041 464336 266093
rect 304048 265967 304054 266019
rect 304106 266007 304112 266019
rect 471376 266007 471382 266019
rect 304106 265979 471382 266007
rect 304106 265967 304112 265979
rect 471376 265967 471382 265979
rect 471434 265967 471440 266019
rect 226384 265893 226390 265945
rect 226442 265933 226448 265945
rect 329584 265933 329590 265945
rect 226442 265905 329590 265933
rect 226442 265893 226448 265905
rect 329584 265893 329590 265905
rect 329642 265893 329648 265945
rect 367024 265893 367030 265945
rect 367082 265933 367088 265945
rect 378832 265933 378838 265945
rect 367082 265905 378838 265933
rect 367082 265893 367088 265905
rect 378832 265893 378838 265905
rect 378890 265893 378896 265945
rect 378928 265893 378934 265945
rect 378986 265933 378992 265945
rect 398800 265933 398806 265945
rect 378986 265905 398806 265933
rect 378986 265893 378992 265905
rect 398800 265893 398806 265905
rect 398858 265893 398864 265945
rect 398896 265893 398902 265945
rect 398954 265933 398960 265945
rect 533200 265933 533206 265945
rect 398954 265905 533206 265933
rect 398954 265893 398960 265905
rect 533200 265893 533206 265905
rect 533258 265893 533264 265945
rect 304720 265819 304726 265871
rect 304778 265859 304784 265871
rect 478576 265859 478582 265871
rect 304778 265831 478582 265859
rect 304778 265819 304784 265831
rect 478576 265819 478582 265831
rect 478634 265819 478640 265871
rect 305584 265745 305590 265797
rect 305642 265785 305648 265797
rect 485680 265785 485686 265797
rect 305642 265757 485686 265785
rect 305642 265745 305648 265757
rect 485680 265745 485686 265757
rect 485738 265745 485744 265797
rect 212464 265671 212470 265723
rect 212522 265711 212528 265723
rect 327856 265711 327862 265723
rect 212522 265683 327862 265711
rect 212522 265671 212528 265683
rect 327856 265671 327862 265683
rect 327914 265671 327920 265723
rect 327952 265671 327958 265723
rect 328010 265711 328016 265723
rect 339088 265711 339094 265723
rect 328010 265683 339094 265711
rect 328010 265671 328016 265683
rect 339088 265671 339094 265683
rect 339146 265671 339152 265723
rect 350704 265671 350710 265723
rect 350762 265711 350768 265723
rect 368368 265711 368374 265723
rect 350762 265683 368374 265711
rect 350762 265671 350768 265683
rect 368368 265671 368374 265683
rect 368426 265671 368432 265723
rect 368560 265671 368566 265723
rect 368618 265711 368624 265723
rect 370672 265711 370678 265723
rect 368618 265683 370678 265711
rect 368618 265671 368624 265683
rect 370672 265671 370678 265683
rect 370730 265671 370736 265723
rect 372898 265683 397694 265711
rect 306736 265597 306742 265649
rect 306794 265637 306800 265649
rect 372898 265637 372926 265683
rect 306794 265609 372926 265637
rect 306794 265597 306800 265609
rect 377200 265597 377206 265649
rect 377258 265637 377264 265649
rect 378928 265637 378934 265649
rect 377258 265609 378934 265637
rect 377258 265597 377264 265609
rect 378928 265597 378934 265609
rect 378986 265597 378992 265649
rect 379024 265597 379030 265649
rect 379082 265637 379088 265649
rect 397552 265637 397558 265649
rect 379082 265609 397558 265637
rect 379082 265597 379088 265609
rect 397552 265597 397558 265609
rect 397610 265597 397616 265649
rect 397666 265637 397694 265683
rect 398800 265671 398806 265723
rect 398858 265711 398864 265723
rect 419248 265711 419254 265723
rect 398858 265683 419254 265711
rect 398858 265671 398864 265683
rect 419248 265671 419254 265683
rect 419306 265671 419312 265723
rect 419344 265671 419350 265723
rect 419402 265711 419408 265723
rect 547600 265711 547606 265723
rect 419402 265683 547606 265711
rect 419402 265671 419408 265683
rect 547600 265671 547606 265683
rect 547658 265671 547664 265723
rect 492880 265637 492886 265649
rect 397666 265609 492886 265637
rect 492880 265597 492886 265609
rect 492938 265597 492944 265649
rect 307312 265523 307318 265575
rect 307370 265563 307376 265575
rect 499888 265563 499894 265575
rect 307370 265535 499894 265563
rect 307370 265523 307376 265535
rect 499888 265523 499894 265535
rect 499946 265523 499952 265575
rect 309328 265449 309334 265501
rect 309386 265489 309392 265501
rect 309386 265461 378878 265489
rect 309386 265449 309392 265461
rect 309904 265375 309910 265427
rect 309962 265415 309968 265427
rect 309962 265387 378302 265415
rect 309962 265375 309968 265387
rect 311632 265301 311638 265353
rect 311690 265341 311696 265353
rect 311690 265313 369662 265341
rect 311690 265301 311696 265313
rect 221680 265227 221686 265279
rect 221738 265267 221744 265279
rect 273136 265267 273142 265279
rect 221738 265239 273142 265267
rect 221738 265227 221744 265239
rect 273136 265227 273142 265239
rect 273194 265227 273200 265279
rect 313264 265227 313270 265279
rect 313322 265267 313328 265279
rect 319312 265267 319318 265279
rect 313322 265239 319318 265267
rect 313322 265227 313328 265239
rect 319312 265227 319318 265239
rect 319370 265227 319376 265279
rect 369328 265267 369334 265279
rect 319522 265239 369334 265267
rect 255664 265153 255670 265205
rect 255722 265193 255728 265205
rect 267856 265193 267862 265205
rect 255722 265165 267862 265193
rect 255722 265153 255728 265165
rect 267856 265153 267862 265165
rect 267914 265153 267920 265205
rect 276496 265153 276502 265205
rect 276554 265193 276560 265205
rect 308080 265193 308086 265205
rect 276554 265165 308086 265193
rect 276554 265153 276560 265165
rect 308080 265153 308086 265165
rect 308138 265153 308144 265205
rect 219568 265079 219574 265131
rect 219626 265119 219632 265131
rect 219626 265091 312926 265119
rect 219626 265079 219632 265091
rect 201424 265005 201430 265057
rect 201482 265045 201488 265057
rect 311920 265045 311926 265057
rect 201482 265017 311926 265045
rect 201482 265005 201488 265017
rect 311920 265005 311926 265017
rect 311978 265005 311984 265057
rect 312898 265045 312926 265091
rect 319408 265079 319414 265131
rect 319466 265119 319472 265131
rect 319522 265119 319550 265239
rect 369328 265227 369334 265239
rect 369386 265227 369392 265279
rect 369634 265267 369662 265313
rect 369712 265301 369718 265353
rect 369770 265341 369776 265353
rect 378160 265341 378166 265353
rect 369770 265313 378166 265341
rect 369770 265301 369776 265313
rect 378160 265301 378166 265313
rect 378218 265301 378224 265353
rect 378274 265341 378302 265387
rect 378352 265375 378358 265427
rect 378410 265415 378416 265427
rect 378736 265415 378742 265427
rect 378410 265387 378742 265415
rect 378410 265375 378416 265387
rect 378736 265375 378742 265387
rect 378794 265375 378800 265427
rect 378850 265415 378878 265461
rect 378928 265449 378934 265501
rect 378986 265489 378992 265501
rect 378986 265461 379838 265489
rect 378986 265449 378992 265461
rect 379696 265415 379702 265427
rect 378850 265387 379702 265415
rect 379696 265375 379702 265387
rect 379754 265375 379760 265427
rect 379600 265341 379606 265353
rect 378274 265313 379606 265341
rect 379600 265301 379606 265313
rect 379658 265301 379664 265353
rect 379810 265341 379838 265461
rect 379888 265449 379894 265501
rect 379946 265489 379952 265501
rect 392944 265489 392950 265501
rect 379946 265461 392950 265489
rect 379946 265449 379952 265461
rect 392944 265449 392950 265461
rect 393002 265449 393008 265501
rect 395728 265449 395734 265501
rect 395786 265489 395792 265501
rect 407056 265489 407062 265501
rect 395786 265461 407062 265489
rect 395786 265449 395792 265461
rect 407056 265449 407062 265461
rect 407114 265449 407120 265501
rect 408208 265449 408214 265501
rect 408266 265489 408272 265501
rect 412816 265489 412822 265501
rect 408266 265461 412822 265489
rect 408266 265449 408272 265461
rect 412816 265449 412822 265461
rect 412874 265449 412880 265501
rect 514288 265489 514294 265501
rect 418978 265461 514294 265489
rect 379984 265375 379990 265427
rect 380042 265415 380048 265427
rect 418978 265415 419006 265461
rect 514288 265449 514294 265461
rect 514346 265449 514352 265501
rect 380042 265387 419006 265415
rect 380042 265375 380048 265387
rect 419056 265375 419062 265427
rect 419114 265415 419120 265427
rect 521392 265415 521398 265427
rect 419114 265387 521398 265415
rect 419114 265375 419120 265387
rect 521392 265375 521398 265387
rect 521450 265375 521456 265427
rect 379810 265313 380126 265341
rect 379408 265267 379414 265279
rect 369634 265239 379414 265267
rect 379408 265227 379414 265239
rect 379466 265227 379472 265279
rect 379984 265227 379990 265279
rect 380042 265227 380048 265279
rect 380098 265267 380126 265313
rect 380176 265301 380182 265353
rect 380234 265341 380240 265353
rect 380234 265313 388766 265341
rect 380234 265301 380240 265313
rect 388738 265267 388766 265313
rect 388816 265301 388822 265353
rect 388874 265341 388880 265353
rect 389584 265341 389590 265353
rect 388874 265313 389590 265341
rect 388874 265301 388880 265313
rect 389584 265301 389590 265313
rect 389642 265301 389648 265353
rect 389776 265301 389782 265353
rect 389834 265341 389840 265353
rect 395728 265341 395734 265353
rect 389834 265313 395734 265341
rect 389834 265301 389840 265313
rect 395728 265301 395734 265313
rect 395786 265301 395792 265353
rect 395920 265301 395926 265353
rect 395978 265341 395984 265353
rect 535600 265341 535606 265353
rect 395978 265313 535606 265341
rect 395978 265301 395984 265313
rect 535600 265301 535606 265313
rect 535658 265301 535664 265353
rect 419056 265267 419062 265279
rect 380098 265239 381278 265267
rect 388738 265239 419062 265267
rect 320272 265153 320278 265205
rect 320330 265193 320336 265205
rect 327280 265193 327286 265205
rect 320330 265165 327286 265193
rect 320330 265153 320336 265165
rect 327280 265153 327286 265165
rect 327338 265153 327344 265205
rect 329392 265153 329398 265205
rect 329450 265193 329456 265205
rect 375952 265193 375958 265205
rect 329450 265165 375958 265193
rect 329450 265153 329456 265165
rect 375952 265153 375958 265165
rect 376010 265153 376016 265205
rect 376048 265153 376054 265205
rect 376106 265193 376112 265205
rect 379504 265193 379510 265205
rect 376106 265165 379510 265193
rect 376106 265153 376112 265165
rect 379504 265153 379510 265165
rect 379562 265153 379568 265205
rect 380002 265193 380030 265227
rect 381136 265193 381142 265205
rect 380002 265165 381142 265193
rect 381136 265153 381142 265165
rect 381194 265153 381200 265205
rect 381250 265193 381278 265239
rect 419056 265227 419062 265239
rect 419114 265227 419120 265279
rect 419152 265227 419158 265279
rect 419210 265267 419216 265279
rect 546352 265267 546358 265279
rect 419210 265239 546358 265267
rect 419210 265227 419216 265239
rect 546352 265227 546358 265239
rect 546410 265227 546416 265279
rect 388528 265193 388534 265205
rect 381250 265165 388534 265193
rect 388528 265153 388534 265165
rect 388586 265153 388592 265205
rect 389008 265153 389014 265205
rect 389066 265193 389072 265205
rect 390448 265193 390454 265205
rect 389066 265165 390454 265193
rect 389066 265153 389072 265165
rect 390448 265153 390454 265165
rect 390506 265153 390512 265205
rect 608176 265193 608182 265205
rect 399106 265165 608182 265193
rect 328432 265119 328438 265131
rect 319466 265091 319550 265119
rect 319618 265091 328438 265119
rect 319466 265079 319472 265091
rect 319618 265045 319646 265091
rect 328432 265079 328438 265091
rect 328490 265079 328496 265131
rect 367120 265119 367126 265131
rect 332626 265091 367126 265119
rect 312418 265017 312830 265045
rect 312898 265017 319646 265045
rect 267760 264931 267766 264983
rect 267818 264971 267824 264983
rect 312418 264971 312446 265017
rect 267818 264943 312446 264971
rect 267818 264931 267824 264943
rect 312688 264931 312694 264983
rect 312746 264931 312752 264983
rect 312802 264971 312830 265017
rect 320560 265005 320566 265057
rect 320618 265045 320624 265057
rect 326224 265045 326230 265057
rect 320618 265017 326230 265045
rect 320618 265005 320624 265017
rect 326224 265005 326230 265017
rect 326282 265005 326288 265057
rect 332626 265045 332654 265091
rect 367120 265079 367126 265091
rect 367178 265079 367184 265131
rect 369058 265091 369278 265119
rect 369058 265045 369086 265091
rect 326530 265017 332654 265045
rect 367138 265017 369086 265045
rect 369250 265045 369278 265091
rect 369328 265079 369334 265131
rect 369386 265119 369392 265131
rect 390256 265119 390262 265131
rect 369386 265091 390262 265119
rect 369386 265079 369392 265091
rect 390256 265079 390262 265091
rect 390314 265079 390320 265131
rect 399106 265119 399134 265165
rect 608176 265153 608182 265165
rect 608234 265153 608240 265205
rect 390370 265091 399134 265119
rect 369250 265017 369374 265045
rect 325072 264971 325078 264983
rect 312802 264943 325078 264971
rect 325072 264931 325078 264943
rect 325130 264931 325136 264983
rect 325186 264943 325502 264971
rect 210640 264857 210646 264909
rect 210698 264897 210704 264909
rect 212464 264897 212470 264909
rect 210698 264869 212470 264897
rect 210698 264857 210704 264869
rect 212464 264857 212470 264869
rect 212522 264857 212528 264909
rect 312706 264897 312734 264931
rect 325186 264897 325214 264943
rect 312706 264869 325214 264897
rect 325474 264897 325502 264943
rect 325744 264931 325750 264983
rect 325802 264971 325808 264983
rect 326530 264971 326558 265017
rect 325802 264943 326558 264971
rect 325802 264931 325808 264943
rect 326704 264931 326710 264983
rect 326762 264931 326768 264983
rect 327280 264931 327286 264983
rect 327338 264931 327344 264983
rect 329392 264931 329398 264983
rect 329450 264931 329456 264983
rect 329488 264931 329494 264983
rect 329546 264971 329552 264983
rect 341008 264971 341014 264983
rect 329546 264943 341014 264971
rect 329546 264931 329552 264943
rect 341008 264931 341014 264943
rect 341066 264931 341072 264983
rect 326722 264897 326750 264931
rect 325474 264869 326750 264897
rect 327298 264897 327326 264931
rect 329410 264897 329438 264931
rect 327298 264869 329438 264897
rect 349840 264857 349846 264909
rect 349898 264897 349904 264909
rect 367138 264897 367166 265017
rect 369346 264971 369374 265017
rect 376432 265005 376438 265057
rect 376490 265045 376496 265057
rect 390370 265045 390398 265091
rect 399376 265079 399382 265131
rect 399434 265119 399440 265131
rect 419152 265119 419158 265131
rect 399434 265091 419158 265119
rect 399434 265079 399440 265091
rect 419152 265079 419158 265091
rect 419210 265079 419216 265131
rect 419248 265079 419254 265131
rect 419306 265119 419312 265131
rect 615376 265119 615382 265131
rect 419306 265091 615382 265119
rect 419306 265079 419312 265091
rect 615376 265079 615382 265091
rect 615434 265079 615440 265131
rect 376490 265017 390398 265045
rect 376490 265005 376496 265017
rect 390448 265005 390454 265057
rect 390506 265045 390512 265057
rect 406960 265045 406966 265057
rect 390506 265017 406966 265045
rect 390506 265005 390512 265017
rect 406960 265005 406966 265017
rect 407018 265005 407024 265057
rect 407056 265005 407062 265057
rect 407114 265045 407120 265057
rect 412720 265045 412726 265057
rect 407114 265017 412726 265045
rect 407114 265005 407120 265017
rect 412720 265005 412726 265017
rect 412778 265005 412784 265057
rect 379024 264971 379030 264983
rect 369346 264943 379030 264971
rect 379024 264931 379030 264943
rect 379082 264931 379088 264983
rect 379120 264931 379126 264983
rect 379178 264971 379184 264983
rect 389776 264971 389782 264983
rect 379178 264943 389782 264971
rect 379178 264931 379184 264943
rect 389776 264931 389782 264943
rect 389834 264931 389840 264983
rect 390256 264931 390262 264983
rect 390314 264971 390320 264983
rect 399376 264971 399382 264983
rect 390314 264943 399382 264971
rect 390314 264931 390320 264943
rect 399376 264931 399382 264943
rect 399434 264931 399440 264983
rect 399856 264931 399862 264983
rect 399914 264971 399920 264983
rect 412624 264971 412630 264983
rect 399914 264943 412630 264971
rect 399914 264931 399920 264943
rect 412624 264931 412630 264943
rect 412682 264931 412688 264983
rect 349898 264869 367166 264897
rect 349898 264857 349904 264869
rect 369040 264857 369046 264909
rect 369098 264897 369104 264909
rect 369712 264897 369718 264909
rect 369098 264869 369718 264897
rect 369098 264857 369104 264869
rect 369712 264857 369718 264869
rect 369770 264857 369776 264909
rect 371536 264857 371542 264909
rect 371594 264897 371600 264909
rect 388048 264897 388054 264909
rect 371594 264869 388054 264897
rect 371594 264857 371600 264869
rect 388048 264857 388054 264869
rect 388106 264857 388112 264909
rect 633616 262159 633622 262171
rect 627874 262131 633622 262159
rect 625840 262045 625846 262097
rect 625898 262085 625904 262097
rect 627874 262085 627902 262131
rect 633616 262119 633622 262131
rect 633674 262119 633680 262171
rect 625898 262057 627902 262085
rect 625898 262045 625904 262057
rect 642256 260491 642262 260543
rect 642314 260531 642320 260543
rect 645712 260531 645718 260543
rect 642314 260503 645718 260531
rect 642314 260491 642320 260503
rect 645712 260491 645718 260503
rect 645770 260491 645776 260543
rect 42544 259677 42550 259729
rect 42602 259717 42608 259729
rect 50512 259717 50518 259729
rect 42602 259689 50518 259717
rect 42602 259677 42608 259689
rect 50512 259677 50518 259689
rect 50570 259677 50576 259729
rect 83536 259307 83542 259359
rect 83594 259347 83600 259359
rect 83594 259319 92222 259347
rect 83594 259307 83600 259319
rect 92194 259199 92222 259319
rect 95056 259199 95062 259211
rect 92194 259171 95062 259199
rect 95056 259159 95062 259171
rect 95114 259159 95120 259211
rect 42640 258937 42646 258989
rect 42698 258977 42704 258989
rect 53392 258977 53398 258989
rect 42698 258949 53398 258977
rect 42698 258937 42704 258949
rect 53392 258937 53398 258949
rect 53450 258937 53456 258989
rect 42544 258197 42550 258249
rect 42602 258237 42608 258249
rect 47440 258237 47446 258249
rect 42602 258209 47446 258237
rect 42602 258197 42608 258209
rect 47440 258197 47446 258209
rect 47498 258197 47504 258249
rect 42256 257753 42262 257805
rect 42314 257793 42320 257805
rect 43120 257793 43126 257805
rect 42314 257765 43126 257793
rect 42314 257753 42320 257765
rect 43120 257753 43126 257765
rect 43178 257753 43184 257805
rect 616336 257753 616342 257805
rect 616394 257793 616400 257805
rect 625840 257793 625846 257805
rect 616394 257765 625846 257793
rect 616394 257753 616400 257765
rect 625840 257753 625846 257765
rect 625898 257753 625904 257805
rect 42544 257161 42550 257213
rect 42602 257201 42608 257213
rect 43216 257201 43222 257213
rect 42602 257173 43222 257201
rect 42602 257161 42608 257173
rect 43216 257161 43222 257173
rect 43274 257161 43280 257213
rect 639280 256347 639286 256399
rect 639338 256387 639344 256399
rect 677008 256387 677014 256399
rect 639338 256359 677014 256387
rect 639338 256347 639344 256359
rect 677008 256347 677014 256359
rect 677066 256347 677072 256399
rect 67600 253387 67606 253439
rect 67658 253427 67664 253439
rect 74896 253427 74902 253439
rect 67658 253399 74902 253427
rect 67658 253387 67664 253399
rect 74896 253387 74902 253399
rect 74954 253387 74960 253439
rect 675184 250945 675190 250997
rect 675242 250985 675248 250997
rect 675376 250985 675382 250997
rect 675242 250957 675382 250985
rect 675242 250945 675248 250957
rect 675376 250945 675382 250957
rect 675434 250945 675440 250997
rect 607696 250575 607702 250627
rect 607754 250615 607760 250627
rect 616336 250615 616342 250627
rect 607754 250587 616342 250615
rect 607754 250575 607760 250587
rect 616336 250575 616342 250587
rect 616394 250575 616400 250627
rect 636496 250575 636502 250627
rect 636554 250615 636560 250627
rect 642256 250615 642262 250627
rect 636554 250587 642262 250615
rect 636554 250575 636560 250587
rect 642256 250575 642262 250587
rect 642314 250575 642320 250627
rect 674512 250353 674518 250405
rect 674570 250393 674576 250405
rect 675184 250393 675190 250405
rect 674570 250365 675190 250393
rect 674570 250353 674576 250365
rect 675184 250353 675190 250365
rect 675242 250353 675248 250405
rect 74896 249317 74902 249369
rect 74954 249357 74960 249369
rect 90640 249357 90646 249369
rect 74954 249329 90646 249357
rect 74954 249317 74960 249329
rect 90640 249317 90646 249329
rect 90698 249317 90704 249369
rect 56176 249243 56182 249295
rect 56234 249283 56240 249295
rect 205552 249283 205558 249295
rect 56234 249255 205558 249283
rect 56234 249243 56240 249255
rect 205552 249243 205558 249255
rect 205610 249243 205616 249295
rect 53776 249169 53782 249221
rect 53834 249209 53840 249221
rect 210736 249209 210742 249221
rect 53834 249181 210742 249209
rect 53834 249169 53840 249181
rect 210736 249169 210742 249181
rect 210794 249169 210800 249221
rect 45040 249095 45046 249147
rect 45098 249135 45104 249147
rect 206896 249135 206902 249147
rect 45098 249107 206902 249135
rect 45098 249095 45104 249107
rect 206896 249095 206902 249107
rect 206954 249095 206960 249147
rect 200080 247689 200086 247741
rect 200138 247729 200144 247741
rect 200138 247701 204446 247729
rect 200138 247689 200144 247701
rect 204418 247655 204446 247701
rect 627856 247689 627862 247741
rect 627914 247729 627920 247741
rect 636496 247729 636502 247741
rect 627914 247701 636502 247729
rect 627914 247689 627920 247701
rect 636496 247689 636502 247701
rect 636554 247689 636560 247741
rect 205264 247655 205270 247667
rect 204418 247627 205270 247655
rect 205264 247615 205270 247627
rect 205322 247615 205328 247667
rect 126544 247319 126550 247371
rect 126602 247359 126608 247371
rect 126602 247331 409022 247359
rect 126602 247319 126608 247331
rect 129520 247245 129526 247297
rect 129578 247285 129584 247297
rect 129578 247257 407006 247285
rect 129578 247245 129584 247257
rect 132304 247171 132310 247223
rect 132362 247211 132368 247223
rect 132362 247183 401918 247211
rect 132362 247171 132368 247183
rect 135184 247097 135190 247149
rect 135242 247137 135248 247149
rect 135242 247109 401822 247137
rect 135242 247097 135248 247109
rect 140944 247023 140950 247075
rect 141002 247063 141008 247075
rect 141002 247035 401726 247063
rect 141002 247023 141008 247035
rect 143920 246949 143926 247001
rect 143978 246989 143984 247001
rect 143978 246961 398270 246989
rect 143978 246949 143984 246961
rect 146704 246875 146710 246927
rect 146762 246915 146768 246927
rect 146762 246887 397886 246915
rect 146762 246875 146768 246887
rect 80464 246801 80470 246853
rect 80522 246841 80528 246853
rect 86512 246841 86518 246853
rect 80522 246813 86518 246841
rect 80522 246801 80528 246813
rect 86512 246801 86518 246813
rect 86570 246801 86576 246853
rect 171280 246801 171286 246853
rect 171338 246841 171344 246853
rect 181360 246841 181366 246853
rect 171338 246813 181366 246841
rect 171338 246801 171344 246813
rect 181360 246801 181366 246813
rect 181418 246801 181424 246853
rect 211696 246801 211702 246853
rect 211754 246841 211760 246853
rect 211754 246813 227966 246841
rect 211754 246801 211760 246813
rect 227938 246779 227966 246813
rect 231778 246813 248222 246841
rect 63280 246727 63286 246779
rect 63338 246767 63344 246779
rect 204592 246767 204598 246779
rect 63338 246739 204598 246767
rect 63338 246727 63344 246739
rect 204592 246727 204598 246739
rect 204650 246727 204656 246779
rect 211888 246727 211894 246779
rect 211946 246767 211952 246779
rect 227440 246767 227446 246779
rect 211946 246739 227446 246767
rect 211946 246727 211952 246739
rect 227440 246727 227446 246739
rect 227498 246727 227504 246779
rect 227920 246727 227926 246779
rect 227978 246727 227984 246779
rect 47632 246653 47638 246705
rect 47690 246693 47696 246705
rect 65008 246693 65014 246705
rect 47690 246665 65014 246693
rect 47690 246653 47696 246665
rect 65008 246653 65014 246665
rect 65066 246653 65072 246705
rect 65200 246653 65206 246705
rect 65258 246693 65264 246705
rect 171280 246693 171286 246705
rect 65258 246665 171286 246693
rect 65258 246653 65264 246665
rect 171280 246653 171286 246665
rect 171338 246653 171344 246705
rect 181360 246653 181366 246705
rect 181418 246693 181424 246705
rect 210928 246693 210934 246705
rect 181418 246665 210934 246693
rect 181418 246653 181424 246665
rect 210928 246653 210934 246665
rect 210986 246653 210992 246705
rect 212080 246653 212086 246705
rect 212138 246693 212144 246705
rect 227056 246693 227062 246705
rect 212138 246665 227062 246693
rect 212138 246653 212144 246665
rect 227056 246653 227062 246665
rect 227114 246653 227120 246705
rect 227824 246653 227830 246705
rect 227882 246693 227888 246705
rect 231778 246693 231806 246813
rect 248194 246779 248222 246813
rect 248290 246813 280382 246841
rect 248290 246779 248318 246813
rect 231856 246727 231862 246779
rect 231914 246767 231920 246779
rect 247888 246767 247894 246779
rect 231914 246739 247894 246767
rect 231914 246727 231920 246739
rect 247888 246727 247894 246739
rect 247946 246727 247952 246779
rect 248176 246727 248182 246779
rect 248234 246727 248240 246779
rect 248272 246727 248278 246779
rect 248330 246727 248336 246779
rect 251920 246727 251926 246779
rect 251978 246767 251984 246779
rect 276880 246767 276886 246779
rect 251978 246739 276886 246767
rect 251978 246727 251984 246739
rect 276880 246727 276886 246739
rect 276938 246727 276944 246779
rect 280354 246767 280382 246813
rect 281218 246813 288446 246841
rect 280816 246767 280822 246779
rect 280354 246739 280822 246767
rect 280816 246727 280822 246739
rect 280874 246727 280880 246779
rect 280912 246727 280918 246779
rect 280970 246767 280976 246779
rect 281218 246767 281246 246813
rect 280970 246739 281246 246767
rect 280970 246727 280976 246739
rect 284944 246727 284950 246779
rect 285002 246767 285008 246779
rect 288304 246767 288310 246779
rect 285002 246739 288310 246767
rect 285002 246727 285008 246739
rect 288304 246727 288310 246739
rect 288362 246727 288368 246779
rect 288418 246767 288446 246813
rect 292258 246813 309374 246841
rect 292258 246779 292286 246813
rect 309346 246779 309374 246813
rect 312130 246813 397790 246841
rect 288688 246767 288694 246779
rect 288418 246739 288694 246767
rect 288688 246727 288694 246739
rect 288746 246727 288752 246779
rect 292240 246727 292246 246779
rect 292298 246727 292304 246779
rect 292354 246739 294686 246767
rect 227882 246665 231806 246693
rect 227882 246653 227888 246665
rect 232144 246653 232150 246705
rect 232202 246693 232208 246705
rect 232202 246665 248414 246693
rect 232202 246653 232208 246665
rect 56080 246579 56086 246631
rect 56138 246619 56144 246631
rect 180976 246619 180982 246631
rect 56138 246591 180982 246619
rect 56138 246579 56144 246591
rect 180976 246579 180982 246591
rect 181034 246579 181040 246631
rect 181264 246579 181270 246631
rect 181322 246619 181328 246631
rect 204784 246619 204790 246631
rect 181322 246591 204790 246619
rect 181322 246579 181328 246591
rect 204784 246579 204790 246591
rect 204842 246579 204848 246631
rect 211792 246579 211798 246631
rect 211850 246619 211856 246631
rect 226480 246619 226486 246631
rect 211850 246591 226486 246619
rect 211850 246579 211856 246591
rect 226480 246579 226486 246591
rect 226538 246579 226544 246631
rect 226960 246579 226966 246631
rect 227018 246619 227024 246631
rect 227018 246591 228254 246619
rect 227018 246579 227024 246591
rect 53488 246505 53494 246557
rect 53546 246545 53552 246557
rect 204496 246545 204502 246557
rect 53546 246517 204502 246545
rect 53546 246505 53552 246517
rect 204496 246505 204502 246517
rect 204554 246505 204560 246557
rect 225328 246505 225334 246557
rect 225386 246545 225392 246557
rect 227824 246545 227830 246557
rect 225386 246517 227830 246545
rect 225386 246505 225392 246517
rect 227824 246505 227830 246517
rect 227882 246505 227888 246557
rect 228226 246545 228254 246591
rect 231376 246579 231382 246631
rect 231434 246619 231440 246631
rect 248176 246619 248182 246631
rect 231434 246591 248182 246619
rect 231434 246579 231440 246591
rect 248176 246579 248182 246591
rect 248234 246579 248240 246631
rect 247312 246545 247318 246557
rect 227938 246517 228158 246545
rect 228226 246517 247318 246545
rect 53200 246431 53206 246483
rect 53258 246471 53264 246483
rect 204688 246471 204694 246483
rect 53258 246443 204694 246471
rect 53258 246431 53264 246443
rect 204688 246431 204694 246443
rect 204746 246431 204752 246483
rect 211984 246431 211990 246483
rect 212042 246471 212048 246483
rect 227938 246471 227966 246517
rect 212042 246443 227966 246471
rect 228130 246471 228158 246517
rect 247312 246505 247318 246517
rect 247370 246505 247376 246557
rect 248386 246545 248414 246665
rect 248578 246665 281150 246693
rect 248578 246545 248606 246665
rect 252112 246579 252118 246631
rect 252170 246619 252176 246631
rect 281122 246619 281150 246665
rect 281296 246653 281302 246705
rect 281354 246693 281360 246705
rect 287536 246693 287542 246705
rect 281354 246665 287542 246693
rect 281354 246653 281360 246665
rect 287536 246653 287542 246665
rect 287594 246653 287600 246705
rect 292354 246693 292382 246739
rect 288322 246665 292382 246693
rect 294658 246693 294686 246739
rect 295696 246727 295702 246779
rect 295754 246767 295760 246779
rect 309232 246767 309238 246779
rect 295754 246739 309238 246767
rect 295754 246727 295760 246739
rect 309232 246727 309238 246739
rect 309290 246727 309296 246779
rect 309328 246727 309334 246779
rect 309386 246727 309392 246779
rect 309424 246727 309430 246779
rect 309482 246767 309488 246779
rect 312130 246767 312158 246813
rect 397762 246779 397790 246813
rect 313744 246767 313750 246779
rect 309482 246739 312158 246767
rect 312226 246739 313750 246767
rect 309482 246727 309488 246739
rect 311728 246693 311734 246705
rect 294658 246665 311734 246693
rect 288322 246619 288350 246665
rect 311728 246653 311734 246665
rect 311786 246653 311792 246705
rect 252170 246591 281054 246619
rect 281122 246591 288350 246619
rect 252170 246579 252176 246591
rect 276976 246545 276982 246557
rect 248386 246517 248606 246545
rect 248722 246517 276982 246545
rect 248722 246471 248750 246517
rect 276976 246505 276982 246517
rect 277034 246505 277040 246557
rect 280912 246545 280918 246557
rect 277186 246517 280918 246545
rect 228130 246443 248750 246471
rect 212042 246431 212048 246443
rect 249040 246431 249046 246483
rect 249098 246471 249104 246483
rect 259120 246471 259126 246483
rect 249098 246443 259126 246471
rect 249098 246431 249104 246443
rect 259120 246431 259126 246443
rect 259178 246431 259184 246483
rect 268816 246431 268822 246483
rect 268874 246471 268880 246483
rect 274096 246471 274102 246483
rect 268874 246443 274102 246471
rect 268874 246431 268880 246443
rect 274096 246431 274102 246443
rect 274154 246431 274160 246483
rect 80464 246357 80470 246409
rect 80522 246397 80528 246409
rect 145840 246397 145846 246409
rect 80522 246369 145846 246397
rect 80522 246357 80528 246369
rect 145840 246357 145846 246369
rect 145898 246357 145904 246409
rect 161296 246357 161302 246409
rect 161354 246397 161360 246409
rect 161354 246369 202814 246397
rect 161354 246357 161360 246369
rect 44752 246283 44758 246335
rect 44810 246323 44816 246335
rect 160912 246323 160918 246335
rect 44810 246295 160918 246323
rect 44810 246283 44816 246295
rect 160912 246283 160918 246295
rect 160970 246283 160976 246335
rect 165520 246283 165526 246335
rect 165578 246323 165584 246335
rect 199600 246323 199606 246335
rect 165578 246295 199606 246323
rect 165578 246283 165584 246295
rect 199600 246283 199606 246295
rect 199658 246283 199664 246335
rect 202786 246323 202814 246369
rect 212176 246357 212182 246409
rect 212234 246397 212240 246409
rect 230896 246397 230902 246409
rect 212234 246369 230902 246397
rect 212234 246357 212240 246369
rect 230896 246357 230902 246369
rect 230954 246357 230960 246409
rect 247792 246357 247798 246409
rect 247850 246397 247856 246409
rect 260752 246397 260758 246409
rect 247850 246369 260758 246397
rect 247850 246357 247856 246369
rect 260752 246357 260758 246369
rect 260810 246357 260816 246409
rect 268048 246397 268054 246409
rect 260866 246369 268054 246397
rect 214192 246323 214198 246335
rect 202786 246295 214198 246323
rect 214192 246283 214198 246295
rect 214250 246283 214256 246335
rect 227920 246283 227926 246335
rect 227978 246323 227984 246335
rect 260866 246323 260894 246369
rect 268048 246357 268054 246369
rect 268106 246357 268112 246409
rect 268624 246357 268630 246409
rect 268682 246397 268688 246409
rect 277186 246397 277214 246517
rect 280912 246505 280918 246517
rect 280970 246505 280976 246557
rect 281026 246545 281054 246591
rect 288400 246579 288406 246631
rect 288458 246619 288464 246631
rect 292240 246619 292246 246631
rect 288458 246591 292246 246619
rect 288458 246579 288464 246591
rect 292240 246579 292246 246591
rect 292298 246579 292304 246631
rect 312226 246619 312254 246739
rect 313744 246727 313750 246739
rect 313802 246727 313808 246779
rect 314032 246727 314038 246779
rect 314090 246767 314096 246779
rect 397264 246767 397270 246779
rect 314090 246739 397270 246767
rect 314090 246727 314096 246739
rect 397264 246727 397270 246739
rect 397322 246727 397328 246779
rect 397744 246727 397750 246779
rect 397802 246727 397808 246779
rect 313936 246653 313942 246705
rect 313994 246693 314000 246705
rect 397360 246693 397366 246705
rect 313994 246665 397366 246693
rect 313994 246653 314000 246665
rect 397360 246653 397366 246665
rect 397418 246653 397424 246705
rect 294658 246591 312254 246619
rect 294658 246545 294686 246591
rect 312304 246579 312310 246631
rect 312362 246619 312368 246631
rect 312362 246591 313502 246619
rect 312362 246579 312368 246591
rect 281026 246517 294686 246545
rect 294832 246505 294838 246557
rect 294890 246545 294896 246557
rect 294890 246517 311294 246545
rect 294890 246505 294896 246517
rect 280816 246431 280822 246483
rect 280874 246471 280880 246483
rect 280874 246443 287966 246471
rect 280874 246431 280880 246443
rect 268682 246369 277214 246397
rect 268682 246357 268688 246369
rect 277360 246357 277366 246409
rect 277418 246397 277424 246409
rect 277418 246369 287678 246397
rect 277418 246357 277424 246369
rect 227978 246295 260894 246323
rect 227978 246283 227984 246295
rect 268240 246283 268246 246335
rect 268298 246323 268304 246335
rect 280816 246323 280822 246335
rect 268298 246295 280822 246323
rect 268298 246283 268304 246295
rect 280816 246283 280822 246295
rect 280874 246283 280880 246335
rect 44560 246209 44566 246261
rect 44618 246249 44624 246261
rect 161008 246249 161014 246261
rect 44618 246221 161014 246249
rect 44618 246209 44624 246221
rect 161008 246209 161014 246221
rect 161066 246209 161072 246261
rect 163696 246209 163702 246261
rect 163754 246249 163760 246261
rect 198736 246249 198742 246261
rect 163754 246221 198742 246249
rect 163754 246209 163760 246221
rect 198736 246209 198742 246221
rect 198794 246209 198800 246261
rect 210256 246209 210262 246261
rect 210314 246249 210320 246261
rect 229264 246249 229270 246261
rect 210314 246221 229270 246249
rect 210314 246209 210320 246221
rect 229264 246209 229270 246221
rect 229322 246209 229328 246261
rect 230896 246209 230902 246261
rect 230954 246249 230960 246261
rect 260848 246249 260854 246261
rect 230954 246221 260854 246249
rect 230954 246209 230960 246221
rect 260848 246209 260854 246221
rect 260906 246209 260912 246261
rect 268528 246209 268534 246261
rect 268586 246249 268592 246261
rect 287650 246249 287678 246369
rect 287938 246323 287966 246443
rect 289168 246431 289174 246483
rect 289226 246471 289232 246483
rect 311152 246471 311158 246483
rect 289226 246443 311158 246471
rect 289226 246431 289232 246443
rect 311152 246431 311158 246443
rect 311210 246431 311216 246483
rect 311266 246471 311294 246517
rect 311728 246505 311734 246557
rect 311786 246545 311792 246557
rect 313474 246545 313502 246591
rect 313744 246579 313750 246631
rect 313802 246619 313808 246631
rect 397858 246619 397886 246887
rect 398242 246779 398270 246961
rect 398224 246727 398230 246779
rect 398282 246727 398288 246779
rect 401698 246693 401726 247035
rect 401794 246915 401822 247109
rect 401890 247063 401918 247183
rect 401890 247035 403262 247063
rect 401794 246887 403070 246915
rect 403042 246779 403070 246887
rect 403024 246727 403030 246779
rect 403082 246727 403088 246779
rect 403234 246767 403262 247035
rect 406978 246779 407006 247257
rect 408994 246779 409022 247331
rect 674320 247245 674326 247297
rect 674378 247285 674384 247297
rect 675184 247285 675190 247297
rect 674378 247257 675190 247285
rect 674378 247245 674384 247257
rect 675184 247245 675190 247257
rect 675242 247245 675248 247297
rect 674800 247171 674806 247223
rect 674858 247211 674864 247223
rect 675088 247211 675094 247223
rect 674858 247183 675094 247211
rect 674858 247171 674864 247183
rect 675088 247171 675094 247183
rect 675146 247171 675152 247223
rect 406096 246767 406102 246779
rect 403234 246739 406102 246767
rect 406096 246727 406102 246739
rect 406154 246727 406160 246779
rect 406960 246727 406966 246779
rect 407018 246727 407024 246779
rect 408976 246727 408982 246779
rect 409034 246727 409040 246779
rect 408304 246693 408310 246705
rect 401698 246665 408310 246693
rect 408304 246653 408310 246665
rect 408362 246653 408368 246705
rect 406576 246619 406582 246631
rect 313802 246591 397790 246619
rect 397858 246591 406582 246619
rect 313802 246579 313808 246591
rect 328912 246545 328918 246557
rect 311786 246517 313406 246545
rect 313474 246517 328918 246545
rect 311786 246505 311792 246517
rect 311266 246443 313310 246471
rect 313282 246409 313310 246443
rect 288688 246357 288694 246409
rect 288746 246397 288752 246409
rect 307504 246397 307510 246409
rect 288746 246369 307510 246397
rect 288746 246357 288752 246369
rect 307504 246357 307510 246369
rect 307562 246357 307568 246409
rect 307696 246357 307702 246409
rect 307754 246397 307760 246409
rect 307984 246397 307990 246409
rect 307754 246369 307990 246397
rect 307754 246357 307760 246369
rect 307984 246357 307990 246369
rect 308042 246357 308048 246409
rect 312304 246397 312310 246409
rect 308098 246369 312310 246397
rect 308098 246323 308126 246369
rect 312304 246357 312310 246369
rect 312362 246357 312368 246409
rect 313264 246357 313270 246409
rect 313322 246357 313328 246409
rect 313378 246397 313406 246517
rect 328912 246505 328918 246517
rect 328970 246505 328976 246557
rect 330640 246505 330646 246557
rect 330698 246545 330704 246557
rect 342736 246545 342742 246557
rect 330698 246517 342742 246545
rect 330698 246505 330704 246517
rect 342736 246505 342742 246517
rect 342794 246505 342800 246557
rect 347248 246505 347254 246557
rect 347306 246545 347312 246557
rect 349648 246545 349654 246557
rect 347306 246517 349654 246545
rect 347306 246505 347312 246517
rect 349648 246505 349654 246517
rect 349706 246505 349712 246557
rect 366448 246505 366454 246557
rect 366506 246545 366512 246557
rect 366506 246517 367358 246545
rect 366506 246505 366512 246517
rect 313648 246431 313654 246483
rect 313706 246471 313712 246483
rect 339856 246471 339862 246483
rect 313706 246443 339862 246471
rect 313706 246431 313712 246443
rect 339856 246431 339862 246443
rect 339914 246431 339920 246483
rect 349072 246471 349078 246483
rect 340066 246443 340286 246471
rect 313936 246397 313942 246409
rect 313378 246369 313942 246397
rect 313936 246357 313942 246369
rect 313994 246357 314000 246409
rect 317200 246357 317206 246409
rect 317258 246397 317264 246409
rect 317488 246397 317494 246409
rect 317258 246369 317494 246397
rect 317258 246357 317264 246369
rect 317488 246357 317494 246369
rect 317546 246357 317552 246409
rect 328432 246357 328438 246409
rect 328490 246397 328496 246409
rect 340066 246397 340094 246443
rect 328490 246369 340094 246397
rect 340258 246397 340286 246443
rect 347458 246443 349078 246471
rect 347248 246397 347254 246409
rect 340258 246369 347254 246397
rect 328490 246357 328496 246369
rect 347248 246357 347254 246369
rect 347306 246357 347312 246409
rect 287938 246295 308126 246323
rect 309328 246283 309334 246335
rect 309386 246323 309392 246335
rect 347458 246323 347486 246443
rect 349072 246431 349078 246443
rect 349130 246431 349136 246483
rect 367216 246471 367222 246483
rect 349858 246443 367222 246471
rect 348592 246357 348598 246409
rect 348650 246397 348656 246409
rect 349858 246397 349886 246443
rect 367216 246431 367222 246443
rect 367274 246431 367280 246483
rect 367330 246471 367358 246517
rect 367408 246505 367414 246557
rect 367466 246545 367472 246557
rect 367984 246545 367990 246557
rect 367466 246517 367990 246545
rect 367466 246505 367472 246517
rect 367984 246505 367990 246517
rect 368042 246505 368048 246557
rect 368464 246505 368470 246557
rect 368522 246545 368528 246557
rect 397648 246545 397654 246557
rect 368522 246517 397654 246545
rect 368522 246505 368528 246517
rect 397648 246505 397654 246517
rect 397706 246505 397712 246557
rect 397762 246545 397790 246591
rect 406576 246579 406582 246591
rect 406634 246579 406640 246631
rect 406384 246545 406390 246557
rect 397762 246517 406390 246545
rect 406384 246505 406390 246517
rect 406442 246505 406448 246557
rect 382864 246471 382870 246483
rect 367330 246443 382870 246471
rect 382864 246431 382870 246443
rect 382922 246431 382928 246483
rect 382960 246431 382966 246483
rect 383018 246471 383024 246483
rect 389392 246471 389398 246483
rect 383018 246443 389398 246471
rect 383018 246431 383024 246443
rect 389392 246431 389398 246443
rect 389450 246431 389456 246483
rect 397744 246431 397750 246483
rect 397802 246471 397808 246483
rect 397802 246443 407870 246471
rect 397802 246431 397808 246443
rect 348650 246369 349886 246397
rect 348650 246357 348656 246369
rect 349936 246357 349942 246409
rect 349994 246397 350000 246409
rect 368464 246397 368470 246409
rect 349994 246369 368470 246397
rect 349994 246357 350000 246369
rect 368464 246357 368470 246369
rect 368522 246357 368528 246409
rect 369520 246357 369526 246409
rect 369578 246397 369584 246409
rect 370672 246397 370678 246409
rect 369578 246369 370678 246397
rect 369578 246357 369584 246369
rect 370672 246357 370678 246369
rect 370730 246357 370736 246409
rect 372976 246357 372982 246409
rect 373034 246397 373040 246409
rect 407728 246397 407734 246409
rect 373034 246369 407734 246397
rect 373034 246357 373040 246369
rect 407728 246357 407734 246369
rect 407786 246357 407792 246409
rect 309386 246295 347486 246323
rect 309386 246283 309392 246295
rect 348208 246283 348214 246335
rect 348266 246323 348272 246335
rect 388912 246323 388918 246335
rect 348266 246295 388918 246323
rect 348266 246283 348272 246295
rect 388912 246283 388918 246295
rect 388970 246283 388976 246335
rect 397840 246283 397846 246335
rect 397898 246323 397904 246335
rect 407344 246323 407350 246335
rect 397898 246295 407350 246323
rect 397898 246283 397904 246295
rect 407344 246283 407350 246295
rect 407402 246283 407408 246335
rect 407842 246323 407870 246443
rect 408112 246357 408118 246409
rect 408170 246397 408176 246409
rect 410512 246397 410518 246409
rect 408170 246369 410518 246397
rect 408170 246357 408176 246369
rect 410512 246357 410518 246369
rect 410570 246357 410576 246409
rect 410800 246323 410806 246335
rect 407842 246295 410806 246323
rect 410800 246283 410806 246295
rect 410858 246283 410864 246335
rect 674896 246283 674902 246335
rect 674954 246283 674960 246335
rect 287920 246249 287926 246261
rect 268586 246221 287486 246249
rect 287650 246221 287926 246249
rect 268586 246209 268592 246221
rect 65008 246135 65014 246187
rect 65066 246175 65072 246187
rect 80464 246175 80470 246187
rect 65066 246147 80470 246175
rect 65066 246135 65072 246147
rect 80464 246135 80470 246147
rect 80522 246135 80528 246187
rect 145840 246135 145846 246187
rect 145898 246175 145904 246187
rect 145898 246147 155582 246175
rect 145898 246135 145904 246147
rect 43408 246061 43414 246113
rect 43466 246101 43472 246113
rect 155554 246101 155582 246147
rect 207280 246135 207286 246187
rect 207338 246175 207344 246187
rect 207338 246147 260606 246175
rect 207338 246135 207344 246147
rect 161296 246101 161302 246113
rect 43466 246073 80414 246101
rect 43466 246061 43472 246073
rect 80386 245953 80414 246073
rect 106594 246073 148382 246101
rect 155554 246073 161302 246101
rect 106594 246027 106622 246073
rect 86434 245999 106622 246027
rect 148354 246027 148382 246073
rect 161296 246061 161302 246073
rect 161354 246061 161360 246113
rect 161488 246061 161494 246113
rect 161546 246101 161552 246113
rect 161546 246073 208766 246101
rect 161546 246061 161552 246073
rect 155536 246027 155542 246039
rect 148354 245999 155542 246027
rect 86434 245953 86462 245999
rect 155536 245987 155542 245999
rect 155594 245987 155600 246039
rect 208738 246027 208766 246073
rect 210160 246061 210166 246113
rect 210218 246101 210224 246113
rect 228304 246101 228310 246113
rect 210218 246073 228310 246101
rect 210218 246061 210224 246073
rect 228304 246061 228310 246073
rect 228362 246061 228368 246113
rect 249136 246061 249142 246113
rect 249194 246101 249200 246113
rect 260368 246101 260374 246113
rect 249194 246073 260374 246101
rect 249194 246061 249200 246073
rect 260368 246061 260374 246073
rect 260426 246061 260432 246113
rect 260578 246101 260606 246147
rect 268144 246135 268150 246187
rect 268202 246175 268208 246187
rect 287344 246175 287350 246187
rect 268202 246147 287350 246175
rect 268202 246135 268208 246147
rect 287344 246135 287350 246147
rect 287402 246135 287408 246187
rect 287458 246175 287486 246221
rect 287920 246209 287926 246221
rect 287978 246209 287984 246261
rect 288016 246209 288022 246261
rect 288074 246249 288080 246261
rect 328240 246249 328246 246261
rect 288074 246221 328246 246249
rect 288074 246209 288080 246221
rect 328240 246209 328246 246221
rect 328298 246209 328304 246261
rect 328336 246209 328342 246261
rect 328394 246249 328400 246261
rect 339952 246249 339958 246261
rect 328394 246221 339958 246249
rect 328394 246209 328400 246221
rect 339952 246209 339958 246221
rect 340010 246209 340016 246261
rect 340144 246209 340150 246261
rect 340202 246249 340208 246261
rect 391216 246249 391222 246261
rect 340202 246221 348350 246249
rect 340202 246209 340208 246221
rect 287824 246175 287830 246187
rect 287458 246147 287830 246175
rect 287824 246135 287830 246147
rect 287882 246135 287888 246187
rect 288112 246135 288118 246187
rect 288170 246175 288176 246187
rect 307696 246175 307702 246187
rect 288170 246147 307702 246175
rect 288170 246135 288176 246147
rect 307696 246135 307702 246147
rect 307754 246135 307760 246187
rect 307888 246135 307894 246187
rect 307946 246175 307952 246187
rect 328144 246175 328150 246187
rect 307946 246147 328150 246175
rect 307946 246135 307952 246147
rect 328144 246135 328150 246147
rect 328202 246135 328208 246187
rect 328258 246147 329054 246175
rect 268816 246101 268822 246113
rect 260578 246073 268822 246101
rect 268816 246061 268822 246073
rect 268874 246061 268880 246113
rect 268912 246061 268918 246113
rect 268970 246101 268976 246113
rect 277744 246101 277750 246113
rect 268970 246073 277750 246101
rect 268970 246061 268976 246073
rect 277744 246061 277750 246073
rect 277802 246061 277808 246113
rect 328258 246101 328286 246147
rect 277858 246073 328286 246101
rect 329026 246101 329054 246147
rect 329680 246135 329686 246187
rect 329738 246175 329744 246187
rect 339664 246175 339670 246187
rect 329738 246147 339670 246175
rect 329738 246135 329744 246147
rect 339664 246135 339670 246147
rect 339722 246135 339728 246187
rect 339760 246135 339766 246187
rect 339818 246175 339824 246187
rect 348208 246175 348214 246187
rect 339818 246147 348214 246175
rect 339818 246135 339824 246147
rect 348208 246135 348214 246147
rect 348266 246135 348272 246187
rect 348322 246175 348350 246221
rect 348610 246221 391222 246249
rect 348400 246175 348406 246187
rect 348322 246147 348406 246175
rect 348400 246135 348406 246147
rect 348458 246135 348464 246187
rect 348496 246135 348502 246187
rect 348554 246175 348560 246187
rect 348610 246175 348638 246221
rect 391216 246209 391222 246221
rect 391274 246209 391280 246261
rect 397264 246209 397270 246261
rect 397322 246249 397328 246261
rect 411184 246249 411190 246261
rect 397322 246221 411190 246249
rect 397322 246209 397328 246221
rect 411184 246209 411190 246221
rect 411242 246209 411248 246261
rect 348554 246147 348638 246175
rect 348554 246135 348560 246147
rect 349360 246135 349366 246187
rect 349418 246175 349424 246187
rect 382960 246175 382966 246187
rect 349418 246147 382966 246175
rect 349418 246135 349424 246147
rect 382960 246135 382966 246147
rect 383018 246135 383024 246187
rect 390178 246147 391646 246175
rect 329026 246073 371870 246101
rect 236176 246027 236182 246039
rect 208738 245999 236182 246027
rect 236176 245987 236182 245999
rect 236234 245987 236240 246039
rect 248272 246027 248278 246039
rect 246178 245999 248278 246027
rect 80386 245925 86462 245953
rect 161008 245913 161014 245965
rect 161066 245953 161072 245965
rect 163696 245953 163702 245965
rect 161066 245925 163702 245953
rect 161066 245913 161072 245925
rect 163696 245913 163702 245925
rect 163754 245913 163760 245965
rect 208720 245913 208726 245965
rect 208778 245953 208784 245965
rect 246178 245953 246206 245999
rect 248272 245987 248278 245999
rect 248330 245987 248336 246039
rect 259120 245987 259126 246039
rect 259178 246027 259184 246039
rect 277858 246027 277886 246073
rect 368080 246027 368086 246039
rect 259178 245999 277886 246027
rect 277954 245999 368086 246027
rect 259178 245987 259184 245999
rect 208778 245925 246206 245953
rect 208778 245913 208784 245925
rect 251728 245913 251734 245965
rect 251786 245953 251792 245965
rect 277360 245953 277366 245965
rect 251786 245925 277366 245953
rect 251786 245913 251792 245925
rect 277360 245913 277366 245925
rect 277418 245913 277424 245965
rect 277552 245913 277558 245965
rect 277610 245953 277616 245965
rect 277954 245953 277982 245999
rect 368080 245987 368086 245999
rect 368138 245987 368144 246039
rect 277610 245925 277982 245953
rect 277610 245913 277616 245925
rect 278032 245913 278038 245965
rect 278090 245953 278096 245965
rect 367504 245953 367510 245965
rect 278090 245925 367510 245953
rect 278090 245913 278096 245925
rect 367504 245913 367510 245925
rect 367562 245913 367568 245965
rect 371842 245953 371870 246073
rect 390178 245953 390206 246147
rect 391618 246101 391646 246147
rect 397360 246135 397366 246187
rect 397418 246175 397424 246187
rect 411760 246175 411766 246187
rect 397418 246147 411766 246175
rect 397418 246135 397424 246147
rect 411760 246135 411766 246147
rect 411818 246135 411824 246187
rect 505840 246101 505846 246113
rect 391618 246073 505846 246101
rect 505840 246061 505846 246073
rect 505898 246061 505904 246113
rect 674914 246101 674942 246283
rect 675280 246101 675286 246113
rect 674914 246073 675286 246101
rect 675280 246061 675286 246073
rect 675338 246061 675344 246113
rect 391216 245987 391222 246039
rect 391274 246027 391280 246039
rect 412336 246027 412342 246039
rect 391274 245999 412342 246027
rect 391274 245987 391280 245999
rect 412336 245987 412342 245999
rect 412394 245987 412400 246039
rect 371842 245925 390206 245953
rect 398224 245913 398230 245965
rect 398282 245953 398288 245965
rect 408112 245953 408118 245965
rect 398282 245925 408118 245953
rect 398282 245913 398288 245925
rect 408112 245913 408118 245925
rect 408170 245913 408176 245965
rect 160912 245839 160918 245891
rect 160970 245879 160976 245891
rect 165520 245879 165526 245891
rect 160970 245851 165526 245879
rect 160970 245839 160976 245851
rect 165520 245839 165526 245851
rect 165578 245839 165584 245891
rect 229264 245839 229270 245891
rect 229322 245879 229328 245891
rect 246256 245879 246262 245891
rect 229322 245851 246262 245879
rect 229322 245839 229328 245851
rect 246256 245839 246262 245851
rect 246314 245839 246320 245891
rect 247888 245839 247894 245891
rect 247946 245879 247952 245891
rect 251920 245879 251926 245891
rect 247946 245851 251926 245879
rect 247946 245839 247952 245851
rect 251920 245839 251926 245851
rect 251978 245839 251984 245891
rect 356272 245879 356278 245891
rect 254050 245851 356278 245879
rect 155536 245765 155542 245817
rect 155594 245805 155600 245817
rect 161488 245805 161494 245817
rect 155594 245777 161494 245805
rect 155594 245765 155600 245777
rect 161488 245765 161494 245777
rect 161546 245765 161552 245817
rect 210352 245765 210358 245817
rect 210410 245805 210416 245817
rect 226960 245805 226966 245817
rect 210410 245777 226966 245805
rect 210410 245765 210416 245777
rect 226960 245765 226966 245777
rect 227018 245765 227024 245817
rect 227440 245765 227446 245817
rect 227498 245805 227504 245817
rect 231856 245805 231862 245817
rect 227498 245777 231862 245805
rect 227498 245765 227504 245777
rect 231856 245765 231862 245777
rect 231914 245765 231920 245817
rect 248176 245765 248182 245817
rect 248234 245805 248240 245817
rect 252112 245805 252118 245817
rect 248234 245777 252118 245805
rect 248234 245765 248240 245777
rect 252112 245765 252118 245777
rect 252170 245765 252176 245817
rect 206896 245691 206902 245743
rect 206954 245731 206960 245743
rect 207280 245731 207286 245743
rect 206954 245703 207286 245731
rect 206954 245691 206960 245703
rect 207280 245691 207286 245703
rect 207338 245691 207344 245743
rect 224848 245691 224854 245743
rect 224906 245731 224912 245743
rect 228112 245731 228118 245743
rect 224906 245703 228118 245731
rect 224906 245691 224912 245703
rect 228112 245691 228118 245703
rect 228170 245691 228176 245743
rect 251344 245691 251350 245743
rect 251402 245731 251408 245743
rect 254050 245731 254078 245851
rect 356272 245839 356278 245851
rect 356330 245839 356336 245891
rect 366832 245839 366838 245891
rect 366890 245879 366896 245891
rect 372976 245879 372982 245891
rect 366890 245851 372982 245879
rect 366890 245839 366896 245851
rect 372976 245839 372982 245851
rect 373034 245839 373040 245891
rect 389392 245839 389398 245891
rect 389450 245879 389456 245891
rect 411376 245879 411382 245891
rect 389450 245851 411382 245879
rect 389450 245839 389456 245851
rect 411376 245839 411382 245851
rect 411434 245839 411440 245891
rect 255088 245765 255094 245817
rect 255146 245805 255152 245817
rect 330640 245805 330646 245817
rect 255146 245777 330646 245805
rect 255146 245765 255152 245777
rect 330640 245765 330646 245777
rect 330698 245765 330704 245817
rect 330736 245765 330742 245817
rect 330794 245805 330800 245817
rect 357136 245805 357142 245817
rect 330794 245777 357142 245805
rect 330794 245765 330800 245777
rect 357136 245765 357142 245777
rect 357194 245765 357200 245817
rect 367984 245765 367990 245817
rect 368042 245805 368048 245817
rect 373456 245805 373462 245817
rect 368042 245777 373462 245805
rect 368042 245765 368048 245777
rect 373456 245765 373462 245777
rect 373514 245765 373520 245817
rect 388912 245765 388918 245817
rect 388970 245805 388976 245817
rect 406000 245805 406006 245817
rect 388970 245777 406006 245805
rect 388970 245765 388976 245777
rect 406000 245765 406006 245777
rect 406058 245765 406064 245817
rect 251402 245703 254078 245731
rect 251402 245691 251408 245703
rect 254128 245691 254134 245743
rect 254186 245731 254192 245743
rect 348496 245731 348502 245743
rect 254186 245703 348502 245731
rect 254186 245691 254192 245703
rect 348496 245691 348502 245703
rect 348554 245691 348560 245743
rect 348592 245691 348598 245743
rect 348650 245731 348656 245743
rect 357424 245731 357430 245743
rect 348650 245703 357430 245731
rect 348650 245691 348656 245703
rect 357424 245691 357430 245703
rect 357482 245691 357488 245743
rect 367216 245691 367222 245743
rect 367274 245731 367280 245743
rect 370192 245731 370198 245743
rect 367274 245703 370198 245731
rect 367274 245691 367280 245703
rect 370192 245691 370198 245703
rect 370250 245691 370256 245743
rect 382864 245691 382870 245743
rect 382922 245731 382928 245743
rect 408208 245731 408214 245743
rect 382922 245703 408214 245731
rect 382922 245691 382928 245703
rect 408208 245691 408214 245703
rect 408266 245691 408272 245743
rect 227056 245617 227062 245669
rect 227114 245657 227120 245669
rect 232144 245657 232150 245669
rect 227114 245629 232150 245657
rect 227114 245617 227120 245629
rect 232144 245617 232150 245629
rect 232202 245617 232208 245669
rect 246448 245617 246454 245669
rect 246506 245657 246512 245669
rect 267472 245657 267478 245669
rect 246506 245629 267478 245657
rect 246506 245617 246512 245629
rect 267472 245617 267478 245629
rect 267530 245617 267536 245669
rect 269008 245617 269014 245669
rect 269066 245657 269072 245669
rect 369232 245657 369238 245669
rect 269066 245629 369238 245657
rect 269066 245617 269072 245629
rect 369232 245617 369238 245629
rect 369290 245617 369296 245669
rect 389008 245617 389014 245669
rect 389066 245657 389072 245669
rect 406768 245657 406774 245669
rect 389066 245629 406774 245657
rect 389066 245617 389072 245629
rect 406768 245617 406774 245629
rect 406826 245617 406832 245669
rect 226480 245543 226486 245595
rect 226538 245583 226544 245595
rect 231376 245583 231382 245595
rect 226538 245555 231382 245583
rect 226538 245543 226544 245555
rect 231376 245543 231382 245555
rect 231434 245543 231440 245595
rect 236176 245543 236182 245595
rect 236234 245583 236240 245595
rect 249040 245583 249046 245595
rect 236234 245555 249046 245583
rect 236234 245543 236240 245555
rect 249040 245543 249046 245555
rect 249098 245543 249104 245595
rect 268432 245543 268438 245595
rect 268490 245583 268496 245595
rect 277648 245583 277654 245595
rect 268490 245555 277654 245583
rect 268490 245543 268496 245555
rect 277648 245543 277654 245555
rect 277706 245543 277712 245595
rect 277744 245543 277750 245595
rect 277802 245583 277808 245595
rect 370960 245583 370966 245595
rect 277802 245555 370966 245583
rect 277802 245543 277808 245555
rect 370960 245543 370966 245555
rect 371018 245543 371024 245595
rect 403024 245543 403030 245595
rect 403082 245583 403088 245595
rect 410320 245583 410326 245595
rect 403082 245555 410326 245583
rect 403082 245543 403088 245555
rect 410320 245543 410326 245555
rect 410378 245543 410384 245595
rect 223120 245469 223126 245521
rect 223178 245509 223184 245521
rect 251728 245509 251734 245521
rect 223178 245481 251734 245509
rect 223178 245469 223184 245481
rect 251728 245469 251734 245481
rect 251786 245469 251792 245521
rect 252400 245469 252406 245521
rect 252458 245509 252464 245521
rect 330736 245509 330742 245521
rect 252458 245481 330742 245509
rect 252458 245469 252464 245481
rect 330736 245469 330742 245481
rect 330794 245469 330800 245521
rect 348496 245509 348502 245521
rect 330850 245481 348502 245509
rect 198832 245395 198838 245447
rect 198890 245435 198896 245447
rect 213136 245435 213142 245447
rect 198890 245407 213142 245435
rect 198890 245395 198896 245407
rect 213136 245395 213142 245407
rect 213194 245395 213200 245447
rect 246160 245395 246166 245447
rect 246218 245435 246224 245447
rect 248368 245435 248374 245447
rect 246218 245407 248374 245435
rect 246218 245395 246224 245407
rect 248368 245395 248374 245407
rect 248426 245395 248432 245447
rect 253360 245395 253366 245447
rect 253418 245435 253424 245447
rect 330850 245435 330878 245481
rect 348496 245469 348502 245481
rect 348554 245469 348560 245521
rect 355792 245509 355798 245521
rect 348610 245481 355798 245509
rect 348610 245435 348638 245481
rect 355792 245469 355798 245481
rect 355850 245469 355856 245521
rect 390256 245509 390262 245521
rect 360034 245481 390262 245509
rect 253418 245407 330878 245435
rect 330946 245407 348638 245435
rect 253418 245395 253424 245407
rect 210160 245321 210166 245373
rect 210218 245361 210224 245373
rect 231856 245361 231862 245373
rect 210218 245333 231862 245361
rect 210218 245321 210224 245333
rect 231856 245321 231862 245333
rect 231914 245321 231920 245373
rect 246256 245321 246262 245373
rect 246314 245361 246320 245373
rect 249136 245361 249142 245373
rect 246314 245333 249142 245361
rect 246314 245321 246320 245333
rect 249136 245321 249142 245333
rect 249194 245321 249200 245373
rect 249616 245321 249622 245373
rect 249674 245361 249680 245373
rect 330946 245361 330974 245407
rect 348688 245395 348694 245447
rect 348746 245435 348752 245447
rect 360034 245435 360062 245481
rect 390256 245469 390262 245481
rect 390314 245469 390320 245521
rect 405904 245469 405910 245521
rect 405962 245509 405968 245521
rect 412144 245509 412150 245521
rect 405962 245481 412150 245509
rect 405962 245469 405968 245481
rect 412144 245469 412150 245481
rect 412202 245469 412208 245521
rect 348746 245407 360062 245435
rect 348746 245395 348752 245407
rect 249674 245333 330974 245361
rect 249674 245321 249680 245333
rect 331024 245321 331030 245373
rect 331082 245361 331088 245373
rect 370096 245361 370102 245373
rect 331082 245333 370102 245361
rect 331082 245321 331088 245333
rect 370096 245321 370102 245333
rect 370154 245321 370160 245373
rect 250288 245247 250294 245299
rect 250346 245287 250352 245299
rect 250346 245259 331166 245287
rect 250346 245247 250352 245259
rect 216592 245173 216598 245225
rect 216650 245213 216656 245225
rect 331024 245213 331030 245225
rect 216650 245185 331030 245213
rect 216650 245173 216656 245185
rect 331024 245173 331030 245185
rect 331082 245173 331088 245225
rect 331138 245213 331166 245259
rect 339664 245247 339670 245299
rect 339722 245287 339728 245299
rect 369904 245287 369910 245299
rect 339722 245259 369910 245287
rect 339722 245247 339728 245259
rect 369904 245247 369910 245259
rect 369962 245247 369968 245299
rect 370192 245247 370198 245299
rect 370250 245287 370256 245299
rect 380176 245287 380182 245299
rect 370250 245259 380182 245287
rect 370250 245247 370256 245259
rect 380176 245247 380182 245259
rect 380234 245247 380240 245299
rect 355888 245213 355894 245225
rect 331138 245185 355894 245213
rect 355888 245173 355894 245185
rect 355946 245173 355952 245225
rect 411472 245213 411478 245225
rect 398818 245185 411478 245213
rect 231856 245099 231862 245151
rect 231914 245139 231920 245151
rect 260272 245139 260278 245151
rect 231914 245111 260278 245139
rect 231914 245099 231920 245111
rect 260272 245099 260278 245111
rect 260330 245099 260336 245151
rect 261808 245099 261814 245151
rect 261866 245139 261872 245151
rect 338416 245139 338422 245151
rect 261866 245111 338422 245139
rect 261866 245099 261872 245111
rect 338416 245099 338422 245111
rect 338474 245099 338480 245151
rect 339472 245099 339478 245151
rect 339530 245139 339536 245151
rect 339530 245111 368990 245139
rect 339530 245099 339536 245111
rect 263440 245025 263446 245077
rect 263498 245065 263504 245077
rect 263498 245037 267614 245065
rect 263498 245025 263504 245037
rect 263824 244951 263830 245003
rect 263882 244991 263888 245003
rect 267472 244991 267478 245003
rect 263882 244963 267478 244991
rect 263882 244951 263888 244963
rect 267472 244951 267478 244963
rect 267530 244951 267536 245003
rect 267586 244991 267614 245037
rect 269488 245025 269494 245077
rect 269546 245065 269552 245077
rect 269546 245037 277886 245065
rect 269546 245025 269552 245037
rect 277552 244991 277558 245003
rect 267586 244963 277558 244991
rect 277552 244951 277558 244963
rect 277610 244951 277616 245003
rect 277858 244991 277886 245037
rect 277936 245025 277942 245077
rect 277994 245065 278000 245077
rect 368962 245065 368990 245111
rect 369904 245099 369910 245151
rect 369962 245139 369968 245151
rect 398704 245139 398710 245151
rect 369962 245111 398710 245139
rect 369962 245099 369968 245111
rect 398704 245099 398710 245111
rect 398762 245099 398768 245151
rect 372016 245065 372022 245077
rect 277994 245037 328574 245065
rect 277994 245025 278000 245037
rect 319696 244991 319702 245003
rect 277858 244963 319702 244991
rect 319696 244951 319702 244963
rect 319754 244951 319760 245003
rect 328546 244991 328574 245037
rect 339778 245037 368894 245065
rect 368962 245037 372022 245065
rect 339778 244991 339806 245037
rect 328546 244963 339806 244991
rect 339952 244951 339958 245003
rect 340010 244991 340016 245003
rect 368866 244991 368894 245037
rect 372016 245025 372022 245037
rect 372074 245025 372080 245077
rect 380176 245025 380182 245077
rect 380234 245065 380240 245077
rect 398818 245065 398846 245185
rect 411472 245173 411478 245185
rect 411530 245173 411536 245225
rect 380234 245037 398846 245065
rect 380234 245025 380240 245037
rect 374032 244991 374038 245003
rect 340010 244963 362846 244991
rect 368866 244963 374038 244991
rect 340010 244951 340016 244963
rect 42544 244877 42550 244929
rect 42602 244917 42608 244929
rect 214288 244917 214294 244929
rect 42602 244889 214294 244917
rect 42602 244877 42608 244889
rect 214288 244877 214294 244889
rect 214346 244877 214352 244929
rect 216496 244877 216502 244929
rect 216554 244917 216560 244929
rect 338128 244917 338134 244929
rect 216554 244889 338134 244917
rect 216554 244877 216560 244889
rect 338128 244877 338134 244889
rect 338186 244877 338192 244929
rect 338416 244877 338422 244929
rect 338474 244917 338480 244929
rect 339472 244917 339478 244929
rect 338474 244889 339478 244917
rect 338474 244877 338480 244889
rect 339472 244877 339478 244889
rect 339530 244877 339536 244929
rect 348880 244877 348886 244929
rect 348938 244917 348944 244929
rect 358000 244917 358006 244929
rect 348938 244889 358006 244917
rect 348938 244877 348944 244889
rect 358000 244877 358006 244889
rect 358058 244877 358064 244929
rect 210064 244803 210070 244855
rect 210122 244843 210128 244855
rect 228592 244843 228598 244855
rect 210122 244815 228598 244843
rect 210122 244803 210128 244815
rect 228592 244803 228598 244815
rect 228650 244803 228656 244855
rect 260272 244803 260278 244855
rect 260330 244843 260336 244855
rect 267952 244843 267958 244855
rect 260330 244815 267958 244843
rect 260330 244803 260336 244815
rect 267952 244803 267958 244815
rect 268010 244803 268016 244855
rect 268048 244803 268054 244855
rect 268106 244843 268112 244855
rect 278032 244843 278038 244855
rect 268106 244815 278038 244843
rect 268106 244803 268112 244815
rect 278032 244803 278038 244815
rect 278090 244803 278096 244855
rect 278128 244803 278134 244855
rect 278186 244843 278192 244855
rect 287248 244843 287254 244855
rect 278186 244815 287254 244843
rect 278186 244803 278192 244815
rect 287248 244803 287254 244815
rect 287306 244803 287312 244855
rect 287344 244803 287350 244855
rect 287402 244843 287408 244855
rect 288784 244843 288790 244855
rect 287402 244815 288790 244843
rect 287402 244803 287408 244815
rect 288784 244803 288790 244815
rect 288842 244803 288848 244855
rect 288880 244803 288886 244855
rect 288938 244843 288944 244855
rect 309424 244843 309430 244855
rect 288938 244815 309430 244843
rect 288938 244803 288944 244815
rect 309424 244803 309430 244815
rect 309482 244803 309488 244855
rect 311824 244803 311830 244855
rect 311882 244843 311888 244855
rect 311882 244815 328574 244843
rect 311882 244803 311888 244815
rect 95056 244729 95062 244781
rect 95114 244769 95120 244781
rect 139984 244769 139990 244781
rect 95114 244741 139990 244769
rect 95114 244729 95120 244741
rect 139984 244729 139990 244741
rect 140042 244729 140048 244781
rect 260944 244729 260950 244781
rect 261002 244769 261008 244781
rect 316816 244769 316822 244781
rect 261002 244741 316822 244769
rect 261002 244729 261008 244741
rect 316816 244729 316822 244741
rect 316874 244729 316880 244781
rect 316912 244729 316918 244781
rect 316970 244769 316976 244781
rect 321232 244769 321238 244781
rect 316970 244741 321238 244769
rect 316970 244729 316976 244741
rect 321232 244729 321238 244741
rect 321290 244729 321296 244781
rect 328546 244769 328574 244815
rect 328624 244803 328630 244855
rect 328682 244843 328688 244855
rect 339568 244843 339574 244855
rect 328682 244815 339574 244843
rect 328682 244803 328688 244815
rect 339568 244803 339574 244815
rect 339626 244803 339632 244855
rect 348688 244843 348694 244855
rect 340066 244815 348694 244843
rect 329680 244769 329686 244781
rect 328546 244741 329686 244769
rect 329680 244729 329686 244741
rect 329738 244729 329744 244781
rect 90640 244655 90646 244707
rect 90698 244695 90704 244707
rect 142480 244695 142486 244707
rect 90698 244667 142486 244695
rect 90698 244655 90704 244667
rect 142480 244655 142486 244667
rect 142538 244655 142544 244707
rect 262864 244655 262870 244707
rect 262922 244695 262928 244707
rect 273040 244695 273046 244707
rect 262922 244667 273046 244695
rect 262922 244655 262928 244667
rect 273040 244655 273046 244667
rect 273098 244655 273104 244707
rect 276016 244655 276022 244707
rect 276074 244695 276080 244707
rect 287440 244695 287446 244707
rect 276074 244667 287446 244695
rect 276074 244655 276080 244667
rect 287440 244655 287446 244667
rect 287498 244655 287504 244707
rect 287920 244655 287926 244707
rect 287978 244695 287984 244707
rect 307312 244695 307318 244707
rect 287978 244667 307318 244695
rect 287978 244655 287984 244667
rect 307312 244655 307318 244667
rect 307370 244655 307376 244707
rect 307408 244655 307414 244707
rect 307466 244695 307472 244707
rect 311824 244695 311830 244707
rect 307466 244667 311830 244695
rect 307466 244655 307472 244667
rect 311824 244655 311830 244667
rect 311882 244655 311888 244707
rect 311920 244655 311926 244707
rect 311978 244695 311984 244707
rect 317008 244695 317014 244707
rect 311978 244667 317014 244695
rect 311978 244655 311984 244667
rect 317008 244655 317014 244667
rect 317066 244655 317072 244707
rect 317104 244655 317110 244707
rect 317162 244695 317168 244707
rect 339952 244695 339958 244707
rect 317162 244667 339958 244695
rect 317162 244655 317168 244667
rect 339952 244655 339958 244667
rect 340010 244655 340016 244707
rect 138160 244581 138166 244633
rect 138218 244621 138224 244633
rect 206992 244621 206998 244633
rect 138218 244593 206998 244621
rect 138218 244581 138224 244593
rect 206992 244581 206998 244593
rect 207050 244581 207056 244633
rect 265936 244581 265942 244633
rect 265994 244621 266000 244633
rect 265994 244593 274046 244621
rect 265994 244581 266000 244593
rect 135280 244507 135286 244559
rect 135338 244547 135344 244559
rect 207088 244547 207094 244559
rect 135338 244519 207094 244547
rect 135338 244507 135344 244519
rect 207088 244507 207094 244519
rect 207146 244507 207152 244559
rect 267472 244507 267478 244559
rect 267530 244547 267536 244559
rect 268048 244547 268054 244559
rect 267530 244519 268054 244547
rect 267530 244507 267536 244519
rect 268048 244507 268054 244519
rect 268106 244507 268112 244559
rect 132400 244433 132406 244485
rect 132458 244473 132464 244485
rect 205168 244473 205174 244485
rect 132458 244445 205174 244473
rect 132458 244433 132464 244445
rect 205168 244433 205174 244445
rect 205226 244433 205232 244485
rect 267952 244433 267958 244485
rect 268010 244473 268016 244485
rect 269200 244473 269206 244485
rect 268010 244445 269206 244473
rect 268010 244433 268016 244445
rect 269200 244433 269206 244445
rect 269258 244433 269264 244485
rect 126640 244359 126646 244411
rect 126698 244399 126704 244411
rect 205552 244399 205558 244411
rect 126698 244371 205558 244399
rect 126698 244359 126704 244371
rect 205552 244359 205558 244371
rect 205610 244359 205616 244411
rect 274018 244399 274046 244593
rect 274096 244581 274102 244633
rect 274154 244621 274160 244633
rect 278032 244621 278038 244633
rect 274154 244593 278038 244621
rect 274154 244581 274160 244593
rect 278032 244581 278038 244593
rect 278090 244581 278096 244633
rect 278128 244581 278134 244633
rect 278186 244621 278192 244633
rect 308944 244621 308950 244633
rect 278186 244593 287390 244621
rect 278186 244581 278192 244593
rect 276880 244507 276886 244559
rect 276938 244547 276944 244559
rect 277744 244547 277750 244559
rect 276938 244519 277750 244547
rect 276938 244507 276944 244519
rect 277744 244507 277750 244519
rect 277802 244507 277808 244559
rect 287362 244547 287390 244593
rect 287650 244593 308950 244621
rect 287650 244547 287678 244593
rect 308944 244581 308950 244593
rect 309002 244581 309008 244633
rect 309232 244581 309238 244633
rect 309290 244621 309296 244633
rect 314032 244621 314038 244633
rect 309290 244593 314038 244621
rect 309290 244581 309296 244593
rect 314032 244581 314038 244593
rect 314090 244581 314096 244633
rect 317218 244593 317390 244621
rect 287362 244519 287678 244547
rect 287824 244507 287830 244559
rect 287882 244547 287888 244559
rect 306640 244547 306646 244559
rect 287882 244519 306646 244547
rect 287882 244507 287888 244519
rect 306640 244507 306646 244519
rect 306698 244507 306704 244559
rect 307504 244507 307510 244559
rect 307562 244547 307568 244559
rect 307562 244519 310910 244547
rect 307562 244507 307568 244519
rect 277840 244433 277846 244485
rect 277898 244473 277904 244485
rect 310768 244473 310774 244485
rect 277898 244445 310774 244473
rect 277898 244433 277904 244445
rect 310768 244433 310774 244445
rect 310826 244433 310832 244485
rect 310882 244473 310910 244519
rect 312016 244507 312022 244559
rect 312074 244547 312080 244559
rect 317218 244547 317246 244593
rect 312074 244519 317246 244547
rect 317362 244547 317390 244593
rect 319600 244581 319606 244633
rect 319658 244621 319664 244633
rect 338320 244621 338326 244633
rect 319658 244593 338326 244621
rect 319658 244581 319664 244593
rect 338320 244581 338326 244593
rect 338378 244581 338384 244633
rect 339568 244581 339574 244633
rect 339626 244621 339632 244633
rect 340066 244621 340094 244815
rect 348688 244803 348694 244815
rect 348746 244803 348752 244855
rect 362818 244843 362846 244963
rect 374032 244951 374038 244963
rect 374090 244951 374096 245003
rect 374608 244843 374614 244855
rect 362818 244815 374614 244843
rect 374608 244803 374614 244815
rect 374666 244803 374672 244855
rect 389296 244769 389302 244781
rect 347266 244741 389302 244769
rect 342544 244655 342550 244707
rect 342602 244695 342608 244707
rect 347266 244695 347294 244741
rect 389296 244729 389302 244741
rect 389354 244729 389360 244781
rect 342602 244667 347294 244695
rect 342602 244655 342608 244667
rect 339626 244593 340094 244621
rect 339626 244581 339632 244593
rect 340144 244581 340150 244633
rect 340202 244621 340208 244633
rect 349936 244621 349942 244633
rect 340202 244593 349942 244621
rect 340202 244581 340208 244593
rect 349936 244581 349942 244593
rect 349994 244581 350000 244633
rect 367888 244547 367894 244559
rect 317362 244519 367894 244547
rect 312074 244507 312080 244519
rect 367888 244507 367894 244519
rect 367946 244507 367952 244559
rect 310882 244445 312062 244473
rect 311920 244399 311926 244411
rect 274018 244371 311926 244399
rect 311920 244359 311926 244371
rect 311978 244359 311984 244411
rect 312034 244399 312062 244445
rect 312400 244433 312406 244485
rect 312458 244473 312464 244485
rect 368752 244473 368758 244485
rect 312458 244445 368758 244473
rect 312458 244433 312464 244445
rect 368752 244433 368758 244445
rect 368810 244433 368816 244485
rect 339856 244399 339862 244411
rect 312034 244371 319742 244399
rect 123760 244285 123766 244337
rect 123818 244325 123824 244337
rect 205360 244325 205366 244337
rect 123818 244297 205366 244325
rect 123818 244285 123824 244297
rect 205360 244285 205366 244297
rect 205418 244285 205424 244337
rect 235120 244285 235126 244337
rect 235178 244325 235184 244337
rect 267184 244325 267190 244337
rect 235178 244297 267190 244325
rect 235178 244285 235184 244297
rect 267184 244285 267190 244297
rect 267242 244285 267248 244337
rect 273040 244285 273046 244337
rect 273098 244325 273104 244337
rect 287728 244325 287734 244337
rect 273098 244297 287734 244325
rect 273098 244285 273104 244297
rect 287728 244285 287734 244297
rect 287786 244285 287792 244337
rect 290032 244285 290038 244337
rect 290090 244325 290096 244337
rect 295696 244325 295702 244337
rect 290090 244297 295702 244325
rect 290090 244285 290096 244297
rect 295696 244285 295702 244297
rect 295754 244285 295760 244337
rect 297424 244285 297430 244337
rect 297482 244325 297488 244337
rect 314896 244325 314902 244337
rect 297482 244297 314902 244325
rect 297482 244285 297488 244297
rect 314896 244285 314902 244297
rect 314954 244285 314960 244337
rect 319600 244325 319606 244337
rect 317122 244297 319606 244325
rect 120880 244211 120886 244263
rect 120938 244251 120944 244263
rect 205648 244251 205654 244263
rect 120938 244223 205654 244251
rect 120938 244211 120944 244223
rect 205648 244211 205654 244223
rect 205706 244211 205712 244263
rect 260752 244211 260758 244263
rect 260810 244251 260816 244263
rect 268144 244251 268150 244263
rect 260810 244223 268150 244251
rect 260810 244211 260816 244223
rect 268144 244211 268150 244223
rect 268202 244211 268208 244263
rect 268240 244211 268246 244263
rect 268298 244251 268304 244263
rect 287440 244251 287446 244263
rect 268298 244223 287446 244251
rect 268298 244211 268304 244223
rect 287440 244211 287446 244223
rect 287498 244211 287504 244263
rect 287920 244211 287926 244263
rect 287978 244251 287984 244263
rect 317122 244251 317150 244297
rect 319600 244285 319606 244297
rect 319658 244285 319664 244337
rect 287978 244223 317150 244251
rect 319714 244251 319742 244371
rect 322594 244371 339862 244399
rect 319792 244285 319798 244337
rect 319850 244325 319856 244337
rect 322594 244325 322622 244371
rect 339856 244359 339862 244371
rect 339914 244359 339920 244411
rect 319850 244297 322622 244325
rect 319850 244285 319856 244297
rect 349360 244251 349366 244263
rect 319714 244223 349366 244251
rect 287978 244211 287984 244223
rect 349360 244211 349366 244223
rect 349418 244211 349424 244263
rect 118000 244137 118006 244189
rect 118058 244177 118064 244189
rect 204976 244177 204982 244189
rect 118058 244149 204982 244177
rect 118058 244137 118064 244149
rect 204976 244137 204982 244149
rect 205034 244137 205040 244189
rect 258352 244137 258358 244189
rect 258410 244177 258416 244189
rect 317200 244177 317206 244189
rect 258410 244149 317206 244177
rect 258410 244137 258416 244149
rect 317200 244137 317206 244149
rect 317258 244137 317264 244189
rect 321232 244137 321238 244189
rect 321290 244177 321296 244189
rect 329296 244177 329302 244189
rect 321290 244149 329302 244177
rect 321290 244137 321296 244149
rect 329296 244137 329302 244149
rect 329354 244137 329360 244189
rect 338128 244137 338134 244189
rect 338186 244177 338192 244189
rect 351568 244177 351574 244189
rect 338186 244149 351574 244177
rect 338186 244137 338192 244149
rect 351568 244137 351574 244149
rect 351626 244137 351632 244189
rect 112240 244063 112246 244115
rect 112298 244103 112304 244115
rect 206608 244103 206614 244115
rect 112298 244075 206614 244103
rect 112298 244063 112304 244075
rect 206608 244063 206614 244075
rect 206666 244063 206672 244115
rect 261136 244063 261142 244115
rect 261194 244103 261200 244115
rect 337552 244103 337558 244115
rect 261194 244075 337558 244103
rect 261194 244063 261200 244075
rect 337552 244063 337558 244075
rect 337610 244063 337616 244115
rect 109360 243989 109366 244041
rect 109418 244029 109424 244041
rect 205744 244029 205750 244041
rect 109418 244001 205750 244029
rect 109418 243989 109424 244001
rect 205744 243989 205750 244001
rect 205802 243989 205808 244041
rect 256336 243989 256342 244041
rect 256394 244029 256400 244041
rect 335344 244029 335350 244041
rect 256394 244001 335350 244029
rect 256394 243989 256400 244001
rect 335344 243989 335350 244001
rect 335402 243989 335408 244041
rect 106480 243915 106486 243967
rect 106538 243955 106544 243967
rect 206512 243955 206518 243967
rect 106538 243927 206518 243955
rect 106538 243915 106544 243927
rect 206512 243915 206518 243927
rect 206570 243915 206576 243967
rect 260080 243915 260086 243967
rect 260138 243955 260144 243967
rect 316816 243955 316822 243967
rect 260138 243927 316822 243955
rect 260138 243915 260144 243927
rect 316816 243915 316822 243927
rect 316874 243915 316880 243967
rect 328240 243915 328246 243967
rect 328298 243955 328304 243967
rect 339760 243955 339766 243967
rect 328298 243927 339766 243955
rect 328298 243915 328304 243927
rect 339760 243915 339766 243927
rect 339818 243915 339824 243967
rect 103600 243841 103606 243893
rect 103658 243881 103664 243893
rect 206320 243881 206326 243893
rect 103658 243853 206326 243881
rect 103658 243841 103664 243853
rect 206320 243841 206326 243853
rect 206378 243841 206384 243893
rect 207184 243841 207190 243893
rect 207242 243881 207248 243893
rect 268048 243881 268054 243893
rect 207242 243853 268054 243881
rect 207242 243841 207248 243853
rect 268048 243841 268054 243853
rect 268106 243841 268112 243893
rect 268144 243841 268150 243893
rect 268202 243881 268208 243893
rect 285232 243881 285238 243893
rect 268202 243853 285238 243881
rect 268202 243841 268208 243853
rect 285232 243841 285238 243853
rect 285290 243841 285296 243893
rect 288112 243841 288118 243893
rect 288170 243881 288176 243893
rect 308080 243881 308086 243893
rect 288170 243853 308086 243881
rect 288170 243841 288176 243853
rect 308080 243841 308086 243853
rect 308138 243841 308144 243893
rect 313360 243841 313366 243893
rect 313418 243881 313424 243893
rect 370288 243881 370294 243893
rect 313418 243853 370294 243881
rect 313418 243841 313424 243853
rect 370288 243841 370294 243853
rect 370346 243841 370352 243893
rect 100720 243767 100726 243819
rect 100778 243807 100784 243819
rect 206416 243807 206422 243819
rect 100778 243779 206422 243807
rect 100778 243767 100784 243779
rect 206416 243767 206422 243779
rect 206474 243767 206480 243819
rect 245392 243767 245398 243819
rect 245450 243807 245456 243819
rect 353680 243807 353686 243819
rect 245450 243779 353686 243807
rect 245450 243767 245456 243779
rect 353680 243767 353686 243779
rect 353738 243767 353744 243819
rect 94960 243693 94966 243745
rect 95018 243733 95024 243745
rect 206224 243733 206230 243745
rect 95018 243705 206230 243733
rect 95018 243693 95024 243705
rect 206224 243693 206230 243705
rect 206282 243693 206288 243745
rect 239344 243693 239350 243745
rect 239402 243733 239408 243745
rect 350800 243733 350806 243745
rect 239402 243705 350806 243733
rect 239402 243693 239408 243705
rect 350800 243693 350806 243705
rect 350858 243693 350864 243745
rect 604816 243693 604822 243745
rect 604874 243733 604880 243745
rect 624880 243733 624886 243745
rect 604874 243705 624886 243733
rect 604874 243693 604880 243705
rect 624880 243693 624886 243705
rect 624938 243693 624944 243745
rect 92080 243619 92086 243671
rect 92138 243659 92144 243671
rect 206032 243659 206038 243671
rect 92138 243631 206038 243659
rect 92138 243619 92144 243631
rect 206032 243619 206038 243631
rect 206090 243619 206096 243671
rect 206800 243619 206806 243671
rect 206858 243659 206864 243671
rect 207184 243659 207190 243671
rect 206858 243631 207190 243659
rect 206858 243619 206864 243631
rect 207184 243619 207190 243631
rect 207242 243619 207248 243671
rect 227056 243619 227062 243671
rect 227114 243659 227120 243671
rect 231664 243659 231670 243671
rect 227114 243631 231670 243659
rect 227114 243619 227120 243631
rect 231664 243619 231670 243631
rect 231722 243619 231728 243671
rect 231760 243619 231766 243671
rect 231818 243659 231824 243671
rect 347344 243659 347350 243671
rect 231818 243631 347350 243659
rect 231818 243619 231824 243631
rect 347344 243619 347350 243631
rect 347402 243619 347408 243671
rect 443536 243619 443542 243671
rect 443594 243659 443600 243671
rect 463600 243659 463606 243671
rect 443594 243631 463606 243659
rect 443594 243619 443600 243631
rect 463600 243619 463606 243631
rect 463658 243619 463664 243671
rect 483856 243619 483862 243671
rect 483914 243659 483920 243671
rect 503920 243659 503926 243671
rect 483914 243631 503926 243659
rect 483914 243619 483920 243631
rect 503920 243619 503926 243631
rect 503978 243619 503984 243671
rect 524176 243619 524182 243671
rect 524234 243659 524240 243671
rect 544240 243659 544246 243671
rect 524234 243631 544246 243659
rect 524234 243619 524240 243631
rect 544240 243619 544246 243631
rect 544298 243619 544304 243671
rect 564496 243619 564502 243671
rect 564554 243659 564560 243671
rect 584560 243659 584566 243671
rect 564554 243631 584566 243659
rect 564554 243619 564560 243631
rect 584560 243619 584566 243631
rect 584618 243619 584624 243671
rect 645136 243619 645142 243671
rect 645194 243659 645200 243671
rect 648016 243659 648022 243671
rect 645194 243631 648022 243659
rect 645194 243619 645200 243631
rect 648016 243619 648022 243631
rect 648074 243619 648080 243671
rect 86320 243545 86326 243597
rect 86378 243585 86384 243597
rect 206704 243585 206710 243597
rect 86378 243557 206710 243585
rect 86378 243545 86384 243557
rect 206704 243545 206710 243557
rect 206762 243545 206768 243597
rect 236272 243545 236278 243597
rect 236330 243585 236336 243597
rect 349264 243585 349270 243597
rect 236330 243557 349270 243585
rect 236330 243545 236336 243557
rect 349264 243545 349270 243557
rect 349322 243545 349328 243597
rect 80560 243471 80566 243523
rect 80618 243511 80624 243523
rect 206800 243511 206806 243523
rect 80618 243483 206806 243511
rect 80618 243471 80624 243483
rect 206800 243471 206806 243483
rect 206858 243471 206864 243523
rect 228496 243471 228502 243523
rect 228554 243511 228560 243523
rect 345616 243511 345622 243523
rect 228554 243483 345622 243511
rect 228554 243471 228560 243483
rect 345616 243471 345622 243483
rect 345674 243471 345680 243523
rect 77680 243397 77686 243449
rect 77738 243437 77744 243449
rect 205936 243437 205942 243449
rect 77738 243409 205942 243437
rect 77738 243397 77744 243409
rect 205936 243397 205942 243409
rect 205994 243397 206000 243449
rect 226768 243397 226774 243449
rect 226826 243437 226832 243449
rect 345136 243437 345142 243449
rect 226826 243409 345142 243437
rect 226826 243397 226832 243409
rect 345136 243397 345142 243409
rect 345194 243397 345200 243449
rect 69040 243323 69046 243375
rect 69098 243363 69104 243375
rect 206128 243363 206134 243375
rect 69098 243335 206134 243363
rect 69098 243323 69104 243335
rect 206128 243323 206134 243335
rect 206186 243323 206192 243375
rect 229744 243323 229750 243375
rect 229802 243363 229808 243375
rect 297808 243363 297814 243375
rect 229802 243335 297814 243363
rect 229802 243323 229808 243335
rect 297808 243323 297814 243335
rect 297866 243323 297872 243375
rect 298192 243363 298198 243375
rect 298114 243335 298198 243363
rect 199600 243249 199606 243301
rect 199658 243289 199664 243301
rect 213520 243289 213526 243301
rect 199658 243261 213526 243289
rect 199658 243249 199664 243261
rect 213520 243249 213526 243261
rect 213578 243249 213584 243301
rect 264784 243249 264790 243301
rect 264842 243289 264848 243301
rect 277840 243289 277846 243301
rect 264842 243261 277846 243289
rect 264842 243249 264848 243261
rect 277840 243249 277846 243261
rect 277898 243249 277904 243301
rect 283216 243249 283222 243301
rect 283274 243289 283280 243301
rect 298114 243289 298142 243335
rect 298192 243323 298198 243335
rect 298250 243323 298256 243375
rect 298480 243323 298486 243375
rect 298538 243323 298544 243375
rect 299440 243323 299446 243375
rect 299498 243363 299504 243375
rect 346384 243363 346390 243375
rect 299498 243335 346390 243363
rect 299498 243323 299504 243335
rect 346384 243323 346390 243335
rect 346442 243323 346448 243375
rect 283274 243261 298142 243289
rect 283274 243249 283280 243261
rect 298288 243249 298294 243301
rect 298346 243289 298352 243301
rect 298498 243289 298526 243323
rect 298346 243261 298526 243289
rect 298346 243249 298352 243261
rect 316912 243249 316918 243301
rect 316970 243289 316976 243301
rect 340720 243289 340726 243301
rect 316970 243261 340726 243289
rect 316970 243249 316976 243261
rect 340720 243249 340726 243261
rect 340778 243249 340784 243301
rect 342736 243249 342742 243301
rect 342794 243289 342800 243301
rect 358384 243289 358390 243301
rect 342794 243261 358390 243289
rect 342794 243249 342800 243261
rect 358384 243249 358390 243261
rect 358442 243249 358448 243301
rect 267376 243175 267382 243227
rect 267434 243215 267440 243227
rect 298576 243215 298582 243227
rect 267434 243187 298582 243215
rect 267434 243175 267440 243187
rect 298576 243175 298582 243187
rect 298634 243175 298640 243227
rect 298672 243175 298678 243227
rect 298730 243215 298736 243227
rect 305104 243215 305110 243227
rect 298730 243187 305110 243215
rect 298730 243175 298736 243187
rect 305104 243175 305110 243187
rect 305162 243175 305168 243227
rect 317200 243175 317206 243227
rect 317258 243215 317264 243227
rect 336304 243215 336310 243227
rect 317258 243187 336310 243215
rect 317258 243175 317264 243187
rect 336304 243175 336310 243187
rect 336362 243175 336368 243227
rect 260368 243101 260374 243153
rect 260426 243141 260432 243153
rect 268624 243141 268630 243153
rect 260426 243113 268630 243141
rect 260426 243101 260432 243113
rect 268624 243101 268630 243113
rect 268682 243101 268688 243153
rect 270832 243101 270838 243153
rect 270890 243141 270896 243153
rect 293104 243141 293110 243153
rect 270890 243113 293110 243141
rect 270890 243101 270896 243113
rect 293104 243101 293110 243113
rect 293162 243101 293168 243153
rect 293392 243101 293398 243153
rect 293450 243141 293456 243153
rect 294352 243141 294358 243153
rect 293450 243113 294358 243141
rect 293450 243101 293456 243113
rect 294352 243101 294358 243113
rect 294410 243101 294416 243153
rect 294562 243113 295646 243141
rect 223504 243027 223510 243079
rect 223562 243067 223568 243079
rect 227344 243067 227350 243079
rect 223562 243039 227350 243067
rect 223562 243027 223568 243039
rect 227344 243027 227350 243039
rect 227402 243027 227408 243079
rect 265264 243027 265270 243079
rect 265322 243067 265328 243079
rect 278128 243067 278134 243079
rect 265322 243039 278134 243067
rect 265322 243027 265328 243039
rect 278128 243027 278134 243039
rect 278186 243027 278192 243079
rect 293776 243067 293782 243079
rect 278914 243039 293782 243067
rect 205264 242953 205270 243005
rect 205322 242993 205328 243005
rect 208528 242993 208534 243005
rect 205322 242965 208534 242993
rect 205322 242953 205328 242965
rect 208528 242953 208534 242965
rect 208586 242953 208592 243005
rect 260848 242953 260854 243005
rect 260906 242993 260912 243005
rect 268528 242993 268534 243005
rect 260906 242965 268534 242993
rect 260906 242953 260912 242965
rect 268528 242953 268534 242965
rect 268586 242953 268592 243005
rect 269872 242953 269878 243005
rect 269930 242993 269936 243005
rect 278914 242993 278942 243039
rect 293776 243027 293782 243039
rect 293834 243027 293840 243079
rect 293872 243027 293878 243079
rect 293930 243067 293936 243079
rect 294448 243067 294454 243079
rect 293930 243039 294454 243067
rect 293930 243027 293936 243039
rect 294448 243027 294454 243039
rect 294506 243027 294512 243079
rect 269930 242965 278942 242993
rect 269930 242953 269936 242965
rect 279088 242953 279094 243005
rect 279146 242993 279152 243005
rect 287536 242993 287542 243005
rect 279146 242965 287542 242993
rect 279146 242953 279152 242965
rect 287536 242953 287542 242965
rect 287594 242953 287600 243005
rect 287728 242953 287734 243005
rect 287786 242993 287792 243005
rect 294562 242993 294590 243113
rect 295618 243067 295646 243113
rect 298864 243101 298870 243153
rect 298922 243141 298928 243153
rect 321328 243141 321334 243153
rect 298922 243113 321334 243141
rect 298922 243101 298928 243113
rect 321328 243101 321334 243113
rect 321386 243101 321392 243153
rect 303376 243067 303382 243079
rect 295618 243039 303382 243067
rect 303376 243027 303382 243039
rect 303434 243027 303440 243079
rect 316816 243027 316822 243079
rect 316874 243067 316880 243079
rect 337072 243067 337078 243079
rect 316874 243039 337078 243067
rect 316874 243027 316880 243039
rect 337072 243027 337078 243039
rect 337130 243027 337136 243079
rect 287786 242965 294590 242993
rect 287786 242953 287792 242965
rect 298576 242953 298582 243005
rect 298634 242993 298640 243005
rect 314320 242993 314326 243005
rect 298634 242965 314326 242993
rect 298634 242953 298640 242965
rect 314320 242953 314326 242965
rect 314378 242953 314384 243005
rect 674608 242953 674614 243005
rect 674666 242993 674672 243005
rect 675376 242993 675382 243005
rect 674666 242965 675382 242993
rect 674666 242953 674672 242965
rect 675376 242953 675382 242965
rect 675434 242953 675440 243005
rect 266032 242879 266038 242931
rect 266090 242919 266096 242931
rect 276016 242919 276022 242931
rect 266090 242891 276022 242919
rect 266090 242879 266096 242891
rect 276016 242879 276022 242891
rect 276074 242879 276080 242931
rect 278032 242879 278038 242931
rect 278090 242919 278096 242931
rect 288304 242919 288310 242931
rect 278090 242891 288310 242919
rect 278090 242879 278096 242891
rect 288304 242879 288310 242891
rect 288362 242879 288368 242931
rect 288592 242879 288598 242931
rect 288650 242919 288656 242931
rect 293392 242919 293398 242931
rect 288650 242891 293398 242919
rect 288650 242879 288656 242891
rect 293392 242879 293398 242891
rect 293450 242879 293456 242931
rect 293584 242879 293590 242931
rect 293642 242919 293648 242931
rect 297904 242919 297910 242931
rect 293642 242891 297910 242919
rect 293642 242879 293648 242891
rect 297904 242879 297910 242891
rect 297962 242879 297968 242931
rect 299440 242919 299446 242931
rect 298402 242891 299446 242919
rect 227824 242805 227830 242857
rect 227882 242845 227888 242857
rect 247792 242845 247798 242857
rect 227882 242817 247798 242845
rect 227882 242805 227888 242817
rect 247792 242805 247798 242817
rect 247850 242805 247856 242857
rect 266608 242805 266614 242857
rect 266666 242845 266672 242857
rect 279088 242845 279094 242857
rect 266666 242817 279094 242845
rect 266666 242805 266672 242817
rect 279088 242805 279094 242817
rect 279146 242805 279152 242857
rect 280816 242805 280822 242857
rect 280874 242845 280880 242857
rect 288880 242845 288886 242857
rect 280874 242817 288886 242845
rect 280874 242805 280880 242817
rect 288880 242805 288886 242817
rect 288938 242805 288944 242857
rect 288976 242805 288982 242857
rect 289034 242845 289040 242857
rect 297424 242845 297430 242857
rect 289034 242817 297430 242845
rect 289034 242805 289040 242817
rect 297424 242805 297430 242817
rect 297482 242805 297488 242857
rect 297808 242805 297814 242857
rect 297866 242845 297872 242857
rect 298402 242845 298430 242891
rect 299440 242879 299446 242891
rect 299498 242879 299504 242931
rect 299632 242879 299638 242931
rect 299690 242919 299696 242931
rect 317392 242919 317398 242931
rect 299690 242891 317398 242919
rect 299690 242879 299696 242891
rect 317392 242879 317398 242891
rect 317450 242879 317456 242931
rect 297866 242817 298430 242845
rect 297866 242805 297872 242817
rect 307696 242805 307702 242857
rect 307754 242845 307760 242857
rect 308272 242845 308278 242857
rect 307754 242817 308278 242845
rect 307754 242805 307760 242817
rect 308272 242805 308278 242817
rect 308330 242805 308336 242857
rect 338128 242805 338134 242857
rect 338186 242845 338192 242857
rect 339184 242845 339190 242857
rect 338186 242817 339190 242845
rect 338186 242805 338192 242817
rect 339184 242805 339190 242817
rect 339242 242805 339248 242857
rect 227056 242731 227062 242783
rect 227114 242771 227120 242783
rect 227632 242771 227638 242783
rect 227114 242743 227638 242771
rect 227114 242731 227120 242743
rect 227632 242731 227638 242743
rect 227690 242731 227696 242783
rect 268048 242731 268054 242783
rect 268106 242771 268112 242783
rect 268106 242743 278270 242771
rect 268106 242731 268112 242743
rect 227344 242657 227350 242709
rect 227402 242697 227408 242709
rect 227728 242697 227734 242709
rect 227402 242669 227734 242697
rect 227402 242657 227408 242669
rect 227728 242657 227734 242669
rect 227786 242657 227792 242709
rect 267760 242657 267766 242709
rect 267818 242697 267824 242709
rect 268240 242697 268246 242709
rect 267818 242669 268246 242697
rect 267818 242657 267824 242669
rect 268240 242657 268246 242669
rect 268298 242657 268304 242709
rect 269680 242657 269686 242709
rect 269738 242697 269744 242709
rect 278128 242697 278134 242709
rect 269738 242669 278134 242697
rect 269738 242657 269744 242669
rect 278128 242657 278134 242669
rect 278186 242657 278192 242709
rect 278242 242697 278270 242743
rect 278320 242731 278326 242783
rect 278378 242771 278384 242783
rect 278378 242743 288158 242771
rect 278378 242731 278384 242743
rect 287536 242697 287542 242709
rect 278242 242669 287542 242697
rect 287536 242657 287542 242669
rect 287594 242657 287600 242709
rect 287632 242657 287638 242709
rect 287690 242697 287696 242709
rect 288016 242697 288022 242709
rect 287690 242669 288022 242697
rect 287690 242657 287696 242669
rect 288016 242657 288022 242669
rect 288074 242657 288080 242709
rect 288130 242697 288158 242743
rect 288208 242731 288214 242783
rect 288266 242771 288272 242783
rect 299632 242771 299638 242783
rect 288266 242743 299638 242771
rect 288266 242731 288272 242743
rect 299632 242731 299638 242743
rect 299690 242731 299696 242783
rect 305776 242731 305782 242783
rect 305834 242771 305840 242783
rect 320368 242771 320374 242783
rect 305834 242743 320374 242771
rect 305834 242731 305840 242743
rect 320368 242731 320374 242743
rect 320426 242731 320432 242783
rect 339856 242731 339862 242783
rect 339914 242771 339920 242783
rect 340240 242771 340246 242783
rect 339914 242743 340246 242771
rect 339914 242731 339920 242743
rect 340240 242731 340246 242743
rect 340298 242731 340304 242783
rect 299536 242697 299542 242709
rect 288130 242669 299542 242697
rect 299536 242657 299542 242669
rect 299594 242657 299600 242709
rect 299728 242657 299734 242709
rect 299786 242697 299792 242709
rect 299786 242669 305918 242697
rect 299786 242657 299792 242669
rect 269200 242583 269206 242635
rect 269258 242623 269264 242635
rect 301264 242623 301270 242635
rect 269258 242595 301270 242623
rect 269258 242583 269264 242595
rect 301264 242583 301270 242595
rect 301322 242583 301328 242635
rect 305776 242583 305782 242635
rect 305834 242583 305840 242635
rect 305890 242623 305918 242669
rect 308080 242657 308086 242709
rect 308138 242697 308144 242709
rect 328720 242697 328726 242709
rect 308138 242669 328726 242697
rect 308138 242657 308144 242669
rect 328720 242657 328726 242669
rect 328778 242657 328784 242709
rect 322576 242623 322582 242635
rect 305890 242595 322582 242623
rect 322576 242583 322582 242595
rect 322634 242583 322640 242635
rect 328336 242583 328342 242635
rect 328394 242623 328400 242635
rect 338800 242623 338806 242635
rect 328394 242595 338806 242623
rect 328394 242583 328400 242595
rect 338800 242583 338806 242595
rect 338858 242583 338864 242635
rect 223984 242509 223990 242561
rect 224042 242549 224048 242561
rect 247312 242549 247318 242561
rect 224042 242521 247318 242549
rect 224042 242509 224048 242521
rect 247312 242509 247318 242521
rect 247370 242509 247376 242561
rect 268144 242509 268150 242561
rect 268202 242549 268208 242561
rect 287728 242549 287734 242561
rect 268202 242521 287734 242549
rect 268202 242509 268208 242521
rect 287728 242509 287734 242521
rect 287786 242509 287792 242561
rect 288112 242509 288118 242561
rect 288170 242549 288176 242561
rect 305794 242549 305822 242583
rect 323440 242549 323446 242561
rect 288170 242521 305822 242549
rect 305890 242521 323446 242549
rect 288170 242509 288176 242521
rect 95056 242435 95062 242487
rect 95114 242475 95120 242487
rect 106576 242475 106582 242487
rect 95114 242447 106582 242475
rect 95114 242435 95120 242447
rect 106576 242435 106582 242447
rect 106634 242435 106640 242487
rect 138256 242435 138262 242487
rect 138314 242475 138320 242487
rect 171376 242475 171382 242487
rect 138314 242447 171382 242475
rect 138314 242435 138320 242447
rect 171376 242435 171382 242447
rect 171434 242435 171440 242487
rect 276976 242435 276982 242487
rect 277034 242475 277040 242487
rect 283984 242475 283990 242487
rect 277034 242447 283990 242475
rect 277034 242435 277040 242447
rect 283984 242435 283990 242447
rect 284042 242435 284048 242487
rect 286480 242435 286486 242487
rect 286538 242475 286544 242487
rect 298000 242475 298006 242487
rect 286538 242447 298006 242475
rect 286538 242435 286544 242447
rect 298000 242435 298006 242447
rect 298058 242435 298064 242487
rect 298096 242435 298102 242487
rect 298154 242475 298160 242487
rect 305890 242475 305918 242521
rect 323440 242509 323446 242521
rect 323498 242509 323504 242561
rect 443536 242509 443542 242561
rect 443594 242549 443600 242561
rect 463600 242549 463606 242561
rect 443594 242521 463606 242549
rect 443594 242509 443600 242521
rect 463600 242509 463606 242521
rect 463658 242509 463664 242561
rect 483856 242509 483862 242561
rect 483914 242549 483920 242561
rect 503920 242549 503926 242561
rect 483914 242521 503926 242549
rect 483914 242509 483920 242521
rect 503920 242509 503926 242521
rect 503978 242509 503984 242561
rect 298154 242447 305918 242475
rect 298154 242435 298160 242447
rect 306640 242435 306646 242487
rect 306698 242475 306704 242487
rect 316912 242475 316918 242487
rect 306698 242447 316918 242475
rect 306698 242435 306704 242447
rect 316912 242435 316918 242447
rect 316970 242435 316976 242487
rect 317008 242435 317014 242487
rect 317066 242475 317072 242487
rect 317488 242475 317494 242487
rect 317066 242447 317494 242475
rect 317066 242435 317072 242447
rect 317488 242435 317494 242447
rect 317546 242435 317552 242487
rect 175696 242361 175702 242413
rect 175754 242401 175760 242413
rect 195760 242401 195766 242413
rect 175754 242373 195766 242401
rect 175754 242361 175760 242373
rect 195760 242361 195766 242373
rect 195818 242361 195824 242413
rect 283696 242361 283702 242413
rect 283754 242401 283760 242413
rect 320176 242401 320182 242413
rect 283754 242373 320182 242401
rect 283754 242361 283760 242373
rect 320176 242361 320182 242373
rect 320234 242361 320240 242413
rect 674128 242361 674134 242413
rect 674186 242401 674192 242413
rect 675376 242401 675382 242413
rect 674186 242373 675382 242401
rect 674186 242361 674192 242373
rect 675376 242361 675382 242373
rect 675434 242361 675440 242413
rect 241936 242287 241942 242339
rect 241994 242327 242000 242339
rect 242320 242327 242326 242339
rect 241994 242299 242326 242327
rect 241994 242287 242000 242299
rect 242320 242287 242326 242299
rect 242378 242287 242384 242339
rect 271888 242287 271894 242339
rect 271946 242327 271952 242339
rect 355216 242327 355222 242339
rect 271946 242299 355222 242327
rect 271946 242287 271952 242299
rect 355216 242287 355222 242299
rect 355274 242287 355280 242339
rect 244432 242213 244438 242265
rect 244490 242253 244496 242265
rect 353008 242253 353014 242265
rect 244490 242225 353014 242253
rect 244490 242213 244496 242225
rect 353008 242213 353014 242225
rect 353066 242213 353072 242265
rect 40048 242139 40054 242191
rect 40106 242179 40112 242191
rect 42256 242179 42262 242191
rect 40106 242151 42262 242179
rect 40106 242139 40112 242151
rect 42256 242139 42262 242151
rect 42314 242139 42320 242191
rect 238288 242139 238294 242191
rect 238346 242179 238352 242191
rect 350032 242179 350038 242191
rect 238346 242151 350038 242179
rect 238346 242139 238352 242151
rect 350032 242139 350038 242151
rect 350090 242139 350096 242191
rect 39952 242065 39958 242117
rect 40010 242105 40016 242117
rect 42928 242105 42934 242117
rect 40010 242077 42934 242105
rect 40010 242065 40016 242077
rect 42928 242065 42934 242077
rect 42986 242065 42992 242117
rect 238960 242065 238966 242117
rect 239018 242105 239024 242117
rect 347824 242105 347830 242117
rect 239018 242077 347830 242105
rect 239018 242065 239024 242077
rect 347824 242065 347830 242077
rect 347882 242065 347888 242117
rect 40144 241991 40150 242043
rect 40202 242031 40208 242043
rect 42544 242031 42550 242043
rect 40202 242003 42550 242031
rect 40202 241991 40208 242003
rect 42544 241991 42550 242003
rect 42602 241991 42608 242043
rect 144016 241991 144022 242043
rect 144074 242031 144080 242043
rect 182800 242031 182806 242043
rect 144074 242003 182806 242031
rect 144074 241991 144080 242003
rect 182800 241991 182806 242003
rect 182858 241991 182864 242043
rect 348592 242031 348598 242043
rect 240994 242003 348598 242031
rect 40240 241917 40246 241969
rect 40298 241957 40304 241969
rect 42352 241957 42358 241969
rect 40298 241929 42358 241957
rect 40298 241917 40304 241929
rect 42352 241917 42358 241929
rect 42410 241917 42416 241969
rect 50320 241917 50326 241969
rect 50378 241957 50384 241969
rect 205840 241957 205846 241969
rect 50378 241929 205846 241957
rect 50378 241917 50384 241929
rect 205840 241917 205846 241929
rect 205898 241917 205904 241969
rect 217552 241843 217558 241895
rect 217610 241883 217616 241895
rect 234448 241883 234454 241895
rect 217610 241855 234454 241883
rect 217610 241843 217616 241855
rect 234448 241843 234454 241855
rect 234506 241843 234512 241895
rect 234544 241843 234550 241895
rect 234602 241883 234608 241895
rect 240994 241883 241022 242003
rect 348592 241991 348598 242003
rect 348650 241991 348656 242043
rect 351760 241957 351766 241969
rect 244354 241929 351766 241957
rect 234602 241855 241022 241883
rect 234602 241843 234608 241855
rect 241072 241843 241078 241895
rect 241130 241883 241136 241895
rect 244354 241883 244382 241929
rect 351760 241917 351766 241929
rect 351818 241917 351824 241969
rect 412048 241917 412054 241969
rect 412106 241957 412112 241969
rect 412240 241957 412246 241969
rect 412106 241929 412246 241957
rect 412106 241917 412112 241929
rect 412240 241917 412246 241929
rect 412298 241917 412304 241969
rect 607696 241957 607702 241969
rect 604834 241929 607702 241957
rect 241130 241855 244382 241883
rect 241130 241843 241136 241855
rect 251824 241843 251830 241895
rect 251882 241883 251888 241895
rect 251882 241855 273086 241883
rect 251882 241843 251888 241855
rect 215440 241769 215446 241821
rect 215498 241809 215504 241821
rect 221392 241809 221398 241821
rect 215498 241781 221398 241809
rect 215498 241769 215504 241781
rect 221392 241769 221398 241781
rect 221450 241769 221456 241821
rect 233488 241769 233494 241821
rect 233546 241809 233552 241821
rect 238960 241809 238966 241821
rect 233546 241781 238966 241809
rect 233546 241769 233552 241781
rect 238960 241769 238966 241781
rect 239018 241769 239024 241821
rect 264304 241769 264310 241821
rect 264362 241809 264368 241821
rect 271984 241809 271990 241821
rect 264362 241781 271990 241809
rect 264362 241769 264368 241781
rect 271984 241769 271990 241781
rect 272042 241769 272048 241821
rect 273058 241809 273086 241855
rect 273136 241843 273142 241895
rect 273194 241883 273200 241895
rect 283888 241883 283894 241895
rect 273194 241855 283894 241883
rect 273194 241843 273200 241855
rect 283888 241843 283894 241855
rect 283946 241843 283952 241895
rect 283984 241843 283990 241895
rect 284042 241883 284048 241895
rect 288592 241883 288598 241895
rect 284042 241855 288598 241883
rect 284042 241843 284048 241855
rect 288592 241843 288598 241855
rect 288650 241843 288656 241895
rect 288688 241843 288694 241895
rect 288746 241883 288752 241895
rect 307888 241883 307894 241895
rect 288746 241855 307894 241883
rect 288746 241843 288752 241855
rect 307888 241843 307894 241855
rect 307946 241843 307952 241895
rect 311728 241843 311734 241895
rect 311786 241883 311792 241895
rect 325168 241883 325174 241895
rect 311786 241855 325174 241883
rect 311786 241843 311792 241855
rect 325168 241843 325174 241855
rect 325226 241843 325232 241895
rect 325264 241843 325270 241895
rect 325322 241883 325328 241895
rect 374416 241883 374422 241895
rect 325322 241855 374422 241883
rect 325322 241843 325328 241855
rect 374416 241843 374422 241855
rect 374474 241843 374480 241895
rect 376048 241843 376054 241895
rect 376106 241883 376112 241895
rect 403216 241883 403222 241895
rect 376106 241855 403222 241883
rect 376106 241843 376112 241855
rect 403216 241843 403222 241855
rect 403274 241843 403280 241895
rect 602896 241843 602902 241895
rect 602954 241883 602960 241895
rect 604834 241883 604862 241929
rect 607696 241917 607702 241929
rect 607754 241917 607760 241969
rect 602954 241855 604862 241883
rect 602954 241843 602960 241855
rect 273616 241809 273622 241821
rect 273058 241781 273622 241809
rect 273616 241769 273622 241781
rect 273674 241769 273680 241821
rect 278224 241769 278230 241821
rect 278282 241809 278288 241821
rect 327952 241809 327958 241821
rect 278282 241781 327958 241809
rect 278282 241769 278288 241781
rect 327952 241769 327958 241781
rect 328010 241769 328016 241821
rect 329296 241769 329302 241821
rect 329354 241809 329360 241821
rect 354544 241809 354550 241821
rect 329354 241781 354550 241809
rect 329354 241769 329360 241781
rect 354544 241769 354550 241781
rect 354602 241769 354608 241821
rect 360592 241769 360598 241821
rect 360650 241809 360656 241821
rect 378640 241809 378646 241821
rect 360650 241781 378646 241809
rect 360650 241769 360656 241781
rect 378640 241769 378646 241781
rect 378698 241769 378704 241821
rect 378736 241769 378742 241821
rect 378794 241809 378800 241821
rect 396400 241809 396406 241821
rect 378794 241781 396406 241809
rect 378794 241769 378800 241781
rect 396400 241769 396406 241781
rect 396458 241769 396464 241821
rect 218704 241695 218710 241747
rect 218762 241735 218768 241747
rect 234352 241735 234358 241747
rect 218762 241707 234358 241735
rect 218762 241695 218768 241707
rect 234352 241695 234358 241707
rect 234410 241695 234416 241747
rect 237424 241695 237430 241747
rect 237482 241735 237488 241747
rect 262192 241735 262198 241747
rect 237482 241707 262198 241735
rect 237482 241695 237488 241707
rect 262192 241695 262198 241707
rect 262250 241695 262256 241747
rect 277648 241695 277654 241747
rect 277706 241735 277712 241747
rect 329968 241735 329974 241747
rect 277706 241707 329974 241735
rect 277706 241695 277712 241707
rect 329968 241695 329974 241707
rect 330026 241695 330032 241747
rect 331024 241695 331030 241747
rect 331082 241735 331088 241747
rect 358288 241735 358294 241747
rect 331082 241707 358294 241735
rect 331082 241695 331088 241707
rect 358288 241695 358294 241707
rect 358346 241695 358352 241747
rect 363184 241695 363190 241747
rect 363242 241735 363248 241747
rect 400144 241735 400150 241747
rect 363242 241707 400150 241735
rect 363242 241695 363248 241707
rect 400144 241695 400150 241707
rect 400202 241695 400208 241747
rect 219280 241621 219286 241673
rect 219338 241661 219344 241673
rect 233776 241661 233782 241673
rect 219338 241633 233782 241661
rect 219338 241621 219344 241633
rect 233776 241621 233782 241633
rect 233834 241621 233840 241673
rect 252784 241621 252790 241673
rect 252842 241661 252848 241673
rect 311728 241661 311734 241673
rect 252842 241633 311734 241661
rect 252842 241621 252848 241633
rect 311728 241621 311734 241633
rect 311786 241621 311792 241673
rect 336496 241661 336502 241673
rect 317410 241633 336502 241661
rect 213904 241547 213910 241599
rect 213962 241587 213968 241599
rect 229168 241587 229174 241599
rect 213962 241559 229174 241587
rect 213962 241547 213968 241559
rect 229168 241547 229174 241559
rect 229226 241547 229232 241599
rect 269296 241547 269302 241599
rect 269354 241587 269360 241599
rect 311632 241587 311638 241599
rect 269354 241559 311638 241587
rect 269354 241547 269360 241559
rect 311632 241547 311638 241559
rect 311690 241547 311696 241599
rect 222544 241473 222550 241525
rect 222602 241513 222608 241525
rect 232528 241513 232534 241525
rect 222602 241485 232534 241513
rect 222602 241473 222608 241485
rect 232528 241473 232534 241485
rect 232586 241473 232592 241525
rect 254992 241473 254998 241525
rect 255050 241513 255056 241525
rect 317410 241513 317438 241633
rect 336496 241621 336502 241633
rect 336554 241621 336560 241673
rect 361552 241621 361558 241673
rect 361610 241661 361616 241673
rect 361610 241633 378590 241661
rect 361610 241621 361616 241633
rect 317872 241547 317878 241599
rect 317930 241587 317936 241599
rect 330160 241587 330166 241599
rect 317930 241559 330166 241587
rect 317930 241547 317936 241559
rect 330160 241547 330166 241559
rect 330218 241547 330224 241599
rect 330256 241547 330262 241599
rect 330314 241587 330320 241599
rect 355696 241587 355702 241599
rect 330314 241559 355702 241587
rect 330314 241547 330320 241559
rect 355696 241547 355702 241559
rect 355754 241547 355760 241599
rect 378562 241587 378590 241633
rect 378640 241621 378646 241673
rect 378698 241661 378704 241673
rect 394096 241661 394102 241673
rect 378698 241633 394102 241661
rect 378698 241621 378704 241633
rect 394096 241621 394102 241633
rect 394154 241621 394160 241673
rect 378736 241587 378742 241599
rect 378562 241559 378742 241587
rect 378736 241547 378742 241559
rect 378794 241547 378800 241599
rect 674992 241547 674998 241599
rect 675050 241587 675056 241599
rect 675472 241587 675478 241599
rect 675050 241559 675478 241587
rect 675050 241547 675056 241559
rect 675472 241547 675478 241559
rect 675530 241547 675536 241599
rect 255050 241485 317438 241513
rect 255050 241473 255056 241485
rect 317488 241473 317494 241525
rect 317546 241513 317552 241525
rect 326896 241513 326902 241525
rect 317546 241485 326902 241513
rect 317546 241473 317552 241485
rect 326896 241473 326902 241485
rect 326954 241473 326960 241525
rect 327184 241473 327190 241525
rect 327242 241513 327248 241525
rect 336112 241513 336118 241525
rect 327242 241485 336118 241513
rect 327242 241473 327248 241485
rect 336112 241473 336118 241485
rect 336170 241473 336176 241525
rect 363760 241473 363766 241525
rect 363818 241513 363824 241525
rect 400720 241513 400726 241525
rect 363818 241485 400726 241513
rect 363818 241473 363824 241485
rect 400720 241473 400726 241485
rect 400778 241473 400784 241525
rect 239152 241399 239158 241451
rect 239210 241439 239216 241451
rect 258544 241439 258550 241451
rect 239210 241411 258550 241439
rect 239210 241399 239216 241411
rect 258544 241399 258550 241411
rect 258602 241399 258608 241451
rect 274096 241399 274102 241451
rect 274154 241439 274160 241451
rect 318256 241439 318262 241451
rect 274154 241411 318262 241439
rect 274154 241399 274160 241411
rect 318256 241399 318262 241411
rect 318314 241399 318320 241451
rect 320464 241399 320470 241451
rect 320522 241439 320528 241451
rect 326992 241439 326998 241451
rect 320522 241411 326998 241439
rect 320522 241399 320528 241411
rect 326992 241399 326998 241411
rect 327050 241399 327056 241451
rect 331504 241399 331510 241451
rect 331562 241439 331568 241451
rect 359344 241439 359350 241451
rect 331562 241411 359350 241439
rect 331562 241399 331568 241411
rect 359344 241399 359350 241411
rect 359402 241399 359408 241451
rect 362320 241399 362326 241451
rect 362378 241439 362384 241451
rect 398416 241439 398422 241451
rect 362378 241411 398422 241439
rect 362378 241399 362384 241411
rect 398416 241399 398422 241411
rect 398474 241399 398480 241451
rect 255952 241325 255958 241377
rect 256010 241365 256016 241377
rect 256010 241337 318206 241365
rect 256010 241325 256016 241337
rect 244720 241251 244726 241303
rect 244778 241291 244784 241303
rect 317488 241291 317494 241303
rect 244778 241263 317494 241291
rect 244778 241251 244784 241263
rect 317488 241251 317494 241263
rect 317546 241251 317552 241303
rect 318178 241291 318206 241337
rect 326704 241325 326710 241377
rect 326762 241365 326768 241377
rect 328912 241365 328918 241377
rect 326762 241337 328918 241365
rect 326762 241325 326768 241337
rect 328912 241325 328918 241337
rect 328970 241325 328976 241377
rect 332272 241325 332278 241377
rect 332330 241365 332336 241377
rect 361072 241365 361078 241377
rect 332330 241337 361078 241365
rect 332330 241325 332336 241337
rect 361072 241325 361078 241337
rect 361130 241325 361136 241377
rect 364144 241325 364150 241377
rect 364202 241365 364208 241377
rect 401872 241365 401878 241377
rect 364202 241337 401878 241365
rect 364202 241325 364208 241337
rect 401872 241325 401878 241337
rect 401930 241325 401936 241377
rect 334480 241291 334486 241303
rect 318178 241263 334486 241291
rect 334480 241251 334486 241263
rect 334538 241251 334544 241303
rect 361936 241251 361942 241303
rect 361994 241291 362000 241303
rect 397456 241291 397462 241303
rect 361994 241263 397462 241291
rect 361994 241251 362000 241263
rect 397456 241251 397462 241263
rect 397514 241251 397520 241303
rect 226288 241177 226294 241229
rect 226346 241217 226352 241229
rect 230704 241217 230710 241229
rect 226346 241189 230710 241217
rect 226346 241177 226352 241189
rect 230704 241177 230710 241189
rect 230762 241177 230768 241229
rect 253744 241177 253750 241229
rect 253802 241217 253808 241229
rect 339376 241217 339382 241229
rect 253802 241189 339382 241217
rect 253802 241177 253808 241189
rect 339376 241177 339382 241189
rect 339434 241177 339440 241229
rect 362416 241177 362422 241229
rect 362474 241217 362480 241229
rect 398992 241217 398998 241229
rect 362474 241189 398998 241217
rect 362474 241177 362480 241189
rect 398992 241177 398998 241189
rect 399050 241177 399056 241229
rect 216688 241103 216694 241155
rect 216746 241143 216752 241155
rect 238384 241143 238390 241155
rect 216746 241115 238390 241143
rect 216746 241103 216752 241115
rect 238384 241103 238390 241115
rect 238442 241103 238448 241155
rect 254224 241103 254230 241155
rect 254282 241143 254288 241155
rect 337840 241143 337846 241155
rect 254282 241115 337846 241143
rect 254282 241103 254288 241115
rect 337840 241103 337846 241115
rect 337898 241103 337904 241155
rect 339664 241103 339670 241155
rect 339722 241143 339728 241155
rect 360496 241143 360502 241155
rect 339722 241115 360502 241143
rect 339722 241103 339728 241115
rect 360496 241103 360502 241115
rect 360554 241103 360560 241155
rect 364528 241103 364534 241155
rect 364586 241143 364592 241155
rect 402736 241143 402742 241155
rect 364586 241115 402742 241143
rect 364586 241103 364592 241115
rect 402736 241103 402742 241115
rect 402794 241103 402800 241155
rect 221488 241029 221494 241081
rect 221546 241069 221552 241081
rect 232912 241069 232918 241081
rect 221546 241041 232918 241069
rect 221546 241029 221552 241041
rect 232912 241029 232918 241041
rect 232970 241029 232976 241081
rect 237520 241029 237526 241081
rect 237578 241069 237584 241081
rect 254608 241069 254614 241081
rect 237578 241041 254614 241069
rect 237578 241029 237584 241041
rect 254608 241029 254614 241041
rect 254666 241029 254672 241081
rect 274480 241029 274486 241081
rect 274538 241069 274544 241081
rect 287632 241069 287638 241081
rect 274538 241041 287638 241069
rect 274538 241029 274544 241041
rect 287632 241029 287638 241041
rect 287690 241029 287696 241081
rect 288304 241029 288310 241081
rect 288362 241069 288368 241081
rect 290032 241069 290038 241081
rect 288362 241041 290038 241069
rect 288362 241029 288368 241041
rect 290032 241029 290038 241041
rect 290090 241029 290096 241081
rect 291952 241029 291958 241081
rect 292010 241069 292016 241081
rect 376144 241069 376150 241081
rect 292010 241041 376150 241069
rect 292010 241029 292016 241041
rect 376144 241029 376150 241041
rect 376202 241029 376208 241081
rect 379216 241029 379222 241081
rect 379274 241069 379280 241081
rect 409264 241069 409270 241081
rect 379274 241041 409270 241069
rect 379274 241029 379280 241041
rect 409264 241029 409270 241041
rect 409322 241029 409328 241081
rect 225232 240955 225238 241007
rect 225290 240995 225296 241007
rect 231184 240995 231190 241007
rect 225290 240967 231190 240995
rect 225290 240955 225296 240967
rect 231184 240955 231190 240967
rect 231242 240955 231248 241007
rect 257680 240955 257686 241007
rect 257738 240995 257744 241007
rect 327856 240995 327862 241007
rect 257738 240967 327862 240995
rect 257738 240955 257744 240967
rect 327856 240955 327862 240967
rect 327914 240955 327920 241007
rect 327952 240955 327958 241007
rect 328010 240995 328016 241007
rect 329584 240995 329590 241007
rect 328010 240967 329590 240995
rect 328010 240955 328016 240967
rect 329584 240955 329590 240967
rect 329642 240955 329648 241007
rect 330736 240955 330742 241007
rect 330794 240995 330800 241007
rect 333616 240995 333622 241007
rect 330794 240967 333622 240995
rect 330794 240955 330800 240967
rect 333616 240955 333622 240967
rect 333674 240955 333680 241007
rect 333712 240955 333718 241007
rect 333770 240995 333776 241007
rect 364336 240995 364342 241007
rect 333770 240967 364342 240995
rect 333770 240955 333776 240967
rect 364336 240955 364342 240967
rect 364394 240955 364400 241007
rect 366352 240955 366358 241007
rect 366410 240995 366416 241007
rect 407152 240995 407158 241007
rect 366410 240967 407158 240995
rect 366410 240955 366416 240967
rect 407152 240955 407158 240967
rect 407210 240955 407216 241007
rect 225424 240881 225430 240933
rect 225482 240921 225488 240933
rect 230896 240921 230902 240933
rect 225482 240893 230902 240921
rect 225482 240881 225488 240893
rect 230896 240881 230902 240893
rect 230954 240881 230960 240933
rect 250672 240921 250678 240933
rect 237586 240893 250678 240921
rect 212752 240807 212758 240859
rect 212810 240847 212816 240859
rect 233296 240847 233302 240859
rect 212810 240819 233302 240847
rect 212810 240807 212816 240819
rect 233296 240807 233302 240819
rect 233354 240807 233360 240859
rect 224080 240733 224086 240785
rect 224138 240773 224144 240785
rect 231568 240773 231574 240785
rect 224138 240745 231574 240773
rect 224138 240733 224144 240745
rect 231568 240733 231574 240745
rect 231626 240733 231632 240785
rect 219280 240659 219286 240711
rect 219338 240699 219344 240711
rect 237586 240699 237614 240893
rect 250672 240881 250678 240893
rect 250730 240881 250736 240933
rect 252304 240881 252310 240933
rect 252362 240921 252368 240933
rect 342640 240921 342646 240933
rect 252362 240893 342646 240921
rect 252362 240881 252368 240893
rect 342640 240881 342646 240893
rect 342698 240881 342704 240933
rect 365008 240881 365014 240933
rect 365066 240921 365072 240933
rect 404464 240921 404470 240933
rect 365066 240893 404470 240921
rect 365066 240881 365072 240893
rect 404464 240881 404470 240893
rect 404522 240881 404528 240933
rect 237808 240807 237814 240859
rect 237866 240847 237872 240859
rect 252880 240847 252886 240859
rect 237866 240819 252886 240847
rect 237866 240807 237872 240819
rect 252880 240807 252886 240819
rect 252938 240807 252944 240859
rect 344176 240847 344182 240859
rect 252994 240819 344182 240847
rect 237712 240733 237718 240785
rect 237770 240773 237776 240785
rect 252016 240773 252022 240785
rect 237770 240745 252022 240773
rect 237770 240733 237776 240745
rect 252016 240733 252022 240745
rect 252074 240733 252080 240785
rect 219338 240671 237614 240699
rect 219338 240659 219344 240671
rect 240304 240659 240310 240711
rect 240362 240699 240368 240711
rect 244144 240699 244150 240711
rect 240362 240671 244150 240699
rect 240362 240659 240368 240671
rect 244144 240659 244150 240671
rect 244202 240659 244208 240711
rect 251536 240659 251542 240711
rect 251594 240699 251600 240711
rect 252994 240699 253022 240819
rect 344176 240807 344182 240819
rect 344234 240807 344240 240859
rect 367216 240807 367222 240859
rect 367274 240847 367280 240859
rect 408880 240847 408886 240859
rect 367274 240819 408886 240847
rect 367274 240807 367280 240819
rect 408880 240807 408886 240819
rect 408938 240807 408944 240859
rect 255472 240733 255478 240785
rect 255530 240773 255536 240785
rect 263344 240773 263350 240785
rect 255530 240745 263350 240773
rect 255530 240733 255536 240745
rect 263344 240733 263350 240745
rect 263402 240733 263408 240785
rect 271024 240733 271030 240785
rect 271082 240773 271088 240785
rect 281392 240773 281398 240785
rect 271082 240745 281398 240773
rect 271082 240733 271088 240745
rect 281392 240733 281398 240745
rect 281450 240733 281456 240785
rect 282256 240733 282262 240785
rect 282314 240773 282320 240785
rect 375760 240773 375766 240785
rect 282314 240745 375766 240773
rect 282314 240733 282320 240745
rect 375760 240733 375766 240745
rect 375818 240733 375824 240785
rect 379600 240733 379606 240785
rect 379658 240773 379664 240785
rect 409936 240773 409942 240785
rect 379658 240745 409942 240773
rect 379658 240733 379664 240745
rect 409936 240733 409942 240745
rect 409994 240733 410000 240785
rect 345712 240699 345718 240711
rect 251594 240671 253022 240699
rect 253090 240671 345718 240699
rect 251594 240659 251600 240671
rect 41776 240585 41782 240637
rect 41834 240585 41840 240637
rect 220240 240585 220246 240637
rect 220298 240625 220304 240637
rect 248656 240625 248662 240637
rect 220298 240597 248662 240625
rect 220298 240585 220304 240597
rect 248656 240585 248662 240597
rect 248714 240585 248720 240637
rect 250576 240585 250582 240637
rect 250634 240625 250640 240637
rect 253090 240625 253118 240671
rect 345712 240659 345718 240671
rect 345770 240659 345776 240711
rect 364624 240659 364630 240711
rect 364682 240699 364688 240711
rect 403408 240699 403414 240711
rect 364682 240671 403414 240699
rect 364682 240659 364688 240671
rect 403408 240659 403414 240671
rect 403466 240659 403472 240711
rect 250634 240597 253118 240625
rect 250634 240585 250640 240597
rect 257872 240585 257878 240637
rect 257930 240625 257936 240637
rect 348304 240625 348310 240637
rect 257930 240597 348310 240625
rect 257930 240585 257936 240597
rect 348304 240585 348310 240597
rect 348362 240585 348368 240637
rect 365392 240585 365398 240637
rect 365450 240625 365456 240637
rect 405136 240625 405142 240637
rect 365450 240597 405142 240625
rect 365450 240585 365456 240597
rect 405136 240585 405142 240597
rect 405194 240585 405200 240637
rect 41794 240415 41822 240585
rect 219664 240511 219670 240563
rect 219722 240551 219728 240563
rect 249808 240551 249814 240563
rect 219722 240523 249814 240551
rect 219722 240511 219728 240523
rect 249808 240511 249814 240523
rect 249866 240511 249872 240563
rect 250192 240511 250198 240563
rect 250250 240551 250256 240563
rect 346288 240551 346294 240563
rect 250250 240523 346294 240551
rect 250250 240511 250256 240523
rect 346288 240511 346294 240523
rect 346346 240511 346352 240563
rect 365968 240511 365974 240563
rect 366026 240551 366032 240563
rect 406096 240551 406102 240563
rect 366026 240523 406102 240551
rect 366026 240511 366032 240523
rect 406096 240511 406102 240523
rect 406154 240511 406160 240563
rect 674704 240511 674710 240563
rect 674762 240551 674768 240563
rect 675472 240551 675478 240563
rect 674762 240523 675478 240551
rect 674762 240511 674768 240523
rect 675472 240511 675478 240523
rect 675530 240511 675536 240563
rect 220432 240437 220438 240489
rect 220490 240477 220496 240489
rect 233392 240477 233398 240489
rect 220490 240449 233398 240477
rect 220490 240437 220496 240449
rect 233392 240437 233398 240449
rect 233450 240437 233456 240489
rect 248080 240477 248086 240489
rect 237586 240449 248086 240477
rect 41776 240363 41782 240415
rect 41834 240363 41840 240415
rect 220624 240363 220630 240415
rect 220682 240403 220688 240415
rect 237586 240403 237614 240449
rect 248080 240437 248086 240449
rect 248138 240437 248144 240489
rect 248368 240437 248374 240489
rect 248426 240477 248432 240489
rect 350224 240477 350230 240489
rect 248426 240449 350230 240477
rect 248426 240437 248432 240449
rect 350224 240437 350230 240449
rect 350282 240437 350288 240489
rect 366736 240437 366742 240489
rect 366794 240477 366800 240489
rect 407824 240477 407830 240489
rect 366794 240449 407830 240477
rect 366794 240437 366800 240449
rect 407824 240437 407830 240449
rect 407882 240437 407888 240489
rect 607600 240437 607606 240489
rect 607658 240477 607664 240489
rect 627760 240477 627766 240489
rect 607658 240449 627766 240477
rect 607658 240437 607664 240449
rect 627760 240437 627766 240449
rect 627818 240437 627824 240489
rect 220682 240375 237614 240403
rect 220682 240363 220688 240375
rect 240880 240363 240886 240415
rect 240938 240403 240944 240415
rect 257680 240403 257686 240415
rect 240938 240375 257686 240403
rect 240938 240363 240944 240375
rect 257680 240363 257686 240375
rect 257738 240363 257744 240415
rect 275344 240363 275350 240415
rect 275402 240403 275408 240415
rect 281104 240403 281110 240415
rect 275402 240375 281110 240403
rect 275402 240363 275408 240375
rect 281104 240363 281110 240375
rect 281162 240363 281168 240415
rect 281392 240363 281398 240415
rect 281450 240403 281456 240415
rect 281450 240375 286238 240403
rect 281450 240363 281456 240375
rect 218800 240289 218806 240341
rect 218858 240329 218864 240341
rect 237712 240329 237718 240341
rect 218858 240301 237718 240329
rect 218858 240289 218864 240301
rect 237712 240289 237718 240301
rect 237770 240289 237776 240341
rect 238960 240289 238966 240341
rect 239018 240329 239024 240341
rect 255472 240329 255478 240341
rect 239018 240301 255478 240329
rect 239018 240289 239024 240301
rect 255472 240289 255478 240301
rect 255530 240289 255536 240341
rect 264400 240329 264406 240341
rect 256162 240301 264406 240329
rect 236560 240215 236566 240267
rect 236618 240255 236624 240267
rect 236618 240227 237950 240255
rect 236618 240215 236624 240227
rect 218416 240141 218422 240193
rect 218474 240181 218480 240193
rect 237808 240181 237814 240193
rect 218474 240153 237814 240181
rect 218474 240141 218480 240153
rect 237808 240141 237814 240153
rect 237866 240141 237872 240193
rect 237922 240181 237950 240227
rect 238864 240215 238870 240267
rect 238922 240255 238928 240267
rect 256162 240255 256190 240301
rect 264400 240289 264406 240301
rect 264458 240289 264464 240341
rect 274000 240289 274006 240341
rect 274058 240329 274064 240341
rect 274058 240301 286142 240329
rect 274058 240289 274064 240301
rect 238922 240227 256190 240255
rect 238922 240215 238928 240227
rect 262000 240215 262006 240267
rect 262058 240255 262064 240267
rect 278224 240255 278230 240267
rect 262058 240227 278230 240255
rect 262058 240215 262064 240227
rect 278224 240215 278230 240227
rect 278282 240215 278288 240267
rect 285616 240255 285622 240267
rect 278338 240227 285622 240255
rect 263920 240181 263926 240193
rect 237922 240153 263926 240181
rect 263920 240141 263926 240153
rect 263978 240141 263984 240193
rect 264016 240141 264022 240193
rect 264074 240181 264080 240193
rect 277648 240181 277654 240193
rect 264074 240153 277654 240181
rect 264074 240141 264080 240153
rect 277648 240141 277654 240153
rect 277706 240141 277712 240193
rect 277744 240141 277750 240193
rect 277802 240181 277808 240193
rect 278338 240181 278366 240227
rect 285616 240215 285622 240227
rect 285674 240215 285680 240267
rect 277802 240153 278366 240181
rect 277802 240141 277808 240153
rect 279472 240141 279478 240193
rect 279530 240181 279536 240193
rect 282160 240181 282166 240193
rect 279530 240153 282166 240181
rect 279530 240141 279536 240153
rect 282160 240141 282166 240153
rect 282218 240141 282224 240193
rect 286114 240181 286142 240301
rect 286210 240255 286238 240375
rect 286864 240363 286870 240415
rect 286922 240403 286928 240415
rect 286922 240375 305054 240403
rect 286922 240363 286928 240375
rect 297040 240329 297046 240341
rect 287266 240301 297046 240329
rect 287266 240255 287294 240301
rect 297040 240289 297046 240301
rect 297098 240289 297104 240341
rect 305026 240329 305054 240375
rect 315568 240363 315574 240415
rect 315626 240403 315632 240415
rect 375088 240403 375094 240415
rect 315626 240375 375094 240403
rect 315626 240363 315632 240375
rect 375088 240363 375094 240375
rect 375146 240363 375152 240415
rect 378256 240363 378262 240415
rect 378314 240403 378320 240415
rect 408304 240403 408310 240415
rect 378314 240375 408310 240403
rect 378314 240363 378320 240375
rect 408304 240363 408310 240375
rect 408362 240363 408368 240415
rect 313168 240329 313174 240341
rect 305026 240301 313174 240329
rect 313168 240289 313174 240301
rect 313226 240289 313232 240341
rect 313648 240289 313654 240341
rect 313706 240329 313712 240341
rect 371824 240329 371830 240341
rect 313706 240301 371830 240329
rect 313706 240289 313712 240301
rect 371824 240289 371830 240301
rect 371882 240289 371888 240341
rect 377776 240289 377782 240341
rect 377834 240329 377840 240341
rect 406672 240329 406678 240341
rect 377834 240301 406678 240329
rect 377834 240289 377840 240301
rect 406672 240289 406678 240301
rect 406730 240289 406736 240341
rect 286210 240227 287294 240255
rect 287440 240215 287446 240267
rect 287498 240255 287504 240267
rect 287824 240255 287830 240267
rect 287498 240227 287830 240255
rect 287498 240215 287504 240227
rect 287824 240215 287830 240227
rect 287882 240215 287888 240267
rect 287920 240215 287926 240267
rect 287978 240255 287984 240267
rect 312592 240255 312598 240267
rect 287978 240227 312598 240255
rect 287978 240215 287984 240227
rect 312592 240215 312598 240227
rect 312650 240215 312656 240267
rect 314608 240215 314614 240267
rect 314666 240255 314672 240267
rect 373552 240255 373558 240267
rect 314666 240227 373558 240255
rect 314666 240215 314672 240227
rect 373552 240215 373558 240227
rect 373610 240215 373616 240267
rect 377200 240215 377206 240267
rect 377258 240255 377264 240267
rect 405520 240255 405526 240267
rect 377258 240227 405526 240255
rect 377258 240215 377264 240227
rect 405520 240215 405526 240227
rect 405578 240215 405584 240267
rect 290704 240181 290710 240193
rect 286114 240153 290710 240181
rect 290704 240141 290710 240153
rect 290762 240141 290768 240193
rect 290800 240141 290806 240193
rect 290858 240181 290864 240193
rect 295408 240181 295414 240193
rect 290858 240153 295414 240181
rect 290858 240141 290864 240153
rect 295408 240141 295414 240153
rect 295466 240141 295472 240193
rect 298192 240141 298198 240193
rect 298250 240181 298256 240193
rect 316048 240181 316054 240193
rect 298250 240153 316054 240181
rect 298250 240141 298256 240153
rect 316048 240141 316054 240153
rect 316106 240141 316112 240193
rect 316144 240141 316150 240193
rect 316202 240181 316208 240193
rect 371344 240181 371350 240193
rect 316202 240153 371350 240181
rect 316202 240141 316208 240153
rect 371344 240141 371350 240153
rect 371402 240141 371408 240193
rect 376432 240141 376438 240193
rect 376490 240181 376496 240193
rect 404080 240181 404086 240193
rect 376490 240153 404086 240181
rect 376490 240141 376496 240153
rect 404080 240141 404086 240153
rect 404138 240141 404144 240193
rect 221776 240067 221782 240119
rect 221834 240107 221840 240119
rect 237520 240107 237526 240119
rect 221834 240079 237526 240107
rect 221834 240067 221840 240079
rect 237520 240067 237526 240079
rect 237578 240067 237584 240119
rect 237904 240067 237910 240119
rect 237962 240107 237968 240119
rect 261616 240107 261622 240119
rect 237962 240079 261622 240107
rect 237962 240067 237968 240079
rect 261616 240067 261622 240079
rect 261674 240067 261680 240119
rect 277456 240067 277462 240119
rect 277514 240107 277520 240119
rect 277514 240079 287582 240107
rect 277514 240067 277520 240079
rect 232336 239993 232342 240045
rect 232394 240033 232400 240045
rect 238192 240033 238198 240045
rect 232394 240005 238198 240033
rect 232394 239993 232400 240005
rect 238192 239993 238198 240005
rect 238250 239993 238256 240045
rect 238288 239993 238294 240045
rect 238346 240033 238352 240045
rect 260656 240033 260662 240045
rect 238346 240005 260662 240033
rect 238346 239993 238352 240005
rect 260656 239993 260662 240005
rect 260714 239993 260720 240045
rect 260752 239993 260758 240045
rect 260810 240033 260816 240045
rect 271888 240033 271894 240045
rect 260810 240005 271894 240033
rect 260810 239993 260816 240005
rect 271888 239993 271894 240005
rect 271946 239993 271952 240045
rect 274672 239993 274678 240045
rect 274730 240033 274736 240045
rect 287344 240033 287350 240045
rect 274730 240005 287350 240033
rect 274730 239993 274736 240005
rect 287344 239993 287350 240005
rect 287402 239993 287408 240045
rect 223216 239919 223222 239971
rect 223274 239959 223280 239971
rect 232144 239959 232150 239971
rect 223274 239931 232150 239959
rect 223274 239919 223280 239931
rect 232144 239919 232150 239931
rect 232202 239919 232208 239971
rect 244624 239919 244630 239971
rect 244682 239959 244688 239971
rect 246064 239959 246070 239971
rect 244682 239931 246070 239959
rect 244682 239919 244688 239931
rect 246064 239919 246070 239931
rect 246122 239919 246128 239971
rect 249712 239919 249718 239971
rect 249770 239959 249776 239971
rect 257872 239959 257878 239971
rect 249770 239931 257878 239959
rect 249770 239919 249776 239931
rect 257872 239919 257878 239931
rect 257930 239919 257936 239971
rect 268720 239919 268726 239971
rect 268778 239959 268784 239971
rect 280144 239959 280150 239971
rect 268778 239931 280150 239959
rect 268778 239919 268784 239931
rect 280144 239919 280150 239931
rect 280202 239919 280208 239971
rect 280240 239919 280246 239971
rect 280298 239959 280304 239971
rect 287554 239959 287582 240079
rect 287824 240067 287830 240119
rect 287882 240107 287888 240119
rect 306640 240107 306646 240119
rect 287882 240079 306646 240107
rect 287882 240067 287888 240079
rect 306640 240067 306646 240079
rect 306698 240067 306704 240119
rect 314224 240067 314230 240119
rect 314282 240107 314288 240119
rect 372400 240107 372406 240119
rect 314282 240079 372406 240107
rect 314282 240067 314288 240079
rect 372400 240067 372406 240079
rect 372458 240067 372464 240119
rect 377008 240067 377014 240119
rect 377066 240107 377072 240119
rect 404944 240107 404950 240119
rect 377066 240079 404950 240107
rect 377066 240067 377072 240079
rect 404944 240067 404950 240079
rect 405002 240067 405008 240119
rect 287632 239993 287638 240045
rect 287690 240033 287696 240045
rect 289456 240033 289462 240045
rect 287690 240005 289462 240033
rect 287690 239993 287696 240005
rect 289456 239993 289462 240005
rect 289514 239993 289520 240045
rect 290512 239993 290518 240045
rect 290570 240033 290576 240045
rect 293392 240033 293398 240045
rect 290570 240005 293398 240033
rect 290570 239993 290576 240005
rect 293392 239993 293398 240005
rect 293450 239993 293456 240045
rect 295696 239993 295702 240045
rect 295754 240033 295760 240045
rect 329104 240033 329110 240045
rect 295754 240005 329110 240033
rect 295754 239993 295760 240005
rect 329104 239993 329110 240005
rect 329162 239993 329168 240045
rect 330064 239993 330070 240045
rect 330122 240033 330128 240045
rect 356560 240033 356566 240045
rect 330122 240005 356566 240033
rect 330122 239993 330128 240005
rect 356560 239993 356566 240005
rect 356618 239993 356624 240045
rect 381808 239993 381814 240045
rect 381866 240033 381872 240045
rect 389872 240033 389878 240045
rect 381866 240005 389878 240033
rect 381866 239993 381872 240005
rect 389872 239993 389878 240005
rect 389930 239993 389936 240045
rect 295600 239959 295606 239971
rect 280298 239931 281630 239959
rect 287554 239931 295606 239959
rect 280298 239919 280304 239931
rect 227152 239845 227158 239897
rect 227210 239885 227216 239897
rect 230320 239885 230326 239897
rect 227210 239857 230326 239885
rect 227210 239845 227216 239857
rect 230320 239845 230326 239857
rect 230378 239845 230384 239897
rect 256432 239845 256438 239897
rect 256490 239885 256496 239897
rect 274096 239885 274102 239897
rect 256490 239857 274102 239885
rect 256490 239845 256496 239857
rect 274096 239845 274102 239857
rect 274154 239845 274160 239897
rect 274192 239845 274198 239897
rect 274250 239885 274256 239897
rect 281488 239885 281494 239897
rect 274250 239857 281494 239885
rect 274250 239845 274256 239857
rect 281488 239845 281494 239857
rect 281546 239845 281552 239897
rect 281602 239885 281630 239931
rect 295600 239919 295606 239931
rect 295658 239919 295664 239971
rect 296080 239919 296086 239971
rect 296138 239959 296144 239971
rect 303664 239959 303670 239971
rect 296138 239931 303670 239959
rect 296138 239919 296144 239931
rect 303664 239919 303670 239931
rect 303722 239919 303728 239971
rect 307792 239919 307798 239971
rect 307850 239959 307856 239971
rect 309808 239959 309814 239971
rect 307850 239931 309814 239959
rect 307850 239919 307856 239931
rect 309808 239919 309814 239931
rect 309866 239919 309872 239971
rect 313744 239919 313750 239971
rect 313802 239959 313808 239971
rect 316144 239959 316150 239971
rect 313802 239931 316150 239959
rect 313802 239919 313808 239931
rect 316144 239919 316150 239931
rect 316202 239919 316208 239971
rect 331696 239959 331702 239971
rect 316258 239931 331702 239959
rect 281602 239857 288062 239885
rect 257200 239771 257206 239823
rect 257258 239811 257264 239823
rect 269296 239811 269302 239823
rect 257258 239783 269302 239811
rect 257258 239771 257264 239783
rect 269296 239771 269302 239783
rect 269354 239771 269360 239823
rect 269392 239771 269398 239823
rect 269450 239811 269456 239823
rect 276304 239811 276310 239823
rect 269450 239783 276310 239811
rect 269450 239771 269456 239783
rect 276304 239771 276310 239783
rect 276362 239771 276368 239823
rect 276688 239771 276694 239823
rect 276746 239811 276752 239823
rect 284464 239811 284470 239823
rect 276746 239783 284470 239811
rect 276746 239771 276752 239783
rect 284464 239771 284470 239783
rect 284522 239771 284528 239823
rect 288034 239811 288062 239857
rect 289456 239845 289462 239897
rect 289514 239885 289520 239897
rect 296656 239885 296662 239897
rect 289514 239857 296662 239885
rect 289514 239845 289520 239857
rect 296656 239845 296662 239857
rect 296714 239845 296720 239897
rect 311632 239845 311638 239897
rect 311690 239885 311696 239897
rect 316258 239885 316286 239931
rect 331696 239919 331702 239931
rect 331754 239919 331760 239971
rect 334480 239919 334486 239971
rect 334538 239959 334544 239971
rect 365872 239959 365878 239971
rect 334538 239931 365878 239959
rect 334538 239919 334544 239931
rect 365872 239919 365878 239931
rect 365930 239919 365936 239971
rect 377872 239919 377878 239971
rect 377930 239959 377936 239971
rect 407536 239959 407542 239971
rect 377930 239931 407542 239959
rect 377930 239919 377936 239931
rect 407536 239919 407542 239931
rect 407594 239919 407600 239971
rect 311690 239857 316286 239885
rect 311690 239845 311696 239857
rect 317776 239845 317782 239897
rect 317834 239885 317840 239897
rect 327952 239885 327958 239897
rect 317834 239857 327958 239885
rect 317834 239845 317840 239857
rect 327952 239845 327958 239857
rect 328010 239845 328016 239897
rect 328240 239845 328246 239897
rect 328298 239885 328304 239897
rect 352432 239885 352438 239897
rect 328298 239857 352438 239885
rect 328298 239845 328304 239857
rect 352432 239845 352438 239857
rect 352490 239845 352496 239897
rect 378640 239845 378646 239897
rect 378698 239885 378704 239897
rect 383824 239885 383830 239897
rect 378698 239857 383830 239885
rect 378698 239845 378704 239857
rect 383824 239845 383830 239857
rect 383882 239845 383888 239897
rect 291664 239811 291670 239823
rect 288034 239783 291670 239811
rect 291664 239771 291670 239783
rect 291722 239771 291728 239823
rect 294448 239771 294454 239823
rect 294506 239811 294512 239823
rect 298192 239811 298198 239823
rect 294506 239783 298198 239811
rect 294506 239771 294512 239783
rect 298192 239771 298198 239783
rect 298250 239771 298256 239823
rect 301840 239771 301846 239823
rect 301898 239811 301904 239823
rect 306640 239811 306646 239823
rect 301898 239783 306646 239811
rect 301898 239771 301904 239783
rect 306640 239771 306646 239783
rect 306698 239771 306704 239823
rect 307888 239771 307894 239823
rect 307946 239811 307952 239823
rect 312112 239811 312118 239823
rect 307946 239783 312118 239811
rect 307946 239771 307952 239783
rect 312112 239771 312118 239783
rect 312170 239771 312176 239823
rect 315184 239771 315190 239823
rect 315242 239811 315248 239823
rect 325264 239811 325270 239823
rect 315242 239783 325270 239811
rect 315242 239771 315248 239783
rect 325264 239771 325270 239783
rect 325322 239771 325328 239823
rect 326224 239771 326230 239823
rect 326282 239811 326288 239823
rect 347920 239811 347926 239823
rect 326282 239783 347926 239811
rect 326282 239771 326288 239783
rect 347920 239771 347926 239783
rect 347978 239771 347984 239823
rect 380560 239771 380566 239823
rect 380618 239811 380624 239823
rect 384880 239811 384886 239823
rect 380618 239783 384886 239811
rect 380618 239771 380624 239783
rect 384880 239771 384886 239783
rect 384938 239771 384944 239823
rect 214480 239697 214486 239749
rect 214538 239737 214544 239749
rect 225136 239737 225142 239749
rect 214538 239709 225142 239737
rect 214538 239697 214544 239709
rect 225136 239697 225142 239709
rect 225194 239697 225200 239749
rect 228016 239697 228022 239749
rect 228074 239737 228080 239749
rect 229936 239737 229942 239749
rect 228074 239709 229942 239737
rect 228074 239697 228080 239709
rect 229936 239697 229942 239709
rect 229994 239697 230000 239749
rect 248560 239697 248566 239749
rect 248618 239737 248624 239749
rect 260752 239737 260758 239749
rect 248618 239709 260758 239737
rect 248618 239697 248624 239709
rect 260752 239697 260758 239709
rect 260810 239697 260816 239749
rect 268240 239697 268246 239749
rect 268298 239737 268304 239749
rect 270928 239737 270934 239749
rect 268298 239709 270934 239737
rect 268298 239697 268304 239709
rect 270928 239697 270934 239709
rect 270986 239697 270992 239749
rect 276208 239697 276214 239749
rect 276266 239737 276272 239749
rect 280528 239737 280534 239749
rect 276266 239709 280534 239737
rect 276266 239697 276272 239709
rect 280528 239697 280534 239709
rect 280586 239697 280592 239749
rect 291376 239697 291382 239749
rect 291434 239737 291440 239749
rect 294736 239737 294742 239749
rect 291434 239709 294742 239737
rect 291434 239697 291440 239709
rect 294736 239697 294742 239709
rect 294794 239697 294800 239749
rect 322672 239697 322678 239749
rect 322730 239737 322736 239749
rect 322730 239709 324830 239737
rect 322730 239697 322736 239709
rect 229072 239623 229078 239675
rect 229130 239663 229136 239675
rect 230224 239663 230230 239675
rect 229130 239635 230230 239663
rect 229130 239623 229136 239635
rect 230224 239623 230230 239635
rect 230282 239623 230288 239675
rect 270256 239623 270262 239675
rect 270314 239663 270320 239675
rect 272272 239663 272278 239675
rect 270314 239635 272278 239663
rect 270314 239623 270320 239635
rect 272272 239623 272278 239635
rect 272330 239623 272336 239675
rect 277744 239663 277750 239675
rect 272386 239635 277750 239663
rect 271792 239549 271798 239601
rect 271850 239589 271856 239601
rect 272386 239589 272414 239635
rect 277744 239623 277750 239635
rect 277802 239623 277808 239675
rect 278032 239623 278038 239675
rect 278090 239663 278096 239675
rect 281776 239663 281782 239675
rect 278090 239635 281782 239663
rect 278090 239623 278096 239635
rect 281776 239623 281782 239635
rect 281834 239623 281840 239675
rect 282160 239623 282166 239675
rect 282218 239663 282224 239675
rect 291184 239663 291190 239675
rect 282218 239635 291190 239663
rect 282218 239623 282224 239635
rect 291184 239623 291190 239635
rect 291242 239623 291248 239675
rect 291472 239623 291478 239675
rect 291530 239663 291536 239675
rect 291530 239635 293150 239663
rect 291530 239623 291536 239635
rect 271850 239561 272414 239589
rect 271850 239549 271856 239561
rect 277648 239549 277654 239601
rect 277706 239589 277712 239601
rect 282928 239589 282934 239601
rect 277706 239561 282934 239589
rect 277706 239549 277712 239561
rect 282928 239549 282934 239561
rect 282986 239549 282992 239601
rect 283024 239549 283030 239601
rect 283082 239589 283088 239601
rect 291376 239589 291382 239601
rect 283082 239561 291382 239589
rect 283082 239549 283088 239561
rect 291376 239549 291382 239561
rect 291434 239549 291440 239601
rect 293122 239589 293150 239635
rect 293200 239623 293206 239675
rect 293258 239663 293264 239675
rect 302800 239663 302806 239675
rect 293258 239635 302806 239663
rect 293258 239623 293264 239635
rect 302800 239623 302806 239635
rect 302858 239623 302864 239675
rect 302992 239623 302998 239675
rect 303050 239663 303056 239675
rect 307600 239663 307606 239675
rect 303050 239635 307606 239663
rect 303050 239623 303056 239635
rect 307600 239623 307606 239635
rect 307658 239623 307664 239675
rect 309520 239623 309526 239675
rect 309578 239663 309584 239675
rect 310288 239663 310294 239675
rect 309578 239635 310294 239663
rect 309578 239623 309584 239635
rect 310288 239623 310294 239635
rect 310346 239623 310352 239675
rect 320848 239623 320854 239675
rect 320906 239663 320912 239675
rect 324688 239663 324694 239675
rect 320906 239635 324694 239663
rect 320906 239623 320912 239635
rect 324688 239623 324694 239635
rect 324746 239623 324752 239675
rect 324802 239663 324830 239709
rect 326992 239697 326998 239749
rect 327050 239737 327056 239749
rect 349552 239737 349558 239749
rect 327050 239709 349558 239737
rect 327050 239697 327056 239709
rect 349552 239697 349558 239709
rect 349610 239697 349616 239749
rect 374800 239697 374806 239749
rect 374858 239737 374864 239749
rect 382672 239737 382678 239749
rect 374858 239709 382678 239737
rect 374858 239697 374864 239709
rect 382672 239697 382678 239709
rect 382730 239697 382736 239749
rect 383536 239737 383542 239749
rect 382786 239709 383542 239737
rect 340912 239663 340918 239675
rect 324802 239635 340918 239663
rect 340912 239623 340918 239635
rect 340970 239623 340976 239675
rect 373840 239623 373846 239675
rect 373898 239663 373904 239675
rect 382786 239663 382814 239709
rect 383536 239697 383542 239709
rect 383594 239697 383600 239749
rect 383632 239697 383638 239749
rect 383690 239737 383696 239749
rect 385552 239737 385558 239749
rect 383690 239709 385558 239737
rect 383690 239697 383696 239709
rect 385552 239697 385558 239709
rect 385610 239697 385616 239749
rect 373898 239635 382814 239663
rect 373898 239623 373904 239635
rect 383152 239623 383158 239675
rect 383210 239663 383216 239675
rect 388144 239663 388150 239675
rect 383210 239635 388150 239663
rect 383210 239623 383216 239635
rect 388144 239623 388150 239635
rect 388202 239623 388208 239675
rect 301840 239589 301846 239601
rect 293122 239561 301846 239589
rect 301840 239549 301846 239561
rect 301898 239549 301904 239601
rect 302512 239549 302518 239601
rect 302570 239589 302576 239601
rect 307216 239589 307222 239601
rect 302570 239561 307222 239589
rect 302570 239549 302576 239561
rect 307216 239549 307222 239561
rect 307274 239549 307280 239601
rect 308848 239549 308854 239601
rect 308906 239589 308912 239601
rect 310192 239589 310198 239601
rect 308906 239561 310198 239589
rect 308906 239549 308912 239561
rect 310192 239549 310198 239561
rect 310250 239549 310256 239601
rect 323056 239549 323062 239601
rect 323114 239589 323120 239601
rect 341296 239589 341302 239601
rect 323114 239561 341302 239589
rect 323114 239549 323120 239561
rect 341296 239549 341302 239561
rect 341354 239549 341360 239601
rect 380080 239549 380086 239601
rect 380138 239589 380144 239601
rect 383728 239589 383734 239601
rect 380138 239561 383734 239589
rect 380138 239549 380144 239561
rect 383728 239549 383734 239561
rect 383786 239549 383792 239601
rect 277072 239475 277078 239527
rect 277130 239515 277136 239527
rect 283792 239515 283798 239527
rect 277130 239487 283798 239515
rect 277130 239475 277136 239487
rect 283792 239475 283798 239487
rect 283850 239475 283856 239527
rect 283888 239475 283894 239527
rect 283946 239515 283952 239527
rect 292144 239515 292150 239527
rect 283946 239487 292150 239515
rect 283946 239475 283952 239487
rect 292144 239475 292150 239487
rect 292202 239475 292208 239527
rect 297808 239475 297814 239527
rect 297866 239515 297872 239527
rect 305008 239515 305014 239527
rect 297866 239487 305014 239515
rect 297866 239475 297872 239487
rect 305008 239475 305014 239487
rect 305066 239475 305072 239527
rect 327376 239475 327382 239527
rect 327434 239515 327440 239527
rect 332944 239515 332950 239527
rect 327434 239487 332950 239515
rect 327434 239475 327440 239487
rect 332944 239475 332950 239487
rect 333002 239475 333008 239527
rect 380848 239475 380854 239527
rect 380906 239515 380912 239527
rect 383056 239515 383062 239527
rect 380906 239487 383062 239515
rect 380906 239475 380912 239487
rect 383056 239475 383062 239487
rect 383114 239475 383120 239527
rect 386608 239515 386614 239527
rect 383170 239487 386614 239515
rect 237136 239401 237142 239453
rect 237194 239441 237200 239453
rect 241840 239441 241846 239453
rect 237194 239413 241846 239441
rect 237194 239401 237200 239413
rect 241840 239401 241846 239413
rect 241898 239401 241904 239453
rect 276208 239401 276214 239453
rect 276266 239441 276272 239453
rect 286000 239441 286006 239453
rect 276266 239413 286006 239441
rect 276266 239401 276272 239413
rect 286000 239401 286006 239413
rect 286058 239401 286064 239453
rect 290800 239441 290806 239453
rect 286114 239413 290806 239441
rect 235504 239327 235510 239379
rect 235562 239367 235568 239379
rect 238672 239367 238678 239379
rect 235562 239339 238678 239367
rect 235562 239327 235568 239339
rect 238672 239327 238678 239339
rect 238730 239327 238736 239379
rect 272464 239327 272470 239379
rect 272522 239367 272528 239379
rect 285520 239367 285526 239379
rect 272522 239339 285526 239367
rect 272522 239327 272528 239339
rect 285520 239327 285526 239339
rect 285578 239327 285584 239379
rect 285616 239327 285622 239379
rect 285674 239367 285680 239379
rect 286114 239367 286142 239413
rect 290800 239401 290806 239413
rect 290858 239401 290864 239453
rect 290896 239401 290902 239453
rect 290954 239441 290960 239453
rect 293296 239441 293302 239453
rect 290954 239413 293302 239441
rect 290954 239401 290960 239413
rect 293296 239401 293302 239413
rect 293354 239401 293360 239453
rect 293392 239401 293398 239453
rect 293450 239441 293456 239453
rect 294448 239441 294454 239453
rect 293450 239413 294454 239441
rect 293450 239401 293456 239413
rect 294448 239401 294454 239413
rect 294506 239401 294512 239453
rect 295984 239401 295990 239453
rect 296042 239441 296048 239453
rect 304144 239441 304150 239453
rect 296042 239413 304150 239441
rect 296042 239401 296048 239413
rect 304144 239401 304150 239413
rect 304202 239401 304208 239453
rect 323440 239401 323446 239453
rect 323498 239441 323504 239453
rect 341968 239441 341974 239453
rect 323498 239413 341974 239441
rect 323498 239401 323504 239413
rect 341968 239401 341974 239413
rect 342026 239401 342032 239453
rect 380080 239401 380086 239453
rect 380138 239441 380144 239453
rect 383170 239441 383198 239487
rect 386608 239475 386614 239487
rect 386666 239475 386672 239527
rect 380138 239413 383198 239441
rect 380138 239401 380144 239413
rect 285674 239339 286142 239367
rect 285674 239327 285680 239339
rect 294256 239327 294262 239379
rect 294314 239367 294320 239379
rect 303568 239367 303574 239379
rect 294314 239339 303574 239367
rect 294314 239327 294320 239339
rect 303568 239327 303574 239339
rect 303626 239327 303632 239379
rect 303664 239327 303670 239379
rect 303722 239367 303728 239379
rect 314800 239367 314806 239379
rect 303722 239339 314806 239367
rect 303722 239327 303728 239339
rect 314800 239327 314806 239339
rect 314858 239327 314864 239379
rect 322192 239327 322198 239379
rect 322250 239367 322256 239379
rect 338896 239367 338902 239379
rect 322250 239339 338902 239367
rect 322250 239327 322256 239339
rect 338896 239327 338902 239339
rect 338954 239327 338960 239379
rect 395824 239367 395830 239379
rect 370546 239339 395830 239367
rect 275728 239253 275734 239305
rect 275786 239293 275792 239305
rect 283024 239293 283030 239305
rect 275786 239265 283030 239293
rect 275786 239253 275792 239265
rect 283024 239253 283030 239265
rect 283082 239253 283088 239305
rect 284080 239293 284086 239305
rect 283330 239265 284086 239293
rect 42544 239179 42550 239231
rect 42602 239219 42608 239231
rect 42602 239191 42782 239219
rect 42602 239179 42608 239191
rect 42448 238883 42454 238935
rect 42506 238923 42512 238935
rect 42754 238923 42782 239191
rect 139984 239179 139990 239231
rect 140042 239219 140048 239231
rect 152464 239219 152470 239231
rect 140042 239191 152470 239219
rect 140042 239179 140048 239191
rect 152464 239179 152470 239191
rect 152522 239179 152528 239231
rect 215920 239179 215926 239231
rect 215978 239219 215984 239231
rect 218896 239219 218902 239231
rect 215978 239191 218902 239219
rect 215978 239179 215984 239191
rect 218896 239179 218902 239191
rect 218954 239179 218960 239231
rect 273424 239179 273430 239231
rect 273482 239219 273488 239231
rect 278800 239219 278806 239231
rect 273482 239191 278806 239219
rect 273482 239179 273488 239191
rect 278800 239179 278806 239191
rect 278858 239179 278864 239231
rect 278896 239179 278902 239231
rect 278954 239219 278960 239231
rect 279664 239219 279670 239231
rect 278954 239191 279670 239219
rect 278954 239179 278960 239191
rect 279664 239179 279670 239191
rect 279722 239179 279728 239231
rect 280432 239179 280438 239231
rect 280490 239219 280496 239231
rect 283330 239219 283358 239265
rect 284080 239253 284086 239265
rect 284138 239253 284144 239305
rect 287344 239253 287350 239305
rect 287402 239293 287408 239305
rect 294352 239293 294358 239305
rect 287402 239265 294358 239293
rect 287402 239253 287408 239265
rect 294352 239253 294358 239265
rect 294410 239253 294416 239305
rect 326608 239253 326614 239305
rect 326666 239293 326672 239305
rect 348976 239293 348982 239305
rect 326666 239265 348982 239293
rect 326666 239253 326672 239265
rect 348976 239253 348982 239265
rect 349034 239253 349040 239305
rect 290896 239219 290902 239231
rect 280490 239191 283358 239219
rect 286690 239191 290902 239219
rect 280490 239179 280496 239191
rect 238480 239105 238486 239157
rect 238538 239145 238544 239157
rect 241648 239145 241654 239157
rect 238538 239117 241654 239145
rect 238538 239105 238544 239117
rect 241648 239105 241654 239117
rect 241706 239105 241712 239157
rect 272656 239105 272662 239157
rect 272714 239145 272720 239157
rect 286690 239145 286718 239191
rect 290896 239179 290902 239191
rect 290954 239179 290960 239231
rect 291280 239179 291286 239231
rect 291338 239219 291344 239231
rect 296560 239219 296566 239231
rect 291338 239191 296566 239219
rect 291338 239179 291344 239191
rect 296560 239179 296566 239191
rect 296618 239179 296624 239231
rect 296656 239179 296662 239231
rect 296714 239219 296720 239231
rect 313840 239219 313846 239231
rect 296714 239191 313846 239219
rect 296714 239179 296720 239191
rect 313840 239179 313846 239191
rect 313898 239179 313904 239231
rect 321232 239179 321238 239231
rect 321290 239219 321296 239231
rect 337168 239219 337174 239231
rect 321290 239191 337174 239219
rect 321290 239179 321296 239191
rect 337168 239179 337174 239191
rect 337226 239179 337232 239231
rect 360976 239179 360982 239231
rect 361034 239219 361040 239231
rect 370546 239219 370574 239339
rect 395824 239327 395830 239339
rect 395882 239327 395888 239379
rect 392080 239293 392086 239305
rect 361034 239191 370574 239219
rect 370690 239265 392086 239293
rect 361034 239179 361040 239191
rect 272714 239117 282398 239145
rect 272714 239105 272720 239117
rect 258640 239031 258646 239083
rect 258698 239071 258704 239083
rect 258928 239071 258934 239083
rect 258698 239043 258934 239071
rect 258698 239031 258704 239043
rect 258928 239031 258934 239043
rect 258986 239031 258992 239083
rect 282256 239071 282262 239083
rect 278338 239043 282262 239071
rect 228112 238957 228118 239009
rect 228170 238997 228176 239009
rect 231952 238997 231958 239009
rect 228170 238969 231958 238997
rect 228170 238957 228176 238969
rect 231952 238957 231958 238969
rect 232010 238957 232016 239009
rect 240112 238957 240118 239009
rect 240170 238997 240176 239009
rect 256816 238997 256822 239009
rect 240170 238969 256822 238997
rect 240170 238957 240176 238969
rect 256816 238957 256822 238969
rect 256874 238957 256880 239009
rect 260368 238957 260374 239009
rect 260426 238997 260432 239009
rect 278338 238997 278366 239043
rect 282256 239031 282262 239043
rect 282314 239031 282320 239083
rect 282370 239071 282398 239117
rect 283426 239117 286718 239145
rect 283426 239071 283454 239117
rect 287056 239105 287062 239157
rect 287114 239145 287120 239157
rect 287114 239117 291134 239145
rect 287114 239105 287120 239117
rect 282370 239043 283454 239071
rect 284080 239031 284086 239083
rect 284138 239071 284144 239083
rect 290800 239071 290806 239083
rect 284138 239043 290806 239071
rect 284138 239031 284144 239043
rect 290800 239031 290806 239043
rect 290858 239031 290864 239083
rect 291106 239071 291134 239117
rect 318256 239105 318262 239157
rect 318314 239145 318320 239157
rect 332752 239145 332758 239157
rect 318314 239117 332758 239145
rect 318314 239105 318320 239117
rect 332752 239105 332758 239117
rect 332810 239105 332816 239157
rect 360208 239105 360214 239157
rect 360266 239145 360272 239157
rect 370690 239145 370718 239265
rect 392080 239253 392086 239265
rect 392138 239253 392144 239305
rect 375664 239179 375670 239231
rect 375722 239219 375728 239231
rect 402352 239219 402358 239231
rect 375722 239191 402358 239219
rect 375722 239179 375728 239191
rect 402352 239179 402358 239191
rect 402410 239179 402416 239231
rect 360266 239117 370718 239145
rect 360266 239105 360272 239117
rect 375184 239105 375190 239157
rect 375242 239145 375248 239157
rect 400624 239145 400630 239157
rect 375242 239117 400630 239145
rect 375242 239105 375248 239117
rect 400624 239105 400630 239117
rect 400682 239105 400688 239157
rect 300016 239071 300022 239083
rect 291106 239043 300022 239071
rect 300016 239031 300022 239043
rect 300074 239031 300080 239083
rect 324400 239031 324406 239083
rect 324458 239071 324464 239083
rect 343696 239071 343702 239083
rect 324458 239043 343702 239071
rect 324458 239031 324464 239043
rect 343696 239031 343702 239043
rect 343754 239031 343760 239083
rect 373360 239031 373366 239083
rect 373418 239071 373424 239083
rect 396880 239071 396886 239083
rect 373418 239043 396886 239071
rect 373418 239031 373424 239043
rect 396880 239031 396886 239043
rect 396938 239031 396944 239083
rect 260426 238969 278366 238997
rect 260426 238957 260432 238969
rect 278416 238957 278422 239009
rect 278474 238997 278480 239009
rect 279376 238997 279382 239009
rect 278474 238969 279382 238997
rect 278474 238957 278480 238969
rect 279376 238957 279382 238969
rect 279434 238957 279440 239009
rect 279472 238957 279478 239009
rect 279530 238997 279536 239009
rect 292240 238997 292246 239009
rect 279530 238969 292246 238997
rect 279530 238957 279536 238969
rect 292240 238957 292246 238969
rect 292298 238957 292304 239009
rect 293968 238957 293974 239009
rect 294026 238997 294032 239009
rect 303184 238997 303190 239009
rect 294026 238969 303190 238997
rect 294026 238957 294032 238969
rect 303184 238957 303190 238969
rect 303242 238957 303248 239009
rect 304720 238957 304726 239009
rect 304778 238997 304784 239009
rect 308176 238997 308182 239009
rect 304778 238969 308182 238997
rect 304778 238957 304784 238969
rect 308176 238957 308182 238969
rect 308234 238957 308240 239009
rect 311632 238957 311638 239009
rect 311690 238997 311696 239009
rect 323632 238997 323638 239009
rect 311690 238969 323638 238997
rect 311690 238957 311696 238969
rect 323632 238957 323638 238969
rect 323690 238957 323696 239009
rect 331312 238997 331318 239009
rect 323746 238969 331318 238997
rect 42506 238895 42782 238923
rect 42506 238883 42512 238895
rect 227728 238883 227734 238935
rect 227786 238923 227792 238935
rect 232816 238923 232822 238935
rect 227786 238895 232822 238923
rect 227786 238883 227792 238895
rect 232816 238883 232822 238895
rect 232874 238883 232880 238935
rect 240496 238883 240502 238935
rect 240554 238923 240560 238935
rect 255664 238923 255670 238935
rect 240554 238895 255670 238923
rect 240554 238883 240560 238895
rect 255664 238883 255670 238895
rect 255722 238883 255728 238935
rect 259984 238883 259990 238935
rect 260042 238923 260048 238935
rect 275248 238923 275254 238935
rect 260042 238895 275254 238923
rect 260042 238883 260048 238895
rect 275248 238883 275254 238895
rect 275306 238883 275312 238935
rect 281680 238883 281686 238935
rect 281738 238923 281744 238935
rect 297424 238923 297430 238935
rect 281738 238895 297430 238923
rect 281738 238883 281744 238895
rect 297424 238883 297430 238895
rect 297482 238883 297488 238935
rect 299056 238883 299062 238935
rect 299114 238923 299120 238935
rect 305776 238923 305782 238935
rect 299114 238895 305782 238923
rect 299114 238883 299120 238895
rect 305776 238883 305782 238895
rect 305834 238883 305840 238935
rect 318544 238883 318550 238935
rect 318602 238923 318608 238935
rect 323746 238923 323774 238969
rect 331312 238957 331318 238969
rect 331370 238957 331376 239009
rect 351088 238957 351094 239009
rect 351146 238997 351152 239009
rect 379024 238997 379030 239009
rect 351146 238969 379030 238997
rect 351146 238957 351152 238969
rect 379024 238957 379030 238969
rect 379082 238957 379088 239009
rect 380464 238957 380470 239009
rect 380522 238997 380528 239009
rect 383152 238997 383158 239009
rect 380522 238969 383158 238997
rect 380522 238957 380528 238969
rect 383152 238957 383158 238969
rect 383210 238957 383216 239009
rect 348400 238923 348406 238935
rect 318602 238895 323774 238923
rect 323842 238895 348406 238923
rect 318602 238883 318608 238895
rect 256816 238809 256822 238861
rect 256874 238849 256880 238861
rect 316240 238849 316246 238861
rect 256874 238821 316246 238849
rect 256874 238809 256880 238821
rect 316240 238809 316246 238821
rect 316298 238809 316304 238861
rect 317392 238809 317398 238861
rect 317450 238849 317456 238861
rect 323728 238849 323734 238861
rect 317450 238821 323734 238849
rect 317450 238809 317456 238821
rect 323728 238809 323734 238821
rect 323786 238809 323792 238861
rect 224560 238735 224566 238787
rect 224618 238775 224624 238787
rect 239440 238775 239446 238787
rect 224618 238747 239446 238775
rect 224618 238735 224624 238747
rect 239440 238735 239446 238747
rect 239498 238735 239504 238787
rect 239536 238735 239542 238787
rect 239594 238775 239600 238787
rect 257392 238775 257398 238787
rect 239594 238747 257398 238775
rect 239594 238735 239600 238747
rect 257392 238735 257398 238747
rect 257450 238735 257456 238787
rect 257776 238735 257782 238787
rect 257834 238775 257840 238787
rect 318160 238775 318166 238787
rect 257834 238747 318166 238775
rect 257834 238735 257840 238747
rect 318160 238735 318166 238747
rect 318218 238735 318224 238787
rect 323842 238775 323870 238895
rect 348400 238883 348406 238895
rect 348458 238883 348464 238935
rect 348496 238883 348502 238935
rect 348554 238923 348560 238935
rect 377296 238923 377302 238935
rect 348554 238895 377302 238923
rect 348554 238883 348560 238895
rect 377296 238883 377302 238895
rect 377354 238883 377360 238935
rect 323920 238809 323926 238861
rect 323978 238849 323984 238861
rect 351088 238849 351094 238861
rect 323978 238821 351094 238849
rect 323978 238809 323984 238821
rect 351088 238809 351094 238821
rect 351146 238809 351152 238861
rect 351184 238809 351190 238861
rect 351242 238849 351248 238861
rect 358768 238849 358774 238861
rect 351242 238821 358774 238849
rect 351242 238809 351248 238821
rect 358768 238809 358774 238821
rect 358826 238809 358832 238861
rect 366832 238809 366838 238861
rect 366890 238849 366896 238861
rect 383344 238849 383350 238861
rect 366890 238821 383350 238849
rect 366890 238809 366896 238821
rect 383344 238809 383350 238821
rect 383402 238809 383408 238861
rect 318370 238747 323870 238775
rect 226288 238661 226294 238713
rect 226346 238701 226352 238713
rect 235600 238701 235606 238713
rect 226346 238673 235606 238701
rect 226346 238661 226352 238673
rect 235600 238661 235606 238673
rect 235658 238661 235664 238713
rect 256240 238661 256246 238713
rect 256298 238701 256304 238713
rect 318256 238701 318262 238713
rect 256298 238673 318262 238701
rect 256298 238661 256304 238673
rect 318256 238661 318262 238673
rect 318314 238661 318320 238713
rect 227248 238587 227254 238639
rect 227306 238627 227312 238639
rect 234064 238627 234070 238639
rect 227306 238599 234070 238627
rect 227306 238587 227312 238599
rect 234064 238587 234070 238599
rect 234122 238587 234128 238639
rect 248944 238587 248950 238639
rect 249002 238627 249008 238639
rect 316336 238627 316342 238639
rect 249002 238599 316342 238627
rect 249002 238587 249008 238599
rect 316336 238587 316342 238599
rect 316394 238587 316400 238639
rect 316432 238587 316438 238639
rect 316490 238627 316496 238639
rect 318370 238627 318398 238747
rect 324208 238735 324214 238787
rect 324266 238775 324272 238787
rect 328816 238775 328822 238787
rect 324266 238747 328822 238775
rect 324266 238735 324272 238747
rect 328816 238735 328822 238747
rect 328874 238735 328880 238787
rect 330640 238735 330646 238787
rect 330698 238775 330704 238787
rect 357232 238775 357238 238787
rect 330698 238747 357238 238775
rect 330698 238735 330704 238747
rect 357232 238735 357238 238747
rect 357290 238735 357296 238787
rect 381424 238735 381430 238787
rect 381482 238775 381488 238787
rect 389200 238775 389206 238787
rect 381482 238747 389206 238775
rect 381482 238735 381488 238747
rect 389200 238735 389206 238747
rect 389258 238735 389264 238787
rect 318640 238661 318646 238713
rect 318698 238701 318704 238713
rect 332176 238701 332182 238713
rect 318698 238673 332182 238701
rect 318698 238661 318704 238673
rect 332176 238661 332182 238673
rect 332234 238661 332240 238713
rect 334096 238661 334102 238713
rect 334154 238701 334160 238713
rect 365296 238701 365302 238713
rect 334154 238673 365302 238701
rect 334154 238661 334160 238673
rect 365296 238661 365302 238673
rect 365354 238661 365360 238713
rect 383152 238661 383158 238713
rect 383210 238701 383216 238713
rect 387568 238701 387574 238713
rect 383210 238673 387574 238701
rect 383210 238661 383216 238673
rect 387568 238661 387574 238673
rect 387626 238661 387632 238713
rect 316490 238599 318398 238627
rect 316490 238587 316496 238599
rect 319024 238587 319030 238639
rect 319082 238627 319088 238639
rect 332368 238627 332374 238639
rect 319082 238599 332374 238627
rect 319082 238587 319088 238599
rect 332368 238587 332374 238599
rect 332426 238587 332432 238639
rect 333616 238587 333622 238639
rect 333674 238627 333680 238639
rect 363280 238627 363286 238639
rect 333674 238599 363286 238627
rect 333674 238587 333680 238599
rect 363280 238587 363286 238599
rect 363338 238587 363344 238639
rect 370384 238587 370390 238639
rect 370442 238627 370448 238639
rect 390352 238627 390358 238639
rect 370442 238599 390358 238627
rect 370442 238587 370448 238599
rect 390352 238587 390358 238599
rect 390410 238587 390416 238639
rect 42160 238513 42166 238565
rect 42218 238553 42224 238565
rect 43024 238553 43030 238565
rect 42218 238525 43030 238553
rect 42218 238513 42224 238525
rect 43024 238513 43030 238525
rect 43082 238513 43088 238565
rect 217072 238513 217078 238565
rect 217130 238553 217136 238565
rect 255184 238553 255190 238565
rect 217130 238525 255190 238553
rect 217130 238513 217136 238525
rect 255184 238513 255190 238525
rect 255242 238513 255248 238565
rect 255568 238513 255574 238565
rect 255626 238553 255632 238565
rect 318064 238553 318070 238565
rect 255626 238525 318070 238553
rect 255626 238513 255632 238525
rect 318064 238513 318070 238525
rect 318122 238513 318128 238565
rect 319600 238513 319606 238565
rect 319658 238553 319664 238565
rect 333424 238553 333430 238565
rect 319658 238525 333430 238553
rect 319658 238513 319664 238525
rect 333424 238513 333430 238525
rect 333482 238513 333488 238565
rect 334864 238513 334870 238565
rect 334922 238553 334928 238565
rect 334922 238525 351422 238553
rect 334922 238513 334928 238525
rect 226864 238439 226870 238491
rect 226922 238479 226928 238491
rect 235024 238479 235030 238491
rect 226922 238451 235030 238479
rect 226922 238439 226928 238451
rect 235024 238439 235030 238451
rect 235082 238439 235088 238491
rect 254128 238439 254134 238491
rect 254186 238479 254192 238491
rect 330928 238479 330934 238491
rect 254186 238451 330934 238479
rect 254186 238439 254192 238451
rect 330928 238439 330934 238451
rect 330986 238439 330992 238491
rect 331120 238439 331126 238491
rect 331178 238479 331184 238491
rect 351184 238479 351190 238491
rect 331178 238451 351190 238479
rect 331178 238439 331184 238451
rect 351184 238439 351190 238451
rect 351242 238439 351248 238491
rect 351394 238479 351422 238525
rect 360880 238513 360886 238565
rect 360938 238553 360944 238565
rect 378352 238553 378358 238565
rect 360938 238525 378358 238553
rect 360938 238513 360944 238525
rect 378352 238513 378358 238525
rect 378410 238513 378416 238565
rect 383056 238513 383062 238565
rect 383114 238553 383120 238565
rect 391408 238553 391414 238565
rect 383114 238525 391414 238553
rect 383114 238513 383120 238525
rect 391408 238513 391414 238525
rect 391466 238513 391472 238565
rect 367024 238479 367030 238491
rect 351394 238451 367030 238479
rect 367024 238439 367030 238451
rect 367082 238439 367088 238491
rect 368464 238439 368470 238491
rect 368522 238479 368528 238491
rect 385936 238479 385942 238491
rect 368522 238451 385942 238479
rect 368522 238439 368528 238451
rect 385936 238439 385942 238451
rect 385994 238439 386000 238491
rect 254608 238365 254614 238417
rect 254666 238405 254672 238417
rect 336976 238405 336982 238417
rect 254666 238377 336982 238405
rect 254666 238365 254672 238377
rect 336976 238365 336982 238377
rect 337034 238365 337040 238417
rect 351376 238365 351382 238417
rect 351434 238405 351440 238417
rect 358864 238405 358870 238417
rect 351434 238377 358870 238405
rect 351434 238365 351440 238377
rect 358864 238365 358870 238377
rect 358922 238365 358928 238417
rect 369424 238365 369430 238417
rect 369482 238405 369488 238417
rect 388816 238405 388822 238417
rect 369482 238377 388822 238405
rect 369482 238365 369488 238377
rect 388816 238365 388822 238377
rect 388874 238365 388880 238417
rect 218032 238291 218038 238343
rect 218090 238331 218096 238343
rect 253456 238331 253462 238343
rect 218090 238303 253462 238331
rect 218090 238291 218096 238303
rect 253456 238291 253462 238303
rect 253514 238291 253520 238343
rect 258544 238291 258550 238343
rect 258602 238331 258608 238343
rect 279472 238331 279478 238343
rect 258602 238303 279478 238331
rect 258602 238291 258608 238303
rect 279472 238291 279478 238303
rect 279530 238291 279536 238343
rect 288112 238291 288118 238343
rect 288170 238331 288176 238343
rect 293680 238331 293686 238343
rect 288170 238303 293686 238331
rect 288170 238291 288176 238303
rect 293680 238291 293686 238303
rect 293738 238291 293744 238343
rect 293776 238291 293782 238343
rect 293834 238331 293840 238343
rect 385264 238331 385270 238343
rect 293834 238303 385270 238331
rect 293834 238291 293840 238303
rect 385264 238291 385270 238303
rect 385322 238291 385328 238343
rect 253360 238217 253366 238269
rect 253418 238257 253424 238269
rect 253418 238229 330878 238257
rect 253418 238217 253424 238229
rect 252400 238143 252406 238195
rect 252458 238183 252464 238195
rect 330850 238183 330878 238229
rect 330928 238217 330934 238269
rect 330986 238257 330992 238269
rect 338704 238257 338710 238269
rect 330986 238229 338710 238257
rect 330986 238217 330992 238229
rect 338704 238217 338710 238229
rect 338762 238217 338768 238269
rect 371632 238217 371638 238269
rect 371690 238257 371696 238269
rect 393616 238257 393622 238269
rect 371690 238229 393622 238257
rect 371690 238217 371696 238229
rect 393616 238217 393622 238229
rect 393674 238217 393680 238269
rect 340432 238183 340438 238195
rect 252458 238155 330782 238183
rect 330850 238155 340438 238183
rect 252458 238143 252464 238155
rect 223216 238069 223222 238121
rect 223274 238109 223280 238121
rect 242608 238109 242614 238121
rect 223274 238081 242614 238109
rect 223274 238069 223280 238081
rect 242608 238069 242614 238081
rect 242666 238069 242672 238121
rect 251920 238069 251926 238121
rect 251978 238109 251984 238121
rect 330754 238109 330782 238155
rect 340432 238143 340438 238155
rect 340490 238143 340496 238195
rect 369808 238143 369814 238195
rect 369866 238183 369872 238195
rect 389680 238183 389686 238195
rect 369866 238155 389686 238183
rect 369866 238143 369872 238155
rect 389680 238143 389686 238155
rect 389738 238143 389744 238195
rect 341488 238109 341494 238121
rect 251978 238081 330686 238109
rect 330754 238081 341494 238109
rect 251978 238069 251984 238081
rect 221872 237995 221878 238047
rect 221930 238035 221936 238047
rect 244816 238035 244822 238047
rect 221930 238007 244822 238035
rect 221930 237995 221936 238007
rect 244816 237995 244822 238007
rect 244874 237995 244880 238047
rect 251152 237995 251158 238047
rect 251210 238035 251216 238047
rect 330544 238035 330550 238047
rect 251210 238007 330550 238035
rect 251210 237995 251216 238007
rect 330544 237995 330550 238007
rect 330602 237995 330608 238047
rect 330658 238035 330686 238081
rect 341488 238069 341494 238081
rect 341546 238069 341552 238121
rect 342736 238069 342742 238121
rect 342794 238109 342800 238121
rect 370000 238109 370006 238121
rect 342794 238081 370006 238109
rect 342794 238069 342800 238081
rect 370000 238069 370006 238081
rect 370058 238069 370064 238121
rect 371152 238069 371158 238121
rect 371210 238109 371216 238121
rect 391888 238109 391894 238121
rect 371210 238081 391894 238109
rect 371210 238069 371216 238081
rect 391888 238069 391894 238081
rect 391946 238069 391952 238121
rect 343504 238035 343510 238047
rect 330658 238007 343510 238035
rect 343504 237995 343510 238007
rect 343562 237995 343568 238047
rect 372016 237995 372022 238047
rect 372074 238035 372080 238047
rect 394192 238035 394198 238047
rect 372074 238007 394198 238035
rect 372074 237995 372080 238007
rect 394192 237995 394198 238007
rect 394250 237995 394256 238047
rect 223312 237921 223318 237973
rect 223370 237961 223376 237973
rect 242128 237961 242134 237973
rect 223370 237933 242134 237961
rect 223370 237921 223376 237933
rect 242128 237921 242134 237933
rect 242186 237921 242192 237973
rect 249808 237921 249814 237973
rect 249866 237961 249872 237973
rect 328432 237961 328438 237973
rect 249866 237933 328438 237961
rect 249866 237921 249872 237933
rect 328432 237921 328438 237933
rect 328490 237921 328496 237973
rect 328528 237921 328534 237973
rect 328586 237961 328592 237973
rect 338224 237961 338230 237973
rect 328586 237933 338230 237961
rect 328586 237921 328592 237933
rect 338224 237921 338230 237933
rect 338282 237921 338288 237973
rect 371248 237921 371254 237973
rect 371306 237961 371312 237973
rect 392464 237961 392470 237973
rect 371306 237933 392470 237961
rect 371306 237921 371312 237933
rect 392464 237921 392470 237933
rect 392522 237921 392528 237973
rect 42160 237847 42166 237899
rect 42218 237887 42224 237899
rect 47536 237887 47542 237899
rect 42218 237859 47542 237887
rect 42218 237847 42224 237859
rect 47536 237847 47542 237859
rect 47594 237847 47600 237899
rect 222832 237847 222838 237899
rect 222890 237887 222896 237899
rect 243760 237887 243766 237899
rect 222890 237859 243766 237887
rect 222890 237847 222896 237859
rect 243760 237847 243766 237859
rect 243818 237847 243824 237899
rect 249328 237847 249334 237899
rect 249386 237887 249392 237899
rect 349168 237887 349174 237899
rect 249386 237859 349174 237887
rect 249386 237847 249392 237859
rect 349168 237847 349174 237859
rect 349226 237847 349232 237899
rect 359824 237847 359830 237899
rect 359882 237887 359888 237899
rect 380944 237887 380950 237899
rect 359882 237859 380950 237887
rect 359882 237847 359888 237859
rect 380944 237847 380950 237859
rect 381002 237847 381008 237899
rect 383056 237847 383062 237899
rect 383114 237887 383120 237899
rect 384400 237887 384406 237899
rect 383114 237859 384406 237887
rect 383114 237847 383120 237859
rect 384400 237847 384406 237859
rect 384458 237847 384464 237899
rect 384496 237847 384502 237899
rect 384554 237887 384560 237899
rect 410992 237887 410998 237899
rect 384554 237859 410998 237887
rect 384554 237847 384560 237859
rect 410992 237847 410998 237859
rect 411050 237847 411056 237899
rect 223696 237773 223702 237825
rect 223754 237813 223760 237825
rect 241552 237813 241558 237825
rect 223754 237785 241558 237813
rect 223754 237773 223760 237785
rect 241552 237773 241558 237785
rect 241610 237773 241616 237825
rect 247120 237773 247126 237825
rect 247178 237813 247184 237825
rect 353968 237813 353974 237825
rect 247178 237785 353974 237813
rect 247178 237773 247184 237785
rect 353968 237773 353974 237785
rect 354026 237773 354032 237825
rect 375568 237773 375574 237825
rect 375626 237813 375632 237825
rect 401200 237813 401206 237825
rect 375626 237785 401206 237813
rect 375626 237773 375632 237785
rect 401200 237773 401206 237785
rect 401258 237773 401264 237825
rect 228496 237699 228502 237751
rect 228554 237739 228560 237751
rect 230800 237739 230806 237751
rect 228554 237711 230806 237739
rect 228554 237699 228560 237711
rect 230800 237699 230806 237711
rect 230858 237699 230864 237751
rect 247600 237699 247606 237751
rect 247658 237739 247664 237751
rect 351952 237739 351958 237751
rect 247658 237711 351958 237739
rect 247658 237699 247664 237711
rect 351952 237699 351958 237711
rect 352010 237699 352016 237751
rect 384400 237699 384406 237751
rect 384458 237739 384464 237751
rect 410608 237739 410614 237751
rect 384458 237711 410614 237739
rect 384458 237699 384464 237711
rect 410608 237699 410614 237711
rect 410666 237699 410672 237751
rect 549232 237699 549238 237751
rect 549290 237739 549296 237751
rect 649360 237739 649366 237751
rect 549290 237711 649366 237739
rect 549290 237699 549296 237711
rect 649360 237699 649366 237711
rect 649418 237699 649424 237751
rect 221488 237625 221494 237677
rect 221546 237665 221552 237677
rect 245872 237665 245878 237677
rect 221546 237637 245878 237665
rect 221546 237625 221552 237637
rect 245872 237625 245878 237637
rect 245930 237625 245936 237677
rect 246160 237625 246166 237677
rect 246218 237665 246224 237677
rect 355024 237665 355030 237677
rect 246218 237637 355030 237665
rect 246218 237625 246224 237637
rect 355024 237625 355030 237637
rect 355082 237625 355088 237677
rect 373456 237625 373462 237677
rect 373514 237665 373520 237677
rect 397936 237665 397942 237677
rect 373514 237637 397942 237665
rect 373514 237625 373520 237637
rect 397936 237625 397942 237637
rect 397994 237625 398000 237677
rect 497488 237625 497494 237677
rect 497546 237665 497552 237677
rect 602896 237665 602902 237677
rect 497546 237637 602902 237665
rect 497546 237625 497552 237637
rect 602896 237625 602902 237637
rect 602954 237625 602960 237677
rect 148336 237551 148342 237603
rect 148394 237591 148400 237603
rect 207184 237591 207190 237603
rect 148394 237563 207190 237591
rect 148394 237551 148400 237563
rect 207184 237551 207190 237563
rect 207242 237591 207248 237603
rect 221968 237591 221974 237603
rect 207242 237563 221974 237591
rect 207242 237551 207248 237563
rect 221968 237551 221974 237563
rect 222026 237551 222032 237603
rect 245776 237551 245782 237603
rect 245834 237591 245840 237603
rect 356176 237591 356182 237603
rect 245834 237563 356182 237591
rect 245834 237551 245840 237563
rect 356176 237551 356182 237563
rect 356234 237551 356240 237603
rect 374224 237551 374230 237603
rect 374282 237591 374288 237603
rect 399664 237591 399670 237603
rect 374282 237563 399670 237591
rect 374282 237551 374288 237563
rect 399664 237551 399670 237563
rect 399722 237551 399728 237603
rect 420592 237551 420598 237603
rect 420650 237591 420656 237603
rect 607600 237591 607606 237603
rect 420650 237563 607606 237591
rect 420650 237551 420656 237563
rect 607600 237551 607606 237563
rect 607658 237551 607664 237603
rect 239056 237477 239062 237529
rect 239114 237517 239120 237529
rect 259120 237517 259126 237529
rect 239114 237489 259126 237517
rect 239114 237477 239120 237489
rect 259120 237477 259126 237489
rect 259178 237477 259184 237529
rect 275248 237477 275254 237529
rect 275306 237517 275312 237529
rect 291952 237517 291958 237529
rect 275306 237489 291958 237517
rect 275306 237477 275312 237489
rect 291952 237477 291958 237489
rect 292010 237477 292016 237529
rect 292048 237477 292054 237529
rect 292106 237517 292112 237529
rect 302416 237517 302422 237529
rect 292106 237489 302422 237517
rect 292106 237477 292112 237489
rect 302416 237477 302422 237489
rect 302474 237477 302480 237529
rect 304048 237477 304054 237529
rect 304106 237517 304112 237529
rect 307984 237517 307990 237529
rect 304106 237489 307990 237517
rect 304106 237477 304112 237489
rect 307984 237477 307990 237489
rect 308042 237477 308048 237529
rect 319984 237477 319990 237529
rect 320042 237517 320048 237529
rect 334384 237517 334390 237529
rect 320042 237489 334390 237517
rect 320042 237477 320048 237489
rect 334384 237477 334390 237489
rect 334442 237477 334448 237529
rect 334498 237489 338462 237517
rect 227344 237403 227350 237455
rect 227402 237443 227408 237455
rect 233584 237443 233590 237455
rect 227402 237415 233590 237443
rect 227402 237403 227408 237415
rect 233584 237403 233590 237415
rect 233642 237403 233648 237455
rect 238768 237403 238774 237455
rect 238826 237443 238832 237455
rect 259408 237443 259414 237455
rect 238826 237415 259414 237443
rect 238826 237403 238832 237415
rect 259408 237403 259414 237415
rect 259466 237403 259472 237455
rect 275440 237403 275446 237455
rect 275498 237443 275504 237455
rect 287152 237443 287158 237455
rect 275498 237415 287158 237443
rect 275498 237403 275504 237415
rect 287152 237403 287158 237415
rect 287210 237403 287216 237455
rect 287248 237403 287254 237455
rect 287306 237443 287312 237455
rect 287920 237443 287926 237455
rect 287306 237415 287926 237443
rect 287306 237403 287312 237415
rect 287920 237403 287926 237415
rect 287978 237403 287984 237455
rect 292528 237443 292534 237455
rect 290242 237415 292534 237443
rect 221008 237329 221014 237381
rect 221066 237369 221072 237381
rect 247216 237369 247222 237381
rect 221066 237341 247222 237369
rect 221066 237329 221072 237341
rect 247216 237329 247222 237341
rect 247274 237329 247280 237381
rect 273232 237329 273238 237381
rect 273290 237369 273296 237381
rect 290242 237369 290270 237415
rect 292528 237403 292534 237415
rect 292586 237403 292592 237455
rect 295312 237403 295318 237455
rect 295370 237443 295376 237455
rect 303664 237443 303670 237455
rect 295370 237415 303670 237443
rect 295370 237403 295376 237415
rect 303664 237403 303670 237415
rect 303722 237403 303728 237455
rect 316048 237403 316054 237455
rect 316106 237443 316112 237455
rect 334498 237443 334526 237489
rect 316106 237415 334526 237443
rect 338434 237443 338462 237489
rect 338512 237477 338518 237529
rect 338570 237517 338576 237529
rect 342736 237517 342742 237529
rect 338570 237489 342742 237517
rect 338570 237477 338576 237489
rect 342736 237477 342742 237489
rect 342794 237477 342800 237529
rect 376624 237517 376630 237529
rect 371746 237489 376630 237517
rect 371746 237443 371774 237489
rect 376624 237477 376630 237489
rect 376682 237477 376688 237529
rect 376720 237477 376726 237529
rect 376778 237517 376784 237529
rect 384592 237517 384598 237529
rect 376778 237489 384598 237517
rect 376778 237477 376784 237489
rect 384592 237477 384598 237489
rect 384650 237477 384656 237529
rect 338434 237415 371774 237443
rect 316106 237403 316112 237415
rect 372592 237403 372598 237455
rect 372650 237443 372656 237455
rect 395344 237443 395350 237455
rect 372650 237415 395350 237443
rect 372650 237403 372656 237415
rect 395344 237403 395350 237415
rect 395402 237403 395408 237455
rect 273290 237341 290270 237369
rect 273290 237329 273296 237341
rect 290320 237329 290326 237381
rect 290378 237369 290384 237381
rect 301456 237369 301462 237381
rect 290378 237341 301462 237369
rect 290378 237329 290384 237341
rect 301456 237329 301462 237341
rect 301514 237329 301520 237381
rect 316816 237329 316822 237381
rect 316874 237369 316880 237381
rect 338512 237369 338518 237381
rect 316874 237341 338518 237369
rect 316874 237329 316880 237341
rect 338512 237329 338518 237341
rect 338570 237329 338576 237381
rect 342832 237329 342838 237381
rect 342890 237369 342896 237381
rect 360880 237369 360886 237381
rect 342890 237341 360886 237369
rect 342890 237329 342896 237341
rect 360880 237329 360886 237341
rect 360938 237329 360944 237381
rect 369040 237329 369046 237381
rect 369098 237369 369104 237381
rect 387664 237369 387670 237381
rect 369098 237341 387670 237369
rect 369098 237329 369104 237341
rect 387664 237329 387670 237341
rect 387722 237329 387728 237381
rect 221104 237255 221110 237307
rect 221162 237295 221168 237307
rect 246544 237295 246550 237307
rect 221162 237267 246550 237295
rect 221162 237255 221168 237267
rect 246544 237255 246550 237267
rect 246602 237255 246608 237307
rect 275824 237255 275830 237307
rect 275882 237295 275888 237307
rect 286576 237295 286582 237307
rect 275882 237267 286582 237295
rect 275882 237255 275888 237267
rect 286576 237255 286582 237267
rect 286634 237255 286640 237307
rect 290608 237295 290614 237307
rect 286690 237267 290614 237295
rect 274000 237181 274006 237233
rect 274058 237221 274064 237233
rect 286690 237221 286718 237267
rect 290608 237255 290614 237267
rect 290666 237255 290672 237307
rect 290704 237255 290710 237307
rect 290762 237295 290768 237307
rect 293968 237295 293974 237307
rect 290762 237267 293974 237295
rect 290762 237255 290768 237267
rect 293968 237255 293974 237267
rect 294026 237255 294032 237307
rect 294064 237255 294070 237307
rect 294122 237295 294128 237307
rect 296464 237295 296470 237307
rect 294122 237267 296470 237295
rect 294122 237255 294128 237267
rect 296464 237255 296470 237267
rect 296522 237255 296528 237307
rect 300208 237255 300214 237307
rect 300266 237295 300272 237307
rect 305872 237295 305878 237307
rect 300266 237267 305878 237295
rect 300266 237255 300272 237267
rect 305872 237255 305878 237267
rect 305930 237255 305936 237307
rect 305968 237255 305974 237307
rect 306026 237295 306032 237307
rect 318448 237295 318454 237307
rect 306026 237267 318454 237295
rect 306026 237255 306032 237267
rect 318448 237255 318454 237267
rect 318506 237255 318512 237307
rect 321808 237255 321814 237307
rect 321866 237295 321872 237307
rect 328528 237295 328534 237307
rect 321866 237267 328534 237295
rect 321866 237255 321872 237267
rect 328528 237255 328534 237267
rect 328586 237255 328592 237307
rect 328720 237255 328726 237307
rect 328778 237295 328784 237307
rect 330736 237295 330742 237307
rect 328778 237267 330742 237295
rect 328778 237255 328784 237267
rect 330736 237255 330742 237267
rect 330794 237255 330800 237307
rect 331792 237255 331798 237307
rect 331850 237295 331856 237307
rect 344752 237295 344758 237307
rect 331850 237267 344758 237295
rect 331850 237255 331856 237267
rect 344752 237255 344758 237267
rect 344810 237255 344816 237307
rect 379984 237255 379990 237307
rect 380042 237295 380048 237307
rect 385360 237295 385366 237307
rect 380042 237267 385366 237295
rect 380042 237255 380048 237267
rect 385360 237255 385366 237267
rect 385418 237255 385424 237307
rect 274058 237193 286718 237221
rect 274058 237181 274064 237193
rect 289264 237181 289270 237233
rect 289322 237221 289328 237233
rect 300976 237221 300982 237233
rect 289322 237193 300982 237221
rect 289322 237181 289328 237193
rect 300976 237181 300982 237193
rect 301034 237181 301040 237233
rect 318160 237181 318166 237233
rect 318218 237221 318224 237233
rect 330832 237221 330838 237233
rect 318218 237193 330838 237221
rect 318218 237181 318224 237193
rect 330832 237181 330838 237193
rect 330890 237181 330896 237233
rect 332848 237181 332854 237233
rect 332906 237221 332912 237233
rect 362224 237221 362230 237233
rect 332906 237193 362230 237221
rect 332906 237181 332912 237193
rect 362224 237181 362230 237193
rect 362282 237181 362288 237233
rect 362800 237181 362806 237233
rect 362858 237221 362864 237233
rect 382288 237221 382294 237233
rect 362858 237193 382294 237221
rect 362858 237181 362864 237193
rect 382288 237181 382294 237193
rect 382346 237181 382352 237233
rect 225520 237107 225526 237159
rect 225578 237147 225584 237159
rect 237328 237147 237334 237159
rect 225578 237119 237334 237147
rect 225578 237107 225584 237119
rect 237328 237107 237334 237119
rect 237386 237107 237392 237159
rect 278512 237107 278518 237159
rect 278570 237147 278576 237159
rect 280720 237147 280726 237159
rect 278570 237119 280726 237147
rect 278570 237107 278576 237119
rect 280720 237107 280726 237119
rect 280778 237107 280784 237159
rect 285808 237107 285814 237159
rect 285866 237147 285872 237159
rect 285866 237119 288350 237147
rect 285866 237107 285872 237119
rect 286384 237033 286390 237085
rect 286442 237073 286448 237085
rect 288322 237073 288350 237119
rect 288400 237107 288406 237159
rect 288458 237147 288464 237159
rect 300592 237147 300598 237159
rect 288458 237119 300598 237147
rect 288458 237107 288464 237119
rect 300592 237107 300598 237119
rect 300650 237107 300656 237159
rect 316240 237107 316246 237159
rect 316298 237147 316304 237159
rect 324112 237147 324118 237159
rect 316298 237119 324118 237147
rect 316298 237107 316304 237119
rect 324112 237107 324118 237119
rect 324170 237107 324176 237159
rect 327856 237107 327862 237159
rect 327914 237147 327920 237159
rect 351472 237147 351478 237159
rect 327914 237119 351478 237147
rect 327914 237107 327920 237119
rect 351472 237107 351478 237119
rect 351530 237107 351536 237159
rect 351568 237107 351574 237159
rect 351626 237147 351632 237159
rect 358768 237147 358774 237159
rect 351626 237119 358774 237147
rect 351626 237107 351632 237119
rect 358768 237107 358774 237119
rect 358826 237107 358832 237159
rect 372976 237107 372982 237159
rect 373034 237147 373040 237159
rect 396208 237147 396214 237159
rect 373034 237119 396214 237147
rect 373034 237107 373040 237119
rect 396208 237107 396214 237119
rect 396266 237107 396272 237159
rect 299536 237073 299542 237085
rect 286442 237045 288254 237073
rect 288322 237045 299542 237073
rect 286442 237033 286448 237045
rect 224080 236959 224086 237011
rect 224138 236999 224144 237011
rect 240400 236999 240406 237011
rect 224138 236971 240406 236999
rect 224138 236959 224144 236971
rect 240400 236959 240406 236971
rect 240458 236959 240464 237011
rect 271888 236959 271894 237011
rect 271946 236999 271952 237011
rect 288112 236999 288118 237011
rect 271946 236971 288118 236999
rect 271946 236959 271952 236971
rect 288112 236959 288118 236971
rect 288170 236959 288176 237011
rect 288226 236999 288254 237045
rect 299536 237033 299542 237045
rect 299594 237033 299600 237085
rect 318256 237033 318262 237085
rect 318314 237073 318320 237085
rect 328720 237073 328726 237085
rect 318314 237045 328726 237073
rect 318314 237033 318320 237045
rect 328720 237033 328726 237045
rect 328778 237033 328784 237085
rect 328816 237033 328822 237085
rect 328874 237073 328880 237085
rect 353488 237073 353494 237085
rect 328874 237045 353494 237073
rect 328874 237033 328880 237045
rect 353488 237033 353494 237045
rect 353546 237033 353552 237085
rect 288226 236971 296798 236999
rect 276784 236885 276790 236937
rect 276842 236925 276848 236937
rect 295216 236925 295222 236937
rect 276842 236897 295222 236925
rect 276842 236885 276848 236897
rect 295216 236885 295222 236897
rect 295274 236885 295280 236937
rect 296770 236925 296798 236971
rect 296848 236959 296854 237011
rect 296906 236999 296912 237011
rect 304432 236999 304438 237011
rect 296906 236971 304438 236999
rect 296906 236959 296912 236971
rect 304432 236959 304438 236971
rect 304490 236959 304496 237011
rect 308002 236971 315518 236999
rect 299632 236925 299638 236937
rect 296770 236897 299638 236925
rect 299632 236885 299638 236897
rect 299690 236885 299696 236937
rect 225040 236811 225046 236863
rect 225098 236851 225104 236863
rect 238576 236851 238582 236863
rect 225098 236823 238582 236851
rect 225098 236811 225104 236823
rect 238576 236811 238582 236823
rect 238634 236811 238640 236863
rect 282736 236811 282742 236863
rect 282794 236851 282800 236863
rect 285232 236851 285238 236863
rect 282794 236823 285238 236851
rect 282794 236811 282800 236823
rect 285232 236811 285238 236823
rect 285290 236811 285296 236863
rect 285904 236811 285910 236863
rect 285962 236851 285968 236863
rect 288976 236851 288982 236863
rect 285962 236823 288982 236851
rect 285962 236811 285968 236823
rect 288976 236811 288982 236823
rect 289034 236811 289040 236863
rect 291760 236811 291766 236863
rect 291818 236851 291824 236863
rect 308002 236851 308030 236971
rect 315490 236925 315518 236971
rect 316336 236959 316342 237011
rect 316394 236999 316400 237011
rect 325840 236999 325846 237011
rect 316394 236971 325846 236999
rect 316394 236959 316400 236971
rect 325840 236959 325846 236971
rect 325898 236959 325904 237011
rect 327472 236959 327478 237011
rect 327530 236999 327536 237011
rect 350704 236999 350710 237011
rect 327530 236971 350710 236999
rect 327530 236959 327536 236971
rect 350704 236959 350710 236971
rect 350762 236959 350768 237011
rect 319312 236925 319318 236937
rect 315490 236897 319318 236925
rect 319312 236885 319318 236897
rect 319370 236885 319376 236937
rect 327088 236885 327094 236937
rect 327146 236925 327152 236937
rect 349744 236925 349750 236937
rect 327146 236897 349750 236925
rect 327146 236885 327152 236897
rect 349744 236885 349750 236897
rect 349802 236885 349808 236937
rect 291818 236823 308030 236851
rect 291818 236811 291824 236823
rect 324784 236811 324790 236863
rect 324842 236851 324848 236863
rect 331792 236851 331798 236863
rect 324842 236823 331798 236851
rect 324842 236811 324848 236823
rect 331792 236811 331798 236823
rect 331850 236811 331856 236863
rect 331888 236811 331894 236863
rect 331946 236851 331952 236863
rect 339664 236851 339670 236863
rect 331946 236823 339670 236851
rect 331946 236811 331952 236823
rect 339664 236811 339670 236823
rect 339722 236811 339728 236863
rect 370768 236811 370774 236863
rect 370826 236851 370832 236863
rect 381136 236851 381142 236863
rect 370826 236823 381142 236851
rect 370826 236811 370832 236823
rect 381136 236811 381142 236823
rect 381194 236811 381200 236863
rect 239056 236737 239062 236789
rect 239114 236777 239120 236789
rect 259120 236777 259126 236789
rect 239114 236749 259126 236777
rect 239114 236737 239120 236749
rect 259120 236737 259126 236749
rect 259178 236737 259184 236789
rect 274864 236737 274870 236789
rect 274922 236777 274928 236789
rect 288496 236777 288502 236789
rect 274922 236749 288502 236777
rect 274922 236737 274928 236749
rect 288496 236737 288502 236749
rect 288554 236737 288560 236789
rect 291664 236737 291670 236789
rect 291722 236777 291728 236789
rect 305968 236777 305974 236789
rect 291722 236749 305974 236777
rect 291722 236737 291728 236749
rect 305968 236737 305974 236749
rect 306026 236737 306032 236789
rect 306448 236737 306454 236789
rect 306506 236777 306512 236789
rect 308944 236777 308950 236789
rect 306506 236749 308950 236777
rect 306506 236737 306512 236749
rect 308944 236737 308950 236749
rect 309002 236737 309008 236789
rect 325648 236737 325654 236789
rect 325706 236777 325712 236789
rect 330448 236777 330454 236789
rect 325706 236749 330454 236777
rect 325706 236737 325712 236749
rect 330448 236737 330454 236749
rect 330506 236737 330512 236789
rect 330544 236737 330550 236789
rect 330602 236777 330608 236789
rect 345232 236777 345238 236789
rect 330602 236749 345238 236777
rect 330602 236737 330608 236749
rect 345232 236737 345238 236749
rect 345290 236737 345296 236789
rect 42160 236663 42166 236715
rect 42218 236703 42224 236715
rect 42352 236703 42358 236715
rect 42218 236675 42358 236703
rect 42218 236663 42224 236675
rect 42352 236663 42358 236675
rect 42410 236663 42416 236715
rect 260752 236663 260758 236715
rect 260810 236703 260816 236715
rect 269488 236703 269494 236715
rect 260810 236675 269494 236703
rect 260810 236663 260816 236675
rect 269488 236663 269494 236675
rect 269546 236663 269552 236715
rect 274096 236663 274102 236715
rect 274154 236703 274160 236715
rect 289744 236703 289750 236715
rect 274154 236675 289750 236703
rect 274154 236663 274160 236675
rect 289744 236663 289750 236675
rect 289802 236663 289808 236715
rect 293488 236663 293494 236715
rect 293546 236703 293552 236715
rect 299728 236703 299734 236715
rect 293546 236675 299734 236703
rect 293546 236663 293552 236675
rect 299728 236663 299734 236675
rect 299786 236663 299792 236715
rect 315376 236703 315382 236715
rect 308866 236675 315382 236703
rect 236464 236589 236470 236641
rect 236522 236629 236528 236641
rect 238864 236629 238870 236641
rect 236522 236601 238870 236629
rect 236522 236589 236528 236601
rect 238864 236589 238870 236601
rect 238922 236589 238928 236641
rect 276400 236589 276406 236641
rect 276458 236629 276464 236641
rect 294832 236629 294838 236641
rect 276458 236601 294838 236629
rect 276458 236589 276464 236601
rect 294832 236589 294838 236601
rect 294890 236589 294896 236641
rect 295792 236589 295798 236641
rect 295850 236629 295856 236641
rect 308866 236629 308894 236675
rect 315376 236663 315382 236675
rect 315434 236663 315440 236715
rect 324016 236663 324022 236715
rect 324074 236703 324080 236715
rect 324074 236675 328478 236703
rect 324074 236663 324080 236675
rect 295850 236601 308894 236629
rect 295850 236589 295856 236601
rect 313648 236589 313654 236641
rect 313706 236629 313712 236641
rect 313840 236629 313846 236641
rect 313706 236601 313846 236629
rect 313706 236589 313712 236601
rect 313840 236589 313846 236601
rect 313898 236589 313904 236641
rect 325264 236589 325270 236641
rect 325322 236629 325328 236641
rect 328336 236629 328342 236641
rect 325322 236601 328342 236629
rect 325322 236589 325328 236601
rect 328336 236589 328342 236601
rect 328394 236589 328400 236641
rect 328450 236629 328478 236675
rect 328528 236663 328534 236715
rect 328586 236703 328592 236715
rect 347440 236703 347446 236715
rect 328586 236675 347446 236703
rect 328586 236663 328592 236675
rect 347440 236663 347446 236675
rect 347498 236663 347504 236715
rect 380176 236663 380182 236715
rect 380234 236703 380240 236715
rect 390160 236703 390166 236715
rect 380234 236675 390166 236703
rect 380234 236663 380240 236675
rect 390160 236663 390166 236675
rect 390218 236663 390224 236715
rect 420496 236663 420502 236715
rect 420554 236703 420560 236715
rect 440560 236703 440566 236715
rect 420554 236675 440566 236703
rect 420554 236663 420560 236675
rect 440560 236663 440566 236675
rect 440618 236663 440624 236715
rect 460816 236663 460822 236715
rect 460874 236703 460880 236715
rect 480880 236703 480886 236715
rect 460874 236675 480886 236703
rect 460874 236663 460880 236675
rect 480880 236663 480886 236675
rect 480938 236663 480944 236715
rect 343024 236629 343030 236641
rect 328450 236601 343030 236629
rect 343024 236589 343030 236601
rect 343082 236589 343088 236641
rect 258160 236515 258166 236567
rect 258218 236555 258224 236567
rect 264016 236555 264022 236567
rect 258218 236527 264022 236555
rect 258218 236515 258224 236527
rect 264016 236515 264022 236527
rect 264074 236515 264080 236567
rect 278704 236515 278710 236567
rect 278762 236555 278768 236567
rect 278762 236527 289214 236555
rect 278762 236515 278768 236527
rect 268336 236441 268342 236493
rect 268394 236481 268400 236493
rect 268394 236453 285182 236481
rect 268394 236441 268400 236453
rect 217456 236367 217462 236419
rect 217514 236407 217520 236419
rect 221776 236407 221782 236419
rect 217514 236379 221782 236407
rect 217514 236367 217520 236379
rect 221776 236367 221782 236379
rect 221834 236367 221840 236419
rect 263056 236367 263062 236419
rect 263114 236407 263120 236419
rect 269008 236407 269014 236419
rect 263114 236379 269014 236407
rect 263114 236367 263120 236379
rect 269008 236367 269014 236379
rect 269066 236367 269072 236419
rect 278416 236367 278422 236419
rect 278474 236407 278480 236419
rect 281200 236407 281206 236419
rect 278474 236379 281206 236407
rect 278474 236367 278480 236379
rect 281200 236367 281206 236379
rect 281258 236367 281264 236419
rect 273520 236293 273526 236345
rect 273578 236333 273584 236345
rect 281584 236333 281590 236345
rect 273578 236305 281590 236333
rect 273578 236293 273584 236305
rect 281584 236293 281590 236305
rect 281642 236293 281648 236345
rect 283312 236293 283318 236345
rect 283370 236333 283376 236345
rect 285040 236333 285046 236345
rect 283370 236305 285046 236333
rect 283370 236293 283376 236305
rect 285040 236293 285046 236305
rect 285098 236293 285104 236345
rect 285154 236333 285182 236453
rect 285232 236367 285238 236419
rect 285290 236407 285296 236419
rect 289186 236407 289214 236527
rect 289264 236515 289270 236567
rect 289322 236555 289328 236567
rect 311440 236555 311446 236567
rect 289322 236527 311446 236555
rect 289322 236515 289328 236527
rect 311440 236515 311446 236527
rect 311498 236515 311504 236567
rect 318064 236515 318070 236567
rect 318122 236555 318128 236567
rect 335632 236555 335638 236567
rect 318122 236527 335638 236555
rect 318122 236515 318128 236527
rect 335632 236515 335638 236527
rect 335690 236515 335696 236567
rect 638032 236515 638038 236567
rect 638090 236555 638096 236567
rect 650512 236555 650518 236567
rect 638090 236527 650518 236555
rect 638090 236515 638096 236527
rect 650512 236515 650518 236527
rect 650570 236515 650576 236567
rect 291280 236441 291286 236493
rect 291338 236481 291344 236493
rect 317584 236481 317590 236493
rect 291338 236453 317590 236481
rect 291338 236441 291344 236453
rect 317584 236441 317590 236453
rect 317642 236441 317648 236493
rect 320368 236441 320374 236493
rect 320426 236481 320432 236493
rect 334960 236481 334966 236493
rect 320426 236453 334966 236481
rect 320426 236441 320432 236453
rect 334960 236441 334966 236453
rect 335018 236441 335024 236493
rect 637552 236441 637558 236493
rect 637610 236481 637616 236493
rect 650224 236481 650230 236493
rect 637610 236453 650230 236481
rect 637610 236441 637616 236453
rect 650224 236441 650230 236453
rect 650282 236441 650288 236493
rect 296176 236407 296182 236419
rect 285290 236379 288830 236407
rect 289186 236379 296182 236407
rect 285290 236367 285296 236379
rect 288112 236333 288118 236345
rect 285154 236305 288118 236333
rect 288112 236293 288118 236305
rect 288170 236293 288176 236345
rect 288802 236333 288830 236379
rect 296176 236367 296182 236379
rect 296234 236367 296240 236419
rect 300784 236367 300790 236419
rect 300842 236407 300848 236419
rect 306256 236407 306262 236419
rect 300842 236379 306262 236407
rect 300842 236367 300848 236379
rect 306256 236367 306262 236379
rect 306314 236367 306320 236419
rect 322480 236367 322486 236419
rect 322538 236407 322544 236419
rect 339856 236407 339862 236419
rect 322538 236379 339862 236407
rect 322538 236367 322544 236379
rect 339856 236367 339862 236379
rect 339914 236367 339920 236419
rect 637936 236367 637942 236419
rect 637994 236407 638000 236419
rect 650320 236407 650326 236419
rect 637994 236379 650326 236407
rect 637994 236367 638000 236379
rect 650320 236367 650326 236379
rect 650378 236367 650384 236419
rect 297808 236333 297814 236345
rect 288802 236305 297814 236333
rect 297808 236293 297814 236305
rect 297866 236293 297872 236345
rect 330448 236293 330454 236345
rect 330506 236333 330512 236345
rect 346960 236333 346966 236345
rect 330506 236305 346966 236333
rect 330506 236293 330512 236305
rect 346960 236293 346966 236305
rect 347018 236293 347024 236345
rect 639184 236293 639190 236345
rect 639242 236333 639248 236345
rect 649840 236333 649846 236345
rect 639242 236305 649846 236333
rect 639242 236293 639248 236305
rect 649840 236293 649846 236305
rect 649898 236293 649904 236345
rect 144016 236219 144022 236271
rect 144074 236259 144080 236271
rect 168400 236259 168406 236271
rect 144074 236231 168406 236259
rect 144074 236219 144080 236231
rect 168400 236219 168406 236231
rect 168458 236219 168464 236271
rect 225904 236219 225910 236271
rect 225962 236259 225968 236271
rect 236752 236259 236758 236271
rect 225962 236231 236758 236259
rect 225962 236219 225968 236231
rect 236752 236219 236758 236231
rect 236810 236219 236816 236271
rect 236944 236219 236950 236271
rect 237002 236259 237008 236271
rect 238960 236259 238966 236271
rect 237002 236231 238966 236259
rect 237002 236219 237008 236231
rect 238960 236219 238966 236231
rect 239018 236219 239024 236271
rect 271408 236219 271414 236271
rect 271466 236259 271472 236271
rect 290704 236259 290710 236271
rect 271466 236231 290710 236259
rect 271466 236219 271472 236231
rect 290704 236219 290710 236231
rect 290762 236219 290768 236271
rect 290800 236219 290806 236271
rect 290858 236259 290864 236271
rect 296944 236259 296950 236271
rect 290858 236231 296950 236259
rect 290858 236219 290864 236231
rect 296944 236219 296950 236231
rect 297002 236219 297008 236271
rect 328336 236219 328342 236271
rect 328394 236259 328400 236271
rect 345904 236259 345910 236271
rect 328394 236231 345910 236259
rect 328394 236219 328400 236231
rect 345904 236219 345910 236231
rect 345962 236219 345968 236271
rect 368944 236219 368950 236271
rect 369002 236259 369008 236271
rect 387088 236259 387094 236271
rect 369002 236231 387094 236259
rect 369002 236219 369008 236231
rect 387088 236219 387094 236231
rect 387146 236219 387152 236271
rect 638800 236219 638806 236271
rect 638858 236259 638864 236271
rect 649648 236259 649654 236271
rect 638858 236231 649654 236259
rect 638858 236219 638864 236231
rect 649648 236219 649654 236231
rect 649706 236219 649712 236271
rect 144112 236145 144118 236197
rect 144170 236185 144176 236197
rect 174160 236185 174166 236197
rect 144170 236157 174166 236185
rect 144170 236145 144176 236157
rect 174160 236145 174166 236157
rect 174218 236145 174224 236197
rect 210256 236145 210262 236197
rect 210314 236185 210320 236197
rect 210736 236185 210742 236197
rect 210314 236157 210742 236185
rect 210314 236145 210320 236157
rect 210736 236145 210742 236157
rect 210794 236185 210800 236197
rect 213040 236185 213046 236197
rect 210794 236157 213046 236185
rect 210794 236145 210800 236157
rect 213040 236145 213046 236157
rect 213098 236145 213104 236197
rect 284368 236145 284374 236197
rect 284426 236185 284432 236197
rect 298768 236185 298774 236197
rect 284426 236157 298774 236185
rect 284426 236145 284432 236157
rect 298768 236145 298774 236157
rect 298826 236145 298832 236197
rect 315952 236145 315958 236197
rect 316010 236185 316016 236197
rect 324208 236185 324214 236197
rect 316010 236157 324214 236185
rect 316010 236145 316016 236157
rect 324208 236145 324214 236157
rect 324266 236145 324272 236197
rect 547120 236145 547126 236197
rect 547178 236185 547184 236197
rect 549232 236185 549238 236197
rect 547178 236157 549238 236185
rect 547178 236145 547184 236157
rect 549232 236145 549238 236157
rect 549290 236145 549296 236197
rect 639760 236145 639766 236197
rect 639818 236185 639824 236197
rect 649936 236185 649942 236197
rect 639818 236157 649942 236185
rect 639818 236145 639824 236157
rect 649936 236145 649942 236157
rect 649994 236145 650000 236197
rect 265648 236071 265654 236123
rect 265706 236111 265712 236123
rect 308368 236111 308374 236123
rect 265706 236083 308374 236111
rect 265706 236071 265712 236083
rect 308368 236071 308374 236083
rect 308426 236071 308432 236123
rect 319696 236071 319702 236123
rect 319754 236111 319760 236123
rect 339760 236111 339766 236123
rect 319754 236083 339766 236111
rect 319754 236071 319760 236083
rect 339760 236071 339766 236083
rect 339818 236071 339824 236123
rect 264880 235997 264886 236049
rect 264938 236037 264944 236049
rect 309904 236037 309910 236049
rect 264938 236009 309910 236037
rect 264938 235997 264944 236009
rect 309904 235997 309910 236009
rect 309962 235997 309968 236049
rect 312976 235997 312982 236049
rect 313034 236037 313040 236049
rect 369616 236037 369622 236049
rect 313034 236009 369622 236037
rect 313034 235997 313040 236009
rect 369616 235997 369622 236009
rect 369674 235997 369680 236049
rect 265072 235923 265078 235975
rect 265130 235963 265136 235975
rect 339376 235963 339382 235975
rect 265130 235935 339382 235963
rect 265130 235923 265136 235935
rect 339376 235923 339382 235935
rect 339434 235923 339440 235975
rect 381904 235923 381910 235975
rect 381962 235963 381968 235975
rect 390928 235963 390934 235975
rect 381962 235935 390934 235963
rect 381962 235923 381968 235935
rect 390928 235923 390934 235935
rect 390986 235923 390992 235975
rect 235696 235849 235702 235901
rect 235754 235889 235760 235901
rect 266128 235889 266134 235901
rect 235754 235861 266134 235889
rect 235754 235849 235760 235861
rect 266128 235849 266134 235861
rect 266186 235849 266192 235901
rect 266800 235849 266806 235901
rect 266858 235889 266864 235901
rect 340336 235889 340342 235901
rect 266858 235861 340342 235889
rect 266858 235849 266864 235861
rect 340336 235849 340342 235861
rect 340394 235849 340400 235901
rect 263728 235775 263734 235827
rect 263786 235815 263792 235827
rect 338896 235815 338902 235827
rect 263786 235787 338902 235815
rect 263786 235775 263792 235787
rect 338896 235775 338902 235787
rect 338954 235775 338960 235827
rect 261904 235701 261910 235753
rect 261962 235741 261968 235753
rect 338128 235741 338134 235753
rect 261962 235713 338134 235741
rect 261962 235701 261968 235713
rect 338128 235701 338134 235713
rect 338186 235701 338192 235753
rect 258928 235627 258934 235679
rect 258986 235667 258992 235679
rect 336688 235667 336694 235679
rect 258986 235639 336694 235667
rect 258986 235627 258992 235639
rect 336688 235627 336694 235639
rect 336746 235627 336752 235679
rect 260560 235553 260566 235605
rect 260618 235593 260624 235605
rect 337168 235593 337174 235605
rect 260618 235565 337174 235593
rect 260618 235553 260624 235565
rect 337168 235553 337174 235565
rect 337226 235553 337232 235605
rect 257296 235479 257302 235531
rect 257354 235519 257360 235531
rect 335920 235519 335926 235531
rect 257354 235491 335926 235519
rect 257354 235479 257360 235491
rect 335920 235479 335926 235491
rect 335978 235479 335984 235531
rect 42160 235405 42166 235457
rect 42218 235445 42224 235457
rect 43120 235445 43126 235457
rect 42218 235417 43126 235445
rect 42218 235405 42224 235417
rect 43120 235405 43126 235417
rect 43178 235405 43184 235457
rect 236080 235405 236086 235457
rect 236138 235445 236144 235457
rect 265456 235445 265462 235457
rect 236138 235417 265462 235445
rect 236138 235405 236144 235417
rect 265456 235405 265462 235417
rect 265514 235405 265520 235457
rect 273616 235405 273622 235457
rect 273674 235445 273680 235457
rect 356656 235445 356662 235457
rect 273674 235417 356662 235445
rect 273674 235405 273680 235417
rect 356656 235405 356662 235417
rect 356714 235405 356720 235457
rect 246064 235331 246070 235383
rect 246122 235371 246128 235383
rect 353584 235371 353590 235383
rect 246122 235343 353590 235371
rect 246122 235331 246128 235343
rect 353584 235331 353590 235343
rect 353642 235331 353648 235383
rect 247792 235257 247798 235309
rect 247850 235297 247856 235309
rect 354832 235297 354838 235309
rect 247850 235269 354838 235297
rect 247850 235257 247856 235269
rect 354832 235257 354838 235269
rect 354890 235257 354896 235309
rect 246352 235183 246358 235235
rect 246410 235223 246416 235235
rect 354352 235223 354358 235235
rect 246410 235195 354358 235223
rect 246410 235183 246416 235195
rect 354352 235183 354358 235195
rect 354410 235183 354416 235235
rect 242032 235109 242038 235161
rect 242090 235149 242096 235161
rect 352144 235149 352150 235161
rect 242090 235121 352150 235149
rect 242090 235109 242096 235121
rect 352144 235109 352150 235121
rect 352202 235109 352208 235161
rect 241840 235035 241846 235087
rect 241898 235075 241904 235087
rect 349936 235075 349942 235087
rect 241898 235047 349942 235075
rect 241898 235035 241904 235047
rect 349936 235035 349942 235047
rect 349994 235035 350000 235087
rect 243280 234961 243286 235013
rect 243338 235001 243344 235013
rect 352624 235001 352630 235013
rect 243338 234973 352630 235001
rect 243338 234961 243344 234973
rect 352624 234961 352630 234973
rect 352682 234961 352688 235013
rect 244144 234887 244150 234939
rect 244202 234927 244208 234939
rect 351376 234927 351382 234939
rect 244202 234899 351382 234927
rect 244202 234887 244208 234899
rect 351376 234887 351382 234899
rect 351434 234887 351440 234939
rect 42160 234813 42166 234865
rect 42218 234853 42224 234865
rect 42928 234853 42934 234865
rect 42218 234825 42934 234853
rect 42218 234813 42224 234825
rect 42928 234813 42934 234825
rect 42986 234813 42992 234865
rect 241648 234813 241654 234865
rect 241706 234853 241712 234865
rect 350416 234853 350422 234865
rect 241706 234825 350422 234853
rect 241706 234813 241712 234825
rect 350416 234813 350422 234825
rect 350474 234813 350480 234865
rect 230608 234739 230614 234791
rect 230666 234779 230672 234791
rect 346960 234779 346966 234791
rect 230666 234751 346966 234779
rect 230666 234739 230672 234751
rect 346960 234739 346966 234751
rect 347018 234739 347024 234791
rect 227920 234665 227926 234717
rect 227978 234705 227984 234717
rect 345520 234705 345526 234717
rect 227978 234677 345526 234705
rect 227978 234665 227984 234677
rect 345520 234665 345526 234677
rect 345578 234665 345584 234717
rect 260848 234591 260854 234643
rect 260906 234631 260912 234643
rect 268432 234631 268438 234643
rect 260906 234603 268438 234631
rect 260906 234591 260912 234603
rect 268432 234591 268438 234603
rect 268490 234591 268496 234643
rect 282448 234591 282454 234643
rect 282506 234631 282512 234643
rect 322768 234631 322774 234643
rect 282506 234603 322774 234631
rect 282506 234591 282512 234603
rect 322768 234591 322774 234603
rect 322826 234591 322832 234643
rect 266992 234517 266998 234569
rect 267050 234557 267056 234569
rect 305680 234557 305686 234569
rect 267050 234529 305686 234557
rect 267050 234517 267056 234529
rect 305680 234517 305686 234529
rect 305738 234517 305744 234569
rect 282832 234443 282838 234495
rect 282890 234483 282896 234495
rect 321904 234483 321910 234495
rect 282890 234455 321910 234483
rect 282890 234443 282896 234455
rect 321904 234443 321910 234455
rect 321962 234443 321968 234495
rect 267472 234369 267478 234421
rect 267530 234409 267536 234421
rect 304240 234409 304246 234421
rect 267530 234381 304246 234409
rect 267530 234369 267536 234381
rect 304240 234369 304246 234381
rect 304298 234369 304304 234421
rect 271600 234295 271606 234347
rect 271658 234335 271664 234347
rect 309424 234335 309430 234347
rect 271658 234307 309430 234335
rect 271658 234295 271664 234307
rect 309424 234295 309430 234307
rect 309482 234295 309488 234347
rect 284656 234221 284662 234273
rect 284714 234261 284720 234273
rect 317968 234261 317974 234273
rect 284714 234233 317974 234261
rect 284714 234221 284720 234233
rect 317968 234221 317974 234233
rect 318026 234221 318032 234273
rect 42064 234147 42070 234199
rect 42122 234187 42128 234199
rect 42448 234187 42454 234199
rect 42122 234159 42454 234187
rect 42122 234147 42128 234159
rect 42448 234147 42454 234159
rect 42506 234147 42512 234199
rect 277264 234147 277270 234199
rect 277322 234187 277328 234199
rect 279760 234187 279766 234199
rect 277322 234159 279766 234187
rect 277322 234147 277328 234159
rect 279760 234147 279766 234159
rect 279818 234147 279824 234199
rect 284272 234147 284278 234199
rect 284330 234187 284336 234199
rect 319120 234187 319126 234199
rect 284330 234159 319126 234187
rect 284330 234147 284336 234159
rect 319120 234147 319126 234159
rect 319178 234147 319184 234199
rect 268816 234073 268822 234125
rect 268874 234113 268880 234125
rect 301936 234113 301942 234125
rect 268874 234085 301942 234113
rect 268874 234073 268880 234085
rect 301936 234073 301942 234085
rect 301994 234073 302000 234125
rect 269584 233999 269590 234051
rect 269642 234039 269648 234051
rect 300304 234039 300310 234051
rect 269642 234011 300310 234039
rect 269642 233999 269648 234011
rect 300304 233999 300310 234011
rect 300362 233999 300368 234051
rect 285136 233925 285142 233977
rect 285194 233965 285200 233977
rect 316528 233965 316534 233977
rect 285194 233937 316534 233965
rect 285194 233925 285200 233937
rect 316528 233925 316534 233937
rect 316586 233925 316592 233977
rect 287344 233851 287350 233903
rect 287402 233891 287408 233903
rect 289264 233891 289270 233903
rect 287402 233863 289270 233891
rect 287402 233851 287408 233863
rect 289264 233851 289270 233863
rect 289322 233851 289328 233903
rect 292528 233851 292534 233903
rect 292586 233891 292592 233903
rect 320560 233891 320566 233903
rect 292586 233863 320566 233891
rect 292586 233851 292592 233863
rect 320560 233851 320566 233863
rect 320618 233851 320624 233903
rect 285040 233777 285046 233829
rect 285098 233817 285104 233829
rect 288208 233817 288214 233829
rect 285098 233789 288214 233817
rect 285098 233777 285104 233789
rect 288208 233777 288214 233789
rect 288266 233777 288272 233829
rect 293104 233777 293110 233829
rect 293162 233817 293168 233829
rect 321424 233817 321430 233829
rect 293162 233789 321430 233817
rect 293162 233777 293168 233789
rect 321424 233777 321430 233789
rect 321482 233777 321488 233829
rect 262336 233703 262342 233755
rect 262394 233743 262400 233755
rect 268912 233743 268918 233755
rect 262394 233715 268918 233743
rect 262394 233703 262400 233715
rect 268912 233703 268918 233715
rect 268970 233703 268976 233755
rect 270064 233703 270070 233755
rect 270122 233743 270128 233755
rect 298576 233743 298582 233755
rect 270122 233715 298582 233743
rect 270122 233703 270128 233715
rect 298576 233703 298582 233715
rect 298634 233703 298640 233755
rect 305584 233703 305590 233755
rect 305642 233743 305648 233755
rect 308704 233743 308710 233755
rect 305642 233715 308710 233743
rect 305642 233703 305648 233715
rect 308704 233703 308710 233715
rect 308762 233703 308768 233755
rect 367936 233703 367942 233755
rect 367994 233743 368000 233755
rect 376720 233743 376726 233755
rect 367994 233715 376726 233743
rect 367994 233703 368000 233715
rect 376720 233703 376726 233715
rect 376778 233703 376784 233755
rect 270640 233629 270646 233681
rect 270698 233669 270704 233681
rect 298480 233669 298486 233681
rect 270698 233641 298486 233669
rect 270698 233629 270704 233641
rect 298480 233629 298486 233641
rect 298538 233629 298544 233681
rect 317008 233669 317014 233681
rect 307906 233641 317014 233669
rect 208144 233555 208150 233607
rect 208202 233595 208208 233607
rect 213520 233595 213526 233607
rect 208202 233567 213526 233595
rect 208202 233555 208208 233567
rect 213520 233555 213526 233567
rect 213578 233555 213584 233607
rect 269104 233555 269110 233607
rect 269162 233595 269168 233607
rect 297040 233595 297046 233607
rect 269162 233567 297046 233595
rect 269162 233555 269168 233567
rect 297040 233555 297046 233567
rect 297098 233555 297104 233607
rect 209968 233481 209974 233533
rect 210026 233521 210032 233533
rect 213136 233521 213142 233533
rect 210026 233493 213142 233521
rect 210026 233481 210032 233493
rect 213136 233481 213142 233493
rect 213194 233481 213200 233533
rect 213904 233481 213910 233533
rect 213962 233481 213968 233533
rect 290896 233481 290902 233533
rect 290954 233521 290960 233533
rect 307906 233521 307934 233641
rect 317008 233629 317014 233641
rect 317066 233629 317072 233681
rect 290954 233493 307934 233521
rect 290954 233481 290960 233493
rect 210064 233407 210070 233459
rect 210122 233447 210128 233459
rect 213922 233447 213950 233481
rect 210122 233419 213950 233447
rect 210122 233407 210128 233419
rect 144016 233259 144022 233311
rect 144074 233299 144080 233311
rect 171280 233299 171286 233311
rect 144074 233271 171286 233299
rect 144074 233259 144080 233271
rect 171280 233259 171286 233271
rect 171338 233259 171344 233311
rect 645520 233185 645526 233237
rect 645578 233225 645584 233237
rect 649744 233225 649750 233237
rect 645578 233197 649750 233225
rect 645578 233185 645584 233197
rect 649744 233185 649750 233197
rect 649802 233185 649808 233237
rect 645232 233111 645238 233163
rect 645290 233151 645296 233163
rect 650416 233151 650422 233163
rect 645290 233123 650422 233151
rect 645290 233111 645296 233123
rect 650416 233111 650422 233123
rect 650474 233111 650480 233163
rect 645328 232963 645334 233015
rect 645386 233003 645392 233015
rect 650128 233003 650134 233015
rect 645386 232975 650134 233003
rect 645386 232963 645392 232975
rect 650128 232963 650134 232975
rect 650186 232963 650192 233015
rect 645136 232889 645142 232941
rect 645194 232929 645200 232941
rect 650608 232929 650614 232941
rect 645194 232901 650614 232929
rect 645194 232889 645200 232901
rect 650608 232889 650614 232901
rect 650666 232889 650672 232941
rect 144016 230521 144022 230573
rect 144074 230561 144080 230573
rect 151120 230561 151126 230573
rect 144074 230533 151126 230561
rect 144074 230521 144080 230533
rect 151120 230521 151126 230533
rect 151178 230521 151184 230573
rect 144112 230447 144118 230499
rect 144170 230487 144176 230499
rect 165520 230487 165526 230499
rect 144170 230459 165526 230487
rect 144170 230447 144176 230459
rect 165520 230447 165526 230459
rect 165578 230447 165584 230499
rect 205744 228153 205750 228205
rect 205802 228193 205808 228205
rect 205936 228193 205942 228205
rect 205802 228165 205942 228193
rect 205802 228153 205808 228165
rect 205936 228153 205942 228165
rect 205994 228153 206000 228205
rect 205264 227857 205270 227909
rect 205322 227897 205328 227909
rect 205648 227897 205654 227909
rect 205322 227869 205654 227897
rect 205322 227857 205328 227869
rect 205648 227857 205654 227869
rect 205706 227857 205712 227909
rect 210256 227783 210262 227835
rect 210314 227783 210320 227835
rect 144016 227709 144022 227761
rect 144074 227749 144080 227761
rect 188560 227749 188566 227761
rect 144074 227721 188566 227749
rect 144074 227709 144080 227721
rect 188560 227709 188566 227721
rect 188618 227709 188624 227761
rect 144112 227635 144118 227687
rect 144170 227675 144176 227687
rect 194320 227675 194326 227687
rect 144170 227647 194326 227675
rect 144170 227635 144176 227647
rect 194320 227635 194326 227647
rect 194378 227635 194384 227687
rect 210274 227613 210302 227783
rect 144208 227561 144214 227613
rect 144266 227601 144272 227613
rect 197200 227601 197206 227613
rect 144266 227573 197206 227601
rect 144266 227561 144272 227573
rect 197200 227561 197206 227573
rect 197258 227561 197264 227613
rect 210256 227561 210262 227613
rect 210314 227561 210320 227613
rect 146800 226377 146806 226429
rect 146858 226417 146864 226429
rect 156880 226417 156886 226429
rect 146858 226389 156886 226417
rect 146858 226377 146864 226389
rect 156880 226377 156886 226389
rect 156938 226377 156944 226429
rect 206608 226417 206614 226429
rect 205762 226389 206614 226417
rect 205762 225973 205790 226389
rect 206608 226377 206614 226389
rect 206666 226377 206672 226429
rect 206320 226229 206326 226281
rect 206378 226269 206384 226281
rect 206608 226269 206614 226281
rect 206378 226241 206614 226269
rect 206378 226229 206384 226241
rect 206608 226229 206614 226241
rect 206666 226229 206672 226281
rect 205840 226155 205846 226207
rect 205898 226195 205904 226207
rect 207088 226195 207094 226207
rect 205898 226167 207094 226195
rect 205898 226155 205904 226167
rect 207088 226155 207094 226167
rect 207146 226155 207152 226207
rect 206032 226081 206038 226133
rect 206090 226121 206096 226133
rect 206320 226121 206326 226133
rect 206090 226093 206326 226121
rect 206090 226081 206096 226093
rect 206320 226081 206326 226093
rect 206378 226081 206384 226133
rect 205840 225973 205846 225985
rect 205762 225945 205846 225973
rect 205840 225933 205846 225945
rect 205898 225933 205904 225985
rect 666832 225045 666838 225097
rect 666890 225085 666896 225097
rect 674704 225085 674710 225097
rect 666890 225057 674710 225085
rect 666890 225045 666896 225057
rect 674704 225045 674710 225057
rect 674762 225045 674768 225097
rect 146128 224675 146134 224727
rect 146186 224715 146192 224727
rect 200080 224715 200086 224727
rect 146186 224687 200086 224715
rect 146186 224675 146192 224687
rect 200080 224675 200086 224687
rect 200138 224675 200144 224727
rect 141040 224601 141046 224653
rect 141098 224641 141104 224653
rect 204496 224641 204502 224653
rect 141098 224613 204502 224641
rect 141098 224601 141104 224613
rect 204496 224601 204502 224613
rect 204554 224601 204560 224653
rect 146416 224527 146422 224579
rect 146474 224567 146480 224579
rect 204592 224567 204598 224579
rect 146474 224539 204598 224567
rect 146474 224527 146480 224539
rect 204592 224527 204598 224539
rect 204650 224527 204656 224579
rect 149680 224453 149686 224505
rect 149738 224493 149744 224505
rect 204688 224493 204694 224505
rect 149738 224465 204694 224493
rect 149738 224453 149744 224465
rect 204688 224453 204694 224465
rect 204746 224453 204752 224505
rect 152560 224379 152566 224431
rect 152618 224419 152624 224431
rect 204784 224419 204790 224431
rect 152618 224391 204790 224419
rect 152618 224379 152624 224391
rect 204784 224379 204790 224391
rect 204842 224379 204848 224431
rect 669520 224305 669526 224357
rect 669578 224345 669584 224357
rect 674416 224345 674422 224357
rect 669578 224317 674422 224345
rect 669578 224305 669584 224317
rect 674416 224305 674422 224317
rect 674474 224305 674480 224357
rect 669616 224009 669622 224061
rect 669674 224049 669680 224061
rect 674704 224049 674710 224061
rect 669674 224021 674710 224049
rect 669674 224009 669680 224021
rect 674704 224009 674710 224021
rect 674762 224009 674768 224061
rect 146704 221937 146710 221989
rect 146762 221977 146768 221989
rect 177040 221977 177046 221989
rect 146762 221949 177046 221977
rect 146762 221937 146768 221949
rect 177040 221937 177046 221949
rect 177098 221937 177104 221989
rect 146800 221863 146806 221915
rect 146858 221903 146864 221915
rect 179920 221903 179926 221915
rect 146858 221875 179926 221903
rect 146858 221863 146864 221875
rect 179920 221863 179926 221875
rect 179978 221863 179984 221915
rect 144400 221789 144406 221841
rect 144458 221829 144464 221841
rect 182896 221829 182902 221841
rect 144458 221801 182902 221829
rect 144458 221789 144464 221801
rect 182896 221789 182902 221801
rect 182954 221789 182960 221841
rect 155440 221715 155446 221767
rect 155498 221755 155504 221767
rect 204496 221755 204502 221767
rect 155498 221727 204502 221755
rect 155498 221715 155504 221727
rect 204496 221715 204502 221727
rect 204554 221715 204560 221767
rect 161200 221641 161206 221693
rect 161258 221681 161264 221693
rect 204592 221681 204598 221693
rect 161258 221653 204598 221681
rect 161258 221641 161264 221653
rect 204592 221641 204598 221653
rect 204650 221641 204656 221693
rect 164080 221567 164086 221619
rect 164138 221607 164144 221619
rect 204688 221607 204694 221619
rect 164138 221579 204694 221607
rect 164138 221567 164144 221579
rect 204688 221567 204694 221579
rect 204746 221567 204752 221619
rect 166960 221493 166966 221545
rect 167018 221533 167024 221545
rect 204784 221533 204790 221545
rect 167018 221505 204790 221533
rect 167018 221493 167024 221505
rect 204784 221493 204790 221505
rect 204842 221493 204848 221545
rect 169840 221419 169846 221471
rect 169898 221459 169904 221471
rect 204880 221459 204886 221471
rect 169898 221431 204886 221459
rect 169898 221419 169904 221431
rect 204880 221419 204886 221431
rect 204938 221419 204944 221471
rect 144400 218903 144406 218955
rect 144458 218943 144464 218955
rect 174256 218943 174262 218955
rect 144458 218915 174262 218943
rect 144458 218903 144464 218915
rect 174256 218903 174262 218915
rect 174314 218903 174320 218955
rect 175600 218829 175606 218881
rect 175658 218869 175664 218881
rect 204496 218869 204502 218881
rect 175658 218841 204502 218869
rect 175658 218829 175664 218841
rect 204496 218829 204502 218841
rect 204554 218829 204560 218881
rect 178480 218755 178486 218807
rect 178538 218795 178544 218807
rect 204592 218795 204598 218807
rect 178538 218767 204598 218795
rect 178538 218755 178544 218767
rect 204592 218755 204598 218767
rect 204650 218755 204656 218807
rect 181360 218681 181366 218733
rect 181418 218721 181424 218733
rect 204688 218721 204694 218733
rect 181418 218693 204694 218721
rect 181418 218681 181424 218693
rect 204688 218681 204694 218693
rect 204746 218681 204752 218733
rect 184240 218607 184246 218659
rect 184298 218647 184304 218659
rect 204784 218647 204790 218659
rect 184298 218619 204790 218647
rect 184298 218607 184304 218619
rect 204784 218607 204790 218619
rect 204842 218607 204848 218659
rect 146800 216535 146806 216587
rect 146858 216575 146864 216587
rect 154000 216575 154006 216587
rect 146858 216547 154006 216575
rect 146858 216535 146864 216547
rect 154000 216535 154006 216547
rect 154058 216535 154064 216587
rect 42736 216313 42742 216365
rect 42794 216353 42800 216365
rect 44944 216353 44950 216365
rect 42794 216325 44950 216353
rect 42794 216313 42800 216325
rect 44944 216313 44950 216325
rect 45002 216313 45008 216365
rect 146224 216091 146230 216143
rect 146282 216131 146288 216143
rect 146282 216103 146366 216131
rect 146282 216091 146288 216103
rect 146338 216069 146366 216103
rect 146320 216017 146326 216069
rect 146378 216017 146384 216069
rect 187120 215943 187126 215995
rect 187178 215983 187184 215995
rect 204496 215983 204502 215995
rect 187178 215955 204502 215983
rect 187178 215943 187184 215955
rect 204496 215943 204502 215955
rect 204554 215943 204560 215995
rect 192880 215869 192886 215921
rect 192938 215909 192944 215921
rect 204592 215909 204598 215921
rect 192938 215881 204598 215909
rect 192938 215869 192944 215881
rect 204592 215869 204598 215881
rect 204650 215869 204656 215921
rect 42736 215721 42742 215773
rect 42794 215761 42800 215773
rect 45136 215761 45142 215773
rect 42794 215733 45142 215761
rect 42794 215721 42800 215733
rect 45136 215721 45142 215733
rect 45194 215721 45200 215773
rect 42736 215203 42742 215255
rect 42794 215243 42800 215255
rect 44848 215243 44854 215255
rect 42794 215215 44854 215243
rect 42794 215203 42800 215215
rect 44848 215203 44854 215215
rect 44906 215203 44912 215255
rect 146800 213205 146806 213257
rect 146858 213245 146864 213257
rect 168496 213245 168502 213257
rect 146858 213217 168502 213245
rect 146858 213205 146864 213217
rect 168496 213205 168502 213217
rect 168554 213205 168560 213257
rect 144400 213131 144406 213183
rect 144458 213171 144464 213183
rect 171376 213171 171382 213183
rect 144458 213143 171382 213171
rect 144458 213131 144464 213143
rect 171376 213131 171382 213143
rect 171434 213131 171440 213183
rect 145264 210245 145270 210297
rect 145322 210285 145328 210297
rect 148240 210285 148246 210297
rect 145322 210257 148246 210285
rect 145322 210245 145328 210257
rect 148240 210245 148246 210257
rect 148298 210245 148304 210297
rect 645616 210245 645622 210297
rect 645674 210285 645680 210297
rect 677008 210285 677014 210297
rect 645674 210257 677014 210285
rect 645674 210245 645680 210257
rect 677008 210245 677014 210257
rect 677066 210245 677072 210297
rect 146608 207433 146614 207485
rect 146666 207473 146672 207485
rect 165616 207473 165622 207485
rect 146666 207445 165622 207473
rect 146666 207433 146672 207445
rect 165616 207433 165622 207445
rect 165674 207433 165680 207485
rect 146800 207359 146806 207411
rect 146858 207399 146864 207411
rect 203056 207399 203062 207411
rect 146858 207371 203062 207399
rect 146858 207359 146864 207371
rect 203056 207359 203062 207371
rect 203114 207359 203120 207411
rect 40240 206767 40246 206819
rect 40298 206807 40304 206819
rect 41776 206807 41782 206819
rect 40298 206779 41782 206807
rect 40298 206767 40304 206779
rect 41776 206767 41782 206779
rect 41834 206767 41840 206819
rect 675472 205953 675478 206005
rect 675530 205953 675536 206005
rect 675490 205783 675518 205953
rect 675472 205731 675478 205783
rect 675530 205731 675536 205783
rect 675184 204991 675190 205043
rect 675242 205031 675248 205043
rect 675472 205031 675478 205043
rect 675242 205003 675478 205031
rect 675242 204991 675248 205003
rect 675472 204991 675478 205003
rect 675530 204991 675536 205043
rect 42736 204399 42742 204451
rect 42794 204439 42800 204451
rect 50320 204439 50326 204451
rect 42794 204411 50326 204439
rect 42794 204399 42800 204411
rect 50320 204399 50326 204411
rect 50378 204399 50384 204451
rect 674896 204399 674902 204451
rect 674954 204439 674960 204451
rect 675376 204439 675382 204451
rect 674954 204411 675382 204439
rect 674954 204399 674960 204411
rect 675376 204399 675382 204411
rect 675434 204399 675440 204451
rect 674992 202179 674998 202231
rect 675050 202219 675056 202231
rect 675280 202219 675286 202231
rect 675050 202191 675286 202219
rect 675050 202179 675056 202191
rect 675280 202179 675286 202191
rect 675338 202179 675344 202231
rect 675088 202031 675094 202083
rect 675146 202071 675152 202083
rect 675280 202071 675286 202083
rect 675146 202043 675286 202071
rect 675146 202031 675152 202043
rect 675280 202031 675286 202043
rect 675338 202031 675344 202083
rect 145840 201661 145846 201713
rect 145898 201701 145904 201713
rect 162640 201701 162646 201713
rect 145898 201673 162646 201701
rect 145898 201661 145904 201673
rect 162640 201661 162646 201673
rect 162698 201661 162704 201713
rect 144016 201587 144022 201639
rect 144074 201627 144080 201639
rect 202960 201627 202966 201639
rect 144074 201599 202966 201627
rect 144074 201587 144080 201599
rect 202960 201587 202966 201599
rect 203018 201587 203024 201639
rect 645904 201587 645910 201639
rect 645962 201627 645968 201639
rect 646096 201627 646102 201639
rect 645962 201599 646102 201627
rect 645962 201587 645968 201599
rect 646096 201587 646102 201599
rect 646154 201587 646160 201639
rect 674224 201291 674230 201343
rect 674282 201331 674288 201343
rect 675376 201331 675382 201343
rect 674282 201303 675382 201331
rect 674282 201291 674288 201303
rect 675376 201291 675382 201303
rect 675434 201291 675440 201343
rect 41968 201069 41974 201121
rect 42026 201109 42032 201121
rect 42352 201109 42358 201121
rect 42026 201081 42358 201109
rect 42026 201069 42032 201081
rect 42352 201069 42358 201081
rect 42410 201069 42416 201121
rect 674800 200329 674806 200381
rect 674858 200369 674864 200381
rect 675280 200369 675286 200381
rect 674858 200341 675286 200369
rect 674858 200329 674864 200341
rect 675280 200329 675286 200341
rect 675338 200329 675344 200381
rect 40144 198997 40150 199049
rect 40202 199037 40208 199049
rect 42160 199037 42166 199049
rect 40202 199009 42166 199037
rect 40202 198997 40208 199009
rect 42160 198997 42166 199009
rect 42218 198997 42224 199049
rect 144016 198923 144022 198975
rect 144074 198963 144080 198975
rect 159760 198963 159766 198975
rect 144074 198935 159766 198963
rect 144074 198923 144080 198935
rect 159760 198923 159766 198935
rect 159818 198923 159824 198975
rect 40048 198849 40054 198901
rect 40106 198889 40112 198901
rect 43120 198889 43126 198901
rect 40106 198861 43126 198889
rect 40106 198849 40112 198861
rect 43120 198849 43126 198861
rect 43178 198849 43184 198901
rect 40240 198701 40246 198753
rect 40298 198741 40304 198753
rect 43120 198741 43126 198753
rect 40298 198713 43126 198741
rect 40298 198701 40304 198713
rect 43120 198701 43126 198713
rect 43178 198701 43184 198753
rect 144496 198701 144502 198753
rect 144554 198741 144560 198753
rect 191440 198741 191446 198753
rect 144554 198713 191446 198741
rect 144554 198701 144560 198713
rect 191440 198701 191446 198713
rect 191498 198701 191504 198753
rect 674704 197739 674710 197791
rect 674762 197779 674768 197791
rect 675376 197779 675382 197791
rect 674762 197751 675382 197779
rect 674762 197739 674768 197751
rect 675376 197739 675382 197751
rect 675434 197739 675440 197791
rect 41776 197369 41782 197421
rect 41834 197369 41840 197421
rect 41794 197199 41822 197369
rect 145072 197221 145078 197273
rect 145130 197261 145136 197273
rect 146224 197261 146230 197273
rect 145130 197233 146230 197261
rect 145130 197221 145136 197233
rect 146224 197221 146230 197233
rect 146282 197221 146288 197273
rect 41776 197147 41782 197199
rect 41834 197147 41840 197199
rect 674512 196999 674518 197051
rect 674570 197039 674576 197051
rect 675472 197039 675478 197051
rect 674570 197011 675478 197039
rect 674570 196999 674576 197011
rect 675472 196999 675478 197011
rect 675530 196999 675536 197051
rect 674608 196555 674614 196607
rect 674666 196595 674672 196607
rect 675376 196595 675382 196607
rect 674666 196567 675382 196595
rect 674666 196555 674672 196567
rect 675376 196555 675382 196567
rect 675434 196555 675440 196607
rect 144688 195815 144694 195867
rect 144746 195855 144752 195867
rect 185680 195855 185686 195867
rect 144746 195827 185686 195855
rect 144746 195815 144752 195827
rect 185680 195815 185686 195827
rect 185738 195815 185744 195867
rect 42160 195297 42166 195349
rect 42218 195337 42224 195349
rect 42352 195337 42358 195349
rect 42218 195309 42358 195337
rect 42218 195297 42224 195309
rect 42352 195297 42358 195309
rect 42410 195297 42416 195349
rect 42064 194483 42070 194535
rect 42122 194523 42128 194535
rect 50416 194523 50422 194535
rect 42122 194495 50422 194523
rect 42122 194483 42128 194495
rect 50416 194483 50422 194495
rect 50474 194483 50480 194535
rect 42064 193447 42070 193499
rect 42122 193487 42128 193499
rect 42928 193487 42934 193499
rect 42122 193459 42934 193487
rect 42122 193447 42128 193459
rect 42928 193447 42934 193459
rect 42986 193447 42992 193499
rect 42928 193299 42934 193351
rect 42986 193339 42992 193351
rect 43216 193339 43222 193351
rect 42986 193311 43222 193339
rect 42986 193299 42992 193311
rect 43216 193299 43222 193311
rect 43274 193299 43280 193351
rect 42160 192189 42166 192241
rect 42218 192229 42224 192241
rect 43024 192229 43030 192241
rect 42218 192201 43030 192229
rect 42218 192189 42224 192201
rect 43024 192189 43030 192201
rect 43082 192189 43088 192241
rect 42064 191449 42070 191501
rect 42122 191489 42128 191501
rect 42352 191489 42358 191501
rect 42122 191461 42358 191489
rect 42122 191449 42128 191461
rect 42352 191449 42358 191461
rect 42410 191449 42416 191501
rect 42160 191005 42166 191057
rect 42218 191045 42224 191057
rect 43120 191045 43126 191057
rect 42218 191017 43126 191045
rect 42218 191005 42224 191017
rect 43120 191005 43126 191017
rect 43178 191005 43184 191057
rect 144304 190191 144310 190243
rect 144362 190231 144368 190243
rect 151216 190231 151222 190243
rect 144362 190203 151222 190231
rect 144362 190191 144368 190203
rect 151216 190191 151222 190203
rect 151274 190191 151280 190243
rect 144016 190117 144022 190169
rect 144074 190157 144080 190169
rect 148432 190157 148438 190169
rect 144074 190129 148438 190157
rect 144074 190117 144080 190129
rect 148432 190117 148438 190129
rect 148490 190117 148496 190169
rect 42256 187897 42262 187949
rect 42314 187937 42320 187949
rect 42928 187937 42934 187949
rect 42314 187909 42934 187937
rect 42314 187897 42320 187909
rect 42928 187897 42934 187909
rect 42986 187897 42992 187949
rect 210256 187379 210262 187431
rect 210314 187379 210320 187431
rect 144016 187231 144022 187283
rect 144074 187271 144080 187283
rect 197296 187271 197302 187283
rect 144074 187243 197302 187271
rect 144074 187231 144080 187243
rect 197296 187231 197302 187243
rect 197354 187231 197360 187283
rect 210274 187135 210302 187379
rect 42160 187083 42166 187135
rect 42218 187123 42224 187135
rect 42832 187123 42838 187135
rect 42218 187095 42838 187123
rect 42218 187083 42224 187095
rect 42832 187083 42838 187095
rect 42890 187083 42896 187135
rect 210256 187083 210262 187135
rect 210314 187083 210320 187135
rect 645712 187083 645718 187135
rect 645770 187123 645776 187135
rect 646096 187123 646102 187135
rect 645770 187095 646102 187123
rect 645770 187083 645776 187095
rect 646096 187083 646102 187095
rect 646154 187083 646160 187135
rect 146320 184567 146326 184619
rect 146378 184607 146384 184619
rect 146800 184607 146806 184619
rect 146378 184579 146806 184607
rect 146378 184567 146384 184579
rect 146800 184567 146806 184579
rect 146858 184567 146864 184619
rect 144016 184345 144022 184397
rect 144074 184385 144080 184397
rect 194416 184385 194422 184397
rect 144074 184357 194422 184385
rect 144074 184345 144080 184357
rect 194416 184345 194422 184357
rect 194474 184345 194480 184397
rect 144208 181533 144214 181585
rect 144266 181573 144272 181585
rect 146608 181573 146614 181585
rect 144266 181545 146614 181573
rect 144266 181533 144272 181545
rect 146608 181533 146614 181545
rect 146666 181533 146672 181585
rect 144016 181459 144022 181511
rect 144074 181499 144080 181511
rect 188656 181499 188662 181511
rect 144074 181471 188662 181499
rect 144074 181459 144080 181471
rect 188656 181459 188662 181471
rect 188714 181459 188720 181511
rect 661072 179313 661078 179365
rect 661130 179353 661136 179365
rect 674416 179353 674422 179365
rect 661130 179325 674422 179353
rect 661130 179313 661136 179325
rect 674416 179313 674422 179325
rect 674474 179313 674480 179365
rect 666640 178795 666646 178847
rect 666698 178835 666704 178847
rect 674416 178835 674422 178847
rect 666698 178807 674422 178835
rect 666698 178795 666704 178807
rect 674416 178795 674422 178807
rect 674474 178795 674480 178847
rect 144112 178647 144118 178699
rect 144170 178687 144176 178699
rect 148528 178687 148534 178699
rect 144170 178659 148534 178687
rect 144170 178647 144176 178659
rect 148528 178647 148534 178659
rect 148586 178647 148592 178699
rect 655216 178647 655222 178699
rect 655274 178687 655280 178699
rect 674704 178687 674710 178699
rect 655274 178659 674710 178687
rect 655274 178647 655280 178659
rect 674704 178647 674710 178659
rect 674762 178647 674768 178699
rect 144016 178573 144022 178625
rect 144074 178613 144080 178625
rect 191536 178613 191542 178625
rect 144074 178585 191542 178613
rect 144074 178573 144080 178585
rect 191536 178573 191542 178585
rect 191594 178573 191600 178625
rect 146512 176131 146518 176183
rect 146570 176171 146576 176183
rect 146992 176171 146998 176183
rect 146570 176143 146998 176171
rect 146570 176131 146576 176143
rect 146992 176131 146998 176143
rect 147050 176131 147056 176183
rect 146224 175983 146230 176035
rect 146282 175983 146288 176035
rect 146242 175813 146270 175983
rect 146224 175761 146230 175813
rect 146282 175761 146288 175813
rect 144016 175687 144022 175739
rect 144074 175727 144080 175739
rect 185776 175727 185782 175739
rect 144074 175699 185782 175727
rect 144074 175687 144080 175699
rect 185776 175687 185782 175699
rect 185834 175687 185840 175739
rect 144496 175613 144502 175665
rect 144554 175653 144560 175665
rect 146800 175653 146806 175665
rect 144554 175625 146806 175653
rect 144554 175613 144560 175625
rect 146800 175613 146806 175625
rect 146858 175613 146864 175665
rect 144112 172875 144118 172927
rect 144170 172915 144176 172927
rect 148624 172915 148630 172927
rect 144170 172887 148630 172915
rect 144170 172875 144176 172887
rect 148624 172875 148630 172887
rect 148682 172875 148688 172927
rect 144016 172801 144022 172853
rect 144074 172841 144080 172853
rect 162736 172841 162742 172853
rect 144074 172813 162742 172841
rect 144074 172801 144080 172813
rect 162736 172801 162742 172813
rect 162794 172801 162800 172853
rect 144112 172727 144118 172779
rect 144170 172767 144176 172779
rect 146704 172767 146710 172779
rect 144170 172739 146710 172767
rect 144170 172727 144176 172739
rect 146704 172727 146710 172739
rect 146762 172727 146768 172779
rect 145072 172579 145078 172631
rect 145130 172619 145136 172631
rect 146704 172619 146710 172631
rect 145130 172591 146710 172619
rect 145130 172579 145136 172591
rect 146704 172579 146710 172591
rect 146762 172579 146768 172631
rect 144016 170211 144022 170263
rect 144074 170251 144080 170263
rect 159856 170251 159862 170263
rect 144074 170223 159862 170251
rect 144074 170211 144080 170223
rect 159856 170211 159862 170223
rect 159914 170211 159920 170263
rect 144016 167251 144022 167303
rect 144074 167291 144080 167303
rect 156976 167291 156982 167303
rect 144074 167263 156982 167291
rect 144074 167251 144080 167263
rect 156976 167251 156982 167263
rect 157034 167251 157040 167303
rect 647056 167251 647062 167303
rect 647114 167291 647120 167303
rect 674416 167291 674422 167303
rect 647114 167263 674422 167291
rect 647114 167251 647120 167263
rect 674416 167251 674422 167263
rect 674474 167251 674480 167303
rect 647824 167177 647830 167229
rect 647882 167217 647888 167229
rect 674608 167217 674614 167229
rect 647882 167189 674614 167217
rect 647882 167177 647888 167189
rect 674608 167177 674614 167189
rect 674666 167177 674672 167229
rect 647920 167103 647926 167155
rect 647978 167143 647984 167155
rect 674704 167143 674710 167155
rect 647978 167115 674710 167143
rect 647978 167103 647984 167115
rect 674704 167103 674710 167115
rect 674762 167103 674768 167155
rect 144880 165549 144886 165601
rect 144938 165589 144944 165601
rect 146800 165589 146806 165601
rect 144938 165561 146806 165589
rect 144938 165549 144944 165561
rect 146800 165549 146806 165561
rect 146858 165549 146864 165601
rect 144688 164143 144694 164195
rect 144746 164183 144752 164195
rect 148720 164183 148726 164195
rect 144746 164155 148726 164183
rect 144746 164143 144752 164155
rect 148720 164143 148726 164155
rect 148778 164143 148784 164195
rect 144688 161257 144694 161309
rect 144746 161297 144752 161309
rect 148816 161297 148822 161309
rect 144746 161269 148822 161297
rect 144746 161257 144752 161269
rect 148816 161257 148822 161269
rect 148874 161257 148880 161309
rect 645712 161257 645718 161309
rect 645770 161297 645776 161309
rect 645904 161297 645910 161309
rect 645770 161269 645910 161297
rect 645770 161257 645776 161269
rect 645904 161257 645910 161269
rect 645962 161257 645968 161309
rect 675568 160961 675574 161013
rect 675626 160961 675632 161013
rect 675760 160961 675766 161013
rect 675818 160961 675824 161013
rect 675586 160791 675614 160961
rect 675568 160739 675574 160791
rect 675626 160739 675632 160791
rect 675778 160051 675806 160961
rect 675760 159999 675766 160051
rect 675818 159999 675824 160051
rect 674032 159407 674038 159459
rect 674090 159447 674096 159459
rect 675376 159447 675382 159459
rect 674090 159419 675382 159447
rect 674090 159407 674096 159419
rect 675376 159407 675382 159419
rect 675434 159407 675440 159459
rect 144688 158445 144694 158497
rect 144746 158485 144752 158497
rect 148912 158485 148918 158497
rect 144746 158457 148918 158485
rect 144746 158445 144752 158457
rect 148912 158445 148918 158457
rect 148970 158445 148976 158497
rect 674800 157705 674806 157757
rect 674858 157745 674864 157757
rect 675472 157745 675478 157757
rect 674858 157717 675478 157745
rect 674858 157705 674864 157717
rect 675472 157705 675478 157717
rect 675530 157705 675536 157757
rect 146128 155781 146134 155833
rect 146186 155821 146192 155833
rect 146704 155821 146710 155833
rect 146186 155793 146710 155821
rect 146186 155781 146192 155793
rect 146704 155781 146710 155793
rect 146762 155781 146768 155833
rect 144112 155707 144118 155759
rect 144170 155747 144176 155759
rect 146416 155747 146422 155759
rect 144170 155719 146422 155747
rect 144170 155707 144176 155719
rect 146416 155707 146422 155719
rect 146474 155707 146480 155759
rect 144496 155633 144502 155685
rect 144554 155673 144560 155685
rect 146704 155673 146710 155685
rect 144554 155645 146710 155673
rect 144554 155633 144560 155645
rect 146704 155633 146710 155645
rect 146762 155633 146768 155685
rect 146896 155633 146902 155685
rect 146954 155673 146960 155685
rect 149008 155673 149014 155685
rect 146954 155645 149014 155673
rect 146954 155633 146960 155645
rect 149008 155633 149014 155645
rect 149066 155633 149072 155685
rect 144688 155559 144694 155611
rect 144746 155599 144752 155611
rect 200176 155599 200182 155611
rect 144746 155571 200182 155599
rect 144746 155559 144752 155571
rect 200176 155559 200182 155571
rect 200234 155559 200240 155611
rect 144688 153117 144694 153169
rect 144746 153157 144752 153169
rect 146704 153157 146710 153169
rect 144746 153129 146710 153157
rect 144746 153117 144752 153129
rect 146704 153117 146710 153129
rect 146762 153117 146768 153169
rect 146800 152747 146806 152799
rect 146858 152787 146864 152799
rect 180016 152787 180022 152799
rect 146858 152759 180022 152787
rect 146858 152747 146864 152759
rect 180016 152747 180022 152759
rect 180074 152747 180080 152799
rect 144496 152673 144502 152725
rect 144554 152713 144560 152725
rect 182992 152713 182998 152725
rect 144554 152685 182998 152713
rect 144554 152673 144560 152685
rect 182992 152673 182998 152685
rect 183050 152673 183056 152725
rect 674320 152599 674326 152651
rect 674378 152639 674384 152651
rect 675376 152639 675382 152651
rect 674378 152611 675382 152639
rect 674378 152599 674384 152611
rect 675376 152599 675382 152611
rect 675434 152599 675440 152651
rect 674512 151489 674518 151541
rect 674570 151529 674576 151541
rect 675376 151529 675382 151541
rect 674570 151501 675382 151529
rect 674570 151489 674576 151501
rect 675376 151489 675382 151501
rect 675434 151489 675440 151541
rect 144496 149861 144502 149913
rect 144554 149901 144560 149913
rect 149104 149901 149110 149913
rect 144554 149873 149110 149901
rect 144554 149861 144560 149873
rect 149104 149861 149110 149873
rect 149162 149861 149168 149913
rect 146800 149787 146806 149839
rect 146858 149827 146864 149839
rect 177136 149827 177142 149839
rect 146858 149799 177142 149827
rect 146858 149787 146864 149799
rect 177136 149787 177142 149799
rect 177194 149787 177200 149839
rect 144496 146975 144502 147027
rect 144554 147015 144560 147027
rect 149200 147015 149206 147027
rect 144554 146987 149206 147015
rect 144554 146975 144560 146987
rect 149200 146975 149206 146987
rect 149258 146975 149264 147027
rect 210256 146975 210262 147027
rect 210314 146975 210320 147027
rect 146800 146901 146806 146953
rect 146858 146941 146864 146953
rect 174352 146941 174358 146953
rect 146858 146913 174358 146941
rect 146858 146901 146864 146913
rect 174352 146901 174358 146913
rect 174410 146901 174416 146953
rect 210274 146583 210302 146975
rect 645712 146901 645718 146953
rect 645770 146941 645776 146953
rect 645770 146913 645854 146941
rect 645770 146901 645776 146913
rect 645826 146879 645854 146913
rect 645808 146827 645814 146879
rect 645866 146827 645872 146879
rect 210256 146531 210262 146583
rect 210314 146531 210320 146583
rect 144496 146383 144502 146435
rect 144554 146423 144560 146435
rect 144688 146423 144694 146435
rect 144554 146395 144694 146423
rect 144554 146383 144560 146395
rect 144688 146383 144694 146395
rect 144746 146383 144752 146435
rect 144112 146235 144118 146287
rect 144170 146275 144176 146287
rect 144688 146275 144694 146287
rect 144170 146247 144694 146275
rect 144170 146235 144176 146247
rect 144688 146235 144694 146247
rect 144746 146235 144752 146287
rect 144016 144015 144022 144067
rect 144074 144055 144080 144067
rect 154096 144055 154102 144067
rect 144074 144027 154102 144055
rect 144074 144015 144080 144027
rect 154096 144015 154102 144027
rect 154154 144015 154160 144067
rect 144016 142535 144022 142587
rect 144074 142575 144080 142587
rect 149296 142575 149302 142587
rect 144074 142547 149302 142575
rect 144074 142535 144080 142547
rect 149296 142535 149302 142547
rect 149354 142535 149360 142587
rect 144016 141129 144022 141181
rect 144074 141169 144080 141181
rect 171472 141169 171478 141181
rect 144074 141141 171478 141169
rect 144074 141129 144080 141141
rect 171472 141129 171478 141141
rect 171530 141129 171536 141181
rect 143728 139723 143734 139775
rect 143786 139763 143792 139775
rect 144496 139763 144502 139775
rect 143786 139735 144502 139763
rect 143786 139723 143792 139735
rect 144496 139723 144502 139735
rect 144554 139723 144560 139775
rect 144304 139575 144310 139627
rect 144362 139615 144368 139627
rect 144496 139615 144502 139627
rect 144362 139587 144502 139615
rect 144362 139575 144368 139587
rect 144496 139575 144502 139587
rect 144554 139575 144560 139627
rect 144304 138391 144310 138443
rect 144362 138431 144368 138443
rect 168592 138431 168598 138443
rect 144362 138403 168598 138431
rect 144362 138391 144368 138403
rect 168592 138391 168598 138403
rect 168650 138391 168656 138443
rect 144016 138243 144022 138295
rect 144074 138283 144080 138295
rect 208720 138283 208726 138295
rect 144074 138255 208726 138283
rect 144074 138243 144080 138255
rect 208720 138243 208726 138255
rect 208778 138243 208784 138295
rect 146992 136023 146998 136075
rect 147050 136063 147056 136075
rect 149392 136063 149398 136075
rect 147050 136035 149398 136063
rect 147050 136023 147056 136035
rect 149392 136023 149398 136035
rect 149450 136023 149456 136075
rect 161200 135579 161206 135631
rect 161258 135619 161264 135631
rect 166960 135619 166966 135631
rect 161258 135591 166966 135619
rect 161258 135579 161264 135591
rect 166960 135579 166966 135591
rect 167018 135579 167024 135631
rect 167056 135579 167062 135631
rect 167114 135619 167120 135631
rect 167114 135591 171326 135619
rect 167114 135579 167120 135591
rect 171298 135545 171326 135591
rect 171298 135517 187166 135545
rect 146704 135357 146710 135409
rect 146762 135397 146768 135409
rect 146896 135397 146902 135409
rect 146762 135369 146902 135397
rect 146762 135357 146768 135369
rect 146896 135357 146902 135369
rect 146954 135357 146960 135409
rect 187138 135397 187166 135517
rect 187138 135369 204926 135397
rect 146128 135283 146134 135335
rect 146186 135323 146192 135335
rect 204898 135323 204926 135369
rect 208816 135323 208822 135335
rect 146186 135295 147038 135323
rect 204898 135295 208822 135323
rect 146186 135283 146192 135295
rect 147010 135261 147038 135295
rect 208816 135283 208822 135295
rect 208874 135283 208880 135335
rect 146992 135209 146998 135261
rect 147050 135209 147056 135261
rect 663760 133581 663766 133633
rect 663818 133621 663824 133633
rect 674416 133621 674422 133633
rect 663818 133593 674422 133621
rect 663818 133581 663824 133593
rect 674416 133581 674422 133593
rect 674474 133581 674480 133633
rect 144016 132915 144022 132967
rect 144074 132955 144080 132967
rect 165712 132955 165718 132967
rect 144074 132927 165718 132955
rect 144074 132915 144080 132927
rect 165712 132915 165718 132927
rect 165770 132915 165776 132967
rect 655312 132767 655318 132819
rect 655370 132807 655376 132819
rect 676912 132807 676918 132819
rect 655370 132779 676918 132807
rect 655370 132767 655376 132779
rect 676912 132767 676918 132779
rect 676970 132767 676976 132819
rect 655120 132619 655126 132671
rect 655178 132659 655184 132671
rect 676816 132659 676822 132671
rect 655178 132631 676822 132659
rect 655178 132619 655184 132631
rect 676816 132619 676822 132631
rect 676874 132619 676880 132671
rect 144304 132545 144310 132597
rect 144362 132585 144368 132597
rect 208912 132585 208918 132597
rect 144362 132557 208918 132585
rect 144362 132545 144368 132557
rect 208912 132545 208918 132557
rect 208970 132545 208976 132597
rect 144016 132471 144022 132523
rect 144074 132511 144080 132523
rect 209008 132511 209014 132523
rect 144074 132483 209014 132511
rect 144074 132471 144080 132483
rect 209008 132471 209014 132483
rect 209066 132471 209072 132523
rect 647728 132471 647734 132523
rect 647786 132511 647792 132523
rect 674416 132511 674422 132523
rect 647786 132483 674422 132511
rect 647786 132471 647792 132483
rect 674416 132471 674422 132483
rect 674474 132471 674480 132523
rect 143920 132397 143926 132449
rect 143978 132437 143984 132449
rect 144304 132437 144310 132449
rect 143978 132409 144310 132437
rect 143978 132397 143984 132409
rect 144304 132397 144310 132409
rect 144362 132397 144368 132449
rect 144112 129659 144118 129711
rect 144170 129699 144176 129711
rect 151504 129699 151510 129711
rect 144170 129671 151510 129699
rect 144170 129659 144176 129671
rect 151504 129659 151510 129671
rect 151562 129659 151568 129711
rect 144016 129585 144022 129637
rect 144074 129625 144080 129637
rect 209104 129625 209110 129637
rect 144074 129597 209110 129625
rect 144074 129585 144080 129597
rect 209104 129585 209110 129597
rect 209162 129585 209168 129637
rect 144016 126995 144022 127047
rect 144074 127035 144080 127047
rect 144074 127007 146846 127035
rect 144074 126995 144080 127007
rect 143920 126847 143926 126899
rect 143978 126887 143984 126899
rect 144496 126887 144502 126899
rect 143978 126859 144502 126887
rect 143978 126847 143984 126859
rect 144496 126847 144502 126859
rect 144554 126847 144560 126899
rect 146818 126813 146846 127007
rect 147088 126847 147094 126899
rect 147146 126887 147152 126899
rect 149488 126887 149494 126899
rect 147146 126859 149494 126887
rect 147146 126847 147152 126859
rect 149488 126847 149494 126859
rect 149546 126847 149552 126899
rect 203152 126813 203158 126825
rect 146818 126785 203158 126813
rect 203152 126773 203158 126785
rect 203210 126773 203216 126825
rect 146704 126699 146710 126751
rect 146762 126739 146768 126751
rect 208624 126739 208630 126751
rect 146762 126711 208630 126739
rect 146762 126699 146768 126711
rect 208624 126699 208630 126711
rect 208682 126699 208688 126751
rect 143728 126625 143734 126677
rect 143786 126665 143792 126677
rect 143920 126665 143926 126677
rect 143786 126637 143926 126665
rect 143786 126625 143792 126637
rect 143920 126625 143926 126637
rect 143978 126625 143984 126677
rect 144688 126625 144694 126677
rect 144746 126665 144752 126677
rect 146128 126665 146134 126677
rect 144746 126637 146134 126665
rect 144746 126625 144752 126637
rect 146128 126625 146134 126637
rect 146186 126625 146192 126677
rect 146416 125737 146422 125789
rect 146474 125777 146480 125789
rect 146704 125777 146710 125789
rect 146474 125749 146710 125777
rect 146474 125737 146480 125749
rect 146704 125737 146710 125749
rect 146762 125737 146768 125789
rect 144592 125367 144598 125419
rect 144650 125407 144656 125419
rect 146416 125407 146422 125419
rect 144650 125379 146422 125407
rect 144650 125367 144656 125379
rect 146416 125367 146422 125379
rect 146474 125367 146480 125419
rect 39856 125293 39862 125345
rect 39914 125333 39920 125345
rect 42448 125333 42454 125345
rect 39914 125305 42454 125333
rect 39914 125293 39920 125305
rect 42448 125293 42454 125305
rect 42506 125293 42512 125345
rect 144112 125219 144118 125271
rect 144170 125259 144176 125271
rect 144592 125259 144598 125271
rect 144170 125231 144598 125259
rect 144170 125219 144176 125231
rect 144592 125219 144598 125231
rect 144650 125219 144656 125271
rect 144400 124627 144406 124679
rect 144458 124667 144464 124679
rect 144688 124667 144694 124679
rect 144458 124639 144694 124667
rect 144458 124627 144464 124639
rect 144688 124627 144694 124639
rect 144746 124627 144752 124679
rect 144016 124479 144022 124531
rect 144074 124519 144080 124531
rect 144400 124519 144406 124531
rect 144074 124491 144406 124519
rect 144074 124479 144080 124491
rect 144400 124479 144406 124491
rect 144458 124479 144464 124531
rect 144016 123961 144022 124013
rect 144074 124001 144080 124013
rect 197392 124001 197398 124013
rect 144074 123973 197398 124001
rect 144074 123961 144080 123973
rect 197392 123961 197398 123973
rect 197450 123961 197456 124013
rect 144112 123887 144118 123939
rect 144170 123927 144176 123939
rect 200272 123927 200278 123939
rect 144170 123899 200278 123927
rect 144170 123887 144176 123899
rect 200272 123887 200278 123899
rect 200330 123887 200336 123939
rect 144112 121519 144118 121571
rect 144170 121559 144176 121571
rect 149584 121559 149590 121571
rect 144170 121531 149590 121559
rect 144170 121519 144176 121531
rect 149584 121519 149590 121531
rect 149642 121519 149648 121571
rect 645712 121223 645718 121275
rect 645770 121263 645776 121275
rect 674704 121263 674710 121275
rect 645770 121235 674710 121263
rect 645770 121223 645776 121235
rect 674704 121223 674710 121235
rect 674762 121223 674768 121275
rect 645424 121149 645430 121201
rect 645482 121189 645488 121201
rect 676912 121189 676918 121201
rect 645482 121161 676918 121189
rect 645482 121149 645488 121161
rect 676912 121149 676918 121161
rect 676970 121149 676976 121201
rect 645712 121075 645718 121127
rect 645770 121115 645776 121127
rect 676816 121115 676822 121127
rect 645770 121087 676822 121115
rect 645770 121075 645776 121087
rect 676816 121075 676822 121087
rect 676874 121075 676880 121127
rect 144016 121001 144022 121053
rect 144074 121041 144080 121053
rect 149680 121041 149686 121053
rect 144074 121013 149686 121041
rect 144074 121001 144080 121013
rect 149680 121001 149686 121013
rect 149738 121001 149744 121053
rect 209296 120927 209302 120979
rect 209354 120967 209360 120979
rect 210256 120967 210262 120979
rect 209354 120939 210262 120967
rect 209354 120927 209360 120939
rect 210256 120927 210262 120939
rect 210314 120927 210320 120979
rect 645904 120927 645910 120979
rect 645962 120967 645968 120979
rect 646096 120967 646102 120979
rect 645962 120939 646102 120967
rect 645962 120927 645968 120939
rect 646096 120927 646102 120939
rect 646154 120927 646160 120979
rect 146896 119003 146902 119055
rect 146954 119043 146960 119055
rect 151312 119043 151318 119055
rect 146954 119015 151318 119043
rect 146954 119003 146960 119015
rect 151312 119003 151318 119015
rect 151370 119003 151376 119055
rect 181456 118485 181462 118537
rect 181514 118525 181520 118537
rect 188752 118525 188758 118537
rect 181514 118497 188758 118525
rect 181514 118485 181520 118497
rect 188752 118485 188758 118497
rect 188810 118485 188816 118537
rect 167152 118337 167158 118389
rect 167210 118377 167216 118389
rect 181456 118377 181462 118389
rect 167210 118349 181462 118377
rect 167210 118337 167216 118349
rect 181456 118337 181462 118349
rect 181514 118337 181520 118389
rect 144016 118263 144022 118315
rect 144074 118303 144080 118315
rect 166960 118303 166966 118315
rect 144074 118275 166966 118303
rect 144074 118263 144080 118275
rect 166960 118263 166966 118275
rect 167018 118263 167024 118315
rect 146704 118229 146710 118241
rect 144034 118201 146710 118229
rect 144034 118167 144062 118201
rect 146704 118189 146710 118201
rect 146762 118189 146768 118241
rect 144016 118115 144022 118167
rect 144074 118115 144080 118167
rect 144112 118115 144118 118167
rect 144170 118155 144176 118167
rect 194512 118155 194518 118167
rect 144170 118127 194518 118155
rect 144170 118115 144176 118127
rect 194512 118115 194518 118127
rect 194570 118115 194576 118167
rect 143920 117967 143926 118019
rect 143978 118007 143984 118019
rect 144112 118007 144118 118019
rect 143978 117979 144118 118007
rect 143978 117967 143984 117979
rect 144112 117967 144118 117979
rect 144170 117967 144176 118019
rect 146896 116635 146902 116687
rect 146954 116675 146960 116687
rect 148048 116675 148054 116687
rect 146954 116647 148054 116675
rect 146954 116635 146960 116647
rect 148048 116635 148054 116647
rect 148106 116635 148112 116687
rect 146896 115895 146902 115947
rect 146954 115935 146960 115947
rect 148144 115935 148150 115947
rect 146954 115907 148150 115935
rect 146954 115895 146960 115907
rect 148144 115895 148150 115907
rect 148202 115895 148208 115947
rect 675184 115377 675190 115429
rect 675242 115417 675248 115429
rect 675472 115417 675478 115429
rect 675242 115389 675478 115417
rect 675242 115377 675248 115389
rect 675472 115377 675478 115389
rect 675530 115377 675536 115429
rect 674800 114785 674806 114837
rect 674858 114825 674864 114837
rect 675376 114825 675382 114837
rect 674858 114797 675382 114825
rect 674858 114785 674864 114797
rect 675376 114785 675382 114797
rect 675434 114785 675440 114837
rect 674512 114119 674518 114171
rect 674570 114159 674576 114171
rect 675376 114159 675382 114171
rect 674570 114131 675382 114159
rect 674570 114119 674576 114131
rect 675376 114119 675382 114131
rect 675434 114119 675440 114171
rect 143824 113231 143830 113283
rect 143882 113271 143888 113283
rect 144112 113271 144118 113283
rect 143882 113243 144118 113271
rect 143882 113231 143888 113243
rect 144112 113231 144118 113243
rect 144170 113231 144176 113283
rect 144016 112639 144022 112691
rect 144074 112679 144080 112691
rect 191632 112679 191638 112691
rect 144074 112651 191638 112679
rect 144074 112639 144080 112651
rect 191632 112639 191638 112651
rect 191690 112639 191696 112691
rect 144112 112417 144118 112469
rect 144170 112457 144176 112469
rect 147952 112457 147958 112469
rect 144170 112429 147958 112457
rect 144170 112417 144176 112429
rect 147952 112417 147958 112429
rect 148010 112417 148016 112469
rect 144016 112343 144022 112395
rect 144074 112383 144080 112395
rect 147856 112383 147862 112395
rect 144074 112355 147862 112383
rect 144074 112343 144080 112355
rect 147856 112343 147862 112355
rect 147914 112343 147920 112395
rect 674320 111825 674326 111877
rect 674378 111865 674384 111877
rect 675088 111865 675094 111877
rect 674378 111837 675094 111865
rect 674378 111825 674384 111837
rect 675088 111825 675094 111837
rect 675146 111825 675152 111877
rect 674608 111307 674614 111359
rect 674666 111347 674672 111359
rect 675088 111347 675094 111359
rect 674666 111319 675094 111347
rect 674666 111307 674672 111319
rect 675088 111307 675094 111319
rect 675146 111307 675152 111359
rect 674704 111159 674710 111211
rect 674762 111199 674768 111211
rect 675376 111199 675382 111211
rect 674762 111171 675382 111199
rect 674762 111159 674768 111171
rect 675376 111159 675382 111171
rect 675434 111159 675440 111211
rect 144112 109531 144118 109583
rect 144170 109571 144176 109583
rect 147760 109571 147766 109583
rect 144170 109543 147766 109571
rect 144170 109531 144176 109543
rect 147760 109531 147766 109543
rect 147818 109531 147824 109583
rect 144016 109457 144022 109509
rect 144074 109497 144080 109509
rect 185872 109497 185878 109509
rect 144074 109469 185878 109497
rect 144074 109457 144080 109469
rect 185872 109457 185878 109469
rect 185930 109457 185936 109509
rect 144112 109383 144118 109435
rect 144170 109423 144176 109435
rect 144592 109423 144598 109435
rect 144170 109395 144598 109423
rect 144170 109383 144176 109395
rect 144592 109383 144598 109395
rect 144650 109383 144656 109435
rect 674992 107533 674998 107585
rect 675050 107573 675056 107585
rect 675376 107573 675382 107585
rect 675050 107545 675382 107573
rect 675050 107533 675056 107545
rect 675376 107533 675382 107545
rect 675434 107533 675440 107585
rect 143632 107163 143638 107215
rect 143690 107203 143696 107215
rect 144112 107203 144118 107215
rect 143690 107175 144118 107203
rect 143690 107163 143696 107175
rect 144112 107163 144118 107175
rect 144170 107163 144176 107215
rect 143728 107089 143734 107141
rect 143786 107129 143792 107141
rect 144400 107129 144406 107141
rect 143786 107101 144406 107129
rect 143786 107089 143792 107101
rect 144400 107089 144406 107101
rect 144458 107089 144464 107141
rect 143824 107015 143830 107067
rect 143882 107015 143888 107067
rect 144112 107015 144118 107067
rect 144170 107055 144176 107067
rect 146128 107055 146134 107067
rect 144170 107027 146134 107055
rect 144170 107015 144176 107027
rect 146128 107015 146134 107027
rect 146186 107015 146192 107067
rect 143842 106981 143870 107015
rect 144400 106981 144406 106993
rect 143842 106953 144406 106981
rect 144400 106941 144406 106953
rect 144458 106941 144464 106993
rect 143824 106867 143830 106919
rect 143882 106907 143888 106919
rect 146416 106907 146422 106919
rect 143882 106879 146422 106907
rect 143882 106867 143888 106879
rect 146416 106867 146422 106879
rect 146474 106867 146480 106919
rect 673936 106867 673942 106919
rect 673994 106907 674000 106919
rect 675472 106907 675478 106919
rect 673994 106879 675478 106907
rect 673994 106867 674000 106879
rect 675472 106867 675478 106879
rect 675530 106867 675536 106919
rect 144592 106833 144598 106845
rect 143938 106805 144598 106833
rect 143938 106611 143966 106805
rect 144592 106793 144598 106805
rect 144650 106793 144656 106845
rect 144016 106719 144022 106771
rect 144074 106759 144080 106771
rect 162832 106759 162838 106771
rect 144074 106731 162838 106759
rect 144074 106719 144080 106731
rect 162832 106719 162838 106731
rect 162890 106719 162896 106771
rect 144016 106611 144022 106623
rect 143938 106583 144022 106611
rect 144016 106571 144022 106583
rect 144074 106571 144080 106623
rect 144688 106571 144694 106623
rect 144746 106611 144752 106623
rect 208528 106611 208534 106623
rect 144746 106583 208534 106611
rect 144746 106571 144752 106583
rect 208528 106571 208534 106583
rect 208586 106571 208592 106623
rect 143728 106497 143734 106549
rect 143786 106537 143792 106549
rect 146704 106537 146710 106549
rect 143786 106509 146710 106537
rect 143786 106497 143792 106509
rect 146704 106497 146710 106509
rect 146762 106497 146768 106549
rect 668176 106497 668182 106549
rect 668234 106537 668240 106549
rect 675088 106537 675094 106549
rect 668234 106509 675094 106537
rect 668234 106497 668240 106509
rect 675088 106497 675094 106509
rect 675146 106497 675152 106549
rect 674224 106349 674230 106401
rect 674282 106389 674288 106401
rect 675376 106389 675382 106401
rect 674282 106361 675382 106389
rect 674282 106349 674288 106361
rect 675376 106349 675382 106361
rect 675434 106349 675440 106401
rect 209296 106275 209302 106327
rect 209354 106315 209360 106327
rect 210160 106315 210166 106327
rect 209354 106287 210166 106315
rect 209354 106275 209360 106287
rect 210160 106275 210166 106287
rect 210218 106275 210224 106327
rect 144208 106127 144214 106179
rect 144266 106167 144272 106179
rect 146416 106167 146422 106179
rect 144266 106139 146422 106167
rect 144266 106127 144272 106139
rect 146416 106127 146422 106139
rect 146474 106127 146480 106179
rect 144016 105979 144022 106031
rect 144074 106019 144080 106031
rect 144208 106019 144214 106031
rect 144074 105991 144214 106019
rect 144074 105979 144080 105991
rect 144208 105979 144214 105991
rect 144266 105979 144272 106031
rect 144112 104869 144118 104921
rect 144170 104909 144176 104921
rect 144592 104909 144598 104921
rect 144170 104881 144598 104909
rect 144170 104869 144176 104881
rect 144592 104869 144598 104881
rect 144650 104869 144656 104921
rect 645424 104499 645430 104551
rect 645482 104539 645488 104551
rect 665200 104539 665206 104551
rect 645482 104511 665206 104539
rect 645482 104499 645488 104511
rect 665200 104499 665206 104511
rect 665258 104499 665264 104551
rect 144016 104351 144022 104403
rect 144074 104391 144080 104403
rect 151408 104391 151414 104403
rect 144074 104363 151414 104391
rect 144074 104351 144080 104363
rect 151408 104351 151414 104363
rect 151466 104351 151472 104403
rect 144016 104203 144022 104255
rect 144074 104243 144080 104255
rect 159952 104243 159958 104255
rect 144074 104215 159958 104243
rect 144074 104203 144080 104215
rect 159952 104203 159958 104215
rect 160010 104203 160016 104255
rect 144112 103685 144118 103737
rect 144170 103725 144176 103737
rect 208432 103725 208438 103737
rect 144170 103697 208438 103725
rect 144170 103685 144176 103697
rect 208432 103685 208438 103697
rect 208490 103685 208496 103737
rect 663184 103685 663190 103737
rect 663242 103725 663248 103737
rect 665104 103725 665110 103737
rect 663242 103697 665110 103725
rect 663242 103685 663248 103697
rect 665104 103685 665110 103697
rect 665162 103685 665168 103737
rect 146992 103611 146998 103663
rect 147050 103651 147056 103663
rect 204496 103651 204502 103663
rect 147050 103623 204502 103651
rect 147050 103611 147056 103623
rect 204496 103611 204502 103623
rect 204554 103611 204560 103663
rect 144688 103537 144694 103589
rect 144746 103577 144752 103589
rect 204592 103577 204598 103589
rect 144746 103549 204598 103577
rect 144746 103537 144752 103549
rect 204592 103537 204598 103549
rect 204650 103537 204656 103589
rect 144400 103463 144406 103515
rect 144458 103503 144464 103515
rect 204688 103503 204694 103515
rect 144458 103475 204694 103503
rect 144458 103463 144464 103475
rect 204688 103463 204694 103475
rect 204746 103463 204752 103515
rect 143632 103315 143638 103367
rect 143690 103355 143696 103367
rect 144400 103355 144406 103367
rect 143690 103327 144406 103355
rect 143690 103315 143696 103327
rect 144400 103315 144406 103327
rect 144458 103315 144464 103367
rect 144016 101539 144022 101591
rect 144074 101579 144080 101591
rect 157072 101579 157078 101591
rect 144074 101551 157078 101579
rect 144074 101539 144080 101551
rect 157072 101539 157078 101551
rect 157130 101539 157136 101591
rect 146128 101391 146134 101443
rect 146186 101431 146192 101443
rect 146320 101431 146326 101443
rect 146186 101403 146326 101431
rect 146186 101391 146192 101403
rect 146320 101391 146326 101403
rect 146378 101391 146384 101443
rect 144112 100799 144118 100851
rect 144170 100839 144176 100851
rect 147664 100839 147670 100851
rect 144170 100811 147670 100839
rect 144170 100799 144176 100811
rect 147664 100799 147670 100811
rect 147722 100799 147728 100851
rect 645808 100799 645814 100851
rect 645866 100839 645872 100851
rect 646096 100839 646102 100851
rect 645866 100811 646102 100839
rect 645866 100799 645872 100811
rect 646096 100799 646102 100811
rect 646154 100799 646160 100851
rect 144208 100725 144214 100777
rect 144266 100765 144272 100777
rect 204880 100765 204886 100777
rect 144266 100737 204886 100765
rect 144266 100725 144272 100737
rect 204880 100725 204886 100737
rect 204938 100725 204944 100777
rect 144016 100651 144022 100703
rect 144074 100691 144080 100703
rect 204784 100691 204790 100703
rect 144074 100663 204790 100691
rect 144074 100651 144080 100663
rect 204784 100651 204790 100663
rect 204842 100651 204848 100703
rect 151120 100577 151126 100629
rect 151178 100617 151184 100629
rect 204592 100617 204598 100629
rect 151178 100589 204598 100617
rect 151178 100577 151184 100589
rect 204592 100577 204598 100589
rect 204650 100577 204656 100629
rect 159760 100503 159766 100555
rect 159818 100543 159824 100555
rect 204688 100543 204694 100555
rect 159818 100515 204694 100543
rect 159818 100503 159824 100515
rect 204688 100503 204694 100515
rect 204746 100503 204752 100555
rect 162640 100429 162646 100481
rect 162698 100469 162704 100481
rect 204496 100469 204502 100481
rect 162698 100441 204502 100469
rect 162698 100429 162704 100441
rect 204496 100429 204502 100441
rect 204554 100429 204560 100481
rect 144016 98061 144022 98113
rect 144074 98101 144080 98113
rect 180112 98101 180118 98113
rect 144074 98073 180118 98101
rect 144074 98061 144080 98073
rect 180112 98061 180118 98073
rect 180170 98061 180176 98113
rect 144112 97987 144118 98039
rect 144170 98027 144176 98039
rect 183088 98027 183094 98039
rect 144170 97999 183094 98027
rect 144170 97987 144176 97999
rect 183088 97987 183094 97999
rect 183146 97987 183152 98039
rect 144208 97913 144214 97965
rect 144266 97953 144272 97965
rect 208336 97953 208342 97965
rect 144266 97925 208342 97953
rect 144266 97913 144272 97925
rect 208336 97913 208342 97925
rect 208394 97913 208400 97965
rect 154000 97839 154006 97891
rect 154058 97879 154064 97891
rect 204784 97879 204790 97891
rect 154058 97851 204790 97879
rect 154058 97839 154064 97851
rect 204784 97839 204790 97851
rect 204842 97839 204848 97891
rect 156880 97765 156886 97817
rect 156938 97805 156944 97817
rect 204496 97805 204502 97817
rect 156938 97777 204502 97805
rect 156938 97765 156944 97777
rect 204496 97765 204502 97777
rect 204554 97765 204560 97817
rect 171376 97691 171382 97743
rect 171434 97731 171440 97743
rect 204688 97731 204694 97743
rect 171434 97703 204694 97731
rect 171434 97691 171440 97703
rect 204688 97691 204694 97703
rect 204746 97691 204752 97743
rect 174256 97617 174262 97669
rect 174314 97657 174320 97669
rect 204592 97657 204598 97669
rect 174314 97629 204598 97657
rect 174314 97617 174320 97629
rect 204592 97617 204598 97629
rect 204650 97617 204656 97669
rect 182896 97543 182902 97595
rect 182954 97583 182960 97595
rect 204496 97583 204502 97595
rect 182954 97555 204502 97583
rect 182954 97543 182960 97555
rect 204496 97543 204502 97555
rect 204554 97543 204560 97595
rect 144016 95101 144022 95153
rect 144074 95141 144080 95153
rect 174448 95141 174454 95153
rect 144074 95113 174454 95141
rect 144074 95101 144080 95113
rect 174448 95101 174454 95113
rect 174506 95101 174512 95153
rect 144112 95027 144118 95079
rect 144170 95067 144176 95079
rect 177232 95067 177238 95079
rect 144170 95039 177238 95067
rect 144170 95027 144176 95039
rect 177232 95027 177238 95039
rect 177290 95027 177296 95079
rect 146704 94879 146710 94931
rect 146762 94919 146768 94931
rect 201712 94919 201718 94931
rect 146762 94891 201718 94919
rect 146762 94879 146768 94891
rect 201712 94879 201718 94891
rect 201770 94879 201776 94931
rect 151216 94805 151222 94857
rect 151274 94845 151280 94857
rect 204784 94845 204790 94857
rect 151274 94817 204790 94845
rect 151274 94805 151280 94817
rect 204784 94805 204790 94817
rect 204842 94805 204848 94857
rect 165616 94731 165622 94783
rect 165674 94771 165680 94783
rect 204496 94771 204502 94783
rect 165674 94743 204502 94771
rect 165674 94731 165680 94743
rect 204496 94731 204502 94743
rect 204554 94731 204560 94783
rect 168496 94657 168502 94709
rect 168554 94697 168560 94709
rect 204592 94697 204598 94709
rect 168554 94669 204598 94697
rect 168554 94657 168560 94669
rect 204592 94657 204598 94669
rect 204650 94657 204656 94709
rect 146416 94583 146422 94635
rect 146474 94623 146480 94635
rect 204688 94623 204694 94635
rect 146474 94595 204694 94623
rect 146474 94583 146480 94595
rect 204688 94583 204694 94595
rect 204746 94583 204752 94635
rect 203056 94435 203062 94487
rect 203114 94475 203120 94487
rect 205264 94475 205270 94487
rect 203114 94447 205270 94475
rect 203114 94435 203120 94447
rect 205264 94435 205270 94447
rect 205322 94435 205328 94487
rect 646384 92659 646390 92711
rect 646442 92699 646448 92711
rect 659824 92699 659830 92711
rect 646442 92671 659830 92699
rect 646442 92659 646448 92671
rect 659824 92659 659830 92671
rect 659882 92659 659888 92711
rect 647536 92585 647542 92637
rect 647594 92625 647600 92637
rect 661744 92625 661750 92637
rect 647594 92597 661750 92625
rect 647594 92585 647600 92597
rect 661744 92585 661750 92597
rect 661802 92585 661808 92637
rect 647152 92511 647158 92563
rect 647210 92551 647216 92563
rect 660688 92551 660694 92563
rect 647210 92523 660694 92551
rect 647210 92511 647216 92523
rect 660688 92511 660694 92523
rect 660746 92511 660752 92563
rect 647824 92437 647830 92489
rect 647882 92477 647888 92489
rect 663088 92477 663094 92489
rect 647882 92449 663094 92477
rect 647882 92437 647888 92449
rect 663088 92437 663094 92449
rect 663146 92437 663152 92489
rect 647728 92289 647734 92341
rect 647786 92329 647792 92341
rect 662512 92329 662518 92341
rect 647786 92301 662518 92329
rect 647786 92289 647792 92301
rect 662512 92289 662518 92301
rect 662570 92289 662576 92341
rect 144112 92215 144118 92267
rect 144170 92255 144176 92267
rect 154000 92255 154006 92267
rect 144170 92227 154006 92255
rect 144170 92215 144176 92227
rect 154000 92215 154006 92227
rect 154058 92215 154064 92267
rect 646096 92215 646102 92267
rect 646154 92255 646160 92267
rect 661168 92255 661174 92267
rect 646154 92227 661174 92255
rect 646154 92215 646160 92227
rect 661168 92215 661174 92227
rect 661226 92215 661232 92267
rect 144016 92141 144022 92193
rect 144074 92181 144080 92193
rect 171376 92181 171382 92193
rect 144074 92153 171382 92181
rect 144074 92141 144080 92153
rect 171376 92141 171382 92153
rect 171434 92141 171440 92193
rect 646672 92141 646678 92193
rect 646730 92181 646736 92193
rect 658864 92181 658870 92193
rect 646730 92153 658870 92181
rect 646730 92141 646736 92153
rect 658864 92141 658870 92153
rect 658922 92141 658928 92193
rect 144400 92067 144406 92119
rect 144458 92107 144464 92119
rect 204496 92107 204502 92119
rect 144458 92079 204502 92107
rect 144458 92067 144464 92079
rect 204496 92067 204502 92079
rect 204554 92067 204560 92119
rect 188656 91993 188662 92045
rect 188714 92033 188720 92045
rect 204688 92033 204694 92045
rect 188714 92005 204694 92033
rect 188714 91993 188720 92005
rect 204688 91993 204694 92005
rect 204746 91993 204752 92045
rect 194416 91919 194422 91971
rect 194474 91959 194480 91971
rect 204592 91959 204598 91971
rect 194474 91931 204598 91959
rect 194474 91919 194480 91931
rect 204592 91919 204598 91931
rect 204650 91919 204656 91971
rect 200176 91845 200182 91897
rect 200234 91885 200240 91897
rect 205360 91885 205366 91897
rect 200234 91857 205366 91885
rect 200234 91845 200240 91857
rect 205360 91845 205366 91857
rect 205418 91845 205424 91897
rect 197296 91771 197302 91823
rect 197354 91811 197360 91823
rect 204496 91811 204502 91823
rect 197354 91783 204502 91811
rect 197354 91771 197360 91783
rect 204496 91771 204502 91783
rect 204554 91771 204560 91823
rect 144016 89403 144022 89455
rect 144074 89443 144080 89455
rect 151120 89443 151126 89455
rect 144074 89415 151126 89443
rect 144074 89403 144080 89415
rect 151120 89403 151126 89415
rect 151178 89403 151184 89455
rect 144112 89329 144118 89381
rect 144170 89369 144176 89381
rect 165616 89369 165622 89381
rect 144170 89341 165622 89369
rect 144170 89329 144176 89341
rect 165616 89329 165622 89341
rect 165674 89329 165680 89381
rect 144208 89255 144214 89307
rect 144266 89295 144272 89307
rect 168496 89295 168502 89307
rect 144266 89267 168502 89295
rect 144266 89255 144272 89267
rect 168496 89255 168502 89267
rect 168554 89255 168560 89307
rect 156976 89181 156982 89233
rect 157034 89221 157040 89233
rect 204880 89221 204886 89233
rect 157034 89193 204886 89221
rect 157034 89181 157040 89193
rect 204880 89181 204886 89193
rect 204938 89181 204944 89233
rect 159856 89107 159862 89159
rect 159914 89147 159920 89159
rect 204784 89147 204790 89159
rect 159914 89119 204790 89147
rect 159914 89107 159920 89119
rect 204784 89107 204790 89119
rect 204842 89107 204848 89159
rect 162736 89033 162742 89085
rect 162794 89073 162800 89085
rect 204688 89073 204694 89085
rect 162794 89045 204694 89073
rect 162794 89033 162800 89045
rect 204688 89033 204694 89045
rect 204746 89033 204752 89085
rect 185776 88959 185782 89011
rect 185834 88999 185840 89011
rect 204592 88999 204598 89011
rect 185834 88971 204598 88999
rect 185834 88959 185840 88971
rect 204592 88959 204598 88971
rect 204650 88959 204656 89011
rect 191536 88885 191542 88937
rect 191594 88925 191600 88937
rect 204496 88925 204502 88937
rect 191594 88897 204502 88925
rect 191594 88885 191600 88897
rect 204496 88885 204502 88897
rect 204554 88885 204560 88937
rect 651376 87331 651382 87383
rect 651434 87371 651440 87383
rect 659344 87371 659350 87383
rect 651434 87343 659350 87371
rect 651434 87331 651440 87343
rect 659344 87331 659350 87343
rect 659402 87331 659408 87383
rect 658000 87297 658006 87309
rect 657058 87269 658006 87297
rect 657058 87161 657086 87269
rect 658000 87257 658006 87269
rect 658058 87257 658064 87309
rect 657040 87109 657046 87161
rect 657098 87109 657104 87161
rect 645424 87035 645430 87087
rect 645482 87075 645488 87087
rect 663280 87075 663286 87087
rect 645482 87047 663286 87075
rect 645482 87035 645488 87047
rect 663280 87035 663286 87047
rect 663338 87035 663344 87087
rect 645712 86961 645718 87013
rect 645770 87001 645776 87013
rect 650992 87001 650998 87013
rect 645770 86973 650998 87001
rect 645770 86961 645776 86973
rect 650992 86961 650998 86973
rect 651050 86961 651056 87013
rect 645712 86813 645718 86865
rect 645770 86853 645776 86865
rect 645904 86853 645910 86865
rect 645770 86825 645910 86853
rect 645770 86813 645776 86825
rect 645904 86813 645910 86825
rect 645962 86813 645968 86865
rect 210160 86739 210166 86791
rect 210218 86739 210224 86791
rect 146128 86443 146134 86495
rect 146186 86483 146192 86495
rect 146320 86483 146326 86495
rect 146186 86455 146326 86483
rect 146186 86443 146192 86455
rect 146320 86443 146326 86455
rect 146378 86443 146384 86495
rect 210178 86483 210206 86739
rect 210256 86483 210262 86495
rect 210178 86455 210262 86483
rect 210256 86443 210262 86455
rect 210314 86443 210320 86495
rect 645424 86443 645430 86495
rect 645482 86483 645488 86495
rect 651088 86483 651094 86495
rect 645482 86455 651094 86483
rect 645482 86443 645488 86455
rect 651088 86443 651094 86455
rect 651146 86443 651152 86495
rect 144400 86369 144406 86421
rect 144458 86409 144464 86421
rect 144592 86409 144598 86421
rect 144458 86381 144598 86409
rect 144458 86369 144464 86381
rect 144592 86369 144598 86381
rect 144650 86369 144656 86421
rect 154096 86369 154102 86421
rect 154154 86409 154160 86421
rect 204880 86409 204886 86421
rect 154154 86381 204886 86409
rect 154154 86369 154160 86381
rect 204880 86369 204886 86381
rect 204938 86369 204944 86421
rect 174352 86295 174358 86347
rect 174410 86335 174416 86347
rect 204784 86335 204790 86347
rect 174410 86307 204790 86335
rect 174410 86295 174416 86307
rect 204784 86295 204790 86307
rect 204842 86295 204848 86347
rect 177136 86221 177142 86273
rect 177194 86261 177200 86273
rect 204688 86261 204694 86273
rect 177194 86233 204694 86261
rect 177194 86221 177200 86233
rect 204688 86221 204694 86233
rect 204746 86221 204752 86273
rect 180016 86147 180022 86199
rect 180074 86187 180080 86199
rect 204592 86187 204598 86199
rect 180074 86159 204598 86187
rect 180074 86147 180080 86159
rect 204592 86147 204598 86159
rect 204650 86147 204656 86199
rect 182992 86073 182998 86125
rect 183050 86113 183056 86125
rect 204496 86113 204502 86125
rect 183050 86085 204502 86113
rect 183050 86073 183056 86085
rect 204496 86073 204502 86085
rect 204554 86073 204560 86125
rect 646288 85185 646294 85237
rect 646346 85225 646352 85237
rect 650896 85225 650902 85237
rect 646346 85197 650902 85225
rect 646346 85185 646352 85197
rect 650896 85185 650902 85197
rect 650954 85185 650960 85237
rect 144016 84963 144022 85015
rect 144074 85003 144080 85015
rect 204496 85003 204502 85015
rect 144074 84975 204502 85003
rect 144074 84963 144080 84975
rect 204496 84963 204502 84975
rect 204554 84963 204560 85015
rect 151504 83483 151510 83535
rect 151562 83523 151568 83535
rect 204784 83523 204790 83535
rect 151562 83495 204790 83523
rect 151562 83483 151568 83495
rect 204784 83483 204790 83495
rect 204842 83483 204848 83535
rect 165712 83409 165718 83461
rect 165770 83449 165776 83461
rect 204688 83449 204694 83461
rect 165770 83421 204694 83449
rect 165770 83409 165776 83421
rect 204688 83409 204694 83421
rect 204746 83409 204752 83461
rect 647920 83409 647926 83461
rect 647978 83449 647984 83461
rect 657040 83449 657046 83461
rect 647978 83421 657046 83449
rect 647978 83409 647984 83421
rect 657040 83409 657046 83421
rect 657098 83409 657104 83461
rect 168592 83335 168598 83387
rect 168650 83375 168656 83387
rect 204592 83375 204598 83387
rect 168650 83347 204598 83375
rect 168650 83335 168656 83347
rect 204592 83335 204598 83347
rect 204650 83335 204656 83387
rect 171472 83261 171478 83313
rect 171530 83301 171536 83313
rect 204496 83301 204502 83313
rect 171530 83273 204502 83301
rect 171530 83261 171536 83273
rect 204496 83261 204502 83273
rect 204554 83261 204560 83313
rect 144016 82077 144022 82129
rect 144074 82117 144080 82129
rect 204496 82117 204502 82129
rect 144074 82089 204502 82117
rect 144074 82077 144080 82089
rect 204496 82077 204502 82089
rect 204554 82077 204560 82129
rect 647920 81855 647926 81907
rect 647978 81895 647984 81907
rect 663280 81895 663286 81907
rect 647978 81867 663286 81895
rect 647978 81855 647984 81867
rect 663280 81855 663286 81867
rect 663338 81855 663344 81907
rect 645904 81781 645910 81833
rect 645962 81821 645968 81833
rect 663376 81821 663382 81833
rect 645962 81793 663382 81821
rect 645962 81781 645968 81793
rect 663376 81781 663382 81793
rect 663434 81781 663440 81833
rect 647632 81633 647638 81685
rect 647690 81673 647696 81685
rect 661072 81673 661078 81685
rect 647690 81645 661078 81673
rect 647690 81633 647696 81645
rect 661072 81633 661078 81645
rect 661130 81633 661136 81685
rect 647920 81263 647926 81315
rect 647978 81303 647984 81315
rect 657520 81303 657526 81315
rect 647978 81275 657526 81303
rect 647978 81263 647984 81275
rect 657520 81263 657526 81275
rect 657578 81263 657584 81315
rect 144016 80819 144022 80871
rect 144074 80859 144080 80871
rect 144400 80859 144406 80871
rect 144074 80831 144406 80859
rect 144074 80819 144080 80831
rect 144400 80819 144406 80831
rect 144458 80819 144464 80871
rect 645712 80745 645718 80797
rect 645770 80785 645776 80797
rect 645770 80757 645854 80785
rect 645770 80745 645776 80757
rect 645826 80723 645854 80757
rect 645808 80671 645814 80723
rect 645866 80671 645872 80723
rect 659440 80671 659446 80723
rect 659498 80711 659504 80723
rect 659536 80711 659542 80723
rect 659498 80683 659542 80711
rect 659498 80671 659504 80683
rect 659536 80671 659542 80683
rect 659594 80671 659600 80723
rect 188752 80597 188758 80649
rect 188810 80637 188816 80649
rect 204592 80637 204598 80649
rect 188810 80609 204598 80637
rect 188810 80597 188816 80609
rect 204592 80597 204598 80609
rect 204650 80597 204656 80649
rect 194512 80523 194518 80575
rect 194570 80563 194576 80575
rect 204496 80563 204502 80575
rect 194570 80535 204502 80563
rect 194570 80523 194576 80535
rect 204496 80523 204502 80535
rect 204554 80523 204560 80575
rect 203152 80449 203158 80501
rect 203210 80489 203216 80501
rect 206896 80489 206902 80501
rect 203210 80461 206902 80489
rect 203210 80449 203216 80461
rect 206896 80449 206902 80461
rect 206954 80449 206960 80501
rect 200272 80375 200278 80427
rect 200330 80415 200336 80427
rect 205456 80415 205462 80427
rect 200330 80387 205462 80415
rect 200330 80375 200336 80387
rect 205456 80375 205462 80387
rect 205514 80375 205520 80427
rect 197392 80301 197398 80353
rect 197450 80341 197456 80353
rect 204688 80341 204694 80353
rect 197450 80313 204694 80341
rect 197450 80301 197456 80313
rect 204688 80301 204694 80313
rect 204746 80301 204752 80353
rect 647920 80153 647926 80205
rect 647978 80193 647984 80205
rect 656944 80193 656950 80205
rect 647978 80165 656950 80193
rect 647978 80153 647984 80165
rect 656944 80153 656950 80165
rect 657002 80153 657008 80205
rect 646096 79117 646102 79169
rect 646154 79157 646160 79169
rect 658864 79157 658870 79169
rect 646154 79129 658870 79157
rect 646154 79117 646160 79129
rect 658864 79117 658870 79129
rect 658922 79117 658928 79169
rect 647824 78673 647830 78725
rect 647882 78713 647888 78725
rect 660688 78713 660694 78725
rect 647882 78685 660694 78713
rect 647882 78673 647888 78685
rect 660688 78673 660694 78685
rect 660746 78673 660752 78725
rect 646864 78599 646870 78651
rect 646922 78639 646928 78651
rect 651184 78639 651190 78651
rect 646922 78611 651190 78639
rect 646922 78599 646928 78611
rect 651184 78599 651190 78611
rect 651242 78599 651248 78651
rect 647920 78303 647926 78355
rect 647978 78343 647984 78355
rect 662512 78343 662518 78355
rect 647978 78315 662518 78343
rect 647978 78303 647984 78315
rect 662512 78303 662518 78315
rect 662570 78303 662576 78355
rect 144112 77859 144118 77911
rect 144170 77899 144176 77911
rect 187216 77899 187222 77911
rect 144170 77871 187222 77899
rect 144170 77859 144176 77871
rect 187216 77859 187222 77871
rect 187274 77859 187280 77911
rect 144016 77785 144022 77837
rect 144074 77825 144080 77837
rect 208240 77825 208246 77837
rect 144074 77797 208246 77825
rect 144074 77785 144080 77797
rect 208240 77785 208246 77797
rect 208298 77785 208304 77837
rect 157072 77711 157078 77763
rect 157130 77751 157136 77763
rect 204976 77751 204982 77763
rect 157130 77723 204982 77751
rect 157130 77711 157136 77723
rect 204976 77711 204982 77723
rect 205034 77711 205040 77763
rect 647344 77711 647350 77763
rect 647402 77751 647408 77763
rect 659440 77751 659446 77763
rect 647402 77723 659446 77751
rect 647402 77711 647408 77723
rect 659440 77711 659446 77723
rect 659498 77711 659504 77763
rect 159952 77637 159958 77689
rect 160010 77677 160016 77689
rect 204880 77677 204886 77689
rect 160010 77649 204886 77677
rect 160010 77637 160016 77649
rect 204880 77637 204886 77649
rect 204938 77637 204944 77689
rect 647920 77637 647926 77689
rect 647978 77677 647984 77689
rect 650992 77677 650998 77689
rect 647978 77649 650998 77677
rect 647978 77637 647984 77649
rect 650992 77637 650998 77649
rect 651050 77637 651056 77689
rect 162832 77563 162838 77615
rect 162890 77603 162896 77615
rect 204784 77603 204790 77615
rect 162890 77575 204790 77603
rect 162890 77563 162896 77575
rect 204784 77563 204790 77575
rect 204842 77563 204848 77615
rect 185872 77489 185878 77541
rect 185930 77529 185936 77541
rect 204688 77529 204694 77541
rect 185930 77501 204694 77529
rect 185930 77489 185936 77501
rect 204688 77489 204694 77501
rect 204746 77489 204752 77541
rect 187216 77415 187222 77467
rect 187274 77455 187280 77467
rect 204496 77455 204502 77467
rect 187274 77427 204502 77455
rect 187274 77415 187280 77427
rect 204496 77415 204502 77427
rect 204554 77415 204560 77467
rect 191632 77341 191638 77393
rect 191690 77381 191696 77393
rect 204592 77381 204598 77393
rect 191690 77353 204598 77381
rect 191690 77341 191696 77353
rect 204592 77341 204598 77353
rect 204650 77341 204656 77393
rect 647920 77267 647926 77319
rect 647978 77307 647984 77319
rect 662896 77307 662902 77319
rect 647978 77279 662902 77307
rect 647978 77267 647984 77279
rect 662896 77267 662902 77279
rect 662954 77267 662960 77319
rect 646480 76897 646486 76949
rect 646538 76937 646544 76949
rect 658288 76937 658294 76949
rect 646538 76909 658294 76937
rect 646538 76897 646544 76909
rect 658288 76897 658294 76909
rect 658346 76897 658352 76949
rect 646480 76749 646486 76801
rect 646538 76789 646544 76801
rect 650896 76789 650902 76801
rect 646538 76761 650902 76789
rect 646538 76749 646544 76761
rect 650896 76749 650902 76761
rect 650954 76749 650960 76801
rect 144208 76379 144214 76431
rect 144266 76419 144272 76431
rect 145456 76419 145462 76431
rect 144266 76391 145462 76419
rect 144266 76379 144272 76391
rect 145456 76379 145462 76391
rect 145514 76379 145520 76431
rect 146032 76305 146038 76357
rect 146090 76345 146096 76357
rect 146800 76345 146806 76357
rect 146090 76317 146806 76345
rect 146090 76305 146096 76317
rect 146800 76305 146806 76317
rect 146858 76305 146864 76357
rect 145552 76157 145558 76209
rect 145610 76197 145616 76209
rect 146512 76197 146518 76209
rect 145610 76169 146518 76197
rect 145610 76157 145616 76169
rect 146512 76157 146518 76169
rect 146570 76157 146576 76209
rect 646864 75565 646870 75617
rect 646922 75605 646928 75617
rect 656848 75605 656854 75617
rect 646922 75577 656854 75605
rect 646922 75565 646928 75577
rect 656848 75565 656854 75577
rect 656906 75565 656912 75617
rect 647920 75269 647926 75321
rect 647978 75309 647984 75321
rect 661744 75309 661750 75321
rect 647978 75281 661750 75309
rect 647978 75269 647984 75281
rect 661744 75269 661750 75281
rect 661802 75269 661808 75321
rect 144016 75047 144022 75099
rect 144074 75087 144080 75099
rect 160528 75087 160534 75099
rect 144074 75059 160534 75087
rect 144074 75047 144080 75059
rect 160528 75047 160534 75059
rect 160586 75047 160592 75099
rect 146896 74973 146902 75025
rect 146954 75013 146960 75025
rect 156880 75013 156886 75025
rect 146954 74985 156886 75013
rect 146954 74973 146960 74985
rect 156880 74973 156886 74985
rect 156938 74973 156944 75025
rect 144112 74899 144118 74951
rect 144170 74939 144176 74951
rect 161584 74939 161590 74951
rect 144170 74911 161590 74939
rect 144170 74899 144176 74911
rect 161584 74899 161590 74911
rect 161642 74899 161648 74951
rect 154000 74825 154006 74877
rect 154058 74865 154064 74877
rect 204880 74865 204886 74877
rect 154058 74837 204886 74865
rect 154058 74825 154064 74837
rect 204880 74825 204886 74837
rect 204938 74825 204944 74877
rect 174448 74751 174454 74803
rect 174506 74791 174512 74803
rect 204784 74791 204790 74803
rect 174506 74763 204790 74791
rect 174506 74751 174512 74763
rect 204784 74751 204790 74763
rect 204842 74751 204848 74803
rect 177232 74677 177238 74729
rect 177290 74717 177296 74729
rect 204688 74717 204694 74729
rect 177290 74689 204694 74717
rect 177290 74677 177296 74689
rect 204688 74677 204694 74689
rect 204746 74677 204752 74729
rect 180112 74603 180118 74655
rect 180170 74643 180176 74655
rect 204592 74643 204598 74655
rect 180170 74615 204598 74643
rect 180170 74603 180176 74615
rect 204592 74603 204598 74615
rect 204650 74603 204656 74655
rect 183088 74529 183094 74581
rect 183146 74569 183152 74581
rect 204496 74569 204502 74581
rect 183146 74541 204502 74569
rect 183146 74529 183152 74541
rect 204496 74529 204502 74541
rect 204554 74529 204560 74581
rect 144112 74233 144118 74285
rect 144170 74273 144176 74285
rect 148336 74273 148342 74285
rect 144170 74245 148342 74273
rect 144170 74233 144176 74245
rect 148336 74233 148342 74245
rect 148394 74233 148400 74285
rect 640720 73419 640726 73471
rect 640778 73459 640784 73471
rect 663184 73459 663190 73471
rect 640778 73431 663190 73459
rect 640778 73419 640784 73431
rect 663184 73419 663190 73431
rect 663242 73419 663248 73471
rect 647920 72679 647926 72731
rect 647978 72719 647984 72731
rect 663280 72719 663286 72731
rect 647978 72691 663286 72719
rect 647978 72679 647984 72691
rect 663280 72679 663286 72691
rect 663338 72679 663344 72731
rect 143824 72605 143830 72657
rect 143882 72645 143888 72657
rect 144112 72645 144118 72657
rect 143882 72617 144118 72645
rect 143882 72605 143888 72617
rect 144112 72605 144118 72617
rect 144170 72605 144176 72657
rect 646960 72605 646966 72657
rect 647018 72645 647024 72657
rect 663472 72645 663478 72657
rect 647018 72617 663478 72645
rect 647018 72605 647024 72617
rect 663472 72605 663478 72617
rect 663530 72605 663536 72657
rect 144592 72457 144598 72509
rect 144650 72497 144656 72509
rect 146512 72497 146518 72509
rect 144650 72469 146518 72497
rect 144650 72457 144656 72469
rect 146512 72457 146518 72469
rect 146570 72457 146576 72509
rect 647824 72235 647830 72287
rect 647882 72275 647888 72287
rect 660112 72275 660118 72287
rect 647882 72247 660118 72275
rect 647882 72235 647888 72247
rect 660112 72235 660118 72247
rect 660170 72235 660176 72287
rect 144016 72013 144022 72065
rect 144074 72053 144080 72065
rect 154576 72053 154582 72065
rect 144074 72025 154582 72053
rect 144074 72013 144080 72025
rect 154576 72013 154582 72025
rect 154634 72013 154640 72065
rect 151120 71939 151126 71991
rect 151178 71979 151184 71991
rect 204784 71979 204790 71991
rect 151178 71951 204790 71979
rect 151178 71939 151184 71951
rect 204784 71939 204790 71951
rect 204842 71939 204848 71991
rect 161584 71865 161590 71917
rect 161642 71905 161648 71917
rect 204880 71905 204886 71917
rect 161642 71877 204886 71905
rect 161642 71865 161648 71877
rect 204880 71865 204886 71877
rect 204938 71865 204944 71917
rect 165616 71791 165622 71843
rect 165674 71831 165680 71843
rect 204688 71831 204694 71843
rect 165674 71803 204694 71831
rect 165674 71791 165680 71803
rect 204688 71791 204694 71803
rect 204746 71791 204752 71843
rect 168496 71717 168502 71769
rect 168554 71757 168560 71769
rect 204592 71757 204598 71769
rect 168554 71729 204598 71757
rect 168554 71717 168560 71729
rect 204592 71717 204598 71729
rect 204650 71717 204656 71769
rect 171376 71643 171382 71695
rect 171434 71683 171440 71695
rect 204496 71683 204502 71695
rect 171434 71655 204502 71683
rect 171434 71643 171440 71655
rect 204496 71643 204502 71655
rect 204554 71643 204560 71695
rect 144016 70829 144022 70881
rect 144074 70869 144080 70881
rect 149776 70869 149782 70881
rect 144074 70841 149782 70869
rect 144074 70829 144080 70841
rect 149776 70829 149782 70841
rect 149834 70829 149840 70881
rect 144016 69127 144022 69179
rect 144074 69167 144080 69179
rect 144074 69139 148094 69167
rect 144074 69127 144080 69139
rect 148066 69093 148094 69139
rect 204880 69093 204886 69105
rect 148066 69065 204886 69093
rect 204880 69053 204886 69065
rect 204938 69053 204944 69105
rect 149776 68979 149782 69031
rect 149834 69019 149840 69031
rect 204784 69019 204790 69031
rect 149834 68991 204790 69019
rect 149834 68979 149840 68991
rect 204784 68979 204790 68991
rect 204842 68979 204848 69031
rect 154576 68905 154582 68957
rect 154634 68945 154640 68957
rect 204688 68945 204694 68957
rect 154634 68917 204694 68945
rect 154634 68905 154640 68917
rect 204688 68905 204694 68917
rect 204746 68905 204752 68957
rect 156880 68831 156886 68883
rect 156938 68871 156944 68883
rect 204592 68871 204598 68883
rect 156938 68843 204598 68871
rect 156938 68831 156944 68843
rect 204592 68831 204598 68843
rect 204650 68831 204656 68883
rect 160528 68757 160534 68809
rect 160586 68797 160592 68809
rect 204496 68797 204502 68809
rect 160586 68769 204502 68797
rect 160586 68757 160592 68769
rect 204496 68757 204502 68769
rect 204554 68757 204560 68809
rect 144016 67351 144022 67403
rect 144074 67391 144080 67403
rect 152656 67391 152662 67403
rect 144074 67363 152662 67391
rect 144074 67351 144080 67363
rect 152656 67351 152662 67363
rect 152714 67351 152720 67403
rect 144592 67203 144598 67255
rect 144650 67243 144656 67255
rect 144650 67215 144734 67243
rect 144650 67203 144656 67215
rect 144706 67033 144734 67215
rect 144688 66981 144694 67033
rect 144746 66981 144752 67033
rect 146128 66833 146134 66885
rect 146186 66873 146192 66885
rect 146704 66873 146710 66885
rect 146186 66845 146710 66873
rect 146186 66833 146192 66845
rect 146704 66833 146710 66845
rect 146762 66833 146768 66885
rect 144016 66685 144022 66737
rect 144074 66725 144080 66737
rect 146704 66725 146710 66737
rect 144074 66697 146710 66725
rect 144074 66685 144080 66697
rect 146704 66685 146710 66697
rect 146762 66685 146768 66737
rect 144208 66503 144214 66515
rect 144034 66475 144214 66503
rect 144034 66293 144062 66475
rect 144208 66463 144214 66475
rect 144266 66463 144272 66515
rect 146512 66315 146518 66367
rect 146570 66355 146576 66367
rect 157648 66355 157654 66367
rect 146570 66327 157654 66355
rect 146570 66315 146576 66327
rect 157648 66315 157654 66327
rect 157706 66315 157712 66367
rect 144016 66241 144022 66293
rect 144074 66241 144080 66293
rect 144208 66241 144214 66293
rect 144266 66281 144272 66293
rect 144266 66253 149822 66281
rect 144266 66241 144272 66253
rect 146320 66167 146326 66219
rect 146378 66207 146384 66219
rect 146800 66207 146806 66219
rect 146378 66179 146806 66207
rect 146378 66167 146384 66179
rect 146800 66167 146806 66179
rect 146858 66167 146864 66219
rect 149794 66207 149822 66253
rect 204688 66207 204694 66219
rect 149794 66179 204694 66207
rect 204688 66167 204694 66179
rect 204746 66167 204752 66219
rect 210256 66167 210262 66219
rect 210314 66167 210320 66219
rect 152656 66093 152662 66145
rect 152714 66133 152720 66145
rect 204496 66133 204502 66145
rect 152714 66105 204502 66133
rect 152714 66093 152720 66105
rect 204496 66093 204502 66105
rect 204554 66093 204560 66145
rect 157648 66019 157654 66071
rect 157706 66059 157712 66071
rect 204592 66059 204598 66071
rect 157706 66031 204598 66059
rect 157706 66019 157712 66031
rect 204592 66019 204598 66031
rect 204650 66019 204656 66071
rect 210274 65997 210302 66167
rect 210256 65945 210262 65997
rect 210314 65945 210320 65997
rect 144016 65575 144022 65627
rect 144074 65615 144080 65627
rect 144208 65615 144214 65627
rect 144074 65587 144214 65615
rect 144074 65575 144080 65587
rect 144208 65575 144214 65587
rect 144266 65575 144272 65627
rect 145456 65131 145462 65183
rect 145514 65171 145520 65183
rect 146512 65171 146518 65183
rect 145514 65143 146518 65171
rect 145514 65131 145520 65143
rect 146512 65131 146518 65143
rect 146570 65131 146576 65183
rect 144976 64983 144982 65035
rect 145034 65023 145040 65035
rect 145456 65023 145462 65035
rect 145034 64995 145462 65023
rect 145034 64983 145040 64995
rect 145456 64983 145462 64995
rect 145514 64983 145520 65035
rect 144016 64835 144022 64887
rect 144074 64875 144080 64887
rect 204496 64875 204502 64887
rect 144074 64847 204502 64875
rect 144074 64835 144080 64847
rect 204496 64835 204502 64847
rect 204554 64835 204560 64887
rect 144880 64761 144886 64813
rect 144938 64801 144944 64813
rect 204592 64801 204598 64813
rect 144938 64773 204598 64801
rect 144938 64761 144944 64773
rect 204592 64761 204598 64773
rect 204650 64761 204656 64813
rect 146896 63355 146902 63407
rect 146954 63395 146960 63407
rect 204496 63395 204502 63407
rect 146954 63367 204502 63395
rect 146954 63355 146960 63367
rect 204496 63355 204502 63367
rect 204554 63355 204560 63407
rect 144016 62171 144022 62223
rect 144074 62211 144080 62223
rect 149776 62211 149782 62223
rect 144074 62183 149782 62211
rect 144074 62171 144080 62183
rect 149776 62171 149782 62183
rect 149834 62171 149840 62223
rect 160528 60765 160534 60817
rect 160586 60805 160592 60817
rect 204592 60805 204598 60817
rect 160586 60777 204598 60805
rect 160586 60765 160592 60777
rect 204592 60765 204598 60777
rect 204650 60765 204656 60817
rect 156304 60691 156310 60743
rect 156362 60731 156368 60743
rect 204688 60731 204694 60743
rect 156362 60703 204694 60731
rect 156362 60691 156368 60703
rect 204688 60691 204694 60703
rect 204746 60691 204752 60743
rect 152656 60617 152662 60669
rect 152714 60657 152720 60669
rect 204496 60657 204502 60669
rect 152714 60629 204502 60657
rect 152714 60617 152720 60629
rect 204496 60617 204502 60629
rect 204554 60617 204560 60669
rect 151120 60543 151126 60595
rect 151178 60583 151184 60595
rect 204880 60583 204886 60595
rect 151178 60555 204886 60583
rect 151178 60543 151184 60555
rect 204880 60543 204886 60555
rect 204938 60543 204944 60595
rect 148336 60469 148342 60521
rect 148394 60509 148400 60521
rect 204784 60509 204790 60521
rect 148394 60481 204790 60509
rect 148394 60469 148400 60481
rect 204784 60469 204790 60481
rect 204842 60469 204848 60521
rect 146896 60395 146902 60447
rect 146954 60435 146960 60447
rect 204496 60435 204502 60447
rect 146954 60407 204502 60435
rect 146954 60395 146960 60407
rect 204496 60395 204502 60407
rect 204554 60395 204560 60447
rect 149776 60321 149782 60373
rect 149834 60361 149840 60373
rect 204688 60361 204694 60373
rect 149834 60333 204694 60361
rect 149834 60321 149840 60333
rect 204688 60321 204694 60333
rect 204746 60321 204752 60373
rect 207760 59951 207766 60003
rect 207818 59991 207824 60003
rect 208720 59991 208726 60003
rect 207818 59963 208726 59991
rect 207818 59951 207824 59963
rect 208720 59951 208726 59963
rect 208778 59951 208784 60003
rect 144016 59581 144022 59633
rect 144074 59621 144080 59633
rect 160528 59621 160534 59633
rect 144074 59593 160534 59621
rect 144074 59581 144080 59593
rect 160528 59581 160534 59593
rect 160586 59581 160592 59633
rect 144016 58989 144022 59041
rect 144074 59029 144080 59041
rect 204592 59029 204598 59041
rect 144074 59001 204598 59029
rect 144074 58989 144080 59001
rect 204592 58989 204598 59001
rect 204650 58989 204656 59041
rect 144016 57065 144022 57117
rect 144074 57105 144080 57117
rect 156304 57105 156310 57117
rect 144074 57077 156310 57105
rect 144074 57065 144080 57077
rect 156304 57065 156310 57077
rect 156362 57065 156368 57117
rect 144016 56473 144022 56525
rect 144074 56513 144080 56525
rect 152656 56513 152662 56525
rect 144074 56485 152662 56513
rect 144074 56473 144080 56485
rect 152656 56473 152662 56485
rect 152714 56473 152720 56525
rect 210160 55215 210166 55267
rect 210218 55215 210224 55267
rect 144016 54623 144022 54675
rect 144074 54663 144080 54675
rect 151120 54663 151126 54675
rect 144074 54635 151126 54663
rect 144074 54623 144080 54635
rect 151120 54623 151126 54635
rect 151178 54623 151184 54675
rect 210178 54441 210206 55215
rect 210178 54413 228542 54441
rect 228514 54305 228542 54413
rect 209488 54253 209494 54305
rect 209546 54293 209552 54305
rect 217168 54293 217174 54305
rect 209546 54265 217174 54293
rect 209546 54253 209552 54265
rect 217168 54253 217174 54265
rect 217226 54253 217232 54305
rect 228496 54253 228502 54305
rect 228554 54253 228560 54305
rect 209968 54179 209974 54231
rect 210026 54219 210032 54231
rect 219184 54219 219190 54231
rect 210026 54191 219190 54219
rect 210026 54179 210032 54191
rect 219184 54179 219190 54191
rect 219242 54179 219248 54231
rect 144016 54105 144022 54157
rect 144074 54145 144080 54157
rect 148336 54145 148342 54157
rect 144074 54117 148342 54145
rect 144074 54105 144080 54117
rect 148336 54105 148342 54117
rect 148394 54105 148400 54157
rect 209296 54105 209302 54157
rect 209354 54145 209360 54157
rect 256048 54145 256054 54157
rect 209354 54117 256054 54145
rect 209354 54105 209360 54117
rect 256048 54105 256054 54117
rect 256106 54105 256112 54157
rect 206992 54031 206998 54083
rect 207050 54071 207056 54083
rect 221392 54071 221398 54083
rect 207050 54043 221398 54071
rect 207050 54031 207056 54043
rect 221392 54031 221398 54043
rect 221450 54031 221456 54083
rect 210832 53957 210838 54009
rect 210890 53997 210896 54009
rect 216976 53997 216982 54009
rect 210890 53969 216982 53997
rect 210890 53957 210896 53969
rect 216976 53957 216982 53969
rect 217034 53957 217040 54009
rect 282160 53923 282166 53935
rect 262114 53895 282166 53923
rect 210256 53809 210262 53861
rect 210314 53849 210320 53861
rect 210314 53821 262046 53849
rect 210314 53809 210320 53821
rect 208048 53735 208054 53787
rect 208106 53775 208112 53787
rect 218176 53775 218182 53787
rect 208106 53747 218182 53775
rect 208106 53735 208112 53747
rect 218176 53735 218182 53747
rect 218234 53735 218240 53787
rect 262018 53775 262046 53821
rect 262114 53775 262142 53895
rect 282160 53883 282166 53895
rect 282218 53883 282224 53935
rect 262018 53747 262142 53775
rect 208336 53661 208342 53713
rect 208394 53701 208400 53713
rect 208394 53673 215822 53701
rect 208394 53661 208400 53673
rect 205648 53587 205654 53639
rect 205706 53627 205712 53639
rect 205706 53599 215630 53627
rect 205706 53587 205712 53599
rect 215602 53565 215630 53599
rect 215794 53565 215822 53673
rect 216976 53661 216982 53713
rect 217034 53701 217040 53713
rect 217034 53673 256286 53701
rect 217034 53661 217040 53673
rect 256258 53627 256286 53673
rect 262114 53673 282206 53701
rect 262114 53627 262142 53673
rect 256258 53599 262142 53627
rect 282178 53627 282206 53673
rect 357424 53627 357430 53639
rect 282178 53599 357430 53627
rect 357424 53587 357430 53599
rect 357482 53587 357488 53639
rect 383152 53587 383158 53639
rect 383210 53627 383216 53639
rect 403120 53627 403126 53639
rect 383210 53599 403126 53627
rect 383210 53587 383216 53599
rect 403120 53587 403126 53599
rect 403178 53587 403184 53639
rect 490960 53627 490966 53639
rect 480994 53599 490966 53627
rect 210352 53513 210358 53565
rect 210410 53553 210416 53565
rect 215248 53553 215254 53565
rect 210410 53525 215254 53553
rect 210410 53513 210416 53525
rect 215248 53513 215254 53525
rect 215306 53513 215312 53565
rect 215584 53513 215590 53565
rect 215642 53513 215648 53565
rect 215776 53513 215782 53565
rect 215834 53513 215840 53565
rect 217168 53513 217174 53565
rect 217226 53553 217232 53565
rect 217456 53553 217462 53565
rect 217226 53525 217462 53553
rect 217226 53513 217232 53525
rect 217456 53513 217462 53525
rect 217514 53513 217520 53565
rect 228496 53513 228502 53565
rect 228554 53553 228560 53565
rect 398320 53553 398326 53565
rect 228554 53525 398326 53553
rect 228554 53513 228560 53525
rect 398320 53513 398326 53525
rect 398378 53513 398384 53565
rect 423568 53513 423574 53565
rect 423626 53553 423632 53565
rect 443344 53553 443350 53565
rect 423626 53525 443350 53553
rect 423626 53513 423632 53525
rect 443344 53513 443350 53525
rect 443402 53513 443408 53565
rect 460816 53513 460822 53565
rect 460874 53553 460880 53565
rect 480994 53553 481022 53599
rect 490960 53587 490966 53599
rect 491018 53587 491024 53639
rect 460874 53525 481022 53553
rect 460874 53513 460880 53525
rect 209200 53439 209206 53491
rect 209258 53479 209264 53491
rect 216352 53479 216358 53491
rect 209258 53451 216358 53479
rect 209258 53439 209264 53451
rect 216352 53439 216358 53451
rect 216410 53439 216416 53491
rect 219664 53479 219670 53491
rect 217282 53451 219670 53479
rect 209392 53365 209398 53417
rect 209450 53405 209456 53417
rect 217282 53405 217310 53451
rect 219664 53439 219670 53451
rect 219722 53439 219728 53491
rect 256240 53439 256246 53491
rect 256298 53479 256304 53491
rect 443440 53479 443446 53491
rect 256298 53451 443446 53479
rect 256298 53439 256304 53451
rect 443440 53439 443446 53451
rect 443498 53439 443504 53491
rect 255952 53405 255958 53417
rect 209450 53377 217310 53405
rect 217378 53377 255958 53405
rect 209450 53365 209456 53377
rect 209776 53291 209782 53343
rect 209834 53331 209840 53343
rect 213424 53331 213430 53343
rect 209834 53303 213430 53331
rect 209834 53291 209840 53303
rect 213424 53291 213430 53303
rect 213482 53291 213488 53343
rect 209680 53217 209686 53269
rect 209738 53257 209744 53269
rect 213712 53257 213718 53269
rect 209738 53229 213718 53257
rect 209738 53217 209744 53229
rect 213712 53217 213718 53229
rect 213770 53217 213776 53269
rect 207280 53143 207286 53195
rect 207338 53183 207344 53195
rect 217378 53183 217406 53377
rect 255952 53365 255958 53377
rect 256010 53365 256016 53417
rect 256144 53365 256150 53417
rect 256202 53405 256208 53417
rect 443344 53405 443350 53417
rect 256202 53377 443350 53405
rect 256202 53365 256208 53377
rect 443344 53365 443350 53377
rect 443402 53365 443408 53417
rect 460816 53365 460822 53417
rect 460874 53365 460880 53417
rect 293680 53291 293686 53343
rect 293738 53331 293744 53343
rect 293738 53303 383102 53331
rect 293738 53291 293744 53303
rect 383074 53269 383102 53303
rect 403408 53291 403414 53343
rect 403466 53331 403472 53343
rect 423376 53331 423382 53343
rect 403466 53303 423382 53331
rect 403466 53291 403472 53303
rect 423376 53291 423382 53303
rect 423434 53291 423440 53343
rect 443632 53291 443638 53343
rect 443690 53331 443696 53343
rect 460834 53331 460862 53365
rect 443690 53303 460862 53331
rect 443690 53291 443696 53303
rect 490960 53291 490966 53343
rect 491018 53331 491024 53343
rect 512272 53331 512278 53343
rect 491018 53303 512278 53331
rect 491018 53291 491024 53303
rect 512272 53291 512278 53303
rect 512330 53291 512336 53343
rect 273616 53257 273622 53269
rect 239074 53229 273622 53257
rect 239074 53183 239102 53229
rect 273616 53217 273622 53229
rect 273674 53217 273680 53269
rect 321040 53257 321046 53269
rect 308290 53229 321046 53257
rect 207338 53155 217406 53183
rect 218914 53155 239102 53183
rect 207338 53143 207344 53155
rect 210736 53069 210742 53121
rect 210794 53109 210800 53121
rect 218914 53109 218942 53155
rect 276400 53109 276406 53121
rect 210794 53081 218942 53109
rect 227218 53081 276406 53109
rect 210794 53069 210800 53081
rect 207088 52995 207094 53047
rect 207146 53035 207152 53047
rect 220336 53035 220342 53047
rect 207146 53007 220342 53035
rect 207146 52995 207152 53007
rect 220336 52995 220342 53007
rect 220394 52995 220400 53047
rect 221392 52995 221398 53047
rect 221450 53035 221456 53047
rect 227218 53035 227246 53081
rect 276400 53069 276406 53081
rect 276458 53069 276464 53121
rect 276592 53069 276598 53121
rect 276650 53109 276656 53121
rect 308290 53109 308318 53229
rect 321040 53217 321046 53229
rect 321098 53217 321104 53269
rect 383056 53217 383062 53269
rect 383114 53217 383120 53269
rect 443728 53217 443734 53269
rect 443786 53257 443792 53269
rect 525904 53257 525910 53269
rect 443786 53229 470846 53257
rect 443786 53217 443792 53229
rect 331120 53143 331126 53195
rect 331178 53183 331184 53195
rect 362704 53183 362710 53195
rect 331178 53155 362710 53183
rect 331178 53143 331184 53155
rect 362704 53143 362710 53155
rect 362762 53143 362768 53195
rect 362992 53143 362998 53195
rect 363050 53183 363056 53195
rect 403120 53183 403126 53195
rect 363050 53155 403126 53183
rect 363050 53143 363056 53155
rect 403120 53143 403126 53155
rect 403178 53143 403184 53195
rect 403312 53143 403318 53195
rect 403370 53183 403376 53195
rect 440656 53183 440662 53195
rect 403370 53155 440662 53183
rect 403370 53143 403376 53155
rect 440656 53143 440662 53155
rect 440714 53143 440720 53195
rect 276650 53081 308318 53109
rect 470818 53109 470846 53229
rect 509890 53229 525910 53257
rect 509890 53109 509918 53229
rect 525904 53217 525910 53229
rect 525962 53217 525968 53269
rect 470818 53081 509918 53109
rect 276650 53069 276656 53081
rect 221450 53007 227246 53035
rect 221450 52995 221456 53007
rect 321040 52995 321046 53047
rect 321098 53035 321104 53047
rect 331120 53035 331126 53047
rect 321098 53007 331126 53035
rect 321098 52995 321104 53007
rect 331120 52995 331126 53007
rect 331178 52995 331184 53047
rect 208144 52921 208150 52973
rect 208202 52961 208208 52973
rect 220048 52961 220054 52973
rect 208202 52933 220054 52961
rect 208202 52921 208208 52933
rect 220048 52921 220054 52933
rect 220106 52921 220112 52973
rect 210160 52847 210166 52899
rect 210218 52887 210224 52899
rect 218896 52887 218902 52899
rect 210218 52859 218902 52887
rect 210218 52847 210224 52859
rect 218896 52847 218902 52859
rect 218954 52847 218960 52899
rect 151408 52699 151414 52751
rect 151466 52739 151472 52751
rect 217264 52739 217270 52751
rect 151466 52711 217270 52739
rect 151466 52699 151472 52711
rect 217264 52699 217270 52711
rect 217322 52699 217328 52751
rect 443344 52551 443350 52603
rect 443402 52591 443408 52603
rect 460720 52591 460726 52603
rect 443402 52563 460726 52591
rect 443402 52551 443408 52563
rect 460720 52551 460726 52563
rect 460778 52551 460784 52603
rect 211888 52477 211894 52529
rect 211946 52517 211952 52529
rect 220912 52517 220918 52529
rect 211946 52489 220918 52517
rect 211946 52477 211952 52489
rect 220912 52477 220918 52489
rect 220970 52477 220976 52529
rect 212176 52329 212182 52381
rect 212234 52369 212240 52381
rect 226960 52369 226966 52381
rect 212234 52341 226966 52369
rect 212234 52329 212240 52341
rect 226960 52329 226966 52341
rect 227018 52329 227024 52381
rect 137488 52255 137494 52307
rect 137546 52295 137552 52307
rect 239056 52295 239062 52307
rect 137546 52267 239062 52295
rect 137546 52255 137552 52267
rect 239056 52255 239062 52267
rect 239114 52255 239120 52307
rect 151312 52181 151318 52233
rect 151370 52221 151376 52233
rect 219856 52221 219862 52233
rect 151370 52193 219862 52221
rect 151370 52181 151376 52193
rect 219856 52181 219862 52193
rect 219914 52181 219920 52233
rect 146704 52107 146710 52159
rect 146762 52147 146768 52159
rect 212176 52147 212182 52159
rect 146762 52119 212182 52147
rect 146762 52107 146768 52119
rect 212176 52107 212182 52119
rect 212234 52107 212240 52159
rect 225712 52147 225718 52159
rect 212290 52119 225718 52147
rect 144400 52033 144406 52085
rect 144458 52073 144464 52085
rect 211888 52073 211894 52085
rect 144458 52045 211894 52073
rect 144458 52033 144464 52045
rect 211888 52033 211894 52045
rect 211946 52033 211952 52085
rect 144592 51959 144598 52011
rect 144650 51999 144656 52011
rect 212290 51999 212318 52119
rect 225712 52107 225718 52119
rect 225770 52107 225776 52159
rect 212368 52033 212374 52085
rect 212426 52073 212432 52085
rect 213424 52073 213430 52085
rect 212426 52045 213430 52073
rect 212426 52033 212432 52045
rect 213424 52033 213430 52045
rect 213482 52033 213488 52085
rect 144650 51971 212318 51999
rect 213346 51971 213566 51999
rect 144650 51959 144656 51971
rect 146416 51885 146422 51937
rect 146474 51925 146480 51937
rect 213346 51925 213374 51971
rect 146474 51897 213374 51925
rect 213538 51925 213566 51971
rect 331120 51959 331126 52011
rect 331178 51999 331184 52011
rect 342544 51999 342550 52011
rect 331178 51971 342550 51999
rect 331178 51959 331184 51971
rect 342544 51959 342550 51971
rect 342602 51959 342608 52011
rect 460816 51959 460822 52011
rect 460874 51999 460880 52011
rect 470800 51999 470806 52011
rect 460874 51971 470806 51999
rect 460874 51959 460880 51971
rect 470800 51959 470806 51971
rect 470858 51959 470864 52011
rect 625936 51959 625942 52011
rect 625994 51999 626000 52011
rect 639664 51999 639670 52011
rect 625994 51971 639670 51999
rect 625994 51959 626000 51971
rect 639664 51959 639670 51971
rect 639722 51959 639728 52011
rect 227536 51925 227542 51937
rect 213538 51897 227542 51925
rect 146474 51885 146480 51897
rect 227536 51885 227542 51897
rect 227594 51885 227600 51937
rect 541360 51925 541366 51937
rect 282274 51897 302366 51925
rect 213424 51811 213430 51863
rect 213482 51851 213488 51863
rect 237424 51851 237430 51863
rect 213482 51823 237430 51851
rect 213482 51811 213488 51823
rect 237424 51811 237430 51823
rect 237482 51811 237488 51863
rect 239056 51811 239062 51863
rect 239114 51851 239120 51863
rect 244144 51851 244150 51863
rect 239114 51823 244150 51851
rect 239114 51811 239120 51823
rect 244144 51811 244150 51823
rect 244202 51811 244208 51863
rect 254416 51811 254422 51863
rect 254474 51851 254480 51863
rect 282274 51851 282302 51897
rect 254474 51823 282302 51851
rect 254474 51811 254480 51823
rect 211216 51737 211222 51789
rect 211274 51777 211280 51789
rect 302338 51777 302366 51897
rect 388738 51897 388862 51925
rect 322576 51811 322582 51863
rect 322634 51851 322640 51863
rect 331120 51851 331126 51863
rect 322634 51823 331126 51851
rect 322634 51811 322640 51823
rect 331120 51811 331126 51823
rect 331178 51811 331184 51863
rect 342736 51811 342742 51863
rect 342794 51851 342800 51863
rect 368464 51851 368470 51863
rect 342794 51823 368470 51851
rect 342794 51811 342800 51823
rect 368464 51811 368470 51823
rect 368522 51811 368528 51863
rect 368560 51811 368566 51863
rect 368618 51851 368624 51863
rect 388738 51851 388766 51897
rect 368618 51823 388766 51851
rect 388834 51851 388862 51897
rect 429058 51897 429182 51925
rect 408880 51851 408886 51863
rect 388834 51823 408886 51851
rect 368618 51811 368624 51823
rect 408880 51811 408886 51823
rect 408938 51811 408944 51863
rect 408976 51811 408982 51863
rect 409034 51851 409040 51863
rect 429058 51851 429086 51897
rect 409034 51823 429086 51851
rect 429154 51851 429182 51897
rect 538594 51897 541366 51925
rect 449200 51851 449206 51863
rect 429154 51823 449206 51851
rect 409034 51811 409040 51823
rect 449200 51811 449206 51823
rect 449258 51811 449264 51863
rect 449296 51811 449302 51863
rect 449354 51851 449360 51863
rect 460816 51851 460822 51863
rect 449354 51823 460822 51851
rect 449354 51811 449360 51823
rect 460816 51811 460822 51823
rect 460874 51811 460880 51863
rect 509776 51811 509782 51863
rect 509834 51851 509840 51863
rect 538594 51851 538622 51897
rect 541360 51885 541366 51897
rect 541418 51885 541424 51937
rect 558736 51925 558742 51937
rect 558658 51897 558742 51925
rect 509834 51823 518366 51851
rect 509834 51811 509840 51823
rect 308080 51777 308086 51789
rect 211274 51749 227486 51777
rect 302338 51749 308086 51777
rect 211274 51737 211280 51749
rect 209872 51663 209878 51715
rect 209930 51703 209936 51715
rect 214096 51703 214102 51715
rect 209930 51675 214102 51703
rect 209930 51663 209936 51675
rect 214096 51663 214102 51675
rect 214154 51663 214160 51715
rect 227458 51703 227486 51749
rect 308080 51737 308086 51749
rect 308138 51737 308144 51789
rect 308176 51737 308182 51789
rect 308234 51777 308240 51789
rect 322480 51777 322486 51789
rect 308234 51749 322486 51777
rect 308234 51737 308240 51749
rect 322480 51737 322486 51749
rect 322538 51737 322544 51789
rect 518338 51777 518366 51823
rect 527362 51823 538622 51851
rect 527362 51777 527390 51823
rect 541456 51811 541462 51863
rect 541514 51851 541520 51863
rect 558658 51851 558686 51897
rect 558736 51885 558742 51897
rect 558794 51885 558800 51937
rect 625090 51897 635006 51925
rect 590320 51851 590326 51863
rect 541514 51823 558686 51851
rect 584578 51823 590326 51851
rect 541514 51811 541520 51823
rect 518338 51749 527390 51777
rect 558832 51737 558838 51789
rect 558890 51777 558896 51789
rect 584578 51777 584606 51823
rect 590320 51811 590326 51823
rect 590378 51811 590384 51863
rect 590416 51811 590422 51863
rect 590474 51851 590480 51863
rect 625090 51851 625118 51897
rect 590474 51823 610526 51851
rect 590474 51811 590480 51823
rect 558890 51749 584606 51777
rect 610498 51777 610526 51823
rect 624898 51823 625118 51851
rect 624898 51777 624926 51823
rect 610498 51749 624926 51777
rect 634978 51777 635006 51897
rect 645520 51777 645526 51789
rect 634978 51749 645526 51777
rect 558890 51737 558896 51749
rect 645520 51737 645526 51749
rect 645578 51737 645584 51789
rect 251920 51703 251926 51715
rect 227458 51675 251926 51703
rect 251920 51663 251926 51675
rect 251978 51663 251984 51715
rect 322384 51703 322390 51715
rect 273538 51675 282110 51703
rect 209584 51589 209590 51641
rect 209642 51629 209648 51641
rect 214480 51629 214486 51641
rect 209642 51601 214486 51629
rect 209642 51589 209648 51601
rect 214480 51589 214486 51601
rect 214538 51589 214544 51641
rect 253552 51589 253558 51641
rect 253610 51629 253616 51641
rect 273538 51629 273566 51675
rect 253610 51601 273566 51629
rect 282082 51629 282110 51675
rect 308290 51675 322390 51703
rect 308080 51629 308086 51641
rect 282082 51601 308086 51629
rect 253610 51589 253616 51601
rect 308080 51589 308086 51601
rect 308138 51589 308144 51641
rect 308176 51589 308182 51641
rect 308234 51629 308240 51641
rect 308290 51629 308318 51675
rect 322384 51663 322390 51675
rect 322442 51663 322448 51715
rect 414640 51703 414646 51715
rect 397282 51675 414646 51703
rect 308234 51601 308318 51629
rect 322690 51601 334142 51629
rect 308234 51589 308240 51601
rect 145360 51515 145366 51567
rect 145418 51555 145424 51567
rect 236752 51555 236758 51567
rect 145418 51527 236758 51555
rect 145418 51515 145424 51527
rect 236752 51515 236758 51527
rect 236810 51515 236816 51567
rect 237424 51515 237430 51567
rect 237482 51555 237488 51567
rect 237482 51527 251294 51555
rect 237482 51515 237488 51527
rect 145936 51441 145942 51493
rect 145994 51481 146000 51493
rect 237136 51481 237142 51493
rect 145994 51453 237142 51481
rect 145994 51441 146000 51453
rect 237136 51441 237142 51453
rect 237194 51441 237200 51493
rect 144784 51367 144790 51419
rect 144842 51407 144848 51419
rect 233584 51407 233590 51419
rect 144842 51379 233590 51407
rect 144842 51367 144848 51379
rect 233584 51367 233590 51379
rect 233642 51367 233648 51419
rect 251266 51407 251294 51527
rect 322384 51515 322390 51567
rect 322442 51555 322448 51567
rect 322690 51555 322718 51601
rect 322442 51527 322718 51555
rect 334114 51555 334142 51601
rect 342736 51589 342742 51641
rect 342794 51629 342800 51641
rect 342794 51601 354206 51629
rect 342794 51589 342800 51601
rect 342640 51555 342646 51567
rect 334114 51527 342646 51555
rect 322442 51515 322448 51527
rect 342640 51515 342646 51527
rect 342698 51515 342704 51567
rect 354178 51555 354206 51601
rect 362992 51589 362998 51641
rect 363050 51629 363056 51641
rect 374416 51629 374422 51641
rect 363050 51601 374422 51629
rect 363050 51589 363056 51601
rect 374416 51589 374422 51601
rect 374474 51589 374480 51641
rect 394480 51589 394486 51641
rect 394538 51629 394544 51641
rect 397282 51629 397310 51675
rect 414640 51663 414646 51675
rect 414698 51663 414704 51715
rect 470800 51663 470806 51715
rect 470858 51703 470864 51715
rect 509680 51703 509686 51715
rect 470858 51675 509686 51703
rect 470858 51663 470864 51675
rect 509680 51663 509686 51675
rect 509738 51663 509744 51715
rect 518320 51663 518326 51715
rect 518378 51703 518384 51715
rect 518378 51675 528158 51703
rect 518378 51663 518384 51675
rect 423280 51629 423286 51641
rect 394538 51601 397310 51629
rect 420514 51601 423286 51629
rect 394538 51589 394544 51601
rect 362800 51555 362806 51567
rect 354178 51527 362806 51555
rect 362800 51515 362806 51527
rect 362858 51515 362864 51567
rect 417520 51515 417526 51567
rect 417578 51555 417584 51567
rect 420514 51555 420542 51601
rect 423280 51589 423286 51601
rect 423338 51589 423344 51641
rect 423376 51589 423382 51641
rect 423434 51629 423440 51641
rect 457936 51629 457942 51641
rect 423434 51601 457942 51629
rect 423434 51589 423440 51601
rect 457936 51589 457942 51601
rect 457994 51589 458000 51641
rect 480880 51589 480886 51641
rect 480938 51629 480944 51641
rect 498256 51629 498262 51641
rect 480938 51601 498262 51629
rect 480938 51589 480944 51601
rect 498256 51589 498262 51601
rect 498314 51589 498320 51641
rect 528130 51629 528158 51675
rect 604720 51663 604726 51715
rect 604778 51703 604784 51715
rect 604778 51675 610430 51703
rect 604778 51663 604784 51675
rect 538576 51629 538582 51641
rect 528130 51601 538582 51629
rect 538576 51589 538582 51601
rect 538634 51589 538640 51641
rect 541456 51589 541462 51641
rect 541514 51629 541520 51641
rect 584656 51629 584662 51641
rect 541514 51601 558686 51629
rect 541514 51589 541520 51601
rect 417578 51527 420542 51555
rect 558658 51555 558686 51601
rect 561442 51601 584662 51629
rect 561442 51555 561470 51601
rect 584656 51589 584662 51601
rect 584714 51589 584720 51641
rect 558658 51527 561470 51555
rect 610402 51555 610430 51675
rect 625936 51629 625942 51641
rect 611938 51601 625942 51629
rect 611938 51555 611966 51601
rect 625936 51589 625942 51601
rect 625994 51589 626000 51641
rect 610402 51527 611966 51555
rect 417578 51515 417584 51527
rect 251920 51441 251926 51493
rect 251978 51481 251984 51493
rect 253456 51481 253462 51493
rect 251978 51453 253462 51481
rect 251978 51441 251984 51453
rect 253456 51441 253462 51453
rect 253514 51441 253520 51493
rect 478000 51441 478006 51493
rect 478058 51481 478064 51493
rect 480880 51481 480886 51493
rect 478058 51453 480886 51481
rect 478058 51441 478064 51453
rect 480880 51441 480886 51453
rect 480938 51441 480944 51493
rect 254416 51407 254422 51419
rect 251266 51379 254422 51407
rect 254416 51367 254422 51379
rect 254474 51367 254480 51419
rect 414640 51367 414646 51419
rect 414698 51407 414704 51419
rect 417520 51407 417526 51419
rect 414698 51379 417526 51407
rect 414698 51367 414704 51379
rect 417520 51367 417526 51379
rect 417578 51367 417584 51419
rect 144976 51293 144982 51345
rect 145034 51333 145040 51345
rect 234544 51333 234550 51345
rect 145034 51305 234550 51333
rect 145034 51293 145040 51305
rect 234544 51293 234550 51305
rect 234602 51293 234608 51345
rect 145648 51219 145654 51271
rect 145706 51259 145712 51271
rect 235312 51259 235318 51271
rect 145706 51231 235318 51259
rect 145706 51219 145712 51231
rect 235312 51219 235318 51231
rect 235370 51219 235376 51271
rect 145840 51145 145846 51197
rect 145898 51185 145904 51197
rect 234928 51185 234934 51197
rect 145898 51157 234934 51185
rect 145898 51145 145904 51157
rect 234928 51145 234934 51157
rect 234986 51145 234992 51197
rect 146224 51071 146230 51123
rect 146282 51111 146288 51123
rect 232336 51111 232342 51123
rect 146282 51083 232342 51111
rect 146282 51071 146288 51083
rect 232336 51071 232342 51083
rect 232394 51071 232400 51123
rect 146800 50997 146806 51049
rect 146858 51037 146864 51049
rect 231952 51037 231958 51049
rect 146858 51009 231958 51037
rect 146858 50997 146864 51009
rect 231952 50997 231958 51009
rect 232010 50997 232016 51049
rect 146608 50923 146614 50975
rect 146666 50963 146672 50975
rect 230992 50963 230998 50975
rect 146666 50935 230998 50963
rect 146666 50923 146672 50935
rect 230992 50923 230998 50935
rect 231050 50923 231056 50975
rect 145552 50849 145558 50901
rect 145610 50889 145616 50901
rect 231376 50889 231382 50901
rect 145610 50861 231382 50889
rect 145610 50849 145616 50861
rect 231376 50849 231382 50861
rect 231434 50849 231440 50901
rect 146032 50775 146038 50827
rect 146090 50815 146096 50827
rect 230512 50815 230518 50827
rect 146090 50787 230518 50815
rect 146090 50775 146096 50787
rect 230512 50775 230518 50787
rect 230570 50775 230576 50827
rect 145072 50701 145078 50753
rect 145130 50741 145136 50753
rect 228304 50741 228310 50753
rect 145130 50713 228310 50741
rect 145130 50701 145136 50713
rect 228304 50701 228310 50713
rect 228362 50701 228368 50753
rect 145456 50627 145462 50679
rect 145514 50667 145520 50679
rect 228688 50667 228694 50679
rect 145514 50639 228694 50667
rect 145514 50627 145520 50639
rect 228688 50627 228694 50639
rect 228746 50627 228752 50679
rect 145264 50553 145270 50605
rect 145322 50593 145328 50605
rect 229744 50593 229750 50605
rect 145322 50565 229750 50593
rect 145322 50553 145328 50565
rect 229744 50553 229750 50565
rect 229802 50553 229808 50605
rect 145168 50479 145174 50531
rect 145226 50519 145232 50531
rect 228784 50519 228790 50531
rect 145226 50491 228790 50519
rect 145226 50479 145232 50491
rect 228784 50479 228790 50491
rect 228842 50479 228848 50531
rect 144496 50405 144502 50457
rect 144554 50445 144560 50457
rect 208048 50445 208054 50457
rect 144554 50417 208054 50445
rect 144554 50405 144560 50417
rect 208048 50405 208054 50417
rect 208106 50405 208112 50457
rect 144112 50331 144118 50383
rect 144170 50371 144176 50383
rect 207952 50371 207958 50383
rect 144170 50343 207958 50371
rect 144170 50331 144176 50343
rect 207952 50331 207958 50343
rect 208010 50331 208016 50383
rect 208240 50331 208246 50383
rect 208298 50371 208304 50383
rect 216112 50371 216118 50383
rect 208298 50343 216118 50371
rect 208298 50331 208304 50343
rect 216112 50331 216118 50343
rect 216170 50331 216176 50383
rect 146128 50257 146134 50309
rect 146186 50297 146192 50309
rect 207856 50297 207862 50309
rect 146186 50269 207862 50297
rect 146186 50257 146192 50269
rect 207856 50257 207862 50269
rect 207914 50257 207920 50309
rect 208432 50257 208438 50309
rect 208490 50297 208496 50309
rect 216880 50297 216886 50309
rect 208490 50269 216886 50297
rect 208490 50257 208496 50269
rect 216880 50257 216886 50269
rect 216938 50257 216944 50309
rect 144304 50183 144310 50235
rect 144362 50223 144368 50235
rect 208336 50223 208342 50235
rect 144362 50195 208342 50223
rect 144362 50183 144368 50195
rect 208336 50183 208342 50195
rect 208394 50183 208400 50235
rect 208528 50183 208534 50235
rect 208586 50223 208592 50235
rect 217648 50223 217654 50235
rect 208586 50195 217654 50223
rect 208586 50183 208592 50195
rect 217648 50183 217654 50195
rect 217706 50183 217712 50235
rect 144208 50109 144214 50161
rect 144266 50149 144272 50161
rect 235792 50149 235798 50161
rect 144266 50121 235798 50149
rect 144266 50109 144272 50121
rect 235792 50109 235798 50121
rect 235850 50109 235856 50161
rect 146512 50035 146518 50087
rect 146570 50075 146576 50087
rect 235408 50075 235414 50087
rect 146570 50047 235414 50075
rect 146570 50035 146576 50047
rect 235408 50035 235414 50047
rect 235466 50035 235472 50087
rect 144688 49961 144694 50013
rect 144746 50001 144752 50013
rect 232720 50001 232726 50013
rect 144746 49973 232726 50001
rect 144746 49961 144752 49973
rect 232720 49961 232726 49973
rect 232778 49961 232784 50013
rect 208048 49887 208054 49939
rect 208106 49927 208112 49939
rect 224944 49927 224950 49939
rect 208106 49899 224950 49927
rect 208106 49887 208112 49899
rect 224944 49887 224950 49899
rect 225002 49887 225008 49939
rect 208336 49813 208342 49865
rect 208394 49853 208400 49865
rect 224272 49853 224278 49865
rect 208394 49825 224278 49853
rect 208394 49813 208400 49825
rect 224272 49813 224278 49825
rect 224330 49813 224336 49865
rect 207952 49739 207958 49791
rect 208010 49779 208016 49791
rect 225328 49779 225334 49791
rect 208010 49751 225334 49779
rect 208010 49739 208016 49751
rect 225328 49739 225334 49751
rect 225386 49739 225392 49791
rect 645808 49779 645814 49791
rect 225442 49751 645814 49779
rect 145744 49665 145750 49717
rect 145802 49705 145808 49717
rect 145802 49677 178622 49705
rect 145802 49665 145808 49677
rect 178594 49631 178622 49677
rect 211600 49665 211606 49717
rect 211658 49705 211664 49717
rect 225442 49705 225470 49751
rect 645808 49739 645814 49751
rect 645866 49739 645872 49791
rect 211658 49677 225470 49705
rect 211658 49665 211664 49677
rect 178594 49603 205886 49631
rect 205858 49557 205886 49603
rect 207856 49591 207862 49643
rect 207914 49631 207920 49643
rect 226576 49631 226582 49643
rect 207914 49603 226582 49631
rect 207914 49591 207920 49603
rect 226576 49591 226582 49603
rect 226634 49591 226640 49643
rect 205858 49529 215870 49557
rect 215842 49495 215870 49529
rect 215824 49443 215830 49495
rect 215882 49443 215888 49495
rect 215920 49443 215926 49495
rect 215978 49483 215984 49495
rect 218800 49483 218806 49495
rect 215978 49455 218806 49483
rect 215978 49443 215984 49455
rect 218800 49443 218806 49455
rect 218858 49443 218864 49495
rect 218800 49295 218806 49347
rect 218858 49335 218864 49347
rect 241168 49335 241174 49347
rect 218858 49307 241174 49335
rect 218858 49295 218864 49307
rect 241168 49295 241174 49307
rect 241226 49295 241232 49347
rect 443440 48999 443446 49051
rect 443498 49039 443504 49051
rect 443498 49011 460862 49039
rect 443498 48999 443504 49011
rect 210064 48925 210070 48977
rect 210122 48965 210128 48977
rect 220720 48965 220726 48977
rect 210122 48937 220726 48965
rect 210122 48925 210128 48937
rect 220720 48925 220726 48937
rect 220778 48925 220784 48977
rect 223696 48925 223702 48977
rect 223754 48965 223760 48977
rect 229648 48965 229654 48977
rect 223754 48937 229654 48965
rect 223754 48925 223760 48937
rect 229648 48925 229654 48937
rect 229706 48925 229712 48977
rect 282352 48925 282358 48977
rect 282410 48965 282416 48977
rect 302416 48965 302422 48977
rect 282410 48937 302422 48965
rect 282410 48925 282416 48937
rect 302416 48925 302422 48937
rect 302474 48925 302480 48977
rect 460834 48965 460862 49011
rect 471376 48965 471382 48977
rect 460834 48937 471382 48965
rect 471376 48925 471382 48937
rect 471434 48925 471440 48977
rect 222256 48851 222262 48903
rect 222314 48891 222320 48903
rect 645136 48891 645142 48903
rect 222314 48863 645142 48891
rect 222314 48851 222320 48863
rect 645136 48851 645142 48863
rect 645194 48851 645200 48903
rect 209008 48777 209014 48829
rect 209066 48817 209072 48829
rect 222064 48817 222070 48829
rect 209066 48789 222070 48817
rect 209066 48777 209072 48789
rect 222064 48777 222070 48789
rect 222122 48777 222128 48829
rect 222928 48777 222934 48829
rect 222986 48817 222992 48829
rect 645232 48817 645238 48829
rect 222986 48789 645238 48817
rect 222986 48777 222992 48789
rect 645232 48777 645238 48789
rect 645290 48777 645296 48829
rect 208624 48703 208630 48755
rect 208682 48743 208688 48755
rect 221680 48743 221686 48755
rect 208682 48715 221686 48743
rect 208682 48703 208688 48715
rect 221680 48703 221686 48715
rect 221738 48703 221744 48755
rect 224080 48703 224086 48755
rect 224138 48743 224144 48755
rect 645328 48743 645334 48755
rect 224138 48715 645334 48743
rect 224138 48703 224144 48715
rect 645328 48703 645334 48715
rect 645386 48703 645392 48755
rect 148240 48629 148246 48681
rect 148298 48669 148304 48681
rect 236368 48669 236374 48681
rect 148298 48641 236374 48669
rect 148298 48629 148304 48641
rect 236368 48629 236374 48641
rect 236426 48629 236432 48681
rect 148816 48555 148822 48607
rect 148874 48595 148880 48607
rect 234160 48595 234166 48607
rect 148874 48567 234166 48595
rect 148874 48555 148880 48567
rect 234160 48555 234166 48567
rect 234218 48555 234224 48607
rect 185680 48481 185686 48533
rect 185738 48521 185744 48533
rect 240208 48521 240214 48533
rect 185738 48493 240214 48521
rect 185738 48481 185744 48493
rect 240208 48481 240214 48493
rect 240266 48481 240272 48533
rect 197200 48407 197206 48459
rect 197258 48447 197264 48459
rect 239824 48447 239830 48459
rect 197258 48419 239830 48447
rect 197258 48407 197264 48419
rect 239824 48407 239830 48419
rect 239882 48407 239888 48459
rect 194320 48333 194326 48385
rect 194378 48373 194384 48385
rect 239728 48373 239734 48385
rect 194378 48345 239734 48373
rect 194378 48333 194384 48345
rect 239728 48333 239734 48345
rect 239786 48333 239792 48385
rect 202960 48259 202966 48311
rect 203018 48299 203024 48311
rect 241552 48299 241558 48311
rect 203018 48271 241558 48299
rect 203018 48259 203024 48271
rect 241552 48259 241558 48271
rect 241610 48259 241616 48311
rect 149296 48185 149302 48237
rect 149354 48225 149360 48237
rect 208528 48225 208534 48237
rect 149354 48197 208534 48225
rect 149354 48185 149360 48197
rect 208528 48185 208534 48197
rect 208586 48185 208592 48237
rect 208912 48185 208918 48237
rect 208970 48225 208976 48237
rect 222448 48225 222454 48237
rect 208970 48197 222454 48225
rect 208970 48185 208976 48197
rect 222448 48185 222454 48197
rect 222506 48185 222512 48237
rect 149392 48111 149398 48163
rect 149450 48151 149456 48163
rect 208624 48151 208630 48163
rect 149450 48123 208630 48151
rect 149450 48111 149456 48123
rect 208624 48111 208630 48123
rect 208682 48111 208688 48163
rect 208816 48111 208822 48163
rect 208874 48151 208880 48163
rect 222736 48151 222742 48163
rect 208874 48123 222742 48151
rect 208874 48111 208880 48123
rect 222736 48111 222742 48123
rect 222794 48111 222800 48163
rect 148048 48037 148054 48089
rect 148106 48077 148112 48089
rect 219472 48077 219478 48089
rect 148106 48049 219478 48077
rect 148106 48037 148112 48049
rect 219472 48037 219478 48049
rect 219530 48037 219536 48089
rect 148144 47963 148150 48015
rect 148202 48003 148208 48015
rect 219088 48003 219094 48015
rect 148202 47975 219094 48003
rect 148202 47963 148208 47975
rect 219088 47963 219094 47975
rect 219146 47963 219152 48015
rect 149488 47889 149494 47941
rect 149546 47929 149552 47941
rect 221296 47929 221302 47941
rect 149546 47901 221302 47929
rect 149546 47889 149552 47901
rect 221296 47889 221302 47901
rect 221354 47889 221360 47941
rect 149584 47815 149590 47867
rect 149642 47855 149648 47867
rect 220528 47855 220534 47867
rect 149642 47827 220534 47855
rect 149642 47815 149648 47827
rect 220528 47815 220534 47827
rect 220586 47815 220592 47867
rect 149680 47741 149686 47793
rect 149738 47781 149744 47793
rect 220240 47781 220246 47793
rect 149738 47753 220246 47781
rect 149738 47741 149744 47753
rect 220240 47741 220246 47753
rect 220298 47741 220304 47793
rect 147664 47667 147670 47719
rect 147722 47707 147728 47719
rect 216496 47707 216502 47719
rect 147722 47679 216502 47707
rect 147722 47667 147728 47679
rect 216496 47667 216502 47679
rect 216554 47667 216560 47719
rect 147760 47593 147766 47645
rect 147818 47633 147824 47645
rect 218032 47633 218038 47645
rect 147818 47605 218038 47633
rect 147818 47593 147824 47605
rect 218032 47593 218038 47605
rect 218090 47593 218096 47645
rect 218512 47593 218518 47645
rect 218570 47633 218576 47645
rect 645616 47633 645622 47645
rect 218570 47605 645622 47633
rect 218570 47593 218576 47605
rect 645616 47593 645622 47605
rect 645674 47593 645680 47645
rect 147952 47519 147958 47571
rect 148010 47559 148016 47571
rect 218704 47559 218710 47571
rect 148010 47531 218710 47559
rect 148010 47519 148016 47531
rect 218704 47519 218710 47531
rect 218762 47519 218768 47571
rect 147856 47445 147862 47497
rect 147914 47485 147920 47497
rect 218320 47485 218326 47497
rect 147914 47457 218326 47485
rect 147914 47445 147920 47457
rect 218320 47445 218326 47457
rect 218378 47445 218384 47497
rect 177040 47371 177046 47423
rect 177098 47411 177104 47423
rect 238000 47411 238006 47423
rect 177098 47383 238006 47411
rect 177098 47371 177104 47383
rect 238000 47371 238006 47383
rect 238058 47371 238064 47423
rect 179920 47297 179926 47349
rect 179978 47337 179984 47349
rect 238576 47337 238582 47349
rect 179978 47309 238582 47337
rect 179978 47297 179984 47309
rect 238576 47297 238582 47309
rect 238634 47297 238640 47349
rect 200080 47223 200086 47275
rect 200138 47263 200144 47275
rect 238960 47263 238966 47275
rect 200138 47235 238966 47263
rect 200138 47223 200144 47235
rect 238960 47223 238966 47235
rect 239018 47223 239024 47275
rect 148912 47149 148918 47201
rect 148970 47189 148976 47201
rect 233296 47189 233302 47201
rect 148970 47161 233302 47189
rect 148970 47149 148976 47161
rect 233296 47149 233302 47161
rect 233354 47149 233360 47201
rect 188560 47075 188566 47127
rect 188618 47115 188624 47127
rect 239344 47115 239350 47127
rect 188618 47087 239350 47115
rect 188618 47075 188624 47087
rect 239344 47075 239350 47087
rect 239402 47075 239408 47127
rect 148528 47001 148534 47053
rect 148586 47041 148592 47053
rect 230896 47041 230902 47053
rect 148586 47013 230902 47041
rect 148586 47001 148592 47013
rect 230896 47001 230902 47013
rect 230954 47001 230960 47053
rect 191440 46927 191446 46979
rect 191498 46967 191504 46979
rect 240784 46967 240790 46979
rect 191498 46939 240790 46967
rect 191498 46927 191504 46939
rect 240784 46927 240790 46939
rect 240842 46927 240848 46979
rect 148720 46853 148726 46905
rect 148778 46893 148784 46905
rect 227920 46893 227926 46905
rect 148778 46865 227926 46893
rect 148778 46853 148784 46865
rect 227920 46853 227926 46865
rect 227978 46853 227984 46905
rect 148432 46779 148438 46831
rect 148490 46819 148496 46831
rect 233104 46819 233110 46831
rect 148490 46791 233110 46819
rect 148490 46779 148496 46791
rect 233104 46779 233110 46791
rect 233162 46779 233168 46831
rect 149200 46705 149206 46757
rect 149258 46745 149264 46757
rect 208432 46745 208438 46757
rect 149258 46717 208438 46745
rect 149258 46705 149264 46717
rect 208432 46705 208438 46717
rect 208490 46705 208496 46757
rect 208720 46705 208726 46757
rect 208778 46745 208784 46757
rect 223504 46745 223510 46757
rect 208778 46717 223510 46745
rect 208778 46705 208784 46717
rect 223504 46705 223510 46717
rect 223562 46705 223568 46757
rect 149008 46631 149014 46683
rect 149066 46671 149072 46683
rect 230128 46671 230134 46683
rect 149066 46643 230134 46671
rect 149066 46631 149072 46643
rect 230128 46631 230134 46643
rect 230186 46631 230192 46683
rect 207760 46557 207766 46609
rect 207818 46597 207824 46609
rect 223888 46597 223894 46609
rect 207818 46569 223894 46597
rect 207818 46557 207824 46569
rect 223888 46557 223894 46569
rect 223946 46557 223952 46609
rect 149104 46483 149110 46535
rect 149162 46523 149168 46535
rect 208336 46523 208342 46535
rect 149162 46495 208342 46523
rect 149162 46483 149168 46495
rect 208336 46483 208342 46495
rect 208394 46483 208400 46535
rect 208624 46483 208630 46535
rect 208682 46523 208688 46535
rect 223120 46523 223126 46535
rect 208682 46495 223126 46523
rect 208682 46483 208688 46495
rect 223120 46483 223126 46495
rect 223178 46483 223184 46535
rect 148624 46409 148630 46461
rect 148682 46449 148688 46461
rect 229168 46449 229174 46461
rect 148682 46421 229174 46449
rect 148682 46409 148688 46421
rect 229168 46409 229174 46421
rect 229226 46409 229232 46461
rect 208528 46335 208534 46387
rect 208586 46375 208592 46387
rect 224656 46375 224662 46387
rect 208586 46347 224662 46375
rect 208586 46335 208592 46347
rect 224656 46335 224662 46347
rect 224714 46335 224720 46387
rect 208432 46261 208438 46313
rect 208490 46301 208496 46313
rect 226096 46301 226102 46313
rect 208490 46273 226102 46301
rect 208490 46261 208496 46273
rect 226096 46261 226102 46273
rect 226154 46261 226160 46313
rect 208336 46187 208342 46239
rect 208394 46227 208400 46239
rect 226480 46227 226486 46239
rect 208394 46199 226486 46227
rect 208394 46187 208400 46199
rect 226480 46187 226486 46199
rect 226538 46187 226544 46239
rect 398320 46113 398326 46165
rect 398378 46153 398384 46165
rect 398378 46125 403262 46153
rect 398378 46113 398384 46125
rect 403234 46079 403262 46125
rect 408880 46079 408886 46091
rect 403234 46051 408886 46079
rect 408880 46039 408886 46051
rect 408938 46039 408944 46091
rect 211408 45299 211414 45351
rect 211466 45339 211472 45351
rect 361744 45339 361750 45351
rect 211466 45311 361750 45339
rect 211466 45299 211472 45311
rect 361744 45299 361750 45311
rect 361802 45299 361808 45351
rect 213232 45225 213238 45277
rect 213290 45265 213296 45277
rect 406096 45265 406102 45277
rect 213290 45237 406102 45265
rect 213290 45225 213296 45237
rect 406096 45225 406102 45237
rect 406154 45225 406160 45277
rect 212848 45151 212854 45203
rect 212906 45191 212912 45203
rect 411568 45191 411574 45203
rect 212906 45163 411574 45191
rect 212906 45151 212912 45163
rect 411568 45151 411574 45163
rect 411626 45151 411632 45203
rect 213904 45077 213910 45129
rect 213962 45117 213968 45129
rect 443920 45117 443926 45129
rect 213962 45089 443926 45117
rect 213962 45077 213968 45089
rect 443920 45077 443926 45089
rect 443978 45077 443984 45129
rect 215056 45003 215062 45055
rect 215114 45043 215120 45055
rect 509680 45043 509686 45055
rect 215114 45015 509686 45043
rect 215114 45003 215120 45015
rect 509680 45003 509686 45015
rect 509738 45003 509744 45055
rect 214672 44929 214678 44981
rect 214730 44969 214736 44981
rect 508240 44969 508246 44981
rect 214730 44941 508246 44969
rect 214730 44929 214736 44941
rect 508240 44929 508246 44941
rect 508298 44929 508304 44981
rect 508240 43227 508246 43279
rect 508298 43267 508304 43279
rect 508298 43239 521534 43267
rect 508298 43227 508304 43239
rect 521506 43205 521534 43239
rect 406096 43153 406102 43205
rect 406154 43193 406160 43205
rect 410992 43193 410998 43205
rect 406154 43165 410998 43193
rect 406154 43153 406160 43165
rect 410992 43153 410998 43165
rect 411050 43153 411056 43205
rect 521488 43153 521494 43205
rect 521546 43153 521552 43205
rect 133648 42783 133654 42835
rect 133706 42823 133712 42835
rect 136528 42823 136534 42835
rect 133706 42795 136534 42823
rect 133706 42783 133712 42795
rect 136528 42783 136534 42795
rect 136586 42783 136592 42835
rect 212464 42339 212470 42391
rect 212522 42379 212528 42391
rect 310096 42379 310102 42391
rect 212522 42351 310102 42379
rect 212522 42339 212528 42351
rect 310096 42339 310102 42351
rect 310154 42339 310160 42391
rect 206896 42117 206902 42169
rect 206954 42157 206960 42169
rect 405232 42157 405238 42169
rect 206954 42129 405238 42157
rect 206954 42117 206960 42129
rect 405232 42117 405238 42129
rect 405290 42117 405296 42169
rect 213616 42043 213622 42095
rect 213674 42083 213680 42095
rect 460048 42083 460054 42095
rect 213674 42055 460054 42083
rect 213674 42043 213680 42055
rect 460048 42043 460054 42055
rect 460106 42043 460112 42095
rect 214288 41969 214294 42021
rect 214346 42009 214352 42021
rect 514864 42009 514870 42021
rect 214346 41981 514870 42009
rect 214346 41969 214352 41981
rect 514864 41969 514870 41981
rect 514922 41969 514928 42021
rect 459184 41525 459190 41577
rect 459242 41565 459248 41577
rect 464194 41565 464222 41786
rect 459242 41537 464222 41565
rect 459242 41525 459248 41537
rect 443920 37381 443926 37433
rect 443978 37421 443984 37433
rect 459184 37421 459190 37433
rect 443978 37393 459190 37421
rect 443978 37381 443984 37393
rect 459184 37381 459190 37393
rect 459242 37381 459248 37433
<< via1 >>
rect 452182 1008113 452234 1008165
rect 472150 1008113 472202 1008165
rect 434998 1008039 435050 1008091
rect 471574 1008039 471626 1008091
rect 434710 1007965 434762 1008017
rect 452182 1007965 452234 1008017
rect 367222 1005449 367274 1005501
rect 383638 1005449 383690 1005501
rect 434614 1005449 434666 1005501
rect 471862 1005449 471914 1005501
rect 434902 1005301 434954 1005353
rect 469366 1005301 469418 1005353
rect 164278 1005227 164330 1005279
rect 172822 1005227 172874 1005279
rect 437494 1005227 437546 1005279
rect 470134 1005227 470186 1005279
rect 218806 1005153 218858 1005205
rect 222646 1005153 222698 1005205
rect 316822 1005153 316874 1005205
rect 331222 1005153 331274 1005205
rect 195286 1003229 195338 1003281
rect 377302 1003229 377354 1003281
rect 434614 1003229 434666 1003281
rect 439126 1003229 439178 1003281
rect 466486 1003229 466538 1003281
rect 519670 1003229 519722 1003281
rect 160438 1003155 160490 1003207
rect 164278 1003155 164330 1003207
rect 209110 1003155 209162 1003207
rect 211798 1003155 211850 1003207
rect 213814 1003155 213866 1003207
rect 357430 1003155 357482 1003207
rect 362518 1003155 362570 1003207
rect 367222 1003155 367274 1003207
rect 428662 1003155 428714 1003207
rect 429526 1003155 429578 1003207
rect 466390 1003155 466442 1003207
rect 502390 1003155 502442 1003207
rect 425398 1003081 425450 1003133
rect 466294 1003081 466346 1003133
rect 428278 1003007 428330 1003059
rect 429142 1003007 429194 1003059
rect 430294 1003007 430346 1003059
rect 434902 1003007 434954 1003059
rect 435382 1003007 435434 1003059
rect 466198 1003007 466250 1003059
rect 501334 1003007 501386 1003059
rect 519766 1003155 519818 1003207
rect 502966 1003007 503018 1003059
rect 519862 1003007 519914 1003059
rect 555382 1003007 555434 1003059
rect 572758 1003007 572810 1003059
rect 161494 1002933 161546 1002985
rect 169942 1002933 169994 1002985
rect 298294 1002933 298346 1002985
rect 312118 1002933 312170 1002985
rect 426070 1002933 426122 1002985
rect 299350 1002859 299402 1002911
rect 308854 1002859 308906 1002911
rect 423862 1002859 423914 1002911
rect 435382 1002859 435434 1002911
rect 299446 1002785 299498 1002837
rect 309334 1002785 309386 1002837
rect 424342 1002785 424394 1002837
rect 429526 1002785 429578 1002837
rect 432022 1002785 432074 1002837
rect 434998 1002785 435050 1002837
rect 439222 1002933 439274 1002985
rect 465526 1002933 465578 1002985
rect 554326 1002933 554378 1002985
rect 573046 1002933 573098 1002985
rect 553750 1002859 553802 1002911
rect 570742 1002859 570794 1002911
rect 439222 1002785 439274 1002837
rect 299254 1002711 299306 1002763
rect 308278 1002711 308330 1002763
rect 358582 1002711 358634 1002763
rect 373366 1002711 373418 1002763
rect 424822 1002711 424874 1002763
rect 439126 1002711 439178 1002763
rect 554902 1002711 554954 1002763
rect 571222 1002711 571274 1002763
rect 358006 1002637 358058 1002689
rect 372502 1002637 372554 1002689
rect 427606 1002637 427658 1002689
rect 435094 1002637 435146 1002689
rect 143926 1002563 143978 1002615
rect 153334 1002563 153386 1002615
rect 429238 1002563 429290 1002615
rect 434710 1002563 434762 1002615
rect 553270 1002563 553322 1002615
rect 572950 1002563 573002 1002615
rect 143734 1002489 143786 1002541
rect 152662 1002489 152714 1002541
rect 361846 1002489 361898 1002541
rect 371542 1002489 371594 1002541
rect 426646 1002489 426698 1002541
rect 435190 1002489 435242 1002541
rect 144022 1002415 144074 1002467
rect 151606 1002415 151658 1002467
rect 427126 1002415 427178 1002467
rect 435286 1002415 435338 1002467
rect 143830 1002341 143882 1002393
rect 151030 1002341 151082 1002393
rect 362902 1002341 362954 1002393
rect 371638 1002341 371690 1002393
rect 429142 1002341 429194 1002393
rect 443542 1002341 443594 1002393
rect 144118 1002267 144170 1002319
rect 175702 1002267 175754 1002319
rect 359062 1002267 359114 1002319
rect 365782 1002267 365834 1002319
rect 489142 1002267 489194 1002319
rect 519094 1002267 519146 1002319
rect 361366 1002193 361418 1002245
rect 379990 1002193 380042 1002245
rect 356374 1001231 356426 1001283
rect 379798 1001231 379850 1001283
rect 357142 1001083 357194 1001135
rect 380086 1001083 380138 1001135
rect 465238 1001009 465290 1001061
rect 472534 1001009 472586 1001061
rect 365782 1000935 365834 1000987
rect 383158 1000935 383210 1000987
rect 506326 1000935 506378 1000987
rect 515542 1000935 515594 1000987
rect 360214 1000861 360266 1000913
rect 383446 1000861 383498 1000913
rect 430966 1000861 431018 1000913
rect 472438 1000861 472490 1000913
rect 359638 1000787 359690 1000839
rect 383254 1000787 383306 1000839
rect 429910 1000787 429962 1000839
rect 472630 1000787 472682 1000839
rect 507862 1000787 507914 1000839
rect 512662 1000787 512714 1000839
rect 552310 1000787 552362 1000839
rect 573142 1000787 573194 1000839
rect 506902 1000639 506954 1000691
rect 512182 1000639 512234 1000691
rect 377302 999825 377354 999877
rect 383350 999825 383402 999877
rect 504694 999825 504746 999877
rect 512086 999825 512138 999877
rect 509686 999751 509738 999803
rect 519958 999751 520010 999803
rect 613462 999751 613514 999803
rect 625846 999751 625898 999803
rect 503638 999677 503690 999729
rect 512278 999677 512330 999729
rect 610582 999677 610634 999729
rect 625558 999677 625610 999729
rect 195478 999603 195530 999655
rect 195190 999455 195242 999507
rect 500758 999603 500810 999655
rect 511990 999603 512042 999655
rect 512086 999603 512138 999655
rect 604246 999603 604298 999655
rect 625654 999603 625706 999655
rect 503638 999529 503690 999581
rect 609046 999529 609098 999581
rect 625462 999529 625514 999581
rect 92662 999381 92714 999433
rect 126646 999381 126698 999433
rect 143734 999381 143786 999433
rect 155542 999381 155594 999433
rect 195094 999381 195146 999433
rect 206902 999381 206954 999433
rect 226006 999455 226058 999507
rect 371542 999455 371594 999507
rect 222934 999381 222986 999433
rect 246550 999381 246602 999433
rect 258358 999381 258410 999433
rect 298198 999381 298250 999433
rect 309910 999381 309962 999433
rect 371638 999381 371690 999433
rect 379894 999381 379946 999433
rect 502006 999455 502058 999507
rect 512086 999455 512138 999507
rect 596182 999455 596234 999507
rect 625846 999455 625898 999507
rect 313750 999307 313802 999359
rect 328342 999307 328394 999359
rect 364534 999307 364586 999359
rect 380374 999307 380426 999359
rect 488950 999381 489002 999433
rect 509686 999381 509738 999433
rect 552982 999381 553034 999433
rect 383542 999307 383594 999359
rect 593302 999381 593354 999433
rect 625750 999381 625802 999433
rect 567382 999307 567434 999359
rect 466294 999233 466346 999285
rect 472054 999233 472106 999285
rect 558838 999233 558890 999285
rect 573718 999233 573770 999285
rect 466486 999011 466538 999063
rect 472246 999011 472298 999063
rect 465526 998937 465578 998989
rect 471958 998937 472010 998989
rect 379990 998863 380042 998915
rect 383062 998863 383114 998915
rect 557206 998789 557258 998841
rect 573910 998789 573962 998841
rect 298390 997901 298442 997953
rect 348886 997901 348938 997953
rect 572758 997901 572810 997953
rect 604246 997901 604298 997953
rect 314806 997827 314858 997879
rect 365206 997827 365258 997879
rect 555958 997827 556010 997879
rect 593302 997827 593354 997879
rect 328342 997753 328394 997805
rect 364534 997753 364586 997805
rect 558166 997753 558218 997805
rect 596182 997753 596234 997805
rect 571222 997679 571274 997731
rect 610582 997679 610634 997731
rect 557782 997605 557834 997657
rect 613462 997605 613514 997657
rect 559414 997531 559466 997583
rect 622006 997531 622058 997583
rect 573142 997457 573194 997509
rect 609046 997457 609098 997509
rect 572950 997383 573002 997435
rect 621910 997383 621962 997435
rect 298102 997087 298154 997139
rect 313750 997087 313802 997139
rect 511990 996717 512042 996769
rect 518326 996717 518378 996769
rect 196822 996643 196874 996695
rect 97942 996495 97994 996547
rect 104662 996495 104714 996547
rect 195766 996495 195818 996547
rect 205174 996495 205226 996547
rect 507478 996569 507530 996621
rect 521302 996569 521354 996621
rect 207958 996495 208010 996547
rect 309910 996495 309962 996547
rect 311542 996495 311594 996547
rect 379894 996495 379946 996547
rect 382966 996495 383018 996547
rect 505750 996495 505802 996547
rect 519190 996495 519242 996547
rect 313174 996421 313226 996473
rect 363958 996421 364010 996473
rect 107542 996273 107594 996325
rect 126742 996273 126794 996325
rect 144214 996273 144266 996325
rect 159190 996199 159242 996251
rect 107926 996051 107978 996103
rect 159766 996051 159818 996103
rect 225238 996347 225290 996399
rect 262486 996347 262538 996399
rect 270646 996347 270698 996399
rect 108982 995977 109034 996029
rect 160438 995977 160490 996029
rect 210166 996051 210218 996103
rect 225238 996051 225290 996103
rect 263062 996125 263114 996177
rect 314806 996125 314858 996177
rect 368662 996125 368714 996177
rect 432406 996125 432458 996177
rect 432502 996125 432554 996177
rect 509590 996125 509642 996177
rect 509974 996125 510026 996177
rect 561046 996125 561098 996177
rect 247510 996051 247562 996103
rect 257782 996051 257834 996103
rect 262006 996051 262058 996103
rect 313174 996051 313226 996103
rect 380374 996051 380426 996103
rect 434998 996051 435050 996103
rect 471574 996051 471626 996103
rect 508918 996051 508970 996103
rect 560182 996051 560234 996103
rect 210646 995977 210698 996029
rect 222646 995977 222698 996029
rect 263254 995977 263306 996029
rect 363958 995977 364010 996029
rect 430966 995977 431018 996029
rect 437494 995977 437546 996029
rect 470134 995977 470186 996029
rect 508342 995977 508394 996029
rect 559606 995977 559658 996029
rect 94966 995903 95018 995955
rect 102838 995903 102890 995955
rect 101206 995829 101258 995881
rect 144022 995903 144074 995955
rect 172822 995903 172874 995955
rect 211798 995903 211850 995955
rect 250486 995903 250538 995955
rect 254518 995903 254570 995955
rect 143926 995829 143978 995881
rect 204022 995829 204074 995881
rect 299446 995903 299498 995955
rect 382966 995903 383018 995955
rect 310294 995829 310346 995881
rect 383350 995829 383402 995881
rect 466390 995903 466442 995955
rect 417526 995829 417578 995881
rect 421558 995829 421610 995881
rect 471958 995903 472010 995955
rect 625462 995903 625514 995955
rect 621910 995829 621962 995881
rect 85942 995755 85994 995807
rect 91510 995755 91562 995807
rect 103990 995755 104042 995807
rect 136822 995755 136874 995807
rect 139318 995755 139370 995807
rect 142966 995755 143018 995807
rect 143734 995755 143786 995807
rect 149590 995755 149642 995807
rect 154870 995755 154922 995807
rect 175702 995755 175754 995807
rect 185206 995755 185258 995807
rect 188854 995755 188906 995807
rect 190582 995755 190634 995807
rect 204694 995755 204746 995807
rect 226006 995755 226058 995807
rect 94966 995681 95018 995733
rect 102454 995681 102506 995733
rect 137974 995681 138026 995733
rect 143830 995681 143882 995733
rect 188086 995681 188138 995733
rect 203062 995681 203114 995733
rect 95062 995607 95114 995659
rect 102358 995607 102410 995659
rect 137398 995607 137450 995659
rect 143638 995607 143690 995659
rect 93526 995533 93578 995585
rect 98038 995533 98090 995585
rect 126742 995533 126794 995585
rect 144214 995607 144266 995659
rect 194422 995607 194474 995659
rect 195094 995607 195146 995659
rect 236470 995755 236522 995807
rect 254902 995755 254954 995807
rect 283702 995755 283754 995807
rect 290614 995755 290666 995807
rect 292534 995755 292586 995807
rect 305494 995755 305546 995807
rect 360886 995755 360938 995807
rect 365782 995755 365834 995807
rect 366742 995755 366794 995807
rect 371638 995755 371690 995807
rect 383638 995755 383690 995807
rect 384406 995755 384458 995807
rect 389398 995755 389450 995807
rect 396694 995755 396746 995807
rect 472630 995755 472682 995807
rect 473302 995755 473354 995807
rect 481366 995755 481418 995807
rect 483862 995755 483914 995807
rect 485686 995755 485738 995807
rect 488950 995755 489002 995807
rect 524086 995755 524138 995807
rect 529846 995755 529898 995807
rect 556534 995755 556586 995807
rect 563254 995755 563306 995807
rect 622006 995755 622058 995807
rect 627862 995755 627914 995807
rect 631510 995755 631562 995807
rect 635830 995755 635882 995807
rect 638806 995755 638858 995807
rect 649942 995755 649994 995807
rect 245686 995681 245738 995733
rect 246550 995681 246602 995733
rect 250390 995681 250442 995733
rect 257110 995681 257162 995733
rect 291190 995681 291242 995733
rect 305974 995681 306026 995733
rect 366166 995681 366218 995733
rect 371734 995681 371786 995733
rect 383446 995681 383498 995733
rect 384982 995681 385034 995733
rect 472534 995681 472586 995733
rect 474070 995681 474122 995733
rect 523990 995681 524042 995733
rect 525334 995681 525386 995733
rect 625846 995681 625898 995733
rect 626518 995681 626570 995733
rect 237238 995607 237290 995659
rect 247606 995607 247658 995659
rect 255958 995607 256010 995659
rect 297334 995607 297386 995659
rect 298198 995607 298250 995659
rect 383254 995607 383306 995659
rect 388054 995607 388106 995659
rect 472438 995607 472490 995659
rect 474646 995607 474698 995659
rect 523894 995607 523946 995659
rect 524758 995607 524810 995659
rect 559606 995607 559658 995659
rect 564598 995607 564650 995659
rect 625750 995607 625802 995659
rect 627094 995607 627146 995659
rect 143830 995533 143882 995585
rect 144118 995533 144170 995585
rect 191926 995533 191978 995585
rect 195190 995533 195242 995585
rect 295414 995533 295466 995585
rect 298294 995533 298346 995585
rect 383158 995533 383210 995585
rect 388822 995533 388874 995585
rect 472150 995533 472202 995585
rect 476374 995533 476426 995585
rect 510262 995533 510314 995585
rect 521398 995533 521450 995585
rect 523798 995533 523850 995585
rect 528982 995533 529034 995585
rect 560182 995533 560234 995585
rect 564502 995533 564554 995585
rect 625654 995533 625706 995585
rect 630166 995533 630218 995585
rect 82294 995459 82346 995511
rect 100726 995459 100778 995511
rect 293686 995459 293738 995511
rect 307606 995459 307658 995511
rect 380086 995459 380138 995511
rect 392374 995459 392426 995511
rect 466198 995459 466250 995511
rect 482710 995459 482762 995511
rect 523606 995459 523658 995511
rect 526102 995459 526154 995511
rect 185110 995385 185162 995437
rect 203638 995385 203690 995437
rect 379798 995385 379850 995437
rect 393718 995385 393770 995437
rect 471862 995385 471914 995437
rect 480982 995385 481034 995437
rect 519190 995385 519242 995437
rect 532246 995459 532298 995511
rect 625558 995459 625610 995511
rect 630934 995459 630986 995511
rect 86326 995311 86378 995363
rect 99766 995311 99818 995363
rect 521302 995311 521354 995363
rect 537382 995311 537434 995363
rect 132118 995237 132170 995289
rect 146806 995237 146858 995289
rect 184150 995237 184202 995289
rect 195766 995237 195818 995289
rect 519094 995237 519146 995289
rect 530566 995237 530618 995289
rect 632374 995237 632426 995289
rect 182998 995163 183050 995215
rect 196822 995163 196874 995215
rect 469462 995163 469514 995215
rect 485974 995163 486026 995215
rect 501814 995163 501866 995215
rect 528214 995163 528266 995215
rect 558934 995163 558986 995215
rect 649366 995163 649418 995215
rect 69142 995089 69194 995141
rect 298390 995089 298442 995141
rect 519958 995089 520010 995141
rect 649750 995089 649802 995141
rect 222934 995015 222986 995067
rect 649654 995015 649706 995067
rect 237430 994941 237482 994993
rect 250486 994941 250538 994993
rect 289270 994793 289322 994845
rect 296662 994793 296714 994845
rect 239446 994053 239498 994105
rect 279286 994053 279338 994105
rect 234934 993905 234986 993957
rect 250390 993905 250442 993957
rect 570742 993905 570794 993957
rect 635254 993905 635306 993957
rect 180502 993831 180554 993883
rect 198646 993831 198698 993883
rect 238678 993831 238730 993883
rect 259030 993831 259082 993883
rect 563254 993831 563306 993883
rect 641014 993831 641066 993883
rect 77686 993757 77738 993809
rect 95062 993757 95114 993809
rect 129334 993757 129386 993809
rect 149590 993757 149642 993809
rect 181366 993757 181418 993809
rect 209782 993757 209834 993809
rect 231478 993757 231530 993809
rect 260086 993757 260138 993809
rect 282838 993757 282890 993809
rect 309910 993757 309962 993809
rect 567382 993757 567434 993809
rect 634870 993757 634922 993809
rect 80182 993683 80234 993735
rect 105334 993683 105386 993735
rect 131830 993683 131882 993735
rect 156598 993683 156650 993735
rect 179830 993683 179882 993735
rect 208726 993683 208778 993735
rect 232534 993683 232586 993735
rect 261046 993683 261098 993735
rect 284374 993683 284426 993735
rect 312790 993683 312842 993735
rect 372502 993683 372554 993735
rect 393046 993683 393098 993735
rect 573046 993683 573098 993735
rect 637366 993683 637418 993735
rect 77302 993609 77354 993661
rect 105910 993609 105962 993661
rect 128470 993609 128522 993661
rect 157270 993609 157322 993661
rect 185398 993609 185450 993661
rect 236758 993609 236810 993661
rect 239446 993609 239498 993661
rect 250486 993609 250538 993661
rect 289270 993609 289322 993661
rect 365782 993609 365834 993661
rect 398806 993609 398858 993661
rect 443542 993609 443594 993661
rect 487798 993609 487850 993661
rect 521398 993609 521450 993661
rect 538966 993609 539018 993661
rect 61846 993535 61898 993587
rect 82582 993535 82634 993587
rect 133942 993535 133994 993587
rect 143830 993535 143882 993587
rect 237430 993535 237482 993587
rect 251350 993535 251402 993587
rect 279286 993535 279338 993587
rect 288118 993535 288170 993587
rect 390166 993535 390218 993587
rect 403126 993535 403178 993587
rect 331222 992573 331274 992625
rect 332566 992573 332618 992625
rect 73366 992055 73418 992107
rect 110134 992055 110186 992107
rect 627670 992055 627722 992107
rect 650038 992055 650090 992107
rect 290902 991759 290954 991811
rect 298966 991759 299018 991811
rect 105814 990501 105866 990553
rect 109558 990501 109610 990553
rect 640534 989909 640586 989961
rect 649846 989909 649898 989961
rect 569878 989539 569930 989591
rect 592438 989539 592490 989591
rect 569974 989465 570026 989517
rect 608758 989465 608810 989517
rect 371638 989391 371690 989443
rect 397846 989391 397898 989443
rect 437782 989391 437834 989443
rect 462742 989391 462794 989443
rect 515638 989391 515690 989443
rect 527638 989391 527690 989443
rect 533686 989391 533738 989443
rect 576310 989391 576362 989443
rect 154486 989317 154538 989369
rect 161686 989317 161738 989369
rect 203158 989317 203210 989369
rect 213334 989317 213386 989369
rect 270742 989317 270794 989369
rect 284278 989317 284330 989369
rect 319606 989317 319658 989369
rect 348502 989317 348554 989369
rect 371542 989317 371594 989369
rect 414070 989317 414122 989369
rect 437878 989317 437930 989369
rect 478966 989317 479018 989369
rect 515542 989317 515594 989369
rect 543766 989317 543818 989369
rect 569782 989317 569834 989369
rect 624982 989317 625034 989369
rect 643318 989317 643370 989369
rect 650134 989317 650186 989369
rect 89590 989243 89642 989295
rect 109366 989243 109418 989295
rect 138262 989243 138314 989295
rect 161494 989243 161546 989295
rect 216022 989243 216074 989295
rect 235606 989243 235658 989295
rect 267958 989243 268010 989295
rect 300502 989243 300554 989295
rect 319702 989243 319754 989295
rect 365398 989243 365450 989295
rect 371734 989243 371786 989295
rect 430294 989243 430346 989295
rect 437974 989243 438026 989295
rect 495190 989243 495242 989295
rect 515734 989243 515786 989295
rect 560086 989243 560138 989295
rect 567286 989243 567338 989295
rect 658102 989243 658154 989295
rect 47638 988281 47690 988333
rect 122038 988281 122090 988333
rect 44758 988207 44810 988259
rect 186934 988207 186986 988259
rect 44854 988133 44906 988185
rect 251830 988133 251882 988185
rect 44950 988059 45002 988111
rect 316726 988059 316778 988111
rect 45046 987985 45098 988037
rect 381622 987985 381674 988037
rect 45142 987911 45194 987963
rect 446518 987911 446570 987963
rect 43126 987837 43178 987889
rect 511414 987837 511466 987889
rect 65110 986727 65162 986779
rect 93526 986727 93578 986779
rect 47542 986653 47594 986705
rect 109174 986653 109226 986705
rect 47734 986579 47786 986631
rect 107926 986579 107978 986631
rect 47446 986505 47498 986557
rect 107542 986505 107594 986557
rect 63286 986431 63338 986483
rect 145366 986431 145418 986483
rect 564502 986431 564554 986483
rect 658006 986431 658058 986483
rect 65206 986357 65258 986409
rect 197206 986357 197258 986409
rect 564598 986357 564650 986409
rect 660886 986357 660938 986409
rect 64918 986135 64970 986187
rect 69046 986135 69098 986187
rect 632374 983693 632426 983745
rect 674518 983693 674570 983745
rect 633046 983619 633098 983671
rect 674134 983619 674186 983671
rect 64822 983545 64874 983597
rect 237430 983545 237482 983597
rect 528214 983545 528266 983597
rect 649558 983545 649610 983597
rect 65014 983471 65066 983523
rect 290806 983471 290858 983523
rect 417526 983471 417578 983523
rect 649462 983471 649514 983523
rect 50518 973481 50570 973533
rect 59446 973481 59498 973533
rect 42166 967265 42218 967317
rect 43126 967265 43178 967317
rect 649654 964749 649706 964801
rect 653782 964749 653834 964801
rect 42166 960975 42218 961027
rect 42454 960975 42506 961027
rect 46102 959051 46154 959103
rect 59542 959051 59594 959103
rect 675190 956979 675242 957031
rect 675478 956979 675530 957031
rect 42070 955203 42122 955255
rect 42838 955203 42890 955255
rect 669526 954685 669578 954737
rect 675382 954685 675434 954737
rect 41782 954611 41834 954663
rect 41782 954389 41834 954441
rect 674134 953945 674186 953997
rect 675478 953945 675530 953997
rect 674038 952021 674090 952073
rect 675478 952021 675530 952073
rect 42550 944621 42602 944673
rect 59542 944621 59594 944673
rect 42550 944177 42602 944229
rect 51862 944177 51914 944229
rect 42550 944029 42602 944081
rect 46102 944029 46154 944081
rect 42550 942993 42602 943045
rect 47542 942993 47594 943045
rect 42550 942845 42602 942897
rect 47734 942845 47786 942897
rect 40342 942327 40394 942379
rect 42550 942327 42602 942379
rect 658102 939515 658154 939567
rect 674422 939515 674474 939567
rect 655318 939367 655370 939419
rect 674518 939367 674570 939419
rect 655222 939219 655274 939271
rect 676822 939219 676874 939271
rect 655126 939071 655178 939123
rect 676918 939071 676970 939123
rect 674134 938923 674186 938975
rect 676918 938923 676970 938975
rect 660886 937961 660938 938013
rect 674422 937961 674474 938013
rect 658006 936259 658058 936311
rect 676822 936259 676874 936311
rect 42550 932115 42602 932167
rect 53206 932115 53258 932167
rect 51862 930487 51914 930539
rect 59542 930487 59594 930539
rect 654454 927453 654506 927505
rect 666742 927453 666794 927505
rect 649654 927379 649706 927431
rect 677014 927379 677066 927431
rect 53398 915835 53450 915887
rect 59542 915835 59594 915887
rect 653974 915835 654026 915887
rect 660982 915835 661034 915887
rect 650230 907103 650282 907155
rect 653782 907103 653834 907155
rect 654454 904365 654506 904417
rect 663958 904365 664010 904417
rect 50326 901479 50378 901531
rect 59542 901479 59594 901531
rect 53494 887123 53546 887175
rect 59542 887123 59594 887175
rect 653974 881277 654026 881329
rect 660886 881277 660938 881329
rect 47542 872619 47594 872671
rect 59542 872619 59594 872671
rect 674614 872619 674666 872671
rect 675382 872619 675434 872671
rect 673366 872101 673418 872153
rect 675478 872101 675530 872153
rect 674230 871657 674282 871709
rect 675094 871657 675146 871709
rect 675382 871657 675434 871709
rect 674902 871435 674954 871487
rect 675190 871435 675242 871487
rect 675382 871435 675434 871487
rect 654454 869807 654506 869859
rect 663766 869807 663818 869859
rect 673270 869141 673322 869193
rect 675478 869141 675530 869193
rect 674326 868327 674378 868379
rect 675382 868327 675434 868379
rect 673174 867809 673226 867861
rect 675382 867809 675434 867861
rect 675094 866477 675146 866529
rect 675382 866477 675434 866529
rect 666646 865293 666698 865345
rect 675382 865293 675434 865345
rect 674518 862925 674570 862977
rect 675382 862925 675434 862977
rect 47446 858263 47498 858315
rect 58582 858263 58634 858315
rect 654166 858263 654218 858315
rect 661078 858263 661130 858315
rect 675094 855747 675146 855799
rect 675478 855747 675530 855799
rect 674902 855599 674954 855651
rect 675574 855599 675626 855651
rect 53302 843833 53354 843885
rect 59542 843833 59594 843885
rect 653974 835175 654026 835227
rect 666838 835175 666890 835227
rect 47734 829477 47786 829529
rect 59542 829477 59594 829529
rect 653974 823705 654026 823757
rect 669910 823705 669962 823757
rect 42550 819265 42602 819317
rect 53494 819265 53546 819317
rect 42838 818525 42890 818577
rect 47542 818525 47594 818577
rect 42550 818229 42602 818281
rect 50326 818229 50378 818281
rect 50422 815047 50474 815099
rect 59542 815047 59594 815099
rect 654454 812161 654506 812213
rect 664054 812161 664106 812213
rect 42550 807425 42602 807477
rect 42838 807425 42890 807477
rect 43126 802541 43178 802593
rect 43414 802541 43466 802593
rect 42070 802393 42122 802445
rect 43126 802393 43178 802445
rect 41974 802023 42026 802075
rect 42454 802023 42506 802075
rect 43318 800617 43370 800669
rect 45142 800617 45194 800669
rect 50326 800617 50378 800669
rect 59542 800617 59594 800669
rect 41878 800173 41930 800225
rect 41878 799951 41930 800003
rect 42838 798323 42890 798375
rect 42934 798323 42986 798375
rect 42166 798101 42218 798153
rect 42742 798027 42794 798079
rect 42070 797287 42122 797339
rect 43318 797287 43370 797339
rect 42166 796251 42218 796303
rect 42742 796251 42794 796303
rect 42166 794993 42218 795045
rect 43030 794993 43082 795045
rect 42166 793143 42218 793195
rect 43126 793143 43178 793195
rect 42166 790627 42218 790679
rect 42742 790627 42794 790679
rect 674710 790553 674762 790605
rect 675478 790553 675530 790605
rect 42166 789887 42218 789939
rect 42838 789887 42890 789939
rect 42166 789443 42218 789495
rect 43414 789443 43466 789495
rect 674998 789221 675050 789273
rect 675574 789221 675626 789273
rect 674230 789147 674282 789199
rect 675094 789147 675146 789199
rect 42166 788777 42218 788829
rect 42454 788777 42506 788829
rect 42166 787001 42218 787053
rect 42934 787001 42986 787053
rect 42166 786409 42218 786461
rect 42742 786409 42794 786461
rect 47542 786261 47594 786313
rect 59542 786261 59594 786313
rect 654070 786261 654122 786313
rect 669718 786261 669770 786313
rect 42070 785595 42122 785647
rect 42838 785595 42890 785647
rect 672310 783449 672362 783501
rect 675382 783449 675434 783501
rect 672886 783079 672938 783131
rect 675094 783079 675146 783131
rect 675478 783079 675530 783131
rect 673462 782931 673514 782983
rect 675382 782931 675434 782983
rect 672502 782487 672554 782539
rect 674998 782487 675050 782539
rect 675478 782487 675530 782539
rect 663862 780489 663914 780541
rect 675094 780489 675146 780541
rect 673078 779749 673130 779801
rect 675382 779749 675434 779801
rect 672214 779305 672266 779357
rect 675478 779305 675530 779357
rect 672982 778565 673034 778617
rect 675382 778565 675434 778617
rect 672694 777603 672746 777655
rect 675478 777603 675530 777655
rect 675094 777011 675146 777063
rect 675382 777011 675434 777063
rect 42742 775901 42794 775953
rect 47734 775901 47786 775953
rect 42742 775309 42794 775361
rect 50422 775309 50474 775361
rect 42742 774791 42794 774843
rect 53302 774791 53354 774843
rect 654070 774717 654122 774769
rect 672406 774717 672458 774769
rect 53494 771831 53546 771883
rect 59542 771831 59594 771883
rect 653974 763247 654026 763299
rect 661174 763247 661226 763299
rect 660982 762877 661034 762929
rect 674422 762877 674474 762929
rect 666742 762285 666794 762337
rect 674422 762285 674474 762337
rect 663958 761989 664010 762041
rect 674614 761989 674666 762041
rect 42838 758585 42890 758637
rect 43030 758585 43082 758637
rect 43030 757623 43082 757675
rect 45046 757623 45098 757675
rect 53686 757475 53738 757527
rect 59542 757475 59594 757527
rect 41590 757327 41642 757379
rect 43510 757327 43562 757379
rect 41686 757253 41738 757305
rect 43414 757253 43466 757305
rect 41878 756957 41930 757009
rect 42070 756957 42122 757009
rect 43318 756957 43370 757009
rect 41878 756735 41930 756787
rect 42838 756661 42890 756713
rect 43222 756661 43274 756713
rect 43030 754219 43082 754271
rect 42166 754071 42218 754123
rect 43030 754071 43082 754123
rect 43222 754071 43274 754123
rect 42070 753035 42122 753087
rect 43126 753035 43178 753087
rect 43126 751777 43178 751829
rect 42934 751703 42986 751755
rect 43414 751629 43466 751681
rect 43702 751629 43754 751681
rect 42070 751111 42122 751163
rect 42934 751111 42986 751163
rect 42166 750371 42218 750423
rect 43030 750371 43082 750423
rect 43030 750223 43082 750275
rect 43510 750223 43562 750275
rect 649750 748817 649802 748869
rect 677014 748817 677066 748869
rect 42166 747263 42218 747315
rect 43126 747263 43178 747315
rect 43030 746967 43082 747019
rect 42166 746893 42218 746945
rect 672886 745931 672938 745983
rect 675094 745931 675146 745983
rect 42166 745635 42218 745687
rect 42934 745635 42986 745687
rect 42454 745487 42506 745539
rect 42934 745487 42986 745539
rect 42166 743785 42218 743837
rect 42934 743785 42986 743837
rect 42070 743193 42122 743245
rect 43126 743193 43178 743245
rect 53590 743045 53642 743097
rect 59542 743045 59594 743097
rect 42166 742601 42218 742653
rect 43030 742601 43082 742653
rect 653974 740159 654026 740211
rect 663958 740159 664010 740211
rect 672502 740159 672554 740211
rect 674710 740159 674762 740211
rect 673174 738087 673226 738139
rect 675094 738087 675146 738139
rect 675478 738087 675530 738139
rect 673366 737865 673418 737917
rect 675382 737865 675434 737917
rect 674710 737643 674762 737695
rect 675382 737643 675434 737695
rect 660982 737273 661034 737325
rect 675094 737273 675146 737325
rect 674614 735423 674666 735475
rect 675478 735423 675530 735475
rect 673270 734757 673322 734809
rect 675382 734757 675434 734809
rect 672790 734387 672842 734439
rect 675382 734387 675434 734439
rect 672886 733573 672938 733625
rect 675478 733573 675530 733625
rect 42838 732685 42890 732737
rect 53494 732685 53546 732737
rect 672598 732315 672650 732367
rect 675478 732315 675530 732367
rect 42838 732093 42890 732145
rect 53686 732093 53738 732145
rect 675094 732019 675146 732071
rect 675382 732019 675434 732071
rect 42838 731797 42890 731849
rect 47542 731797 47594 731849
rect 674614 731501 674666 731553
rect 674806 731501 674858 731553
rect 674518 730465 674570 730517
rect 675478 730465 675530 730517
rect 47542 728615 47594 728667
rect 59542 728615 59594 728667
rect 674038 728615 674090 728667
rect 675478 728615 675530 728667
rect 663766 718033 663818 718085
rect 674614 718033 674666 718085
rect 660886 717589 660938 717641
rect 674614 717589 674666 717641
rect 43126 717219 43178 717271
rect 43798 717219 43850 717271
rect 654262 717145 654314 717197
rect 666934 717145 666986 717197
rect 43126 717071 43178 717123
rect 44950 717071 45002 717123
rect 661078 716997 661130 717049
rect 674614 716997 674666 717049
rect 674614 715665 674666 715717
rect 674806 715665 674858 715717
rect 50422 714259 50474 714311
rect 59542 714259 59594 714311
rect 41494 714185 41546 714237
rect 43510 714185 43562 714237
rect 41590 714111 41642 714163
rect 43606 714111 43658 714163
rect 41686 714037 41738 714089
rect 43414 714037 43466 714089
rect 41878 713815 41930 713867
rect 41974 713815 42026 713867
rect 43222 713815 43274 713867
rect 41878 713519 41930 713571
rect 42070 711669 42122 711721
rect 43318 711669 43370 711721
rect 43222 711595 43274 711647
rect 43126 711373 43178 711425
rect 43414 711595 43466 711647
rect 43318 711373 43370 711425
rect 674326 711299 674378 711351
rect 674518 711299 674570 711351
rect 42166 710855 42218 710907
rect 43414 710855 43466 710907
rect 42166 709893 42218 709945
rect 43126 709893 43178 709945
rect 672310 709893 672362 709945
rect 674614 709893 674666 709945
rect 674422 709301 674474 709353
rect 674614 709301 674666 709353
rect 672694 709153 672746 709205
rect 674422 709153 674474 709205
rect 672214 708635 672266 708687
rect 674422 708635 674474 708687
rect 672982 707007 673034 707059
rect 674422 707007 674474 707059
rect 42166 706711 42218 706763
rect 43798 706711 43850 706763
rect 43222 706563 43274 706615
rect 43222 706341 43274 706393
rect 674710 705601 674762 705653
rect 674998 705601 675050 705653
rect 42166 704269 42218 704321
rect 42742 704269 42794 704321
rect 42742 704121 42794 704173
rect 43606 704121 43658 704173
rect 42070 703677 42122 703729
rect 43030 703677 43082 703729
rect 42166 702863 42218 702915
rect 43126 702863 43178 702915
rect 43126 702715 43178 702767
rect 43510 702715 43562 702767
rect 649846 702715 649898 702767
rect 677014 702715 677066 702767
rect 42166 702271 42218 702323
rect 42742 702271 42794 702323
rect 42070 700421 42122 700473
rect 43126 700421 43178 700473
rect 42166 700051 42218 700103
rect 42454 700051 42506 700103
rect 42454 699829 42506 699881
rect 59542 699829 59594 699881
rect 672694 699829 672746 699881
rect 673174 699829 673226 699881
rect 42166 699163 42218 699215
rect 43030 699163 43082 699215
rect 654454 694057 654506 694109
rect 669814 694057 669866 694109
rect 672694 692947 672746 692999
rect 675478 692947 675530 692999
rect 672310 692873 672362 692925
rect 675382 692873 675434 692925
rect 674614 692651 674666 692703
rect 675382 692651 675434 692703
rect 674806 690653 674858 690705
rect 675478 690653 675530 690705
rect 673078 689765 673130 689817
rect 675382 689765 675434 689817
rect 42838 689469 42890 689521
rect 50422 689469 50474 689521
rect 672982 689321 673034 689373
rect 675382 689321 675434 689373
rect 42454 688581 42506 688633
rect 47542 688581 47594 688633
rect 673174 688581 673226 688633
rect 675478 688581 675530 688633
rect 674710 687323 674762 687375
rect 675478 687323 675530 687375
rect 669622 686213 669674 686265
rect 675382 686213 675434 686265
rect 47542 685473 47594 685525
rect 59542 685473 59594 685525
rect 673942 685473 673994 685525
rect 675478 685473 675530 685525
rect 675478 683623 675530 683675
rect 675478 683327 675530 683379
rect 43414 673855 43466 673907
rect 44854 673855 44906 673907
rect 674710 673041 674762 673093
rect 674998 673041 675050 673093
rect 669910 672893 669962 672945
rect 674710 672893 674762 672945
rect 666838 672301 666890 672353
rect 674710 672301 674762 672353
rect 664054 671857 664106 671909
rect 674710 671857 674762 671909
rect 50422 671043 50474 671095
rect 59542 671043 59594 671095
rect 654454 671043 654506 671095
rect 661078 671043 661130 671095
rect 41686 670969 41738 671021
rect 42166 670969 42218 671021
rect 43702 670969 43754 671021
rect 674326 670969 674378 671021
rect 674710 670969 674762 671021
rect 41494 670821 41546 670873
rect 43414 670821 43466 670873
rect 43510 670747 43562 670799
rect 41974 670599 42026 670651
rect 42070 670599 42122 670651
rect 43126 670599 43178 670651
rect 41974 670303 42026 670355
rect 43030 670229 43082 670281
rect 43318 670229 43370 670281
rect 42454 670081 42506 670133
rect 43030 670081 43082 670133
rect 43030 668897 43082 668949
rect 42166 668527 42218 668579
rect 42838 668453 42890 668505
rect 43318 668453 43370 668505
rect 42166 667861 42218 667913
rect 43606 667861 43658 667913
rect 42166 666677 42218 666729
rect 42838 666677 42890 666729
rect 42838 666529 42890 666581
rect 43414 666529 43466 666581
rect 42166 665345 42218 665397
rect 43126 665345 43178 665397
rect 43126 665197 43178 665249
rect 43510 665197 43562 665249
rect 672790 665197 672842 665249
rect 673846 665197 673898 665249
rect 672598 664161 672650 664213
rect 674710 664161 674762 664213
rect 42742 663495 42794 663547
rect 42166 663347 42218 663399
rect 42742 663347 42794 663399
rect 43702 663347 43754 663399
rect 672886 662311 672938 662363
rect 673846 662311 673898 662363
rect 42070 661053 42122 661105
rect 42838 661053 42890 661105
rect 42166 659869 42218 659921
rect 42742 659869 42794 659921
rect 650038 659499 650090 659551
rect 674710 659499 674762 659551
rect 42166 659203 42218 659255
rect 43126 659203 43178 659255
rect 674422 658463 674474 658515
rect 675478 658463 675530 658515
rect 42070 657353 42122 657405
rect 42454 657353 42506 657405
rect 42934 656687 42986 656739
rect 59542 656687 59594 656739
rect 42166 656613 42218 656665
rect 43126 656613 43178 656665
rect 672694 653727 672746 653779
rect 674518 653727 674570 653779
rect 673270 648251 673322 648303
rect 675382 648251 675434 648303
rect 654262 648029 654314 648081
rect 664054 648029 664106 648081
rect 673750 648029 673802 648081
rect 675382 648029 675434 648081
rect 673366 647067 673418 647119
rect 674518 647067 674570 647119
rect 675382 647067 675434 647119
rect 675382 646401 675434 646453
rect 674806 646327 674858 646379
rect 674518 645883 674570 645935
rect 674998 645883 675050 645935
rect 42934 645217 42986 645269
rect 50422 645217 50474 645269
rect 42454 645069 42506 645121
rect 59542 645069 59594 645121
rect 672790 644551 672842 644603
rect 675478 644551 675530 644603
rect 672502 644033 672554 644085
rect 675478 644033 675530 644085
rect 672886 643367 672938 643419
rect 675382 643367 675434 643419
rect 672694 642257 672746 642309
rect 675478 642257 675530 642309
rect 673942 642109 673994 642161
rect 674134 642109 674186 642161
rect 666742 641073 666794 641125
rect 675478 641073 675530 641125
rect 674806 638187 674858 638239
rect 675478 638187 675530 638239
rect 43126 627975 43178 628027
rect 43702 627975 43754 628027
rect 43510 627901 43562 627953
rect 44758 627901 44810 627953
rect 43030 627827 43082 627879
rect 43414 627827 43466 627879
rect 50422 627827 50474 627879
rect 59542 627827 59594 627879
rect 674422 627827 674474 627879
rect 675094 627827 675146 627879
rect 41686 627679 41738 627731
rect 43030 627679 43082 627731
rect 672406 627679 672458 627731
rect 674422 627679 674474 627731
rect 42166 627605 42218 627657
rect 43126 627605 43178 627657
rect 41878 627383 41930 627435
rect 42070 627383 42122 627435
rect 43126 627383 43178 627435
rect 669718 627309 669770 627361
rect 674902 627309 674954 627361
rect 41878 627161 41930 627213
rect 661174 626569 661226 626621
rect 674422 626569 674474 626621
rect 670966 625459 671018 625511
rect 674422 625459 674474 625511
rect 42166 625311 42218 625363
rect 42934 625311 42986 625363
rect 42934 625163 42986 625215
rect 43222 625163 43274 625215
rect 42166 624645 42218 624697
rect 43510 624645 43562 624697
rect 42166 622203 42218 622255
rect 43414 622203 43466 622255
rect 654358 622203 654410 622255
rect 672598 622203 672650 622255
rect 671926 622129 671978 622181
rect 676918 622129 676970 622181
rect 672022 622055 672074 622107
rect 676822 622055 676874 622107
rect 42166 621611 42218 621663
rect 43126 621611 43178 621663
rect 42070 620871 42122 620923
rect 42934 620871 42986 620923
rect 42166 620353 42218 620405
rect 43030 620353 43082 620405
rect 672982 618429 673034 618481
rect 674422 618429 674474 618481
rect 672310 617837 672362 617889
rect 674422 617837 674474 617889
rect 673078 617541 673130 617593
rect 674710 617541 674762 617593
rect 42166 617171 42218 617223
rect 43702 617171 43754 617223
rect 42166 615987 42218 616039
rect 42454 615987 42506 616039
rect 42166 614137 42218 614189
rect 43126 614137 43178 614189
rect 42838 613471 42890 613523
rect 59542 613471 59594 613523
rect 649942 613471 649994 613523
rect 677110 613471 677162 613523
rect 654358 613397 654410 613449
rect 669526 613397 669578 613449
rect 673366 613397 673418 613449
rect 674998 613397 675050 613449
rect 675094 612139 675146 612191
rect 675478 612139 675530 612191
rect 671830 604073 671882 604125
rect 675478 604073 675530 604125
rect 673558 603259 673610 603311
rect 675382 603259 675434 603311
rect 42166 603111 42218 603163
rect 42838 603111 42890 603163
rect 672118 602815 672170 602867
rect 674998 602815 675050 602867
rect 675478 602815 675530 602867
rect 673366 602667 673418 602719
rect 675382 602667 675434 602719
rect 672310 602445 672362 602497
rect 675094 602445 675146 602497
rect 675382 602445 675434 602497
rect 42742 602223 42794 602275
rect 51862 602223 51914 602275
rect 663766 601927 663818 601979
rect 674422 601927 674474 601979
rect 42838 601853 42890 601905
rect 59542 601853 59594 601905
rect 673078 599781 673130 599833
rect 675382 599781 675434 599833
rect 672982 599263 673034 599315
rect 675382 599263 675434 599315
rect 654454 599041 654506 599093
rect 672406 599041 672458 599093
rect 673174 598375 673226 598427
rect 675478 598375 675530 598427
rect 672214 597117 672266 597169
rect 675478 597117 675530 597169
rect 674422 596821 674474 596873
rect 675382 596821 675434 596873
rect 654454 587497 654506 587549
rect 666838 587497 666890 587549
rect 671926 587497 671978 587549
rect 676822 587497 676874 587549
rect 51862 585943 51914 585995
rect 59542 585943 59594 585995
rect 43126 584685 43178 584737
rect 47638 584685 47690 584737
rect 41494 584463 41546 584515
rect 43222 584463 43274 584515
rect 41782 584241 41834 584293
rect 43414 584241 43466 584293
rect 41878 584167 41930 584219
rect 41878 583945 41930 583997
rect 42838 583797 42890 583849
rect 43318 583797 43370 583849
rect 663958 582021 664010 582073
rect 674422 582021 674474 582073
rect 655222 581947 655274 581999
rect 674614 581947 674666 581999
rect 666934 581577 666986 581629
rect 674614 581577 674666 581629
rect 43030 581503 43082 581555
rect 43318 581503 43370 581555
rect 42070 581429 42122 581481
rect 43126 581429 43178 581481
rect 670966 580837 671018 580889
rect 674422 580837 674474 580889
rect 671926 579135 671978 579187
rect 673846 579135 673898 579187
rect 42166 578987 42218 579039
rect 43030 578987 43082 579039
rect 43030 578839 43082 578891
rect 43414 578839 43466 578891
rect 42166 577137 42218 577189
rect 43126 577137 43178 577189
rect 654454 576027 654506 576079
rect 669910 576027 669962 576079
rect 672694 575953 672746 576005
rect 673846 575953 673898 576005
rect 672502 573585 672554 573637
rect 673846 573585 673898 573637
rect 42166 573437 42218 573489
rect 43030 573437 43082 573489
rect 672790 573067 672842 573119
rect 673846 573067 673898 573119
rect 42166 572623 42218 572675
rect 42934 572623 42986 572675
rect 672886 571587 672938 571639
rect 674422 571587 674474 571639
rect 42166 570995 42218 571047
rect 43126 570995 43178 571047
rect 42934 570255 42986 570307
rect 59542 570255 59594 570307
rect 42070 569663 42122 569715
rect 43126 569663 43178 569715
rect 650134 567369 650186 567421
rect 677014 567369 677066 567421
rect 654454 567295 654506 567347
rect 666646 567295 666698 567347
rect 672310 564409 672362 564461
rect 675094 564409 675146 564461
rect 672118 564335 672170 564387
rect 674998 564335 675050 564387
rect 674230 559525 674282 559577
rect 675382 559525 675434 559577
rect 43030 559303 43082 559355
rect 48886 559303 48938 559355
rect 42838 558859 42890 558911
rect 59542 558859 59594 558911
rect 674710 558045 674762 558097
rect 675382 558045 675434 558097
rect 674998 557823 675050 557875
rect 675382 557823 675434 557875
rect 673750 557601 673802 557653
rect 675478 557601 675530 557653
rect 675094 557083 675146 557135
rect 675478 557083 675530 557135
rect 660886 555825 660938 555877
rect 674998 555825 675050 555877
rect 674422 555233 674474 555285
rect 675478 555233 675530 555285
rect 673270 553753 673322 553805
rect 675478 553753 675530 553805
rect 672886 553161 672938 553213
rect 675382 553161 675434 553213
rect 654454 552939 654506 552991
rect 666646 552939 666698 552991
rect 674326 551903 674378 551955
rect 675478 551903 675530 551955
rect 674998 551607 675050 551659
rect 675382 551607 675434 551659
rect 674518 550053 674570 550105
rect 675478 550053 675530 550105
rect 674614 548203 674666 548255
rect 675478 548203 675530 548255
rect 48886 544651 48938 544703
rect 59542 544651 59594 544703
rect 41878 544207 41930 544259
rect 42934 544207 42986 544259
rect 43030 541469 43082 541521
rect 50518 541469 50570 541521
rect 654454 541469 654506 541521
rect 669718 541469 669770 541521
rect 41590 541247 41642 541299
rect 43606 541247 43658 541299
rect 42070 541173 42122 541225
rect 43222 541173 43274 541225
rect 42454 541099 42506 541151
rect 41974 540951 42026 541003
rect 42454 540951 42506 541003
rect 42166 540729 42218 540781
rect 42070 538879 42122 538931
rect 42934 538879 42986 538931
rect 42934 538731 42986 538783
rect 43222 538731 43274 538783
rect 42166 538139 42218 538191
rect 43030 538139 43082 538191
rect 669814 537177 669866 537229
rect 674806 537177 674858 537229
rect 661078 536585 661130 536637
rect 674806 536585 674858 536637
rect 671926 536141 671978 536193
rect 674806 536141 674858 536193
rect 42070 535771 42122 535823
rect 43126 535771 43178 535823
rect 655126 535771 655178 535823
rect 676822 535771 676874 535823
rect 43126 535623 43178 535675
rect 43606 535623 43658 535675
rect 42166 535031 42218 535083
rect 42934 535031 42986 535083
rect 42166 530887 42218 530939
rect 43030 530887 43082 530939
rect 42070 530221 42122 530273
rect 42454 530221 42506 530273
rect 43126 530147 43178 530199
rect 42454 530073 42506 530125
rect 43318 529999 43370 530051
rect 43702 529999 43754 530051
rect 43030 529925 43082 529977
rect 59542 529925 59594 529977
rect 654070 529925 654122 529977
rect 672502 529925 672554 529977
rect 671830 529851 671882 529903
rect 673654 529851 673706 529903
rect 43126 529481 43178 529533
rect 42934 529333 42986 529385
rect 43126 529333 43178 529385
rect 42454 529185 42506 529237
rect 42934 529185 42986 529237
rect 42838 528889 42890 528941
rect 672214 529037 672266 529089
rect 674806 529037 674858 529089
rect 672982 528445 673034 528497
rect 674806 528445 674858 528497
rect 42166 527631 42218 527683
rect 42934 527631 42986 527683
rect 42070 527039 42122 527091
rect 43126 527039 43178 527091
rect 42166 526447 42218 526499
rect 42838 526447 42890 526499
rect 677206 525929 677258 525981
rect 677398 525929 677450 525981
rect 650230 524301 650282 524353
rect 677014 524301 677066 524353
rect 41878 519787 41930 519839
rect 43030 519787 43082 519839
rect 654454 519269 654506 519321
rect 663862 519269 663914 519321
rect 53974 515495 54026 515547
rect 59542 515495 59594 515547
rect 43126 509723 43178 509775
rect 43318 509723 43370 509775
rect 654454 506911 654506 506963
rect 663862 506911 663914 506963
rect 47734 501139 47786 501191
rect 59542 501139 59594 501191
rect 654358 495367 654410 495419
rect 661174 495367 661226 495419
rect 664054 493221 664106 493273
rect 675094 493221 675146 493273
rect 655318 492481 655370 492533
rect 674902 492481 674954 492533
rect 672598 492407 672650 492459
rect 673846 492407 673898 492459
rect 44758 486709 44810 486761
rect 58582 486709 58634 486761
rect 654262 483823 654314 483875
rect 666934 483823 666986 483875
rect 672886 483749 672938 483801
rect 673846 483749 673898 483801
rect 650326 479457 650378 479509
rect 677014 479457 677066 479509
rect 44854 472353 44906 472405
rect 59542 472353 59594 472405
rect 654454 472205 654506 472257
rect 660982 472205 661034 472257
rect 43318 469393 43370 469445
rect 43606 469393 43658 469445
rect 50518 457923 50570 457975
rect 59542 457923 59594 457975
rect 654454 457923 654506 457975
rect 660982 457923 661034 457975
rect 43222 449265 43274 449317
rect 43606 449265 43658 449317
rect 654358 446379 654410 446431
rect 669814 446379 669866 446431
rect 53878 443567 53930 443619
rect 59542 443567 59594 443619
rect 654454 434909 654506 434961
rect 663958 434909 664010 434961
rect 42838 432245 42890 432297
rect 53974 432245 54026 432297
rect 42550 431949 42602 432001
rect 47734 431949 47786 432001
rect 47638 429137 47690 429189
rect 59542 429137 59594 429189
rect 654454 426177 654506 426229
rect 669622 426177 669674 426229
rect 42934 423365 42986 423417
rect 43702 423365 43754 423417
rect 40246 420479 40298 420531
rect 41782 420479 41834 420531
rect 42454 417593 42506 417645
rect 56182 417593 56234 417645
rect 39958 415891 40010 415943
rect 42454 415891 42506 415943
rect 40054 415373 40106 415425
rect 43126 415373 43178 415425
rect 40150 414707 40202 414759
rect 43030 414707 43082 414759
rect 45046 414707 45098 414759
rect 58390 414707 58442 414759
rect 41782 413375 41834 413427
rect 41782 413153 41834 413205
rect 653878 411821 653930 411873
rect 669526 411821 669578 411873
rect 42454 411377 42506 411429
rect 43222 411377 43274 411429
rect 42166 410933 42218 410985
rect 42550 410933 42602 410985
rect 42166 409675 42218 409727
rect 42550 409675 42602 409727
rect 42166 409453 42218 409505
rect 42358 409453 42410 409505
rect 42358 409305 42410 409357
rect 42934 409305 42986 409357
rect 43318 409083 43370 409135
rect 43030 409009 43082 409061
rect 42166 408195 42218 408247
rect 42358 408195 42410 408247
rect 42070 407455 42122 407507
rect 43126 407455 43178 407507
rect 42166 407011 42218 407063
rect 42934 407011 42986 407063
rect 42550 406049 42602 406101
rect 53398 406049 53450 406101
rect 672406 406049 672458 406101
rect 673846 406049 673898 406101
rect 666838 405457 666890 405509
rect 674710 405457 674762 405509
rect 669910 404421 669962 404473
rect 674710 404421 674762 404473
rect 42166 403163 42218 403215
rect 43030 403163 43082 403215
rect 43318 403163 43370 403215
rect 42934 403089 42986 403141
rect 673366 400425 673418 400477
rect 676918 400425 676970 400477
rect 56278 400351 56330 400403
rect 57622 400351 57674 400403
rect 654454 400351 654506 400403
rect 666838 400351 666890 400403
rect 673750 400351 673802 400403
rect 677206 400351 677258 400403
rect 650422 391767 650474 391819
rect 677110 391767 677162 391819
rect 42358 389325 42410 389377
rect 44854 389325 44906 389377
rect 654454 388807 654506 388859
rect 669622 388807 669674 388859
rect 42646 388733 42698 388785
rect 50518 388733 50570 388785
rect 42646 387993 42698 388045
rect 44758 387993 44810 388045
rect 675382 386365 675434 386417
rect 675382 386143 675434 386195
rect 44950 385921 45002 385973
rect 59254 385921 59306 385973
rect 675190 385403 675242 385455
rect 675478 385403 675530 385455
rect 675094 384811 675146 384863
rect 675382 384811 675434 384863
rect 674902 384663 674954 384715
rect 675094 384663 675146 384715
rect 674134 383109 674186 383161
rect 675286 383109 675338 383161
rect 674230 382443 674282 382495
rect 675478 382443 675530 382495
rect 654454 380075 654506 380127
rect 666742 380075 666794 380127
rect 674806 378151 674858 378203
rect 675382 378151 675434 378203
rect 674518 377559 674570 377611
rect 675382 377559 675434 377611
rect 674614 376893 674666 376945
rect 675478 376893 675530 376945
rect 42646 376523 42698 376575
rect 44758 376523 44810 376575
rect 673942 375709 673994 375761
rect 675478 375709 675530 375761
rect 40054 374303 40106 374355
rect 43126 374303 43178 374355
rect 40246 373637 40298 373689
rect 42838 373637 42890 373689
rect 39958 371565 40010 371617
rect 43318 371565 43370 371617
rect 47734 371565 47786 371617
rect 59542 371565 59594 371617
rect 42742 370455 42794 370507
rect 43222 370455 43274 370507
rect 42166 369937 42218 369989
rect 42358 369937 42410 369989
rect 42358 369789 42410 369841
rect 42838 369789 42890 369841
rect 42934 369493 42986 369545
rect 43126 369493 43178 369545
rect 43222 369197 43274 369249
rect 43414 369197 43466 369249
rect 42070 368087 42122 368139
rect 43126 368087 43178 368139
rect 43222 368087 43274 368139
rect 43222 367865 43274 367917
rect 42070 367347 42122 367399
rect 47446 367347 47498 367399
rect 42070 366237 42122 366289
rect 42934 366237 42986 366289
rect 654454 365793 654506 365845
rect 661078 365793 661130 365845
rect 42166 364979 42218 365031
rect 42838 364979 42890 365031
rect 42070 364239 42122 364291
rect 43030 364239 43082 364291
rect 42166 363795 42218 363847
rect 42358 363795 42410 363847
rect 42166 360095 42218 360147
rect 43126 360095 43178 360147
rect 669718 360021 669770 360073
rect 674422 360021 674474 360073
rect 666646 359725 666698 359777
rect 674710 359725 674762 359777
rect 672502 358985 672554 359037
rect 674422 358985 674474 359037
rect 47446 357135 47498 357187
rect 59542 357135 59594 357187
rect 42838 345887 42890 345939
rect 47638 345887 47690 345939
rect 650518 345591 650570 345643
rect 677014 345591 677066 345643
rect 42838 345369 42890 345421
rect 45046 345369 45098 345421
rect 42838 344777 42890 344829
rect 53878 344777 53930 344829
rect 50518 342779 50570 342831
rect 58390 342779 58442 342831
rect 654454 342705 654506 342757
rect 666646 342705 666698 342757
rect 675190 340929 675242 340981
rect 675478 340929 675530 340981
rect 674998 340781 675050 340833
rect 675190 340781 675242 340833
rect 674902 339523 674954 339575
rect 675382 339523 675434 339575
rect 674326 336563 674378 336615
rect 675382 336563 675434 336615
rect 673942 333529 673994 333581
rect 675382 333529 675434 333581
rect 674038 332715 674090 332767
rect 675382 332715 675434 332767
rect 654454 332271 654506 332323
rect 663766 332271 663818 332323
rect 43222 332197 43274 332249
rect 45046 332197 45098 332249
rect 674134 332197 674186 332249
rect 675478 332197 675530 332249
rect 674518 331753 674570 331805
rect 675382 331753 675434 331805
rect 40150 329533 40202 329585
rect 43030 329533 43082 329585
rect 40054 329311 40106 329363
rect 43126 329311 43178 329363
rect 53398 328349 53450 328401
rect 57814 328349 57866 328401
rect 41782 327017 41834 327069
rect 42262 326943 42314 326995
rect 42934 326943 42986 326995
rect 41782 326721 41834 326773
rect 42070 324871 42122 324923
rect 42838 324871 42890 324923
rect 42166 324131 42218 324183
rect 50326 324131 50378 324183
rect 42166 323095 42218 323147
rect 43126 323095 43178 323147
rect 42070 321763 42122 321815
rect 42550 321763 42602 321815
rect 42166 321023 42218 321075
rect 43030 321023 43082 321075
rect 42262 318729 42314 318781
rect 42838 318729 42890 318781
rect 42070 316879 42122 316931
rect 42934 316879 42986 316931
rect 661174 315029 661226 315081
rect 674422 315029 674474 315081
rect 663862 314733 663914 314785
rect 674710 314733 674762 314785
rect 666934 313993 666986 314045
rect 674422 313993 674474 314045
rect 44854 313919 44906 313971
rect 58006 313919 58058 313971
rect 42838 302671 42890 302723
rect 44950 302671 45002 302723
rect 650614 302597 650666 302649
rect 674422 302597 674474 302649
rect 42454 302301 42506 302353
rect 47734 302301 47786 302353
rect 42838 301635 42890 301687
rect 56278 301635 56330 301687
rect 44950 299563 45002 299615
rect 59446 299563 59498 299615
rect 674902 295419 674954 295471
rect 675094 295419 675146 295471
rect 674038 294753 674090 294805
rect 675094 294753 675146 294805
rect 654550 293791 654602 293843
rect 663766 293791 663818 293843
rect 674806 293495 674858 293547
rect 675094 293495 675146 293547
rect 674326 292903 674378 292955
rect 675382 292903 675434 292955
rect 674710 291719 674762 291771
rect 675094 291719 675146 291771
rect 674518 291645 674570 291697
rect 675190 291645 675242 291697
rect 42838 290091 42890 290143
rect 47638 290091 47690 290143
rect 673942 289425 673994 289477
rect 675382 289425 675434 289477
rect 674998 288537 675050 288589
rect 675478 288537 675530 288589
rect 674422 287723 674474 287775
rect 675382 287723 675434 287775
rect 674134 287205 674186 287257
rect 675478 287205 675530 287257
rect 674230 286761 674282 286813
rect 675382 286761 675434 286813
rect 39958 285355 40010 285407
rect 43318 285355 43370 285407
rect 40054 285281 40106 285333
rect 43126 285281 43178 285333
rect 40150 285207 40202 285259
rect 43030 285207 43082 285259
rect 40246 285133 40298 285185
rect 42934 285133 42986 285185
rect 45142 285133 45194 285185
rect 58102 285133 58154 285185
rect 654070 284763 654122 284815
rect 660886 284763 660938 284815
rect 42166 282913 42218 282965
rect 42454 282913 42506 282965
rect 42166 281729 42218 281781
rect 42358 281729 42410 281781
rect 42166 281063 42218 281115
rect 53590 281063 53642 281115
rect 42166 279879 42218 279931
rect 42934 279879 42986 279931
rect 42934 279731 42986 279783
rect 43318 279731 43370 279783
rect 64822 278547 64874 278599
rect 67222 278547 67274 278599
rect 268150 278547 268202 278599
rect 293782 278547 293834 278599
rect 299542 278547 299594 278599
rect 330166 278547 330218 278599
rect 332758 278547 332810 278599
rect 348790 278547 348842 278599
rect 350326 278547 350378 278599
rect 380662 278547 380714 278599
rect 255190 278473 255242 278525
rect 287254 278473 287306 278525
rect 233782 278399 233834 278451
rect 267766 278399 267818 278451
rect 267862 278399 267914 278451
rect 268150 278399 268202 278451
rect 293782 278399 293834 278451
rect 299734 278399 299786 278451
rect 293206 278325 293258 278377
rect 299542 278325 299594 278377
rect 335542 278473 335594 278525
rect 380854 278547 380906 278599
rect 381238 278547 381290 278599
rect 390262 278547 390314 278599
rect 393814 278547 393866 278599
rect 300406 278399 300458 278451
rect 383062 278473 383114 278525
rect 440662 278473 440714 278525
rect 489622 278473 489674 278525
rect 495382 278473 495434 278525
rect 501334 278473 501386 278525
rect 625078 278473 625130 278525
rect 631030 278473 631082 278525
rect 300310 278325 300362 278377
rect 380278 278325 380330 278377
rect 380662 278325 380714 278377
rect 381910 278325 381962 278377
rect 397462 278399 397514 278451
rect 417430 278399 417482 278451
rect 525526 278399 525578 278451
rect 551254 278399 551306 278451
rect 610486 278399 610538 278451
rect 610774 278399 610826 278451
rect 389014 278325 389066 278377
rect 290806 278251 290858 278303
rect 364150 278251 364202 278303
rect 365782 278251 365834 278303
rect 368854 278251 368906 278303
rect 378262 278251 378314 278303
rect 387766 278251 387818 278303
rect 396694 278251 396746 278303
rect 440662 278251 440714 278303
rect 440758 278251 440810 278303
rect 490198 278251 490250 278303
rect 294742 278177 294794 278229
rect 299542 278177 299594 278229
rect 299830 278177 299882 278229
rect 396214 278177 396266 278229
rect 240982 278103 241034 278155
rect 266038 278029 266090 278081
rect 299926 278103 299978 278155
rect 331318 278103 331370 278155
rect 352918 278103 352970 278155
rect 299830 278029 299882 278081
rect 300406 278029 300458 278081
rect 334390 278029 334442 278081
rect 353494 278029 353546 278081
rect 369622 278103 369674 278155
rect 380182 278103 380234 278155
rect 380662 278103 380714 278155
rect 390166 278103 390218 278155
rect 390262 278103 390314 278155
rect 636502 278103 636554 278155
rect 223126 277955 223178 278007
rect 299494 277955 299546 278007
rect 299638 277955 299690 278007
rect 300310 277955 300362 278007
rect 329110 277955 329162 278007
rect 355510 277955 355562 278007
rect 415318 278029 415370 278081
rect 64918 277881 64970 277933
rect 184342 277881 184394 277933
rect 291478 277881 291530 277933
rect 356950 277881 357002 277933
rect 422326 277955 422378 278007
rect 436630 277881 436682 277933
rect 42166 277807 42218 277859
rect 43126 277807 43178 277859
rect 288406 277807 288458 277859
rect 342742 277807 342794 277859
rect 356854 277807 356906 277859
rect 450838 277807 450890 277859
rect 289942 277733 289994 277785
rect 357046 277733 357098 277785
rect 358774 277733 358826 277785
rect 465238 277733 465290 277785
rect 295798 277659 295850 277711
rect 403606 277659 403658 277711
rect 296470 277585 296522 277637
rect 410806 277585 410858 277637
rect 297526 277511 297578 277563
rect 417910 277511 417962 277563
rect 292054 277437 292106 277489
rect 375094 277437 375146 277489
rect 375190 277437 375242 277489
rect 385174 277437 385226 277489
rect 42070 277363 42122 277415
rect 43030 277363 43082 277415
rect 247894 277363 247946 277415
rect 332182 277363 332234 277415
rect 363766 277363 363818 277415
rect 378742 277363 378794 277415
rect 378838 277363 378890 277415
rect 486838 277363 486890 277415
rect 298198 277289 298250 277341
rect 425014 277289 425066 277341
rect 299062 277215 299114 277267
rect 432214 277215 432266 277267
rect 314710 277141 314762 277193
rect 328054 277141 328106 277193
rect 328150 277141 328202 277193
rect 460726 277141 460778 277193
rect 225238 277067 225290 277119
rect 273622 277067 273674 277119
rect 300214 277067 300266 277119
rect 439318 277067 439370 277119
rect 301270 276993 301322 277045
rect 338806 276993 338858 277045
rect 364822 276993 364874 277045
rect 378646 276993 378698 277045
rect 378742 276993 378794 277045
rect 504694 276993 504746 277045
rect 300790 276919 300842 276971
rect 446518 276919 446570 276971
rect 289270 276845 289322 276897
rect 350038 276845 350090 276897
rect 376630 276845 376682 276897
rect 378550 276845 378602 276897
rect 378646 276845 378698 276897
rect 515446 276845 515498 276897
rect 301846 276771 301898 276823
rect 453526 276771 453578 276823
rect 215734 276697 215786 276749
rect 314710 276697 314762 276749
rect 208534 276623 208586 276675
rect 327382 276697 327434 276749
rect 349174 276697 349226 276749
rect 366934 276697 366986 276749
rect 367030 276697 367082 276749
rect 518998 276697 519050 276749
rect 324982 276623 325034 276675
rect 365782 276623 365834 276675
rect 197878 276549 197930 276601
rect 325846 276549 325898 276601
rect 325942 276549 325994 276601
rect 328150 276549 328202 276601
rect 361558 276549 361610 276601
rect 378838 276623 378890 276675
rect 378934 276623 378986 276675
rect 114646 276475 114698 276527
rect 322102 276475 322154 276527
rect 230614 276401 230666 276453
rect 327190 276475 327242 276527
rect 351094 276475 351146 276527
rect 366934 276475 366986 276527
rect 379030 276549 379082 276601
rect 386998 276549 387050 276601
rect 390166 276623 390218 276675
rect 554710 276623 554762 276675
rect 611830 276549 611882 276601
rect 325462 276401 325514 276453
rect 372022 276401 372074 276453
rect 372118 276401 372170 276453
rect 378454 276401 378506 276453
rect 401206 276475 401258 276527
rect 642262 276475 642314 276527
rect 649558 276475 649610 276527
rect 379030 276401 379082 276453
rect 379606 276401 379658 276453
rect 398902 276401 398954 276453
rect 243766 276327 243818 276379
rect 434518 276327 434570 276379
rect 231958 276253 232010 276305
rect 338230 276253 338282 276305
rect 346486 276253 346538 276305
rect 365590 276253 365642 276305
rect 372214 276253 372266 276305
rect 382966 276253 383018 276305
rect 383062 276253 383114 276305
rect 232342 276179 232394 276231
rect 341782 276179 341834 276231
rect 348406 276179 348458 276231
rect 379894 276179 379946 276231
rect 379990 276179 380042 276231
rect 384982 276179 385034 276231
rect 385174 276253 385226 276305
rect 565462 276253 565514 276305
rect 572470 276179 572522 276231
rect 244726 276105 244778 276157
rect 441718 276105 441770 276157
rect 245398 276031 245450 276083
rect 448822 276031 448874 276083
rect 246358 275957 246410 276009
rect 455926 275957 455978 276009
rect 233494 275883 233546 275935
rect 348982 275883 349034 275935
rect 369526 275883 369578 275935
rect 384886 275883 384938 275935
rect 384982 275883 385034 275935
rect 579670 275883 579722 275935
rect 247414 275809 247466 275861
rect 463126 275809 463178 275861
rect 227446 275735 227498 275787
rect 298966 275735 299018 275787
rect 311542 275735 311594 275787
rect 532150 275735 532202 275787
rect 248086 275661 248138 275713
rect 470230 275661 470282 275713
rect 234070 275587 234122 275639
rect 356086 275587 356138 275639
rect 364246 275587 364298 275639
rect 378742 275587 378794 275639
rect 378838 275587 378890 275639
rect 601078 275587 601130 275639
rect 249142 275513 249194 275565
rect 477430 275513 477482 275565
rect 42262 275439 42314 275491
rect 42934 275439 42986 275491
rect 196726 275439 196778 275491
rect 270262 275439 270314 275491
rect 322582 275439 322634 275491
rect 564214 275439 564266 275491
rect 235030 275365 235082 275417
rect 363190 275365 363242 275417
rect 368566 275365 368618 275417
rect 372982 275365 373034 275417
rect 375574 275365 375626 275417
rect 378838 275365 378890 275417
rect 378934 275365 378986 275417
rect 379990 275365 380042 275417
rect 380950 275365 381002 275417
rect 235990 275291 236042 275343
rect 370294 275291 370346 275343
rect 372598 275291 372650 275343
rect 384598 275291 384650 275343
rect 384790 275365 384842 275417
rect 622486 275365 622538 275417
rect 398806 275291 398858 275343
rect 398902 275291 398954 275343
rect 633142 275291 633194 275343
rect 200182 275217 200234 275269
rect 270838 275217 270890 275269
rect 284950 275217 285002 275269
rect 314422 275217 314474 275269
rect 316630 275217 316682 275269
rect 571318 275217 571370 275269
rect 228022 275143 228074 275195
rect 306070 275143 306122 275195
rect 316918 275143 316970 275195
rect 578518 275143 578570 275195
rect 236758 275069 236810 275121
rect 377494 275069 377546 275121
rect 377686 275069 377738 275121
rect 397462 275069 397514 275121
rect 398806 275069 398858 275121
rect 647542 275069 647594 275121
rect 229078 274995 229130 275047
rect 313270 274995 313322 275047
rect 317974 274995 318026 275047
rect 585622 274995 585674 275047
rect 242998 274921 243050 274973
rect 427414 274921 427466 274973
rect 258550 274847 258602 274899
rect 333142 274847 333194 274899
rect 368086 274847 368138 274899
rect 378646 274847 378698 274899
rect 378742 274847 378794 274899
rect 384790 274847 384842 274899
rect 384886 274847 384938 274899
rect 551062 274847 551114 274899
rect 242230 274773 242282 274825
rect 420214 274773 420266 274825
rect 241078 274699 241130 274751
rect 413206 274699 413258 274751
rect 223030 274625 223082 274677
rect 263350 274625 263402 274677
rect 269206 274625 269258 274677
rect 334486 274625 334538 274677
rect 370966 274625 371018 274677
rect 375190 274625 375242 274677
rect 375958 274625 376010 274677
rect 378358 274625 378410 274677
rect 378646 274625 378698 274677
rect 540406 274625 540458 274677
rect 240502 274551 240554 274603
rect 406006 274551 406058 274603
rect 239350 274477 239402 274529
rect 398614 274477 398666 274529
rect 238486 274403 238538 274455
rect 372790 274403 372842 274455
rect 372886 274403 372938 274455
rect 378646 274403 378698 274455
rect 379030 274403 379082 274455
rect 398902 274403 398954 274455
rect 237814 274329 237866 274381
rect 372598 274329 372650 274381
rect 372982 274329 373034 274381
rect 381622 274329 381674 274381
rect 382774 274329 382826 274381
rect 400054 274329 400106 274381
rect 408982 274329 409034 274381
rect 449302 274329 449354 274381
rect 226294 274255 226346 274307
rect 291862 274255 291914 274307
rect 297814 274255 297866 274307
rect 337942 274255 337994 274307
rect 358294 274255 358346 274307
rect 378646 274255 378698 274307
rect 378742 274255 378794 274307
rect 383542 274255 383594 274307
rect 385078 274255 385130 274307
rect 390550 274255 390602 274307
rect 184342 274181 184394 274233
rect 200086 274181 200138 274233
rect 207382 274181 207434 274233
rect 271318 274181 271370 274233
rect 271414 274181 271466 274233
rect 214582 274107 214634 274159
rect 272470 274107 272522 274159
rect 276406 274181 276458 274233
rect 335638 274181 335690 274233
rect 364342 274181 364394 274233
rect 511894 274255 511946 274307
rect 645718 274255 645770 274307
rect 649462 274255 649514 274307
rect 398902 274181 398954 274233
rect 408982 274181 409034 274233
rect 449302 274181 449354 274233
rect 469462 274181 469514 274233
rect 225430 274033 225482 274085
rect 284662 274033 284714 274085
rect 225238 273959 225290 274011
rect 281110 273959 281162 274011
rect 287062 274107 287114 274159
rect 337078 274107 337130 274159
rect 360502 274107 360554 274159
rect 479734 274107 479786 274159
rect 286678 274033 286730 274085
rect 328726 274033 328778 274085
rect 360022 274033 360074 274085
rect 476182 274033 476234 274085
rect 239446 273885 239498 273937
rect 275254 273885 275306 273937
rect 304918 273959 304970 274011
rect 338902 273959 338954 274011
rect 374326 273959 374378 274011
rect 352246 273885 352298 273937
rect 365878 273885 365930 273937
rect 370294 273885 370346 273937
rect 378550 273959 378602 274011
rect 378646 273959 378698 274011
rect 461974 273959 462026 274011
rect 469462 273959 469514 274011
rect 508342 273959 508394 274011
rect 375670 273885 375722 273937
rect 383446 273885 383498 273937
rect 383542 273885 383594 273937
rect 558262 273885 558314 273937
rect 232438 273811 232490 273863
rect 274678 273811 274730 273863
rect 308854 273811 308906 273863
rect 229750 273737 229802 273789
rect 320086 273737 320138 273789
rect 356182 273811 356234 273863
rect 444118 273811 444170 273863
rect 365110 273737 365162 273789
rect 365206 273737 365258 273789
rect 382390 273737 382442 273789
rect 382486 273737 382538 273789
rect 383158 273737 383210 273789
rect 383254 273737 383306 273789
rect 391702 273737 391754 273789
rect 403126 273737 403178 273789
rect 417334 273737 417386 273789
rect 231766 273663 231818 273715
rect 325462 273663 325514 273715
rect 354454 273663 354506 273715
rect 429814 273663 429866 273715
rect 262678 273589 262730 273641
rect 365782 273589 365834 273641
rect 365878 273589 365930 273641
rect 411958 273589 412010 273641
rect 67222 273515 67274 273567
rect 79030 273515 79082 273567
rect 153814 273515 153866 273567
rect 163126 273515 163178 273567
rect 165814 273515 165866 273567
rect 166966 273515 167018 273567
rect 170518 273515 170570 273567
rect 172726 273515 172778 273567
rect 174070 273515 174122 273567
rect 175510 273515 175562 273567
rect 177622 273515 177674 273567
rect 178390 273515 178442 273567
rect 180022 273515 180074 273567
rect 181366 273515 181418 273567
rect 184726 273515 184778 273567
rect 187030 273515 187082 273567
rect 198646 273515 198698 273567
rect 212374 273515 212426 273567
rect 257878 273515 257930 273567
rect 282454 273515 282506 273567
rect 315382 273515 315434 273567
rect 322582 273515 322634 273567
rect 322678 273515 322730 273567
rect 325270 273515 325322 273567
rect 325462 273515 325514 273567
rect 334582 273515 334634 273567
rect 340630 273515 340682 273567
rect 343510 273515 343562 273567
rect 344662 273515 344714 273567
rect 347734 273515 347786 273567
rect 356950 273515 357002 273567
rect 367894 273515 367946 273567
rect 374134 273515 374186 273567
rect 378070 273515 378122 273567
rect 378358 273515 378410 273567
rect 396214 273515 396266 273567
rect 397366 273515 397418 273567
rect 595126 273515 595178 273567
rect 91990 273441 92042 273493
rect 206038 273441 206090 273493
rect 224566 273441 224618 273493
rect 271510 273441 271562 273493
rect 271606 273441 271658 273493
rect 279478 273441 279530 273493
rect 281206 273441 281258 273493
rect 285814 273441 285866 273493
rect 285910 273441 285962 273493
rect 310870 273441 310922 273493
rect 314518 273441 314570 273493
rect 557014 273441 557066 273493
rect 146518 273367 146570 273419
rect 151126 273367 151178 273419
rect 161014 273367 161066 273419
rect 394582 273367 394634 273419
rect 144406 273293 144458 273345
rect 146806 273293 146858 273345
rect 157462 273293 157514 273345
rect 404086 273367 404138 273419
rect 158614 273219 158666 273271
rect 161206 273219 161258 273271
rect 163126 273219 163178 273271
rect 403990 273293 404042 273345
rect 394870 273219 394922 273271
rect 408214 273219 408266 273271
rect 128950 273145 129002 273197
rect 146518 273145 146570 273197
rect 95638 273071 95690 273123
rect 100726 273071 100778 273123
rect 132502 273071 132554 273123
rect 147862 273145 147914 273197
rect 147958 273145 148010 273197
rect 149686 273145 149738 273197
rect 151414 273145 151466 273197
rect 152566 273145 152618 273197
rect 152662 273145 152714 273197
rect 155350 273145 155402 273197
rect 156214 273145 156266 273197
rect 158326 273145 158378 273197
rect 159862 273145 159914 273197
rect 161110 273145 161162 273197
rect 162166 273145 162218 273197
rect 164086 273145 164138 273197
rect 164182 273145 164234 273197
rect 378454 273145 378506 273197
rect 146710 273071 146762 273123
rect 377974 273071 378026 273123
rect 143158 272997 143210 273049
rect 400630 273145 400682 273197
rect 130102 272923 130154 272975
rect 132406 272923 132458 272975
rect 133558 272923 133610 272975
rect 135286 272923 135338 272975
rect 139606 272923 139658 272975
rect 399670 273071 399722 273123
rect 378742 272997 378794 273049
rect 398614 272997 398666 273049
rect 65878 272849 65930 272901
rect 198646 272849 198698 272901
rect 198742 272849 198794 272901
rect 211606 272849 211658 272901
rect 220822 272849 220874 272901
rect 245494 272849 245546 272901
rect 267862 272849 267914 272901
rect 270358 272849 270410 272901
rect 270454 272849 270506 272901
rect 271414 272849 271466 272901
rect 271510 272849 271562 272901
rect 277558 272849 277610 272901
rect 278806 272849 278858 272901
rect 280054 272849 280106 272901
rect 280726 272849 280778 272901
rect 282358 272849 282410 272901
rect 282454 272849 282506 272901
rect 378262 272849 378314 272901
rect 101494 272775 101546 272827
rect 103606 272775 103658 272827
rect 105046 272775 105098 272827
rect 106486 272775 106538 272827
rect 115798 272775 115850 272827
rect 118006 272775 118058 272827
rect 119350 272775 119402 272827
rect 120886 272775 120938 272827
rect 122902 272775 122954 272827
rect 123766 272775 123818 272827
rect 124150 272775 124202 272827
rect 126550 272775 126602 272827
rect 127702 272775 127754 272827
rect 129526 272775 129578 272827
rect 131254 272775 131306 272827
rect 132310 272775 132362 272827
rect 137206 272775 137258 272827
rect 138166 272775 138218 272827
rect 142006 272775 142058 272827
rect 143926 272775 143978 272827
rect 146710 272775 146762 272827
rect 378646 272849 378698 272901
rect 398038 272923 398090 272975
rect 378934 272849 378986 272901
rect 380758 272849 380810 272901
rect 380854 272849 380906 272901
rect 643894 272849 643946 272901
rect 135958 272701 136010 272753
rect 146614 272701 146666 272753
rect 147862 272701 147914 272753
rect 378838 272775 378890 272827
rect 151126 272627 151178 272679
rect 387574 272701 387626 272753
rect 391414 272775 391466 272827
rect 412246 272775 412298 272827
rect 596182 272775 596234 272827
rect 598486 272775 598538 272827
rect 378742 272627 378794 272679
rect 380374 272627 380426 272679
rect 380758 272627 380810 272679
rect 381334 272627 381386 272679
rect 381622 272627 381674 272679
rect 386422 272627 386474 272679
rect 386518 272627 386570 272679
rect 387862 272627 387914 272679
rect 397270 272701 397322 272753
rect 398806 272627 398858 272679
rect 612982 272627 613034 272679
rect 125302 272553 125354 272605
rect 378358 272553 378410 272605
rect 378550 272553 378602 272605
rect 391894 272553 391946 272605
rect 394582 272553 394634 272605
rect 396886 272553 396938 272605
rect 397366 272553 397418 272605
rect 591574 272553 591626 272605
rect 121750 272479 121802 272531
rect 380278 272479 380330 272531
rect 380374 272479 380426 272531
rect 402358 272479 402410 272531
rect 118102 272405 118154 272457
rect 394198 272405 394250 272457
rect 394294 272405 394346 272457
rect 584374 272405 584426 272457
rect 84886 272331 84938 272383
rect 86326 272331 86378 272383
rect 111094 272331 111146 272383
rect 107446 272257 107498 272309
rect 378550 272257 378602 272309
rect 103894 272183 103946 272235
rect 390934 272257 390986 272309
rect 392470 272331 392522 272383
rect 587926 272331 587978 272383
rect 392566 272257 392618 272309
rect 393814 272257 393866 272309
rect 573718 272257 573770 272309
rect 378742 272183 378794 272235
rect 378934 272183 378986 272235
rect 379990 272183 380042 272235
rect 381430 272183 381482 272235
rect 381526 272183 381578 272235
rect 382486 272183 382538 272235
rect 382678 272183 382730 272235
rect 541558 272183 541610 272235
rect 67030 272109 67082 272161
rect 213238 272109 213290 272161
rect 221014 272109 221066 272161
rect 249046 272109 249098 272161
rect 258358 272109 258410 272161
rect 552310 272109 552362 272161
rect 89590 272035 89642 272087
rect 92086 272035 92138 272087
rect 145558 272035 145610 272087
rect 146710 272035 146762 272087
rect 150262 272035 150314 272087
rect 164182 272035 164234 272087
rect 164566 272035 164618 272087
rect 405910 272035 405962 272087
rect 99190 271961 99242 272013
rect 198742 271961 198794 272013
rect 198838 271961 198890 272013
rect 212182 271961 212234 272013
rect 224086 271961 224138 272013
rect 267958 271961 268010 272013
rect 268054 271961 268106 272013
rect 278998 271961 279050 272013
rect 285526 271961 285578 272013
rect 321526 271961 321578 272013
rect 321622 271961 321674 272013
rect 329782 271961 329834 272013
rect 336982 271961 337034 272013
rect 343030 271961 343082 272013
rect 347926 271961 347978 272013
rect 358486 271961 358538 272013
rect 365782 271961 365834 272013
rect 380182 271961 380234 272013
rect 380278 271961 380330 272013
rect 395254 271961 395306 272013
rect 396886 271961 396938 272013
rect 398710 271961 398762 272013
rect 398806 271961 398858 272013
rect 618838 271961 618890 272013
rect 172918 271887 172970 271939
rect 175606 271887 175658 271939
rect 176470 271887 176522 271939
rect 178486 271887 178538 271939
rect 171670 271739 171722 271791
rect 407542 271887 407594 271939
rect 409654 271887 409706 271939
rect 433462 271887 433514 271939
rect 633622 271887 633674 271939
rect 642262 271887 642314 271939
rect 100726 271591 100778 271643
rect 175318 271665 175370 271717
rect 394870 271813 394922 271865
rect 394966 271813 395018 271865
rect 406678 271813 406730 271865
rect 121174 271591 121226 271643
rect 156886 271591 156938 271643
rect 120982 271443 121034 271495
rect 177046 271443 177098 271495
rect 102646 271369 102698 271421
rect 156886 271369 156938 271421
rect 178870 271591 178922 271643
rect 409270 271739 409322 271791
rect 182422 271665 182474 271717
rect 403174 271665 403226 271717
rect 185974 271591 186026 271643
rect 403030 271591 403082 271643
rect 189526 271517 189578 271569
rect 403126 271517 403178 271569
rect 403318 271517 403370 271569
rect 195766 271443 195818 271495
rect 206614 271443 206666 271495
rect 209782 271443 209834 271495
rect 198838 271369 198890 271421
rect 113494 271295 113546 271347
rect 212086 271369 212138 271421
rect 223702 271443 223754 271495
rect 267862 271443 267914 271495
rect 267958 271443 268010 271495
rect 274006 271443 274058 271495
rect 275158 271443 275210 271495
rect 279670 271443 279722 271495
rect 283798 271443 283850 271495
rect 307318 271443 307370 271495
rect 313654 271443 313706 271495
rect 321622 271443 321674 271495
rect 216118 271369 216170 271421
rect 220342 271369 220394 271421
rect 241846 271369 241898 271421
rect 246646 271369 246698 271421
rect 116950 271221 117002 271273
rect 211894 271295 211946 271347
rect 213334 271295 213386 271347
rect 216694 271295 216746 271347
rect 219766 271295 219818 271347
rect 238294 271295 238346 271347
rect 199126 271221 199178 271273
rect 214966 271221 215018 271273
rect 253750 271369 253802 271421
rect 277270 271369 277322 271421
rect 282742 271369 282794 271421
rect 296662 271369 296714 271421
rect 312118 271369 312170 271421
rect 333334 271443 333386 271495
rect 333430 271443 333482 271495
rect 342646 271443 342698 271495
rect 345718 271443 345770 271495
rect 358390 271443 358442 271495
rect 358486 271443 358538 271495
rect 374422 271443 374474 271495
rect 374710 271443 374762 271495
rect 403222 271443 403274 271495
rect 459286 271517 459338 271569
rect 479446 271517 479498 271569
rect 499606 271517 499658 271569
rect 518326 271517 518378 271569
rect 593974 271443 594026 271495
rect 324118 271369 324170 271421
rect 325558 271369 325610 271421
rect 329974 271369 330026 271421
rect 341974 271369 342026 271421
rect 347446 271369 347498 271421
rect 372694 271369 372746 271421
rect 374038 271369 374090 271421
rect 590326 271369 590378 271421
rect 264502 271295 264554 271347
rect 278518 271295 278570 271347
rect 282934 271295 282986 271347
rect 300118 271295 300170 271347
rect 308182 271295 308234 271347
rect 319414 271295 319466 271347
rect 320374 271295 320426 271347
rect 325654 271295 325706 271347
rect 120502 271147 120554 271199
rect 211798 271147 211850 271199
rect 219286 271147 219338 271199
rect 234646 271147 234698 271199
rect 109846 271073 109898 271125
rect 201526 271073 201578 271125
rect 202582 271073 202634 271125
rect 215446 271073 215498 271125
rect 218902 271073 218954 271125
rect 231190 271073 231242 271125
rect 283414 271221 283466 271273
rect 303670 271221 303722 271273
rect 308470 271221 308522 271273
rect 339382 271295 339434 271347
rect 276406 271147 276458 271199
rect 284470 271147 284522 271199
rect 285910 271147 285962 271199
rect 319126 271147 319178 271199
rect 340918 271221 340970 271273
rect 345334 271295 345386 271347
rect 347254 271295 347306 271347
rect 346390 271221 346442 271273
rect 362038 271221 362090 271273
rect 268726 271073 268778 271125
rect 270454 271073 270506 271125
rect 292534 271073 292586 271125
rect 106294 270999 106346 271051
rect 191446 270999 191498 271051
rect 193078 270999 193130 271051
rect 269878 270999 269930 271051
rect 282166 270999 282218 271051
rect 293014 270999 293066 271051
rect 302518 270999 302570 271051
rect 315958 271073 316010 271125
rect 322006 271073 322058 271125
rect 322774 271073 322826 271125
rect 329494 271073 329546 271125
rect 329686 271073 329738 271125
rect 345238 271147 345290 271199
rect 354838 271147 354890 271199
rect 366166 271295 366218 271347
rect 370390 271295 370442 271347
rect 370486 271295 370538 271347
rect 403414 271295 403466 271347
rect 413206 271295 413258 271347
rect 559414 271295 559466 271347
rect 365110 271221 365162 271273
rect 381526 271221 381578 271273
rect 381910 271221 381962 271273
rect 409654 271221 409706 271273
rect 433462 271221 433514 271273
rect 459286 271221 459338 271273
rect 479446 271221 479498 271273
rect 499606 271221 499658 271273
rect 518326 271221 518378 271273
rect 543958 271221 544010 271273
rect 369142 271147 369194 271199
rect 369238 271147 369290 271199
rect 373654 271147 373706 271199
rect 374422 271147 374474 271199
rect 376246 271147 376298 271199
rect 376342 271147 376394 271199
rect 378070 271147 378122 271199
rect 378166 271147 378218 271199
rect 395062 271147 395114 271199
rect 395446 271147 395498 271199
rect 534454 271147 534506 271199
rect 333334 271073 333386 271125
rect 336694 271073 336746 271125
rect 191926 270925 191978 270977
rect 213814 270925 213866 270977
rect 218710 270925 218762 270977
rect 227638 270925 227690 270977
rect 257302 270925 257354 270977
rect 277462 270925 277514 270977
rect 281686 270925 281738 270977
rect 289462 270925 289514 270977
rect 294262 270925 294314 270977
rect 308182 270925 308234 270977
rect 320278 270999 320330 271051
rect 322102 270999 322154 271051
rect 393622 271073 393674 271125
rect 394486 271073 394538 271125
rect 580918 271073 580970 271125
rect 336886 270999 336938 271051
rect 383062 270999 383114 271051
rect 383158 270999 383210 271051
rect 510646 270999 510698 271051
rect 322678 270925 322730 270977
rect 322966 270925 323018 270977
rect 324886 270925 324938 270977
rect 326326 270925 326378 270977
rect 341494 270925 341546 270977
rect 344758 270925 344810 270977
rect 351286 270925 351338 270977
rect 363862 270925 363914 270977
rect 371542 270925 371594 270977
rect 373462 270925 373514 270977
rect 388630 270925 388682 270977
rect 388726 270925 388778 270977
rect 545206 270925 545258 270977
rect 168118 270851 168170 270903
rect 394966 270851 395018 270903
rect 395062 270851 395114 270903
rect 401302 270851 401354 270903
rect 403414 270851 403466 270903
rect 413206 270851 413258 270903
rect 177046 270777 177098 270829
rect 68182 270703 68234 270755
rect 69046 270703 69098 270755
rect 75382 270703 75434 270755
rect 77686 270703 77738 270755
rect 188374 270703 188426 270755
rect 190006 270703 190058 270755
rect 190774 270703 190826 270755
rect 192886 270703 192938 270755
rect 195478 270777 195530 270829
rect 214486 270777 214538 270829
rect 218230 270777 218282 270829
rect 223990 270777 224042 270829
rect 260950 270777 261002 270829
rect 277942 270777 277994 270829
rect 314806 270777 314858 270829
rect 319702 270777 319754 270829
rect 322006 270777 322058 270829
rect 340438 270777 340490 270829
rect 342742 270777 342794 270829
rect 359638 270777 359690 270829
rect 362038 270777 362090 270829
rect 365206 270777 365258 270829
rect 365302 270777 365354 270829
rect 367030 270777 367082 270829
rect 367126 270777 367178 270829
rect 369238 270777 369290 270829
rect 370678 270777 370730 270829
rect 373558 270777 373610 270829
rect 373654 270777 373706 270829
rect 376150 270777 376202 270829
rect 377590 270777 377642 270829
rect 378838 270777 378890 270829
rect 378934 270777 378986 270829
rect 386902 270777 386954 270829
rect 388054 270777 388106 270829
rect 395446 270777 395498 270829
rect 398902 270777 398954 270829
rect 404950 270777 405002 270829
rect 195766 270703 195818 270755
rect 206230 270703 206282 270755
rect 215542 270703 215594 270755
rect 217558 270703 217610 270755
rect 220438 270703 220490 270755
rect 250198 270703 250250 270755
rect 276790 270703 276842 270755
rect 317494 270703 317546 270755
rect 392086 270703 392138 270755
rect 394486 270703 394538 270755
rect 570166 270703 570218 270755
rect 230230 270629 230282 270681
rect 310294 270629 310346 270681
rect 310390 270629 310442 270681
rect 325654 270629 325706 270681
rect 328342 270629 328394 270681
rect 329686 270629 329738 270681
rect 329782 270629 329834 270681
rect 549910 270629 549962 270681
rect 231286 270555 231338 270607
rect 328534 270555 328586 270607
rect 328630 270555 328682 270607
rect 332278 270555 332330 270607
rect 336694 270555 336746 270607
rect 339862 270555 339914 270607
rect 348310 270555 348362 270607
rect 352726 270555 352778 270607
rect 358486 270555 358538 270607
rect 370678 270555 370730 270607
rect 370774 270555 370826 270607
rect 373462 270555 373514 270607
rect 373558 270555 373610 270607
rect 379126 270555 379178 270607
rect 379798 270555 379850 270607
rect 388726 270555 388778 270607
rect 388822 270555 388874 270607
rect 561814 270555 561866 270607
rect 623062 270555 623114 270607
rect 641494 270555 641546 270607
rect 203830 270481 203882 270533
rect 270934 270481 270986 270533
rect 307798 270481 307850 270533
rect 503542 270481 503594 270533
rect 544438 270481 544490 270533
rect 564406 270481 564458 270533
rect 244150 270407 244202 270459
rect 438070 270407 438122 270459
rect 440662 270407 440714 270459
rect 460726 270407 460778 270459
rect 469174 270407 469226 270459
rect 469654 270407 469706 270459
rect 232822 270333 232874 270385
rect 328342 270333 328394 270385
rect 328534 270333 328586 270385
rect 331126 270333 331178 270385
rect 338998 270333 339050 270385
rect 352438 270333 352490 270385
rect 355606 270333 355658 270385
rect 373846 270333 373898 270385
rect 375094 270333 375146 270385
rect 379030 270333 379082 270385
rect 379222 270333 379274 270385
rect 568918 270333 568970 270385
rect 245302 270259 245354 270311
rect 332566 270259 332618 270311
rect 339190 270259 339242 270311
rect 233974 270185 234026 270237
rect 338998 270185 339050 270237
rect 357622 270185 357674 270237
rect 366166 270185 366218 270237
rect 367510 270185 367562 270237
rect 378838 270185 378890 270237
rect 445270 270259 445322 270311
rect 469078 270259 469130 270311
rect 469558 270259 469610 270311
rect 379318 270185 379370 270237
rect 576118 270185 576170 270237
rect 245878 270111 245930 270163
rect 348310 270111 348362 270163
rect 352726 270111 352778 270163
rect 452374 270111 452426 270163
rect 469366 270111 469418 270163
rect 469558 270111 469610 270163
rect 234550 270037 234602 270089
rect 342742 270037 342794 270089
rect 363094 270037 363146 270089
rect 378934 270037 378986 270089
rect 379126 270037 379178 270089
rect 98038 269963 98090 270015
rect 100726 269963 100778 270015
rect 140758 269963 140810 270015
rect 141046 269963 141098 270015
rect 194326 269963 194378 270015
rect 314038 269963 314090 270015
rect 314422 269963 314474 270015
rect 325462 269963 325514 270015
rect 325558 269963 325610 270015
rect 371446 269963 371498 270015
rect 375766 269963 375818 270015
rect 387382 269963 387434 270015
rect 387574 270037 387626 270089
rect 583222 270037 583274 270089
rect 669814 270037 669866 270089
rect 674422 270037 674474 270089
rect 586774 269963 586826 270015
rect 79030 269889 79082 269941
rect 83446 269889 83498 269941
rect 247030 269889 247082 269941
rect 459574 269889 459626 269941
rect 469462 269889 469514 269941
rect 488278 269889 488330 269941
rect 226966 269815 227018 269867
rect 295414 269815 295466 269867
rect 310294 269815 310346 269867
rect 323350 269815 323402 269867
rect 323446 269815 323498 269867
rect 325558 269815 325610 269867
rect 325654 269815 325706 269867
rect 524950 269815 525002 269867
rect 235702 269741 235754 269793
rect 366454 269741 366506 269793
rect 366550 269741 366602 269793
rect 379030 269741 379082 269793
rect 379126 269741 379178 269793
rect 597526 269741 597578 269793
rect 660982 269741 661034 269793
rect 674710 269741 674762 269793
rect 247606 269667 247658 269719
rect 466582 269667 466634 269719
rect 248566 269593 248618 269645
rect 473782 269593 473834 269645
rect 236278 269519 236330 269571
rect 358486 269519 358538 269571
rect 358582 269519 358634 269571
rect 387286 269519 387338 269571
rect 387382 269519 387434 269571
rect 604630 269519 604682 269571
rect 227542 269445 227594 269497
rect 302614 269445 302666 269497
rect 312598 269445 312650 269497
rect 542806 269445 542858 269497
rect 249622 269371 249674 269423
rect 480982 269371 481034 269423
rect 228502 269297 228554 269349
rect 309718 269297 309770 269349
rect 313846 269297 313898 269349
rect 553462 269297 553514 269349
rect 221494 269223 221546 269275
rect 251254 269223 251306 269275
rect 251350 269223 251402 269275
rect 495190 269223 495242 269275
rect 243286 269149 243338 269201
rect 431062 269149 431114 269201
rect 663958 269149 664010 269201
rect 674710 269149 674762 269201
rect 242614 269075 242666 269127
rect 423862 269075 423914 269127
rect 241558 269001 241610 269053
rect 416662 269001 416714 269053
rect 428950 269001 429002 269053
rect 429238 269001 429290 269053
rect 229558 268927 229610 268979
rect 313942 268927 313994 268979
rect 314038 268927 314090 268979
rect 325174 268927 325226 268979
rect 325270 268927 325322 268979
rect 327094 268927 327146 268979
rect 327190 268927 327242 268979
rect 336406 268927 336458 268979
rect 351766 268927 351818 268979
rect 378358 268927 378410 268979
rect 240886 268853 240938 268905
rect 378742 268927 378794 268979
rect 387574 268927 387626 268979
rect 388630 268927 388682 268979
rect 388918 268927 388970 268979
rect 390166 268927 390218 268979
rect 395446 268927 395498 268979
rect 398806 268927 398858 268979
rect 536854 268927 536906 268979
rect 409558 268853 409610 268905
rect 225814 268779 225866 268831
rect 288214 268779 288266 268831
rect 313942 268779 313994 268831
rect 316438 268779 316490 268831
rect 317686 268779 317738 268831
rect 371446 268779 371498 268831
rect 371542 268779 371594 268831
rect 372982 268779 373034 268831
rect 373366 268779 373418 268831
rect 378742 268779 378794 268831
rect 379030 268779 379082 268831
rect 529750 268779 529802 268831
rect 240022 268705 240074 268757
rect 378646 268705 378698 268757
rect 378838 268705 378890 268757
rect 398806 268705 398858 268757
rect 403222 268705 403274 268757
rect 403990 268705 404042 268757
rect 210934 268631 210986 268683
rect 271990 268631 272042 268683
rect 272758 268631 272810 268683
rect 334966 268631 335018 268683
rect 348598 268631 348650 268683
rect 373078 268631 373130 268683
rect 373174 268631 373226 268683
rect 377014 268631 377066 268683
rect 377110 268631 377162 268683
rect 526102 268631 526154 268683
rect 238870 268557 238922 268609
rect 372982 268557 373034 268609
rect 238294 268483 238346 268535
rect 371062 268483 371114 268535
rect 371350 268483 371402 268535
rect 378550 268557 378602 268609
rect 378646 268557 378698 268609
rect 402454 268557 402506 268609
rect 403702 268557 403754 268609
rect 409942 268557 409994 268609
rect 373174 268483 373226 268535
rect 382390 268483 382442 268535
rect 382486 268483 382538 268535
rect 395350 268483 395402 268535
rect 395446 268483 395498 268535
rect 408118 268483 408170 268535
rect 237142 268409 237194 268461
rect 357622 268409 357674 268461
rect 357718 268409 357770 268461
rect 358582 268409 358634 268461
rect 366358 268409 366410 268461
rect 377110 268409 377162 268461
rect 377206 268409 377258 268461
rect 390454 268409 390506 268461
rect 403702 268409 403754 268461
rect 406102 268409 406154 268461
rect 499414 268409 499466 268461
rect 502006 268409 502058 268461
rect 218038 268335 218090 268387
rect 272662 268335 272714 268387
rect 283510 268335 283562 268387
rect 336502 268335 336554 268387
rect 357238 268335 357290 268387
rect 358870 268335 358922 268387
rect 359446 268335 359498 268387
rect 378646 268335 378698 268387
rect 378934 268335 378986 268387
rect 501142 268335 501194 268387
rect 228790 268261 228842 268313
rect 274198 268261 274250 268313
rect 290614 268261 290666 268313
rect 337462 268261 337514 268313
rect 353974 268261 354026 268313
rect 222550 268187 222602 268239
rect 259702 268187 259754 268239
rect 260086 268187 260138 268239
rect 355606 268187 355658 268239
rect 358390 268187 358442 268239
rect 360982 268261 361034 268313
rect 483286 268261 483338 268313
rect 223222 268113 223274 268165
rect 266806 268113 266858 268165
rect 287062 268113 287114 268165
rect 235894 268039 235946 268091
rect 274870 268039 274922 268091
rect 294550 268039 294602 268091
rect 315958 268039 316010 268091
rect 221974 267965 222026 268017
rect 256150 267965 256202 268017
rect 286006 267965 286058 268017
rect 316150 267965 316202 268017
rect 316534 268113 316586 268165
rect 337846 268113 337898 268165
rect 426262 268187 426314 268239
rect 499318 268187 499370 268239
rect 499798 268187 499850 268239
rect 370870 268113 370922 268165
rect 372502 268113 372554 268165
rect 378550 268113 378602 268165
rect 378646 268113 378698 268165
rect 468982 268113 469034 268165
rect 316438 268039 316490 268091
rect 322966 268039 323018 268091
rect 323062 268039 323114 268091
rect 326902 268039 326954 268091
rect 326998 268039 327050 268091
rect 324502 267965 324554 268017
rect 324598 267965 324650 268017
rect 328630 267965 328682 268017
rect 329014 268039 329066 268091
rect 348598 268039 348650 268091
rect 336118 267965 336170 268017
rect 336214 267965 336266 268017
rect 371542 268039 371594 268091
rect 371638 268039 371690 268091
rect 387190 268039 387242 268091
rect 387286 268039 387338 268091
rect 454774 268039 454826 268091
rect 355702 267965 355754 268017
rect 440470 267965 440522 268017
rect 243094 267891 243146 267943
rect 275734 267891 275786 267943
rect 285046 267891 285098 267943
rect 317782 267891 317834 267943
rect 322390 267891 322442 267943
rect 326806 267891 326858 267943
rect 326902 267891 326954 267943
rect 65014 267817 65066 267869
rect 67606 267817 67658 267869
rect 258550 267817 258602 267869
rect 358390 267817 358442 267869
rect 377782 267891 377834 267943
rect 378358 267891 378410 267943
rect 358870 267817 358922 267869
rect 371638 267817 371690 267869
rect 372982 267817 373034 267869
rect 377302 267817 377354 267869
rect 377494 267817 377546 267869
rect 378454 267817 378506 267869
rect 379318 267891 379370 267943
rect 386518 267891 386570 267943
rect 388726 267891 388778 267943
rect 390358 267891 390410 267943
rect 390454 267891 390506 267943
rect 413398 267891 413450 267943
rect 390166 267817 390218 267869
rect 390262 267817 390314 267869
rect 413302 267817 413354 267869
rect 204982 267743 205034 267795
rect 312694 267743 312746 267795
rect 319414 267743 319466 267795
rect 322390 267743 322442 267795
rect 322486 267743 322538 267795
rect 621238 267743 621290 267795
rect 276214 267669 276266 267721
rect 298006 267669 298058 267721
rect 287734 267595 287786 267647
rect 297814 267595 297866 267647
rect 279958 267521 280010 267573
rect 326710 267669 326762 267721
rect 326806 267669 326858 267721
rect 376054 267669 376106 267721
rect 378454 267669 378506 267721
rect 379318 267669 379370 267721
rect 379414 267669 379466 267721
rect 389110 267669 389162 267721
rect 389206 267669 389258 267721
rect 414358 267669 414410 267721
rect 298390 267595 298442 267647
rect 327958 267595 328010 267647
rect 311926 267521 311978 267573
rect 320566 267521 320618 267573
rect 321526 267521 321578 267573
rect 377206 267595 377258 267647
rect 377302 267595 377354 267647
rect 382486 267595 382538 267647
rect 383062 267595 383114 267647
rect 385462 267595 385514 267647
rect 387190 267595 387242 267647
rect 389014 267595 389066 267647
rect 390358 267595 390410 267647
rect 399862 267595 399914 267647
rect 403030 267595 403082 267647
rect 410998 267595 411050 267647
rect 328630 267521 328682 267573
rect 138358 267447 138410 267499
rect 140950 267447 141002 267499
rect 290326 267447 290378 267499
rect 338326 267447 338378 267499
rect 353302 267521 353354 267573
rect 419062 267521 419114 267573
rect 357238 267447 357290 267499
rect 357334 267447 357386 267499
rect 368278 267447 368330 267499
rect 368374 267447 368426 267499
rect 377686 267447 377738 267499
rect 377782 267447 377834 267499
rect 378934 267447 378986 267499
rect 379030 267447 379082 267499
rect 382774 267447 382826 267499
rect 389014 267447 389066 267499
rect 390262 267447 390314 267499
rect 395638 267447 395690 267499
rect 398710 267447 398762 267499
rect 398806 267447 398858 267499
rect 421462 267447 421514 267499
rect 288790 267373 288842 267425
rect 346582 267373 346634 267425
rect 355030 267373 355082 267425
rect 433366 267373 433418 267425
rect 291670 267299 291722 267351
rect 363862 267299 363914 267351
rect 368278 267299 368330 267351
rect 378646 267299 378698 267351
rect 379510 267299 379562 267351
rect 383062 267299 383114 267351
rect 387862 267299 387914 267351
rect 629686 267299 629738 267351
rect 289462 267225 289514 267277
rect 353686 267225 353738 267277
rect 356566 267225 356618 267277
rect 447670 267225 447722 267277
rect 293590 267151 293642 267203
rect 379030 267151 379082 267203
rect 379126 267151 379178 267203
rect 387862 267151 387914 267203
rect 388534 267151 388586 267203
rect 419350 267151 419402 267203
rect 262390 267077 262442 267129
rect 333910 267077 333962 267129
rect 351286 267077 351338 267129
rect 357334 267077 357386 267129
rect 357814 267077 357866 267129
rect 458326 267077 458378 267129
rect 295318 267003 295370 267055
rect 378742 267003 378794 267055
rect 378838 267003 378890 267055
rect 398902 267003 398954 267055
rect 403126 267003 403178 267055
rect 411958 267003 412010 267055
rect 295990 266929 296042 266981
rect 389014 266929 389066 266981
rect 389110 266929 389162 266981
rect 404758 266929 404810 266981
rect 408214 266929 408266 266981
rect 408694 266929 408746 266981
rect 251158 266855 251210 266907
rect 332374 266855 332426 266907
rect 359830 266855 359882 266907
rect 472630 266855 472682 266907
rect 296854 266781 296906 266833
rect 389206 266781 389258 266833
rect 389302 266781 389354 266833
rect 412918 266781 412970 266833
rect 298006 266707 298058 266759
rect 398806 266707 398858 266759
rect 398998 266707 399050 266759
rect 408214 266707 408266 266759
rect 408406 266707 408458 266759
rect 413302 266707 413354 266759
rect 298582 266633 298634 266685
rect 428662 266633 428714 266685
rect 244246 266559 244298 266611
rect 331702 266559 331754 266611
rect 338326 266559 338378 266611
rect 360790 266559 360842 266611
rect 362230 266559 362282 266611
rect 494038 266559 494090 266611
rect 237430 266485 237482 266537
rect 330646 266485 330698 266537
rect 362710 266485 362762 266537
rect 497590 266485 497642 266537
rect 299734 266411 299786 266463
rect 435670 266411 435722 266463
rect 300310 266337 300362 266389
rect 442870 266337 442922 266389
rect 521590 266337 521642 266389
rect 523510 266337 523562 266389
rect 301270 266263 301322 266315
rect 449974 266263 450026 266315
rect 230038 266189 230090 266241
rect 329974 266189 330026 266241
rect 365974 266189 366026 266241
rect 522550 266189 522602 266241
rect 302326 266115 302378 266167
rect 457174 266115 457226 266167
rect 302998 266041 303050 266093
rect 464278 266041 464330 266093
rect 304054 265967 304106 266019
rect 471382 265967 471434 266019
rect 226390 265893 226442 265945
rect 329590 265893 329642 265945
rect 367030 265893 367082 265945
rect 378838 265893 378890 265945
rect 378934 265893 378986 265945
rect 398806 265893 398858 265945
rect 398902 265893 398954 265945
rect 533206 265893 533258 265945
rect 304726 265819 304778 265871
rect 478582 265819 478634 265871
rect 305590 265745 305642 265797
rect 485686 265745 485738 265797
rect 212470 265671 212522 265723
rect 327862 265671 327914 265723
rect 327958 265671 328010 265723
rect 339094 265671 339146 265723
rect 350710 265671 350762 265723
rect 368374 265671 368426 265723
rect 368566 265671 368618 265723
rect 370678 265671 370730 265723
rect 306742 265597 306794 265649
rect 377206 265597 377258 265649
rect 378934 265597 378986 265649
rect 379030 265597 379082 265649
rect 397558 265597 397610 265649
rect 398806 265671 398858 265723
rect 419254 265671 419306 265723
rect 419350 265671 419402 265723
rect 547606 265671 547658 265723
rect 492886 265597 492938 265649
rect 307318 265523 307370 265575
rect 499894 265523 499946 265575
rect 309334 265449 309386 265501
rect 309910 265375 309962 265427
rect 311638 265301 311690 265353
rect 221686 265227 221738 265279
rect 273142 265227 273194 265279
rect 313270 265227 313322 265279
rect 319318 265227 319370 265279
rect 255670 265153 255722 265205
rect 267862 265153 267914 265205
rect 276502 265153 276554 265205
rect 308086 265153 308138 265205
rect 219574 265079 219626 265131
rect 201430 265005 201482 265057
rect 311926 265005 311978 265057
rect 319414 265079 319466 265131
rect 369334 265227 369386 265279
rect 369718 265301 369770 265353
rect 378166 265301 378218 265353
rect 378358 265375 378410 265427
rect 378742 265375 378794 265427
rect 378934 265449 378986 265501
rect 379702 265375 379754 265427
rect 379606 265301 379658 265353
rect 379894 265449 379946 265501
rect 392950 265449 393002 265501
rect 395734 265449 395786 265501
rect 407062 265449 407114 265501
rect 408214 265449 408266 265501
rect 412822 265449 412874 265501
rect 379990 265375 380042 265427
rect 514294 265449 514346 265501
rect 419062 265375 419114 265427
rect 521398 265375 521450 265427
rect 379414 265227 379466 265279
rect 379990 265227 380042 265279
rect 380182 265301 380234 265353
rect 388822 265301 388874 265353
rect 389590 265301 389642 265353
rect 389782 265301 389834 265353
rect 395734 265301 395786 265353
rect 395926 265301 395978 265353
rect 535606 265301 535658 265353
rect 320278 265153 320330 265205
rect 327286 265153 327338 265205
rect 329398 265153 329450 265205
rect 375958 265153 376010 265205
rect 376054 265153 376106 265205
rect 379510 265153 379562 265205
rect 381142 265153 381194 265205
rect 419062 265227 419114 265279
rect 419158 265227 419210 265279
rect 546358 265227 546410 265279
rect 388534 265153 388586 265205
rect 389014 265153 389066 265205
rect 390454 265153 390506 265205
rect 328438 265079 328490 265131
rect 267766 264931 267818 264983
rect 312694 264931 312746 264983
rect 320566 265005 320618 265057
rect 326230 265005 326282 265057
rect 367126 265079 367178 265131
rect 369334 265079 369386 265131
rect 390262 265079 390314 265131
rect 608182 265153 608234 265205
rect 325078 264931 325130 264983
rect 210646 264857 210698 264909
rect 212470 264857 212522 264909
rect 325750 264931 325802 264983
rect 326710 264931 326762 264983
rect 327286 264931 327338 264983
rect 329398 264931 329450 264983
rect 329494 264931 329546 264983
rect 341014 264931 341066 264983
rect 349846 264857 349898 264909
rect 376438 265005 376490 265057
rect 399382 265079 399434 265131
rect 419158 265079 419210 265131
rect 419254 265079 419306 265131
rect 615382 265079 615434 265131
rect 390454 265005 390506 265057
rect 406966 265005 407018 265057
rect 407062 265005 407114 265057
rect 412726 265005 412778 265057
rect 379030 264931 379082 264983
rect 379126 264931 379178 264983
rect 389782 264931 389834 264983
rect 390262 264931 390314 264983
rect 399382 264931 399434 264983
rect 399862 264931 399914 264983
rect 412630 264931 412682 264983
rect 369046 264857 369098 264909
rect 369718 264857 369770 264909
rect 371542 264857 371594 264909
rect 388054 264857 388106 264909
rect 625846 262045 625898 262097
rect 633622 262119 633674 262171
rect 642262 260491 642314 260543
rect 645718 260491 645770 260543
rect 42550 259677 42602 259729
rect 50518 259677 50570 259729
rect 83542 259307 83594 259359
rect 95062 259159 95114 259211
rect 42646 258937 42698 258989
rect 53398 258937 53450 258989
rect 42550 258197 42602 258249
rect 47446 258197 47498 258249
rect 42262 257753 42314 257805
rect 43126 257753 43178 257805
rect 616342 257753 616394 257805
rect 625846 257753 625898 257805
rect 42550 257161 42602 257213
rect 43222 257161 43274 257213
rect 639286 256347 639338 256399
rect 677014 256347 677066 256399
rect 67606 253387 67658 253439
rect 74902 253387 74954 253439
rect 675190 250945 675242 250997
rect 675382 250945 675434 250997
rect 607702 250575 607754 250627
rect 616342 250575 616394 250627
rect 636502 250575 636554 250627
rect 642262 250575 642314 250627
rect 674518 250353 674570 250405
rect 675190 250353 675242 250405
rect 74902 249317 74954 249369
rect 90646 249317 90698 249369
rect 56182 249243 56234 249295
rect 205558 249243 205610 249295
rect 53782 249169 53834 249221
rect 210742 249169 210794 249221
rect 45046 249095 45098 249147
rect 206902 249095 206954 249147
rect 200086 247689 200138 247741
rect 627862 247689 627914 247741
rect 636502 247689 636554 247741
rect 205270 247615 205322 247667
rect 126550 247319 126602 247371
rect 129526 247245 129578 247297
rect 132310 247171 132362 247223
rect 135190 247097 135242 247149
rect 140950 247023 141002 247075
rect 143926 246949 143978 247001
rect 146710 246875 146762 246927
rect 80470 246801 80522 246853
rect 86518 246801 86570 246853
rect 171286 246801 171338 246853
rect 181366 246801 181418 246853
rect 211702 246801 211754 246853
rect 63286 246727 63338 246779
rect 204598 246727 204650 246779
rect 211894 246727 211946 246779
rect 227446 246727 227498 246779
rect 227926 246727 227978 246779
rect 47638 246653 47690 246705
rect 65014 246653 65066 246705
rect 65206 246653 65258 246705
rect 171286 246653 171338 246705
rect 181366 246653 181418 246705
rect 210934 246653 210986 246705
rect 212086 246653 212138 246705
rect 227062 246653 227114 246705
rect 227830 246653 227882 246705
rect 231862 246727 231914 246779
rect 247894 246727 247946 246779
rect 248182 246727 248234 246779
rect 248278 246727 248330 246779
rect 251926 246727 251978 246779
rect 276886 246727 276938 246779
rect 280822 246727 280874 246779
rect 280918 246727 280970 246779
rect 284950 246727 285002 246779
rect 288310 246727 288362 246779
rect 288694 246727 288746 246779
rect 292246 246727 292298 246779
rect 232150 246653 232202 246705
rect 56086 246579 56138 246631
rect 180982 246579 181034 246631
rect 181270 246579 181322 246631
rect 204790 246579 204842 246631
rect 211798 246579 211850 246631
rect 226486 246579 226538 246631
rect 226966 246579 227018 246631
rect 53494 246505 53546 246557
rect 204502 246505 204554 246557
rect 225334 246505 225386 246557
rect 227830 246505 227882 246557
rect 231382 246579 231434 246631
rect 248182 246579 248234 246631
rect 53206 246431 53258 246483
rect 204694 246431 204746 246483
rect 211990 246431 212042 246483
rect 247318 246505 247370 246557
rect 252118 246579 252170 246631
rect 281302 246653 281354 246705
rect 287542 246653 287594 246705
rect 295702 246727 295754 246779
rect 309238 246727 309290 246779
rect 309334 246727 309386 246779
rect 309430 246727 309482 246779
rect 311734 246653 311786 246705
rect 276982 246505 277034 246557
rect 249046 246431 249098 246483
rect 259126 246431 259178 246483
rect 268822 246431 268874 246483
rect 274102 246431 274154 246483
rect 80470 246357 80522 246409
rect 145846 246357 145898 246409
rect 161302 246357 161354 246409
rect 44758 246283 44810 246335
rect 160918 246283 160970 246335
rect 165526 246283 165578 246335
rect 199606 246283 199658 246335
rect 212182 246357 212234 246409
rect 230902 246357 230954 246409
rect 247798 246357 247850 246409
rect 260758 246357 260810 246409
rect 214198 246283 214250 246335
rect 227926 246283 227978 246335
rect 268054 246357 268106 246409
rect 268630 246357 268682 246409
rect 280918 246505 280970 246557
rect 288406 246579 288458 246631
rect 292246 246579 292298 246631
rect 313750 246727 313802 246779
rect 314038 246727 314090 246779
rect 397270 246727 397322 246779
rect 397750 246727 397802 246779
rect 313942 246653 313994 246705
rect 397366 246653 397418 246705
rect 312310 246579 312362 246631
rect 294838 246505 294890 246557
rect 280822 246431 280874 246483
rect 277366 246357 277418 246409
rect 268246 246283 268298 246335
rect 280822 246283 280874 246335
rect 44566 246209 44618 246261
rect 161014 246209 161066 246261
rect 163702 246209 163754 246261
rect 198742 246209 198794 246261
rect 210262 246209 210314 246261
rect 229270 246209 229322 246261
rect 230902 246209 230954 246261
rect 260854 246209 260906 246261
rect 268534 246209 268586 246261
rect 289174 246431 289226 246483
rect 311158 246431 311210 246483
rect 311734 246505 311786 246557
rect 313750 246579 313802 246631
rect 398230 246727 398282 246779
rect 403030 246727 403082 246779
rect 674326 247245 674378 247297
rect 675190 247245 675242 247297
rect 674806 247171 674858 247223
rect 675094 247171 675146 247223
rect 406102 246727 406154 246779
rect 406966 246727 407018 246779
rect 408982 246727 409034 246779
rect 408310 246653 408362 246705
rect 288694 246357 288746 246409
rect 307510 246357 307562 246409
rect 307702 246357 307754 246409
rect 307990 246357 308042 246409
rect 312310 246357 312362 246409
rect 313270 246357 313322 246409
rect 328918 246505 328970 246557
rect 330646 246505 330698 246557
rect 342742 246505 342794 246557
rect 347254 246505 347306 246557
rect 349654 246505 349706 246557
rect 366454 246505 366506 246557
rect 313654 246431 313706 246483
rect 339862 246431 339914 246483
rect 313942 246357 313994 246409
rect 317206 246357 317258 246409
rect 317494 246357 317546 246409
rect 328438 246357 328490 246409
rect 347254 246357 347306 246409
rect 309334 246283 309386 246335
rect 349078 246431 349130 246483
rect 348598 246357 348650 246409
rect 367222 246431 367274 246483
rect 367414 246505 367466 246557
rect 367990 246505 368042 246557
rect 368470 246505 368522 246557
rect 397654 246505 397706 246557
rect 406582 246579 406634 246631
rect 406390 246505 406442 246557
rect 382870 246431 382922 246483
rect 382966 246431 383018 246483
rect 389398 246431 389450 246483
rect 397750 246431 397802 246483
rect 349942 246357 349994 246409
rect 368470 246357 368522 246409
rect 369526 246357 369578 246409
rect 370678 246357 370730 246409
rect 372982 246357 373034 246409
rect 407734 246357 407786 246409
rect 348214 246283 348266 246335
rect 388918 246283 388970 246335
rect 397846 246283 397898 246335
rect 407350 246283 407402 246335
rect 408118 246357 408170 246409
rect 410518 246357 410570 246409
rect 410806 246283 410858 246335
rect 674902 246283 674954 246335
rect 65014 246135 65066 246187
rect 80470 246135 80522 246187
rect 145846 246135 145898 246187
rect 43414 246061 43466 246113
rect 207286 246135 207338 246187
rect 161302 246061 161354 246113
rect 161494 246061 161546 246113
rect 155542 245987 155594 246039
rect 210166 246061 210218 246113
rect 228310 246061 228362 246113
rect 249142 246061 249194 246113
rect 260374 246061 260426 246113
rect 268150 246135 268202 246187
rect 287350 246135 287402 246187
rect 287926 246209 287978 246261
rect 288022 246209 288074 246261
rect 328246 246209 328298 246261
rect 328342 246209 328394 246261
rect 339958 246209 340010 246261
rect 340150 246209 340202 246261
rect 287830 246135 287882 246187
rect 288118 246135 288170 246187
rect 307702 246135 307754 246187
rect 307894 246135 307946 246187
rect 328150 246135 328202 246187
rect 268822 246061 268874 246113
rect 268918 246061 268970 246113
rect 277750 246061 277802 246113
rect 329686 246135 329738 246187
rect 339670 246135 339722 246187
rect 339766 246135 339818 246187
rect 348214 246135 348266 246187
rect 348406 246135 348458 246187
rect 348502 246135 348554 246187
rect 391222 246209 391274 246261
rect 397270 246209 397322 246261
rect 411190 246209 411242 246261
rect 349366 246135 349418 246187
rect 382966 246135 383018 246187
rect 236182 245987 236234 246039
rect 161014 245913 161066 245965
rect 163702 245913 163754 245965
rect 208726 245913 208778 245965
rect 248278 245987 248330 246039
rect 259126 245987 259178 246039
rect 251734 245913 251786 245965
rect 277366 245913 277418 245965
rect 277558 245913 277610 245965
rect 368086 245987 368138 246039
rect 278038 245913 278090 245965
rect 367510 245913 367562 245965
rect 397366 246135 397418 246187
rect 411766 246135 411818 246187
rect 505846 246061 505898 246113
rect 675286 246061 675338 246113
rect 391222 245987 391274 246039
rect 412342 245987 412394 246039
rect 398230 245913 398282 245965
rect 408118 245913 408170 245965
rect 160918 245839 160970 245891
rect 165526 245839 165578 245891
rect 229270 245839 229322 245891
rect 246262 245839 246314 245891
rect 247894 245839 247946 245891
rect 251926 245839 251978 245891
rect 155542 245765 155594 245817
rect 161494 245765 161546 245817
rect 210358 245765 210410 245817
rect 226966 245765 227018 245817
rect 227446 245765 227498 245817
rect 231862 245765 231914 245817
rect 248182 245765 248234 245817
rect 252118 245765 252170 245817
rect 206902 245691 206954 245743
rect 207286 245691 207338 245743
rect 224854 245691 224906 245743
rect 228118 245691 228170 245743
rect 251350 245691 251402 245743
rect 356278 245839 356330 245891
rect 366838 245839 366890 245891
rect 372982 245839 373034 245891
rect 389398 245839 389450 245891
rect 411382 245839 411434 245891
rect 255094 245765 255146 245817
rect 330646 245765 330698 245817
rect 330742 245765 330794 245817
rect 357142 245765 357194 245817
rect 367990 245765 368042 245817
rect 373462 245765 373514 245817
rect 388918 245765 388970 245817
rect 406006 245765 406058 245817
rect 254134 245691 254186 245743
rect 348502 245691 348554 245743
rect 348598 245691 348650 245743
rect 357430 245691 357482 245743
rect 367222 245691 367274 245743
rect 370198 245691 370250 245743
rect 382870 245691 382922 245743
rect 408214 245691 408266 245743
rect 227062 245617 227114 245669
rect 232150 245617 232202 245669
rect 246454 245617 246506 245669
rect 267478 245617 267530 245669
rect 269014 245617 269066 245669
rect 369238 245617 369290 245669
rect 389014 245617 389066 245669
rect 406774 245617 406826 245669
rect 226486 245543 226538 245595
rect 231382 245543 231434 245595
rect 236182 245543 236234 245595
rect 249046 245543 249098 245595
rect 268438 245543 268490 245595
rect 277654 245543 277706 245595
rect 277750 245543 277802 245595
rect 370966 245543 371018 245595
rect 403030 245543 403082 245595
rect 410326 245543 410378 245595
rect 223126 245469 223178 245521
rect 251734 245469 251786 245521
rect 252406 245469 252458 245521
rect 330742 245469 330794 245521
rect 198838 245395 198890 245447
rect 213142 245395 213194 245447
rect 246166 245395 246218 245447
rect 248374 245395 248426 245447
rect 253366 245395 253418 245447
rect 348502 245469 348554 245521
rect 355798 245469 355850 245521
rect 210166 245321 210218 245373
rect 231862 245321 231914 245373
rect 246262 245321 246314 245373
rect 249142 245321 249194 245373
rect 249622 245321 249674 245373
rect 348694 245395 348746 245447
rect 390262 245469 390314 245521
rect 405910 245469 405962 245521
rect 412150 245469 412202 245521
rect 331030 245321 331082 245373
rect 370102 245321 370154 245373
rect 250294 245247 250346 245299
rect 216598 245173 216650 245225
rect 331030 245173 331082 245225
rect 339670 245247 339722 245299
rect 369910 245247 369962 245299
rect 370198 245247 370250 245299
rect 380182 245247 380234 245299
rect 355894 245173 355946 245225
rect 231862 245099 231914 245151
rect 260278 245099 260330 245151
rect 261814 245099 261866 245151
rect 338422 245099 338474 245151
rect 339478 245099 339530 245151
rect 263446 245025 263498 245077
rect 263830 244951 263882 245003
rect 267478 244951 267530 245003
rect 269494 245025 269546 245077
rect 277558 244951 277610 245003
rect 277942 245025 277994 245077
rect 369910 245099 369962 245151
rect 398710 245099 398762 245151
rect 319702 244951 319754 245003
rect 339958 244951 340010 245003
rect 372022 245025 372074 245077
rect 380182 245025 380234 245077
rect 411478 245173 411530 245225
rect 42550 244877 42602 244929
rect 214294 244877 214346 244929
rect 216502 244877 216554 244929
rect 338134 244877 338186 244929
rect 338422 244877 338474 244929
rect 339478 244877 339530 244929
rect 348886 244877 348938 244929
rect 358006 244877 358058 244929
rect 210070 244803 210122 244855
rect 228598 244803 228650 244855
rect 260278 244803 260330 244855
rect 267958 244803 268010 244855
rect 268054 244803 268106 244855
rect 278038 244803 278090 244855
rect 278134 244803 278186 244855
rect 287254 244803 287306 244855
rect 287350 244803 287402 244855
rect 288790 244803 288842 244855
rect 288886 244803 288938 244855
rect 309430 244803 309482 244855
rect 311830 244803 311882 244855
rect 95062 244729 95114 244781
rect 139990 244729 140042 244781
rect 260950 244729 261002 244781
rect 316822 244729 316874 244781
rect 316918 244729 316970 244781
rect 321238 244729 321290 244781
rect 328630 244803 328682 244855
rect 339574 244803 339626 244855
rect 329686 244729 329738 244781
rect 90646 244655 90698 244707
rect 142486 244655 142538 244707
rect 262870 244655 262922 244707
rect 273046 244655 273098 244707
rect 276022 244655 276074 244707
rect 287446 244655 287498 244707
rect 287926 244655 287978 244707
rect 307318 244655 307370 244707
rect 307414 244655 307466 244707
rect 311830 244655 311882 244707
rect 311926 244655 311978 244707
rect 317014 244655 317066 244707
rect 317110 244655 317162 244707
rect 339958 244655 340010 244707
rect 138166 244581 138218 244633
rect 206998 244581 207050 244633
rect 265942 244581 265994 244633
rect 135286 244507 135338 244559
rect 207094 244507 207146 244559
rect 267478 244507 267530 244559
rect 268054 244507 268106 244559
rect 132406 244433 132458 244485
rect 205174 244433 205226 244485
rect 267958 244433 268010 244485
rect 269206 244433 269258 244485
rect 126646 244359 126698 244411
rect 205558 244359 205610 244411
rect 274102 244581 274154 244633
rect 278038 244581 278090 244633
rect 278134 244581 278186 244633
rect 276886 244507 276938 244559
rect 277750 244507 277802 244559
rect 308950 244581 309002 244633
rect 309238 244581 309290 244633
rect 314038 244581 314090 244633
rect 287830 244507 287882 244559
rect 306646 244507 306698 244559
rect 307510 244507 307562 244559
rect 277846 244433 277898 244485
rect 310774 244433 310826 244485
rect 312022 244507 312074 244559
rect 319606 244581 319658 244633
rect 338326 244581 338378 244633
rect 339574 244581 339626 244633
rect 348694 244803 348746 244855
rect 374038 244951 374090 245003
rect 374614 244803 374666 244855
rect 342550 244655 342602 244707
rect 389302 244729 389354 244781
rect 340150 244581 340202 244633
rect 349942 244581 349994 244633
rect 367894 244507 367946 244559
rect 311926 244359 311978 244411
rect 312406 244433 312458 244485
rect 368758 244433 368810 244485
rect 123766 244285 123818 244337
rect 205366 244285 205418 244337
rect 235126 244285 235178 244337
rect 267190 244285 267242 244337
rect 273046 244285 273098 244337
rect 287734 244285 287786 244337
rect 290038 244285 290090 244337
rect 295702 244285 295754 244337
rect 297430 244285 297482 244337
rect 314902 244285 314954 244337
rect 120886 244211 120938 244263
rect 205654 244211 205706 244263
rect 260758 244211 260810 244263
rect 268150 244211 268202 244263
rect 268246 244211 268298 244263
rect 287446 244211 287498 244263
rect 287926 244211 287978 244263
rect 319606 244285 319658 244337
rect 319798 244285 319850 244337
rect 339862 244359 339914 244411
rect 349366 244211 349418 244263
rect 118006 244137 118058 244189
rect 204982 244137 205034 244189
rect 258358 244137 258410 244189
rect 317206 244137 317258 244189
rect 321238 244137 321290 244189
rect 329302 244137 329354 244189
rect 338134 244137 338186 244189
rect 351574 244137 351626 244189
rect 112246 244063 112298 244115
rect 206614 244063 206666 244115
rect 261142 244063 261194 244115
rect 337558 244063 337610 244115
rect 109366 243989 109418 244041
rect 205750 243989 205802 244041
rect 256342 243989 256394 244041
rect 335350 243989 335402 244041
rect 106486 243915 106538 243967
rect 206518 243915 206570 243967
rect 260086 243915 260138 243967
rect 316822 243915 316874 243967
rect 328246 243915 328298 243967
rect 339766 243915 339818 243967
rect 103606 243841 103658 243893
rect 206326 243841 206378 243893
rect 207190 243841 207242 243893
rect 268054 243841 268106 243893
rect 268150 243841 268202 243893
rect 285238 243841 285290 243893
rect 288118 243841 288170 243893
rect 308086 243841 308138 243893
rect 313366 243841 313418 243893
rect 370294 243841 370346 243893
rect 100726 243767 100778 243819
rect 206422 243767 206474 243819
rect 245398 243767 245450 243819
rect 353686 243767 353738 243819
rect 94966 243693 95018 243745
rect 206230 243693 206282 243745
rect 239350 243693 239402 243745
rect 350806 243693 350858 243745
rect 604822 243693 604874 243745
rect 624886 243693 624938 243745
rect 92086 243619 92138 243671
rect 206038 243619 206090 243671
rect 206806 243619 206858 243671
rect 207190 243619 207242 243671
rect 227062 243619 227114 243671
rect 231670 243619 231722 243671
rect 231766 243619 231818 243671
rect 347350 243619 347402 243671
rect 443542 243619 443594 243671
rect 463606 243619 463658 243671
rect 483862 243619 483914 243671
rect 503926 243619 503978 243671
rect 524182 243619 524234 243671
rect 544246 243619 544298 243671
rect 564502 243619 564554 243671
rect 584566 243619 584618 243671
rect 645142 243619 645194 243671
rect 648022 243619 648074 243671
rect 86326 243545 86378 243597
rect 206710 243545 206762 243597
rect 236278 243545 236330 243597
rect 349270 243545 349322 243597
rect 80566 243471 80618 243523
rect 206806 243471 206858 243523
rect 228502 243471 228554 243523
rect 345622 243471 345674 243523
rect 77686 243397 77738 243449
rect 205942 243397 205994 243449
rect 226774 243397 226826 243449
rect 345142 243397 345194 243449
rect 69046 243323 69098 243375
rect 206134 243323 206186 243375
rect 229750 243323 229802 243375
rect 297814 243323 297866 243375
rect 199606 243249 199658 243301
rect 213526 243249 213578 243301
rect 264790 243249 264842 243301
rect 277846 243249 277898 243301
rect 283222 243249 283274 243301
rect 298198 243323 298250 243375
rect 298486 243323 298538 243375
rect 299446 243323 299498 243375
rect 346390 243323 346442 243375
rect 298294 243249 298346 243301
rect 316918 243249 316970 243301
rect 340726 243249 340778 243301
rect 342742 243249 342794 243301
rect 358390 243249 358442 243301
rect 267382 243175 267434 243227
rect 298582 243175 298634 243227
rect 298678 243175 298730 243227
rect 305110 243175 305162 243227
rect 317206 243175 317258 243227
rect 336310 243175 336362 243227
rect 260374 243101 260426 243153
rect 268630 243101 268682 243153
rect 270838 243101 270890 243153
rect 293110 243101 293162 243153
rect 293398 243101 293450 243153
rect 294358 243101 294410 243153
rect 223510 243027 223562 243079
rect 227350 243027 227402 243079
rect 265270 243027 265322 243079
rect 278134 243027 278186 243079
rect 205270 242953 205322 243005
rect 208534 242953 208586 243005
rect 260854 242953 260906 243005
rect 268534 242953 268586 243005
rect 269878 242953 269930 243005
rect 293782 243027 293834 243079
rect 293878 243027 293930 243079
rect 294454 243027 294506 243079
rect 279094 242953 279146 243005
rect 287542 242953 287594 243005
rect 287734 242953 287786 243005
rect 298870 243101 298922 243153
rect 321334 243101 321386 243153
rect 303382 243027 303434 243079
rect 316822 243027 316874 243079
rect 337078 243027 337130 243079
rect 298582 242953 298634 243005
rect 314326 242953 314378 243005
rect 674614 242953 674666 243005
rect 675382 242953 675434 243005
rect 266038 242879 266090 242931
rect 276022 242879 276074 242931
rect 278038 242879 278090 242931
rect 288310 242879 288362 242931
rect 288598 242879 288650 242931
rect 293398 242879 293450 242931
rect 293590 242879 293642 242931
rect 297910 242879 297962 242931
rect 227830 242805 227882 242857
rect 247798 242805 247850 242857
rect 266614 242805 266666 242857
rect 279094 242805 279146 242857
rect 280822 242805 280874 242857
rect 288886 242805 288938 242857
rect 288982 242805 289034 242857
rect 297430 242805 297482 242857
rect 297814 242805 297866 242857
rect 299446 242879 299498 242931
rect 299638 242879 299690 242931
rect 317398 242879 317450 242931
rect 307702 242805 307754 242857
rect 308278 242805 308330 242857
rect 338134 242805 338186 242857
rect 339190 242805 339242 242857
rect 227062 242731 227114 242783
rect 227638 242731 227690 242783
rect 268054 242731 268106 242783
rect 227350 242657 227402 242709
rect 227734 242657 227786 242709
rect 267766 242657 267818 242709
rect 268246 242657 268298 242709
rect 269686 242657 269738 242709
rect 278134 242657 278186 242709
rect 278326 242731 278378 242783
rect 287542 242657 287594 242709
rect 287638 242657 287690 242709
rect 288022 242657 288074 242709
rect 288214 242731 288266 242783
rect 299638 242731 299690 242783
rect 305782 242731 305834 242783
rect 320374 242731 320426 242783
rect 339862 242731 339914 242783
rect 340246 242731 340298 242783
rect 299542 242657 299594 242709
rect 299734 242657 299786 242709
rect 269206 242583 269258 242635
rect 301270 242583 301322 242635
rect 305782 242583 305834 242635
rect 308086 242657 308138 242709
rect 328726 242657 328778 242709
rect 322582 242583 322634 242635
rect 328342 242583 328394 242635
rect 338806 242583 338858 242635
rect 223990 242509 224042 242561
rect 247318 242509 247370 242561
rect 268150 242509 268202 242561
rect 287734 242509 287786 242561
rect 288118 242509 288170 242561
rect 95062 242435 95114 242487
rect 106582 242435 106634 242487
rect 138262 242435 138314 242487
rect 171382 242435 171434 242487
rect 276982 242435 277034 242487
rect 283990 242435 284042 242487
rect 286486 242435 286538 242487
rect 298006 242435 298058 242487
rect 298102 242435 298154 242487
rect 323446 242509 323498 242561
rect 443542 242509 443594 242561
rect 463606 242509 463658 242561
rect 483862 242509 483914 242561
rect 503926 242509 503978 242561
rect 306646 242435 306698 242487
rect 316918 242435 316970 242487
rect 317014 242435 317066 242487
rect 317494 242435 317546 242487
rect 175702 242361 175754 242413
rect 195766 242361 195818 242413
rect 283702 242361 283754 242413
rect 320182 242361 320234 242413
rect 674134 242361 674186 242413
rect 675382 242361 675434 242413
rect 241942 242287 241994 242339
rect 242326 242287 242378 242339
rect 271894 242287 271946 242339
rect 355222 242287 355274 242339
rect 244438 242213 244490 242265
rect 353014 242213 353066 242265
rect 40054 242139 40106 242191
rect 42262 242139 42314 242191
rect 238294 242139 238346 242191
rect 350038 242139 350090 242191
rect 39958 242065 40010 242117
rect 42934 242065 42986 242117
rect 238966 242065 239018 242117
rect 347830 242065 347882 242117
rect 40150 241991 40202 242043
rect 42550 241991 42602 242043
rect 144022 241991 144074 242043
rect 182806 241991 182858 242043
rect 40246 241917 40298 241969
rect 42358 241917 42410 241969
rect 50326 241917 50378 241969
rect 205846 241917 205898 241969
rect 217558 241843 217610 241895
rect 234454 241843 234506 241895
rect 234550 241843 234602 241895
rect 348598 241991 348650 242043
rect 241078 241843 241130 241895
rect 351766 241917 351818 241969
rect 412054 241917 412106 241969
rect 412246 241917 412298 241969
rect 251830 241843 251882 241895
rect 215446 241769 215498 241821
rect 221398 241769 221450 241821
rect 233494 241769 233546 241821
rect 238966 241769 239018 241821
rect 264310 241769 264362 241821
rect 271990 241769 272042 241821
rect 273142 241843 273194 241895
rect 283894 241843 283946 241895
rect 283990 241843 284042 241895
rect 288598 241843 288650 241895
rect 288694 241843 288746 241895
rect 307894 241843 307946 241895
rect 311734 241843 311786 241895
rect 325174 241843 325226 241895
rect 325270 241843 325322 241895
rect 374422 241843 374474 241895
rect 376054 241843 376106 241895
rect 403222 241843 403274 241895
rect 602902 241843 602954 241895
rect 607702 241917 607754 241969
rect 273622 241769 273674 241821
rect 278230 241769 278282 241821
rect 327958 241769 328010 241821
rect 329302 241769 329354 241821
rect 354550 241769 354602 241821
rect 360598 241769 360650 241821
rect 378646 241769 378698 241821
rect 378742 241769 378794 241821
rect 396406 241769 396458 241821
rect 218710 241695 218762 241747
rect 234358 241695 234410 241747
rect 237430 241695 237482 241747
rect 262198 241695 262250 241747
rect 277654 241695 277706 241747
rect 329974 241695 330026 241747
rect 331030 241695 331082 241747
rect 358294 241695 358346 241747
rect 363190 241695 363242 241747
rect 400150 241695 400202 241747
rect 219286 241621 219338 241673
rect 233782 241621 233834 241673
rect 252790 241621 252842 241673
rect 311734 241621 311786 241673
rect 213910 241547 213962 241599
rect 229174 241547 229226 241599
rect 269302 241547 269354 241599
rect 311638 241547 311690 241599
rect 222550 241473 222602 241525
rect 232534 241473 232586 241525
rect 254998 241473 255050 241525
rect 336502 241621 336554 241673
rect 361558 241621 361610 241673
rect 317878 241547 317930 241599
rect 330166 241547 330218 241599
rect 330262 241547 330314 241599
rect 355702 241547 355754 241599
rect 378646 241621 378698 241673
rect 394102 241621 394154 241673
rect 378742 241547 378794 241599
rect 674998 241547 675050 241599
rect 675478 241547 675530 241599
rect 317494 241473 317546 241525
rect 326902 241473 326954 241525
rect 327190 241473 327242 241525
rect 336118 241473 336170 241525
rect 363766 241473 363818 241525
rect 400726 241473 400778 241525
rect 239158 241399 239210 241451
rect 258550 241399 258602 241451
rect 274102 241399 274154 241451
rect 318262 241399 318314 241451
rect 320470 241399 320522 241451
rect 326998 241399 327050 241451
rect 331510 241399 331562 241451
rect 359350 241399 359402 241451
rect 362326 241399 362378 241451
rect 398422 241399 398474 241451
rect 255958 241325 256010 241377
rect 244726 241251 244778 241303
rect 317494 241251 317546 241303
rect 326710 241325 326762 241377
rect 328918 241325 328970 241377
rect 332278 241325 332330 241377
rect 361078 241325 361130 241377
rect 364150 241325 364202 241377
rect 401878 241325 401930 241377
rect 334486 241251 334538 241303
rect 361942 241251 361994 241303
rect 397462 241251 397514 241303
rect 226294 241177 226346 241229
rect 230710 241177 230762 241229
rect 253750 241177 253802 241229
rect 339382 241177 339434 241229
rect 362422 241177 362474 241229
rect 398998 241177 399050 241229
rect 216694 241103 216746 241155
rect 238390 241103 238442 241155
rect 254230 241103 254282 241155
rect 337846 241103 337898 241155
rect 339670 241103 339722 241155
rect 360502 241103 360554 241155
rect 364534 241103 364586 241155
rect 402742 241103 402794 241155
rect 221494 241029 221546 241081
rect 232918 241029 232970 241081
rect 237526 241029 237578 241081
rect 254614 241029 254666 241081
rect 274486 241029 274538 241081
rect 287638 241029 287690 241081
rect 288310 241029 288362 241081
rect 290038 241029 290090 241081
rect 291958 241029 292010 241081
rect 376150 241029 376202 241081
rect 379222 241029 379274 241081
rect 409270 241029 409322 241081
rect 225238 240955 225290 241007
rect 231190 240955 231242 241007
rect 257686 240955 257738 241007
rect 327862 240955 327914 241007
rect 327958 240955 328010 241007
rect 329590 240955 329642 241007
rect 330742 240955 330794 241007
rect 333622 240955 333674 241007
rect 333718 240955 333770 241007
rect 364342 240955 364394 241007
rect 366358 240955 366410 241007
rect 407158 240955 407210 241007
rect 225430 240881 225482 240933
rect 230902 240881 230954 240933
rect 212758 240807 212810 240859
rect 233302 240807 233354 240859
rect 224086 240733 224138 240785
rect 231574 240733 231626 240785
rect 219286 240659 219338 240711
rect 250678 240881 250730 240933
rect 252310 240881 252362 240933
rect 342646 240881 342698 240933
rect 365014 240881 365066 240933
rect 404470 240881 404522 240933
rect 237814 240807 237866 240859
rect 252886 240807 252938 240859
rect 237718 240733 237770 240785
rect 252022 240733 252074 240785
rect 240310 240659 240362 240711
rect 244150 240659 244202 240711
rect 251542 240659 251594 240711
rect 344182 240807 344234 240859
rect 367222 240807 367274 240859
rect 408886 240807 408938 240859
rect 255478 240733 255530 240785
rect 263350 240733 263402 240785
rect 271030 240733 271082 240785
rect 281398 240733 281450 240785
rect 282262 240733 282314 240785
rect 375766 240733 375818 240785
rect 379606 240733 379658 240785
rect 409942 240733 409994 240785
rect 41782 240585 41834 240637
rect 220246 240585 220298 240637
rect 248662 240585 248714 240637
rect 250582 240585 250634 240637
rect 345718 240659 345770 240711
rect 364630 240659 364682 240711
rect 403414 240659 403466 240711
rect 257878 240585 257930 240637
rect 348310 240585 348362 240637
rect 365398 240585 365450 240637
rect 405142 240585 405194 240637
rect 219670 240511 219722 240563
rect 249814 240511 249866 240563
rect 250198 240511 250250 240563
rect 346294 240511 346346 240563
rect 365974 240511 366026 240563
rect 406102 240511 406154 240563
rect 674710 240511 674762 240563
rect 675478 240511 675530 240563
rect 220438 240437 220490 240489
rect 233398 240437 233450 240489
rect 41782 240363 41834 240415
rect 220630 240363 220682 240415
rect 248086 240437 248138 240489
rect 248374 240437 248426 240489
rect 350230 240437 350282 240489
rect 366742 240437 366794 240489
rect 407830 240437 407882 240489
rect 607606 240437 607658 240489
rect 627766 240437 627818 240489
rect 240886 240363 240938 240415
rect 257686 240363 257738 240415
rect 275350 240363 275402 240415
rect 281110 240363 281162 240415
rect 281398 240363 281450 240415
rect 218806 240289 218858 240341
rect 237718 240289 237770 240341
rect 238966 240289 239018 240341
rect 255478 240289 255530 240341
rect 236566 240215 236618 240267
rect 218422 240141 218474 240193
rect 237814 240141 237866 240193
rect 238870 240215 238922 240267
rect 264406 240289 264458 240341
rect 274006 240289 274058 240341
rect 262006 240215 262058 240267
rect 278230 240215 278282 240267
rect 263926 240141 263978 240193
rect 264022 240141 264074 240193
rect 277654 240141 277706 240193
rect 277750 240141 277802 240193
rect 285622 240215 285674 240267
rect 279478 240141 279530 240193
rect 282166 240141 282218 240193
rect 286870 240363 286922 240415
rect 297046 240289 297098 240341
rect 315574 240363 315626 240415
rect 375094 240363 375146 240415
rect 378262 240363 378314 240415
rect 408310 240363 408362 240415
rect 313174 240289 313226 240341
rect 313654 240289 313706 240341
rect 371830 240289 371882 240341
rect 377782 240289 377834 240341
rect 406678 240289 406730 240341
rect 287446 240215 287498 240267
rect 287830 240215 287882 240267
rect 287926 240215 287978 240267
rect 312598 240215 312650 240267
rect 314614 240215 314666 240267
rect 373558 240215 373610 240267
rect 377206 240215 377258 240267
rect 405526 240215 405578 240267
rect 290710 240141 290762 240193
rect 290806 240141 290858 240193
rect 295414 240141 295466 240193
rect 298198 240141 298250 240193
rect 316054 240141 316106 240193
rect 316150 240141 316202 240193
rect 371350 240141 371402 240193
rect 376438 240141 376490 240193
rect 404086 240141 404138 240193
rect 221782 240067 221834 240119
rect 237526 240067 237578 240119
rect 237910 240067 237962 240119
rect 261622 240067 261674 240119
rect 277462 240067 277514 240119
rect 232342 239993 232394 240045
rect 238198 239993 238250 240045
rect 238294 239993 238346 240045
rect 260662 239993 260714 240045
rect 260758 239993 260810 240045
rect 271894 239993 271946 240045
rect 274678 239993 274730 240045
rect 287350 239993 287402 240045
rect 223222 239919 223274 239971
rect 232150 239919 232202 239971
rect 244630 239919 244682 239971
rect 246070 239919 246122 239971
rect 249718 239919 249770 239971
rect 257878 239919 257930 239971
rect 268726 239919 268778 239971
rect 280150 239919 280202 239971
rect 280246 239919 280298 239971
rect 287830 240067 287882 240119
rect 306646 240067 306698 240119
rect 314230 240067 314282 240119
rect 372406 240067 372458 240119
rect 377014 240067 377066 240119
rect 404950 240067 405002 240119
rect 287638 239993 287690 240045
rect 289462 239993 289514 240045
rect 290518 239993 290570 240045
rect 293398 239993 293450 240045
rect 295702 239993 295754 240045
rect 329110 239993 329162 240045
rect 330070 239993 330122 240045
rect 356566 239993 356618 240045
rect 381814 239993 381866 240045
rect 389878 239993 389930 240045
rect 227158 239845 227210 239897
rect 230326 239845 230378 239897
rect 256438 239845 256490 239897
rect 274102 239845 274154 239897
rect 274198 239845 274250 239897
rect 281494 239845 281546 239897
rect 295606 239919 295658 239971
rect 296086 239919 296138 239971
rect 303670 239919 303722 239971
rect 307798 239919 307850 239971
rect 309814 239919 309866 239971
rect 313750 239919 313802 239971
rect 316150 239919 316202 239971
rect 257206 239771 257258 239823
rect 269302 239771 269354 239823
rect 269398 239771 269450 239823
rect 276310 239771 276362 239823
rect 276694 239771 276746 239823
rect 284470 239771 284522 239823
rect 289462 239845 289514 239897
rect 296662 239845 296714 239897
rect 311638 239845 311690 239897
rect 331702 239919 331754 239971
rect 334486 239919 334538 239971
rect 365878 239919 365930 239971
rect 377878 239919 377930 239971
rect 407542 239919 407594 239971
rect 317782 239845 317834 239897
rect 327958 239845 328010 239897
rect 328246 239845 328298 239897
rect 352438 239845 352490 239897
rect 378646 239845 378698 239897
rect 383830 239845 383882 239897
rect 291670 239771 291722 239823
rect 294454 239771 294506 239823
rect 298198 239771 298250 239823
rect 301846 239771 301898 239823
rect 306646 239771 306698 239823
rect 307894 239771 307946 239823
rect 312118 239771 312170 239823
rect 315190 239771 315242 239823
rect 325270 239771 325322 239823
rect 326230 239771 326282 239823
rect 347926 239771 347978 239823
rect 380566 239771 380618 239823
rect 384886 239771 384938 239823
rect 214486 239697 214538 239749
rect 225142 239697 225194 239749
rect 228022 239697 228074 239749
rect 229942 239697 229994 239749
rect 248566 239697 248618 239749
rect 260758 239697 260810 239749
rect 268246 239697 268298 239749
rect 270934 239697 270986 239749
rect 276214 239697 276266 239749
rect 280534 239697 280586 239749
rect 291382 239697 291434 239749
rect 294742 239697 294794 239749
rect 322678 239697 322730 239749
rect 229078 239623 229130 239675
rect 230230 239623 230282 239675
rect 270262 239623 270314 239675
rect 272278 239623 272330 239675
rect 271798 239549 271850 239601
rect 277750 239623 277802 239675
rect 278038 239623 278090 239675
rect 281782 239623 281834 239675
rect 282166 239623 282218 239675
rect 291190 239623 291242 239675
rect 291478 239623 291530 239675
rect 277654 239549 277706 239601
rect 282934 239549 282986 239601
rect 283030 239549 283082 239601
rect 291382 239549 291434 239601
rect 293206 239623 293258 239675
rect 302806 239623 302858 239675
rect 302998 239623 303050 239675
rect 307606 239623 307658 239675
rect 309526 239623 309578 239675
rect 310294 239623 310346 239675
rect 320854 239623 320906 239675
rect 324694 239623 324746 239675
rect 326998 239697 327050 239749
rect 349558 239697 349610 239749
rect 374806 239697 374858 239749
rect 382678 239697 382730 239749
rect 340918 239623 340970 239675
rect 373846 239623 373898 239675
rect 383542 239697 383594 239749
rect 383638 239697 383690 239749
rect 385558 239697 385610 239749
rect 383158 239623 383210 239675
rect 388150 239623 388202 239675
rect 301846 239549 301898 239601
rect 302518 239549 302570 239601
rect 307222 239549 307274 239601
rect 308854 239549 308906 239601
rect 310198 239549 310250 239601
rect 323062 239549 323114 239601
rect 341302 239549 341354 239601
rect 380086 239549 380138 239601
rect 383734 239549 383786 239601
rect 277078 239475 277130 239527
rect 283798 239475 283850 239527
rect 283894 239475 283946 239527
rect 292150 239475 292202 239527
rect 297814 239475 297866 239527
rect 305014 239475 305066 239527
rect 327382 239475 327434 239527
rect 332950 239475 333002 239527
rect 380854 239475 380906 239527
rect 383062 239475 383114 239527
rect 237142 239401 237194 239453
rect 241846 239401 241898 239453
rect 276214 239401 276266 239453
rect 286006 239401 286058 239453
rect 235510 239327 235562 239379
rect 238678 239327 238730 239379
rect 272470 239327 272522 239379
rect 285526 239327 285578 239379
rect 285622 239327 285674 239379
rect 290806 239401 290858 239453
rect 290902 239401 290954 239453
rect 293302 239401 293354 239453
rect 293398 239401 293450 239453
rect 294454 239401 294506 239453
rect 295990 239401 296042 239453
rect 304150 239401 304202 239453
rect 323446 239401 323498 239453
rect 341974 239401 342026 239453
rect 380086 239401 380138 239453
rect 386614 239475 386666 239527
rect 294262 239327 294314 239379
rect 303574 239327 303626 239379
rect 303670 239327 303722 239379
rect 314806 239327 314858 239379
rect 322198 239327 322250 239379
rect 338902 239327 338954 239379
rect 275734 239253 275786 239305
rect 283030 239253 283082 239305
rect 42550 239179 42602 239231
rect 42454 238883 42506 238935
rect 139990 239179 140042 239231
rect 152470 239179 152522 239231
rect 215926 239179 215978 239231
rect 218902 239179 218954 239231
rect 273430 239179 273482 239231
rect 278806 239179 278858 239231
rect 278902 239179 278954 239231
rect 279670 239179 279722 239231
rect 280438 239179 280490 239231
rect 284086 239253 284138 239305
rect 287350 239253 287402 239305
rect 294358 239253 294410 239305
rect 326614 239253 326666 239305
rect 348982 239253 349034 239305
rect 238486 239105 238538 239157
rect 241654 239105 241706 239157
rect 272662 239105 272714 239157
rect 290902 239179 290954 239231
rect 291286 239179 291338 239231
rect 296566 239179 296618 239231
rect 296662 239179 296714 239231
rect 313846 239179 313898 239231
rect 321238 239179 321290 239231
rect 337174 239179 337226 239231
rect 360982 239179 361034 239231
rect 395830 239327 395882 239379
rect 258646 239031 258698 239083
rect 258934 239031 258986 239083
rect 228118 238957 228170 239009
rect 231958 238957 232010 239009
rect 240118 238957 240170 239009
rect 256822 238957 256874 239009
rect 260374 238957 260426 239009
rect 282262 239031 282314 239083
rect 287062 239105 287114 239157
rect 284086 239031 284138 239083
rect 290806 239031 290858 239083
rect 318262 239105 318314 239157
rect 332758 239105 332810 239157
rect 360214 239105 360266 239157
rect 392086 239253 392138 239305
rect 375670 239179 375722 239231
rect 402358 239179 402410 239231
rect 375190 239105 375242 239157
rect 400630 239105 400682 239157
rect 300022 239031 300074 239083
rect 324406 239031 324458 239083
rect 343702 239031 343754 239083
rect 373366 239031 373418 239083
rect 396886 239031 396938 239083
rect 278422 238957 278474 239009
rect 279382 238957 279434 239009
rect 279478 238957 279530 239009
rect 292246 238957 292298 239009
rect 293974 238957 294026 239009
rect 303190 238957 303242 239009
rect 304726 238957 304778 239009
rect 308182 238957 308234 239009
rect 311638 238957 311690 239009
rect 323638 238957 323690 239009
rect 227734 238883 227786 238935
rect 232822 238883 232874 238935
rect 240502 238883 240554 238935
rect 255670 238883 255722 238935
rect 259990 238883 260042 238935
rect 275254 238883 275306 238935
rect 281686 238883 281738 238935
rect 297430 238883 297482 238935
rect 299062 238883 299114 238935
rect 305782 238883 305834 238935
rect 318550 238883 318602 238935
rect 331318 238957 331370 239009
rect 351094 238957 351146 239009
rect 379030 238957 379082 239009
rect 380470 238957 380522 239009
rect 383158 238957 383210 239009
rect 256822 238809 256874 238861
rect 316246 238809 316298 238861
rect 317398 238809 317450 238861
rect 323734 238809 323786 238861
rect 224566 238735 224618 238787
rect 239446 238735 239498 238787
rect 239542 238735 239594 238787
rect 257398 238735 257450 238787
rect 257782 238735 257834 238787
rect 318166 238735 318218 238787
rect 348406 238883 348458 238935
rect 348502 238883 348554 238935
rect 377302 238883 377354 238935
rect 323926 238809 323978 238861
rect 351094 238809 351146 238861
rect 351190 238809 351242 238861
rect 358774 238809 358826 238861
rect 366838 238809 366890 238861
rect 383350 238809 383402 238861
rect 226294 238661 226346 238713
rect 235606 238661 235658 238713
rect 256246 238661 256298 238713
rect 318262 238661 318314 238713
rect 227254 238587 227306 238639
rect 234070 238587 234122 238639
rect 248950 238587 249002 238639
rect 316342 238587 316394 238639
rect 316438 238587 316490 238639
rect 324214 238735 324266 238787
rect 328822 238735 328874 238787
rect 330646 238735 330698 238787
rect 357238 238735 357290 238787
rect 381430 238735 381482 238787
rect 389206 238735 389258 238787
rect 318646 238661 318698 238713
rect 332182 238661 332234 238713
rect 334102 238661 334154 238713
rect 365302 238661 365354 238713
rect 383158 238661 383210 238713
rect 387574 238661 387626 238713
rect 319030 238587 319082 238639
rect 332374 238587 332426 238639
rect 333622 238587 333674 238639
rect 363286 238587 363338 238639
rect 370390 238587 370442 238639
rect 390358 238587 390410 238639
rect 42166 238513 42218 238565
rect 43030 238513 43082 238565
rect 217078 238513 217130 238565
rect 255190 238513 255242 238565
rect 255574 238513 255626 238565
rect 318070 238513 318122 238565
rect 319606 238513 319658 238565
rect 333430 238513 333482 238565
rect 334870 238513 334922 238565
rect 226870 238439 226922 238491
rect 235030 238439 235082 238491
rect 254134 238439 254186 238491
rect 330934 238439 330986 238491
rect 331126 238439 331178 238491
rect 351190 238439 351242 238491
rect 360886 238513 360938 238565
rect 378358 238513 378410 238565
rect 383062 238513 383114 238565
rect 391414 238513 391466 238565
rect 367030 238439 367082 238491
rect 368470 238439 368522 238491
rect 385942 238439 385994 238491
rect 254614 238365 254666 238417
rect 336982 238365 337034 238417
rect 351382 238365 351434 238417
rect 358870 238365 358922 238417
rect 369430 238365 369482 238417
rect 388822 238365 388874 238417
rect 218038 238291 218090 238343
rect 253462 238291 253514 238343
rect 258550 238291 258602 238343
rect 279478 238291 279530 238343
rect 288118 238291 288170 238343
rect 293686 238291 293738 238343
rect 293782 238291 293834 238343
rect 385270 238291 385322 238343
rect 253366 238217 253418 238269
rect 252406 238143 252458 238195
rect 330934 238217 330986 238269
rect 338710 238217 338762 238269
rect 371638 238217 371690 238269
rect 393622 238217 393674 238269
rect 223222 238069 223274 238121
rect 242614 238069 242666 238121
rect 251926 238069 251978 238121
rect 340438 238143 340490 238195
rect 369814 238143 369866 238195
rect 389686 238143 389738 238195
rect 221878 237995 221930 238047
rect 244822 237995 244874 238047
rect 251158 237995 251210 238047
rect 330550 237995 330602 238047
rect 341494 238069 341546 238121
rect 342742 238069 342794 238121
rect 370006 238069 370058 238121
rect 371158 238069 371210 238121
rect 391894 238069 391946 238121
rect 343510 237995 343562 238047
rect 372022 237995 372074 238047
rect 394198 237995 394250 238047
rect 223318 237921 223370 237973
rect 242134 237921 242186 237973
rect 249814 237921 249866 237973
rect 328438 237921 328490 237973
rect 328534 237921 328586 237973
rect 338230 237921 338282 237973
rect 371254 237921 371306 237973
rect 392470 237921 392522 237973
rect 42166 237847 42218 237899
rect 47542 237847 47594 237899
rect 222838 237847 222890 237899
rect 243766 237847 243818 237899
rect 249334 237847 249386 237899
rect 349174 237847 349226 237899
rect 359830 237847 359882 237899
rect 380950 237847 381002 237899
rect 383062 237847 383114 237899
rect 384406 237847 384458 237899
rect 384502 237847 384554 237899
rect 410998 237847 411050 237899
rect 223702 237773 223754 237825
rect 241558 237773 241610 237825
rect 247126 237773 247178 237825
rect 353974 237773 354026 237825
rect 375574 237773 375626 237825
rect 401206 237773 401258 237825
rect 228502 237699 228554 237751
rect 230806 237699 230858 237751
rect 247606 237699 247658 237751
rect 351958 237699 352010 237751
rect 384406 237699 384458 237751
rect 410614 237699 410666 237751
rect 549238 237699 549290 237751
rect 649366 237699 649418 237751
rect 221494 237625 221546 237677
rect 245878 237625 245930 237677
rect 246166 237625 246218 237677
rect 355030 237625 355082 237677
rect 373462 237625 373514 237677
rect 397942 237625 397994 237677
rect 497494 237625 497546 237677
rect 602902 237625 602954 237677
rect 148342 237551 148394 237603
rect 207190 237551 207242 237603
rect 221974 237551 222026 237603
rect 245782 237551 245834 237603
rect 356182 237551 356234 237603
rect 374230 237551 374282 237603
rect 399670 237551 399722 237603
rect 420598 237551 420650 237603
rect 607606 237551 607658 237603
rect 239062 237477 239114 237529
rect 259126 237477 259178 237529
rect 275254 237477 275306 237529
rect 291958 237477 292010 237529
rect 292054 237477 292106 237529
rect 302422 237477 302474 237529
rect 304054 237477 304106 237529
rect 307990 237477 308042 237529
rect 319990 237477 320042 237529
rect 334390 237477 334442 237529
rect 227350 237403 227402 237455
rect 233590 237403 233642 237455
rect 238774 237403 238826 237455
rect 259414 237403 259466 237455
rect 275446 237403 275498 237455
rect 287158 237403 287210 237455
rect 287254 237403 287306 237455
rect 287926 237403 287978 237455
rect 221014 237329 221066 237381
rect 247222 237329 247274 237381
rect 273238 237329 273290 237381
rect 292534 237403 292586 237455
rect 295318 237403 295370 237455
rect 303670 237403 303722 237455
rect 316054 237403 316106 237455
rect 338518 237477 338570 237529
rect 342742 237477 342794 237529
rect 376630 237477 376682 237529
rect 376726 237477 376778 237529
rect 384598 237477 384650 237529
rect 372598 237403 372650 237455
rect 395350 237403 395402 237455
rect 290326 237329 290378 237381
rect 301462 237329 301514 237381
rect 316822 237329 316874 237381
rect 338518 237329 338570 237381
rect 342838 237329 342890 237381
rect 360886 237329 360938 237381
rect 369046 237329 369098 237381
rect 387670 237329 387722 237381
rect 221110 237255 221162 237307
rect 246550 237255 246602 237307
rect 275830 237255 275882 237307
rect 286582 237255 286634 237307
rect 274006 237181 274058 237233
rect 290614 237255 290666 237307
rect 290710 237255 290762 237307
rect 293974 237255 294026 237307
rect 294070 237255 294122 237307
rect 296470 237255 296522 237307
rect 300214 237255 300266 237307
rect 305878 237255 305930 237307
rect 305974 237255 306026 237307
rect 318454 237255 318506 237307
rect 321814 237255 321866 237307
rect 328534 237255 328586 237307
rect 328726 237255 328778 237307
rect 330742 237255 330794 237307
rect 331798 237255 331850 237307
rect 344758 237255 344810 237307
rect 379990 237255 380042 237307
rect 385366 237255 385418 237307
rect 289270 237181 289322 237233
rect 300982 237181 301034 237233
rect 318166 237181 318218 237233
rect 330838 237181 330890 237233
rect 332854 237181 332906 237233
rect 362230 237181 362282 237233
rect 362806 237181 362858 237233
rect 382294 237181 382346 237233
rect 225526 237107 225578 237159
rect 237334 237107 237386 237159
rect 278518 237107 278570 237159
rect 280726 237107 280778 237159
rect 285814 237107 285866 237159
rect 286390 237033 286442 237085
rect 288406 237107 288458 237159
rect 300598 237107 300650 237159
rect 316246 237107 316298 237159
rect 324118 237107 324170 237159
rect 327862 237107 327914 237159
rect 351478 237107 351530 237159
rect 351574 237107 351626 237159
rect 358774 237107 358826 237159
rect 372982 237107 373034 237159
rect 396214 237107 396266 237159
rect 224086 236959 224138 237011
rect 240406 236959 240458 237011
rect 271894 236959 271946 237011
rect 288118 236959 288170 237011
rect 299542 237033 299594 237085
rect 318262 237033 318314 237085
rect 328726 237033 328778 237085
rect 328822 237033 328874 237085
rect 353494 237033 353546 237085
rect 276790 236885 276842 236937
rect 295222 236885 295274 236937
rect 296854 236959 296906 237011
rect 304438 236959 304490 237011
rect 299638 236885 299690 236937
rect 225046 236811 225098 236863
rect 238582 236811 238634 236863
rect 282742 236811 282794 236863
rect 285238 236811 285290 236863
rect 285910 236811 285962 236863
rect 288982 236811 289034 236863
rect 291766 236811 291818 236863
rect 316342 236959 316394 237011
rect 325846 236959 325898 237011
rect 327478 236959 327530 237011
rect 350710 236959 350762 237011
rect 319318 236885 319370 236937
rect 327094 236885 327146 236937
rect 349750 236885 349802 236937
rect 324790 236811 324842 236863
rect 331798 236811 331850 236863
rect 331894 236811 331946 236863
rect 339670 236811 339722 236863
rect 370774 236811 370826 236863
rect 381142 236811 381194 236863
rect 239062 236737 239114 236789
rect 259126 236737 259178 236789
rect 274870 236737 274922 236789
rect 288502 236737 288554 236789
rect 291670 236737 291722 236789
rect 305974 236737 306026 236789
rect 306454 236737 306506 236789
rect 308950 236737 309002 236789
rect 325654 236737 325706 236789
rect 330454 236737 330506 236789
rect 330550 236737 330602 236789
rect 345238 236737 345290 236789
rect 42166 236663 42218 236715
rect 42358 236663 42410 236715
rect 260758 236663 260810 236715
rect 269494 236663 269546 236715
rect 274102 236663 274154 236715
rect 289750 236663 289802 236715
rect 293494 236663 293546 236715
rect 299734 236663 299786 236715
rect 236470 236589 236522 236641
rect 238870 236589 238922 236641
rect 276406 236589 276458 236641
rect 294838 236589 294890 236641
rect 295798 236589 295850 236641
rect 315382 236663 315434 236715
rect 324022 236663 324074 236715
rect 313654 236589 313706 236641
rect 313846 236589 313898 236641
rect 325270 236589 325322 236641
rect 328342 236589 328394 236641
rect 328534 236663 328586 236715
rect 347446 236663 347498 236715
rect 380182 236663 380234 236715
rect 390166 236663 390218 236715
rect 420502 236663 420554 236715
rect 440566 236663 440618 236715
rect 460822 236663 460874 236715
rect 480886 236663 480938 236715
rect 343030 236589 343082 236641
rect 258166 236515 258218 236567
rect 264022 236515 264074 236567
rect 278710 236515 278762 236567
rect 268342 236441 268394 236493
rect 217462 236367 217514 236419
rect 221782 236367 221834 236419
rect 263062 236367 263114 236419
rect 269014 236367 269066 236419
rect 278422 236367 278474 236419
rect 281206 236367 281258 236419
rect 273526 236293 273578 236345
rect 281590 236293 281642 236345
rect 283318 236293 283370 236345
rect 285046 236293 285098 236345
rect 285238 236367 285290 236419
rect 289270 236515 289322 236567
rect 311446 236515 311498 236567
rect 318070 236515 318122 236567
rect 335638 236515 335690 236567
rect 638038 236515 638090 236567
rect 650518 236515 650570 236567
rect 291286 236441 291338 236493
rect 317590 236441 317642 236493
rect 320374 236441 320426 236493
rect 334966 236441 335018 236493
rect 637558 236441 637610 236493
rect 650230 236441 650282 236493
rect 288118 236293 288170 236345
rect 296182 236367 296234 236419
rect 300790 236367 300842 236419
rect 306262 236367 306314 236419
rect 322486 236367 322538 236419
rect 339862 236367 339914 236419
rect 637942 236367 637994 236419
rect 650326 236367 650378 236419
rect 297814 236293 297866 236345
rect 330454 236293 330506 236345
rect 346966 236293 347018 236345
rect 639190 236293 639242 236345
rect 649846 236293 649898 236345
rect 144022 236219 144074 236271
rect 168406 236219 168458 236271
rect 225910 236219 225962 236271
rect 236758 236219 236810 236271
rect 236950 236219 237002 236271
rect 238966 236219 239018 236271
rect 271414 236219 271466 236271
rect 290710 236219 290762 236271
rect 290806 236219 290858 236271
rect 296950 236219 297002 236271
rect 328342 236219 328394 236271
rect 345910 236219 345962 236271
rect 368950 236219 369002 236271
rect 387094 236219 387146 236271
rect 638806 236219 638858 236271
rect 649654 236219 649706 236271
rect 144118 236145 144170 236197
rect 174166 236145 174218 236197
rect 210262 236145 210314 236197
rect 210742 236145 210794 236197
rect 213046 236145 213098 236197
rect 284374 236145 284426 236197
rect 298774 236145 298826 236197
rect 315958 236145 316010 236197
rect 324214 236145 324266 236197
rect 547126 236145 547178 236197
rect 549238 236145 549290 236197
rect 639766 236145 639818 236197
rect 649942 236145 649994 236197
rect 265654 236071 265706 236123
rect 308374 236071 308426 236123
rect 319702 236071 319754 236123
rect 339766 236071 339818 236123
rect 264886 235997 264938 236049
rect 309910 235997 309962 236049
rect 312982 235997 313034 236049
rect 369622 235997 369674 236049
rect 265078 235923 265130 235975
rect 339382 235923 339434 235975
rect 381910 235923 381962 235975
rect 390934 235923 390986 235975
rect 235702 235849 235754 235901
rect 266134 235849 266186 235901
rect 266806 235849 266858 235901
rect 340342 235849 340394 235901
rect 263734 235775 263786 235827
rect 338902 235775 338954 235827
rect 261910 235701 261962 235753
rect 338134 235701 338186 235753
rect 258934 235627 258986 235679
rect 336694 235627 336746 235679
rect 260566 235553 260618 235605
rect 337174 235553 337226 235605
rect 257302 235479 257354 235531
rect 335926 235479 335978 235531
rect 42166 235405 42218 235457
rect 43126 235405 43178 235457
rect 236086 235405 236138 235457
rect 265462 235405 265514 235457
rect 273622 235405 273674 235457
rect 356662 235405 356714 235457
rect 246070 235331 246122 235383
rect 353590 235331 353642 235383
rect 247798 235257 247850 235309
rect 354838 235257 354890 235309
rect 246358 235183 246410 235235
rect 354358 235183 354410 235235
rect 242038 235109 242090 235161
rect 352150 235109 352202 235161
rect 241846 235035 241898 235087
rect 349942 235035 349994 235087
rect 243286 234961 243338 235013
rect 352630 234961 352682 235013
rect 244150 234887 244202 234939
rect 351382 234887 351434 234939
rect 42166 234813 42218 234865
rect 42934 234813 42986 234865
rect 241654 234813 241706 234865
rect 350422 234813 350474 234865
rect 230614 234739 230666 234791
rect 346966 234739 347018 234791
rect 227926 234665 227978 234717
rect 345526 234665 345578 234717
rect 260854 234591 260906 234643
rect 268438 234591 268490 234643
rect 282454 234591 282506 234643
rect 322774 234591 322826 234643
rect 266998 234517 267050 234569
rect 305686 234517 305738 234569
rect 282838 234443 282890 234495
rect 321910 234443 321962 234495
rect 267478 234369 267530 234421
rect 304246 234369 304298 234421
rect 271606 234295 271658 234347
rect 309430 234295 309482 234347
rect 284662 234221 284714 234273
rect 317974 234221 318026 234273
rect 42070 234147 42122 234199
rect 42454 234147 42506 234199
rect 277270 234147 277322 234199
rect 279766 234147 279818 234199
rect 284278 234147 284330 234199
rect 319126 234147 319178 234199
rect 268822 234073 268874 234125
rect 301942 234073 301994 234125
rect 269590 233999 269642 234051
rect 300310 233999 300362 234051
rect 285142 233925 285194 233977
rect 316534 233925 316586 233977
rect 287350 233851 287402 233903
rect 289270 233851 289322 233903
rect 292534 233851 292586 233903
rect 320566 233851 320618 233903
rect 285046 233777 285098 233829
rect 288214 233777 288266 233829
rect 293110 233777 293162 233829
rect 321430 233777 321482 233829
rect 262342 233703 262394 233755
rect 268918 233703 268970 233755
rect 270070 233703 270122 233755
rect 298582 233703 298634 233755
rect 305590 233703 305642 233755
rect 308710 233703 308762 233755
rect 367942 233703 367994 233755
rect 376726 233703 376778 233755
rect 270646 233629 270698 233681
rect 298486 233629 298538 233681
rect 208150 233555 208202 233607
rect 213526 233555 213578 233607
rect 269110 233555 269162 233607
rect 297046 233555 297098 233607
rect 209974 233481 210026 233533
rect 213142 233481 213194 233533
rect 213910 233481 213962 233533
rect 290902 233481 290954 233533
rect 317014 233629 317066 233681
rect 210070 233407 210122 233459
rect 144022 233259 144074 233311
rect 171286 233259 171338 233311
rect 645526 233185 645578 233237
rect 649750 233185 649802 233237
rect 645238 233111 645290 233163
rect 650422 233111 650474 233163
rect 645334 232963 645386 233015
rect 650134 232963 650186 233015
rect 645142 232889 645194 232941
rect 650614 232889 650666 232941
rect 144022 230521 144074 230573
rect 151126 230521 151178 230573
rect 144118 230447 144170 230499
rect 165526 230447 165578 230499
rect 205750 228153 205802 228205
rect 205942 228153 205994 228205
rect 205270 227857 205322 227909
rect 205654 227857 205706 227909
rect 210262 227783 210314 227835
rect 144022 227709 144074 227761
rect 188566 227709 188618 227761
rect 144118 227635 144170 227687
rect 194326 227635 194378 227687
rect 144214 227561 144266 227613
rect 197206 227561 197258 227613
rect 210262 227561 210314 227613
rect 146806 226377 146858 226429
rect 156886 226377 156938 226429
rect 206614 226377 206666 226429
rect 206326 226229 206378 226281
rect 206614 226229 206666 226281
rect 205846 226155 205898 226207
rect 207094 226155 207146 226207
rect 206038 226081 206090 226133
rect 206326 226081 206378 226133
rect 205846 225933 205898 225985
rect 666838 225045 666890 225097
rect 674710 225045 674762 225097
rect 146134 224675 146186 224727
rect 200086 224675 200138 224727
rect 141046 224601 141098 224653
rect 204502 224601 204554 224653
rect 146422 224527 146474 224579
rect 204598 224527 204650 224579
rect 149686 224453 149738 224505
rect 204694 224453 204746 224505
rect 152566 224379 152618 224431
rect 204790 224379 204842 224431
rect 669526 224305 669578 224357
rect 674422 224305 674474 224357
rect 669622 224009 669674 224061
rect 674710 224009 674762 224061
rect 146710 221937 146762 221989
rect 177046 221937 177098 221989
rect 146806 221863 146858 221915
rect 179926 221863 179978 221915
rect 144406 221789 144458 221841
rect 182902 221789 182954 221841
rect 155446 221715 155498 221767
rect 204502 221715 204554 221767
rect 161206 221641 161258 221693
rect 204598 221641 204650 221693
rect 164086 221567 164138 221619
rect 204694 221567 204746 221619
rect 166966 221493 167018 221545
rect 204790 221493 204842 221545
rect 169846 221419 169898 221471
rect 204886 221419 204938 221471
rect 144406 218903 144458 218955
rect 174262 218903 174314 218955
rect 175606 218829 175658 218881
rect 204502 218829 204554 218881
rect 178486 218755 178538 218807
rect 204598 218755 204650 218807
rect 181366 218681 181418 218733
rect 204694 218681 204746 218733
rect 184246 218607 184298 218659
rect 204790 218607 204842 218659
rect 146806 216535 146858 216587
rect 154006 216535 154058 216587
rect 42742 216313 42794 216365
rect 44950 216313 45002 216365
rect 146230 216091 146282 216143
rect 146326 216017 146378 216069
rect 187126 215943 187178 215995
rect 204502 215943 204554 215995
rect 192886 215869 192938 215921
rect 204598 215869 204650 215921
rect 42742 215721 42794 215773
rect 45142 215721 45194 215773
rect 42742 215203 42794 215255
rect 44854 215203 44906 215255
rect 146806 213205 146858 213257
rect 168502 213205 168554 213257
rect 144406 213131 144458 213183
rect 171382 213131 171434 213183
rect 145270 210245 145322 210297
rect 148246 210245 148298 210297
rect 645622 210245 645674 210297
rect 677014 210245 677066 210297
rect 146614 207433 146666 207485
rect 165622 207433 165674 207485
rect 146806 207359 146858 207411
rect 203062 207359 203114 207411
rect 40246 206767 40298 206819
rect 41782 206767 41834 206819
rect 675478 205953 675530 206005
rect 675478 205731 675530 205783
rect 675190 204991 675242 205043
rect 675478 204991 675530 205043
rect 42742 204399 42794 204451
rect 50326 204399 50378 204451
rect 674902 204399 674954 204451
rect 675382 204399 675434 204451
rect 674998 202179 675050 202231
rect 675286 202179 675338 202231
rect 675094 202031 675146 202083
rect 675286 202031 675338 202083
rect 145846 201661 145898 201713
rect 162646 201661 162698 201713
rect 144022 201587 144074 201639
rect 202966 201587 203018 201639
rect 645910 201587 645962 201639
rect 646102 201587 646154 201639
rect 674230 201291 674282 201343
rect 675382 201291 675434 201343
rect 41974 201069 42026 201121
rect 42358 201069 42410 201121
rect 674806 200329 674858 200381
rect 675286 200329 675338 200381
rect 40150 198997 40202 199049
rect 42166 198997 42218 199049
rect 144022 198923 144074 198975
rect 159766 198923 159818 198975
rect 40054 198849 40106 198901
rect 43126 198849 43178 198901
rect 40246 198701 40298 198753
rect 43126 198701 43178 198753
rect 144502 198701 144554 198753
rect 191446 198701 191498 198753
rect 674710 197739 674762 197791
rect 675382 197739 675434 197791
rect 41782 197369 41834 197421
rect 145078 197221 145130 197273
rect 146230 197221 146282 197273
rect 41782 197147 41834 197199
rect 674518 196999 674570 197051
rect 675478 196999 675530 197051
rect 674614 196555 674666 196607
rect 675382 196555 675434 196607
rect 144694 195815 144746 195867
rect 185686 195815 185738 195867
rect 42166 195297 42218 195349
rect 42358 195297 42410 195349
rect 42070 194483 42122 194535
rect 50422 194483 50474 194535
rect 42070 193447 42122 193499
rect 42934 193447 42986 193499
rect 42934 193299 42986 193351
rect 43222 193299 43274 193351
rect 42166 192189 42218 192241
rect 43030 192189 43082 192241
rect 42070 191449 42122 191501
rect 42358 191449 42410 191501
rect 42166 191005 42218 191057
rect 43126 191005 43178 191057
rect 144310 190191 144362 190243
rect 151222 190191 151274 190243
rect 144022 190117 144074 190169
rect 148438 190117 148490 190169
rect 42262 187897 42314 187949
rect 42934 187897 42986 187949
rect 210262 187379 210314 187431
rect 144022 187231 144074 187283
rect 197302 187231 197354 187283
rect 42166 187083 42218 187135
rect 42838 187083 42890 187135
rect 210262 187083 210314 187135
rect 645718 187083 645770 187135
rect 646102 187083 646154 187135
rect 146326 184567 146378 184619
rect 146806 184567 146858 184619
rect 144022 184345 144074 184397
rect 194422 184345 194474 184397
rect 144214 181533 144266 181585
rect 146614 181533 146666 181585
rect 144022 181459 144074 181511
rect 188662 181459 188714 181511
rect 661078 179313 661130 179365
rect 674422 179313 674474 179365
rect 666646 178795 666698 178847
rect 674422 178795 674474 178847
rect 144118 178647 144170 178699
rect 148534 178647 148586 178699
rect 655222 178647 655274 178699
rect 674710 178647 674762 178699
rect 144022 178573 144074 178625
rect 191542 178573 191594 178625
rect 146518 176131 146570 176183
rect 146998 176131 147050 176183
rect 146230 175983 146282 176035
rect 146230 175761 146282 175813
rect 144022 175687 144074 175739
rect 185782 175687 185834 175739
rect 144502 175613 144554 175665
rect 146806 175613 146858 175665
rect 144118 172875 144170 172927
rect 148630 172875 148682 172927
rect 144022 172801 144074 172853
rect 162742 172801 162794 172853
rect 144118 172727 144170 172779
rect 146710 172727 146762 172779
rect 145078 172579 145130 172631
rect 146710 172579 146762 172631
rect 144022 170211 144074 170263
rect 159862 170211 159914 170263
rect 144022 167251 144074 167303
rect 156982 167251 157034 167303
rect 647062 167251 647114 167303
rect 674422 167251 674474 167303
rect 647830 167177 647882 167229
rect 674614 167177 674666 167229
rect 647926 167103 647978 167155
rect 674710 167103 674762 167155
rect 144886 165549 144938 165601
rect 146806 165549 146858 165601
rect 144694 164143 144746 164195
rect 148726 164143 148778 164195
rect 144694 161257 144746 161309
rect 148822 161257 148874 161309
rect 645718 161257 645770 161309
rect 645910 161257 645962 161309
rect 675574 160961 675626 161013
rect 675766 160961 675818 161013
rect 675574 160739 675626 160791
rect 675766 159999 675818 160051
rect 674038 159407 674090 159459
rect 675382 159407 675434 159459
rect 144694 158445 144746 158497
rect 148918 158445 148970 158497
rect 674806 157705 674858 157757
rect 675478 157705 675530 157757
rect 146134 155781 146186 155833
rect 146710 155781 146762 155833
rect 144118 155707 144170 155759
rect 146422 155707 146474 155759
rect 144502 155633 144554 155685
rect 146710 155633 146762 155685
rect 146902 155633 146954 155685
rect 149014 155633 149066 155685
rect 144694 155559 144746 155611
rect 200182 155559 200234 155611
rect 144694 153117 144746 153169
rect 146710 153117 146762 153169
rect 146806 152747 146858 152799
rect 180022 152747 180074 152799
rect 144502 152673 144554 152725
rect 182998 152673 183050 152725
rect 674326 152599 674378 152651
rect 675382 152599 675434 152651
rect 674518 151489 674570 151541
rect 675382 151489 675434 151541
rect 144502 149861 144554 149913
rect 149110 149861 149162 149913
rect 146806 149787 146858 149839
rect 177142 149787 177194 149839
rect 144502 146975 144554 147027
rect 149206 146975 149258 147027
rect 210262 146975 210314 147027
rect 146806 146901 146858 146953
rect 174358 146901 174410 146953
rect 645718 146901 645770 146953
rect 645814 146827 645866 146879
rect 210262 146531 210314 146583
rect 144502 146383 144554 146435
rect 144694 146383 144746 146435
rect 144118 146235 144170 146287
rect 144694 146235 144746 146287
rect 144022 144015 144074 144067
rect 154102 144015 154154 144067
rect 144022 142535 144074 142587
rect 149302 142535 149354 142587
rect 144022 141129 144074 141181
rect 171478 141129 171530 141181
rect 143734 139723 143786 139775
rect 144502 139723 144554 139775
rect 144310 139575 144362 139627
rect 144502 139575 144554 139627
rect 144310 138391 144362 138443
rect 168598 138391 168650 138443
rect 144022 138243 144074 138295
rect 208726 138243 208778 138295
rect 146998 136023 147050 136075
rect 149398 136023 149450 136075
rect 161206 135579 161258 135631
rect 166966 135579 167018 135631
rect 167062 135579 167114 135631
rect 146710 135357 146762 135409
rect 146902 135357 146954 135409
rect 146134 135283 146186 135335
rect 208822 135283 208874 135335
rect 146998 135209 147050 135261
rect 663766 133581 663818 133633
rect 674422 133581 674474 133633
rect 144022 132915 144074 132967
rect 165718 132915 165770 132967
rect 655318 132767 655370 132819
rect 676918 132767 676970 132819
rect 655126 132619 655178 132671
rect 676822 132619 676874 132671
rect 144310 132545 144362 132597
rect 208918 132545 208970 132597
rect 144022 132471 144074 132523
rect 209014 132471 209066 132523
rect 647734 132471 647786 132523
rect 674422 132471 674474 132523
rect 143926 132397 143978 132449
rect 144310 132397 144362 132449
rect 144118 129659 144170 129711
rect 151510 129659 151562 129711
rect 144022 129585 144074 129637
rect 209110 129585 209162 129637
rect 144022 126995 144074 127047
rect 143926 126847 143978 126899
rect 144502 126847 144554 126899
rect 147094 126847 147146 126899
rect 149494 126847 149546 126899
rect 203158 126773 203210 126825
rect 146710 126699 146762 126751
rect 208630 126699 208682 126751
rect 143734 126625 143786 126677
rect 143926 126625 143978 126677
rect 144694 126625 144746 126677
rect 146134 126625 146186 126677
rect 146422 125737 146474 125789
rect 146710 125737 146762 125789
rect 144598 125367 144650 125419
rect 146422 125367 146474 125419
rect 39862 125293 39914 125345
rect 42454 125293 42506 125345
rect 144118 125219 144170 125271
rect 144598 125219 144650 125271
rect 144406 124627 144458 124679
rect 144694 124627 144746 124679
rect 144022 124479 144074 124531
rect 144406 124479 144458 124531
rect 144022 123961 144074 124013
rect 197398 123961 197450 124013
rect 144118 123887 144170 123939
rect 200278 123887 200330 123939
rect 144118 121519 144170 121571
rect 149590 121519 149642 121571
rect 645718 121223 645770 121275
rect 674710 121223 674762 121275
rect 645430 121149 645482 121201
rect 676918 121149 676970 121201
rect 645718 121075 645770 121127
rect 676822 121075 676874 121127
rect 144022 121001 144074 121053
rect 149686 121001 149738 121053
rect 209302 120927 209354 120979
rect 210262 120927 210314 120979
rect 645910 120927 645962 120979
rect 646102 120927 646154 120979
rect 146902 119003 146954 119055
rect 151318 119003 151370 119055
rect 181462 118485 181514 118537
rect 188758 118485 188810 118537
rect 167158 118337 167210 118389
rect 181462 118337 181514 118389
rect 144022 118263 144074 118315
rect 166966 118263 167018 118315
rect 146710 118189 146762 118241
rect 144022 118115 144074 118167
rect 144118 118115 144170 118167
rect 194518 118115 194570 118167
rect 143926 117967 143978 118019
rect 144118 117967 144170 118019
rect 146902 116635 146954 116687
rect 148054 116635 148106 116687
rect 146902 115895 146954 115947
rect 148150 115895 148202 115947
rect 675190 115377 675242 115429
rect 675478 115377 675530 115429
rect 674806 114785 674858 114837
rect 675382 114785 675434 114837
rect 674518 114119 674570 114171
rect 675382 114119 675434 114171
rect 143830 113231 143882 113283
rect 144118 113231 144170 113283
rect 144022 112639 144074 112691
rect 191638 112639 191690 112691
rect 144118 112417 144170 112469
rect 147958 112417 148010 112469
rect 144022 112343 144074 112395
rect 147862 112343 147914 112395
rect 674326 111825 674378 111877
rect 675094 111825 675146 111877
rect 674614 111307 674666 111359
rect 675094 111307 675146 111359
rect 674710 111159 674762 111211
rect 675382 111159 675434 111211
rect 144118 109531 144170 109583
rect 147766 109531 147818 109583
rect 144022 109457 144074 109509
rect 185878 109457 185930 109509
rect 144118 109383 144170 109435
rect 144598 109383 144650 109435
rect 674998 107533 675050 107585
rect 675382 107533 675434 107585
rect 143638 107163 143690 107215
rect 144118 107163 144170 107215
rect 143734 107089 143786 107141
rect 144406 107089 144458 107141
rect 143830 107015 143882 107067
rect 144118 107015 144170 107067
rect 146134 107015 146186 107067
rect 144406 106941 144458 106993
rect 143830 106867 143882 106919
rect 146422 106867 146474 106919
rect 673942 106867 673994 106919
rect 675478 106867 675530 106919
rect 144598 106793 144650 106845
rect 144022 106719 144074 106771
rect 162838 106719 162890 106771
rect 144022 106571 144074 106623
rect 144694 106571 144746 106623
rect 208534 106571 208586 106623
rect 143734 106497 143786 106549
rect 146710 106497 146762 106549
rect 668182 106497 668234 106549
rect 675094 106497 675146 106549
rect 674230 106349 674282 106401
rect 675382 106349 675434 106401
rect 209302 106275 209354 106327
rect 210166 106275 210218 106327
rect 144214 106127 144266 106179
rect 146422 106127 146474 106179
rect 144022 105979 144074 106031
rect 144214 105979 144266 106031
rect 144118 104869 144170 104921
rect 144598 104869 144650 104921
rect 645430 104499 645482 104551
rect 665206 104499 665258 104551
rect 144022 104351 144074 104403
rect 151414 104351 151466 104403
rect 144022 104203 144074 104255
rect 159958 104203 160010 104255
rect 144118 103685 144170 103737
rect 208438 103685 208490 103737
rect 663190 103685 663242 103737
rect 665110 103685 665162 103737
rect 146998 103611 147050 103663
rect 204502 103611 204554 103663
rect 144694 103537 144746 103589
rect 204598 103537 204650 103589
rect 144406 103463 144458 103515
rect 204694 103463 204746 103515
rect 143638 103315 143690 103367
rect 144406 103315 144458 103367
rect 144022 101539 144074 101591
rect 157078 101539 157130 101591
rect 146134 101391 146186 101443
rect 146326 101391 146378 101443
rect 144118 100799 144170 100851
rect 147670 100799 147722 100851
rect 645814 100799 645866 100851
rect 646102 100799 646154 100851
rect 144214 100725 144266 100777
rect 204886 100725 204938 100777
rect 144022 100651 144074 100703
rect 204790 100651 204842 100703
rect 151126 100577 151178 100629
rect 204598 100577 204650 100629
rect 159766 100503 159818 100555
rect 204694 100503 204746 100555
rect 162646 100429 162698 100481
rect 204502 100429 204554 100481
rect 144022 98061 144074 98113
rect 180118 98061 180170 98113
rect 144118 97987 144170 98039
rect 183094 97987 183146 98039
rect 144214 97913 144266 97965
rect 208342 97913 208394 97965
rect 154006 97839 154058 97891
rect 204790 97839 204842 97891
rect 156886 97765 156938 97817
rect 204502 97765 204554 97817
rect 171382 97691 171434 97743
rect 204694 97691 204746 97743
rect 174262 97617 174314 97669
rect 204598 97617 204650 97669
rect 182902 97543 182954 97595
rect 204502 97543 204554 97595
rect 144022 95101 144074 95153
rect 174454 95101 174506 95153
rect 144118 95027 144170 95079
rect 177238 95027 177290 95079
rect 146710 94879 146762 94931
rect 201718 94879 201770 94931
rect 151222 94805 151274 94857
rect 204790 94805 204842 94857
rect 165622 94731 165674 94783
rect 204502 94731 204554 94783
rect 168502 94657 168554 94709
rect 204598 94657 204650 94709
rect 146422 94583 146474 94635
rect 204694 94583 204746 94635
rect 203062 94435 203114 94487
rect 205270 94435 205322 94487
rect 646390 92659 646442 92711
rect 659830 92659 659882 92711
rect 647542 92585 647594 92637
rect 661750 92585 661802 92637
rect 647158 92511 647210 92563
rect 660694 92511 660746 92563
rect 647830 92437 647882 92489
rect 663094 92437 663146 92489
rect 647734 92289 647786 92341
rect 662518 92289 662570 92341
rect 144118 92215 144170 92267
rect 154006 92215 154058 92267
rect 646102 92215 646154 92267
rect 661174 92215 661226 92267
rect 144022 92141 144074 92193
rect 171382 92141 171434 92193
rect 646678 92141 646730 92193
rect 658870 92141 658922 92193
rect 144406 92067 144458 92119
rect 204502 92067 204554 92119
rect 188662 91993 188714 92045
rect 204694 91993 204746 92045
rect 194422 91919 194474 91971
rect 204598 91919 204650 91971
rect 200182 91845 200234 91897
rect 205366 91845 205418 91897
rect 197302 91771 197354 91823
rect 204502 91771 204554 91823
rect 144022 89403 144074 89455
rect 151126 89403 151178 89455
rect 144118 89329 144170 89381
rect 165622 89329 165674 89381
rect 144214 89255 144266 89307
rect 168502 89255 168554 89307
rect 156982 89181 157034 89233
rect 204886 89181 204938 89233
rect 159862 89107 159914 89159
rect 204790 89107 204842 89159
rect 162742 89033 162794 89085
rect 204694 89033 204746 89085
rect 185782 88959 185834 89011
rect 204598 88959 204650 89011
rect 191542 88885 191594 88937
rect 204502 88885 204554 88937
rect 651382 87331 651434 87383
rect 659350 87331 659402 87383
rect 658006 87257 658058 87309
rect 657046 87109 657098 87161
rect 645430 87035 645482 87087
rect 663286 87035 663338 87087
rect 645718 86961 645770 87013
rect 650998 86961 651050 87013
rect 645718 86813 645770 86865
rect 645910 86813 645962 86865
rect 210166 86739 210218 86791
rect 146134 86443 146186 86495
rect 146326 86443 146378 86495
rect 210262 86443 210314 86495
rect 645430 86443 645482 86495
rect 651094 86443 651146 86495
rect 144406 86369 144458 86421
rect 144598 86369 144650 86421
rect 154102 86369 154154 86421
rect 204886 86369 204938 86421
rect 174358 86295 174410 86347
rect 204790 86295 204842 86347
rect 177142 86221 177194 86273
rect 204694 86221 204746 86273
rect 180022 86147 180074 86199
rect 204598 86147 204650 86199
rect 182998 86073 183050 86125
rect 204502 86073 204554 86125
rect 646294 85185 646346 85237
rect 650902 85185 650954 85237
rect 144022 84963 144074 85015
rect 204502 84963 204554 85015
rect 151510 83483 151562 83535
rect 204790 83483 204842 83535
rect 165718 83409 165770 83461
rect 204694 83409 204746 83461
rect 647926 83409 647978 83461
rect 657046 83409 657098 83461
rect 168598 83335 168650 83387
rect 204598 83335 204650 83387
rect 171478 83261 171530 83313
rect 204502 83261 204554 83313
rect 144022 82077 144074 82129
rect 204502 82077 204554 82129
rect 647926 81855 647978 81907
rect 663286 81855 663338 81907
rect 645910 81781 645962 81833
rect 663382 81781 663434 81833
rect 647638 81633 647690 81685
rect 661078 81633 661130 81685
rect 647926 81263 647978 81315
rect 657526 81263 657578 81315
rect 144022 80819 144074 80871
rect 144406 80819 144458 80871
rect 645718 80745 645770 80797
rect 645814 80671 645866 80723
rect 659446 80671 659498 80723
rect 659542 80671 659594 80723
rect 188758 80597 188810 80649
rect 204598 80597 204650 80649
rect 194518 80523 194570 80575
rect 204502 80523 204554 80575
rect 203158 80449 203210 80501
rect 206902 80449 206954 80501
rect 200278 80375 200330 80427
rect 205462 80375 205514 80427
rect 197398 80301 197450 80353
rect 204694 80301 204746 80353
rect 647926 80153 647978 80205
rect 656950 80153 657002 80205
rect 646102 79117 646154 79169
rect 658870 79117 658922 79169
rect 647830 78673 647882 78725
rect 660694 78673 660746 78725
rect 646870 78599 646922 78651
rect 651190 78599 651242 78651
rect 647926 78303 647978 78355
rect 662518 78303 662570 78355
rect 144118 77859 144170 77911
rect 187222 77859 187274 77911
rect 144022 77785 144074 77837
rect 208246 77785 208298 77837
rect 157078 77711 157130 77763
rect 204982 77711 205034 77763
rect 647350 77711 647402 77763
rect 659446 77711 659498 77763
rect 159958 77637 160010 77689
rect 204886 77637 204938 77689
rect 647926 77637 647978 77689
rect 650998 77637 651050 77689
rect 162838 77563 162890 77615
rect 204790 77563 204842 77615
rect 185878 77489 185930 77541
rect 204694 77489 204746 77541
rect 187222 77415 187274 77467
rect 204502 77415 204554 77467
rect 191638 77341 191690 77393
rect 204598 77341 204650 77393
rect 647926 77267 647978 77319
rect 662902 77267 662954 77319
rect 646486 76897 646538 76949
rect 658294 76897 658346 76949
rect 646486 76749 646538 76801
rect 650902 76749 650954 76801
rect 144214 76379 144266 76431
rect 145462 76379 145514 76431
rect 146038 76305 146090 76357
rect 146806 76305 146858 76357
rect 145558 76157 145610 76209
rect 146518 76157 146570 76209
rect 646870 75565 646922 75617
rect 656854 75565 656906 75617
rect 647926 75269 647978 75321
rect 661750 75269 661802 75321
rect 144022 75047 144074 75099
rect 160534 75047 160586 75099
rect 146902 74973 146954 75025
rect 156886 74973 156938 75025
rect 144118 74899 144170 74951
rect 161590 74899 161642 74951
rect 154006 74825 154058 74877
rect 204886 74825 204938 74877
rect 174454 74751 174506 74803
rect 204790 74751 204842 74803
rect 177238 74677 177290 74729
rect 204694 74677 204746 74729
rect 180118 74603 180170 74655
rect 204598 74603 204650 74655
rect 183094 74529 183146 74581
rect 204502 74529 204554 74581
rect 144118 74233 144170 74285
rect 148342 74233 148394 74285
rect 640726 73419 640778 73471
rect 663190 73419 663242 73471
rect 647926 72679 647978 72731
rect 663286 72679 663338 72731
rect 143830 72605 143882 72657
rect 144118 72605 144170 72657
rect 646966 72605 647018 72657
rect 663478 72605 663530 72657
rect 144598 72457 144650 72509
rect 146518 72457 146570 72509
rect 647830 72235 647882 72287
rect 660118 72235 660170 72287
rect 144022 72013 144074 72065
rect 154582 72013 154634 72065
rect 151126 71939 151178 71991
rect 204790 71939 204842 71991
rect 161590 71865 161642 71917
rect 204886 71865 204938 71917
rect 165622 71791 165674 71843
rect 204694 71791 204746 71843
rect 168502 71717 168554 71769
rect 204598 71717 204650 71769
rect 171382 71643 171434 71695
rect 204502 71643 204554 71695
rect 144022 70829 144074 70881
rect 149782 70829 149834 70881
rect 144022 69127 144074 69179
rect 204886 69053 204938 69105
rect 149782 68979 149834 69031
rect 204790 68979 204842 69031
rect 154582 68905 154634 68957
rect 204694 68905 204746 68957
rect 156886 68831 156938 68883
rect 204598 68831 204650 68883
rect 160534 68757 160586 68809
rect 204502 68757 204554 68809
rect 144022 67351 144074 67403
rect 152662 67351 152714 67403
rect 144598 67203 144650 67255
rect 144694 66981 144746 67033
rect 146134 66833 146186 66885
rect 146710 66833 146762 66885
rect 144022 66685 144074 66737
rect 146710 66685 146762 66737
rect 144214 66463 144266 66515
rect 146518 66315 146570 66367
rect 157654 66315 157706 66367
rect 144022 66241 144074 66293
rect 144214 66241 144266 66293
rect 146326 66167 146378 66219
rect 146806 66167 146858 66219
rect 204694 66167 204746 66219
rect 210262 66167 210314 66219
rect 152662 66093 152714 66145
rect 204502 66093 204554 66145
rect 157654 66019 157706 66071
rect 204598 66019 204650 66071
rect 210262 65945 210314 65997
rect 144022 65575 144074 65627
rect 144214 65575 144266 65627
rect 145462 65131 145514 65183
rect 146518 65131 146570 65183
rect 144982 64983 145034 65035
rect 145462 64983 145514 65035
rect 144022 64835 144074 64887
rect 204502 64835 204554 64887
rect 144886 64761 144938 64813
rect 204598 64761 204650 64813
rect 146902 63355 146954 63407
rect 204502 63355 204554 63407
rect 144022 62171 144074 62223
rect 149782 62171 149834 62223
rect 160534 60765 160586 60817
rect 204598 60765 204650 60817
rect 156310 60691 156362 60743
rect 204694 60691 204746 60743
rect 152662 60617 152714 60669
rect 204502 60617 204554 60669
rect 151126 60543 151178 60595
rect 204886 60543 204938 60595
rect 148342 60469 148394 60521
rect 204790 60469 204842 60521
rect 146902 60395 146954 60447
rect 204502 60395 204554 60447
rect 149782 60321 149834 60373
rect 204694 60321 204746 60373
rect 207766 59951 207818 60003
rect 208726 59951 208778 60003
rect 144022 59581 144074 59633
rect 160534 59581 160586 59633
rect 144022 58989 144074 59041
rect 204598 58989 204650 59041
rect 144022 57065 144074 57117
rect 156310 57065 156362 57117
rect 144022 56473 144074 56525
rect 152662 56473 152714 56525
rect 210166 55215 210218 55267
rect 144022 54623 144074 54675
rect 151126 54623 151178 54675
rect 209494 54253 209546 54305
rect 217174 54253 217226 54305
rect 228502 54253 228554 54305
rect 209974 54179 210026 54231
rect 219190 54179 219242 54231
rect 144022 54105 144074 54157
rect 148342 54105 148394 54157
rect 209302 54105 209354 54157
rect 256054 54105 256106 54157
rect 206998 54031 207050 54083
rect 221398 54031 221450 54083
rect 210838 53957 210890 54009
rect 216982 53957 217034 54009
rect 210262 53809 210314 53861
rect 208054 53735 208106 53787
rect 218182 53735 218234 53787
rect 282166 53883 282218 53935
rect 208342 53661 208394 53713
rect 205654 53587 205706 53639
rect 216982 53661 217034 53713
rect 357430 53587 357482 53639
rect 383158 53587 383210 53639
rect 403126 53587 403178 53639
rect 210358 53513 210410 53565
rect 215254 53513 215306 53565
rect 215590 53513 215642 53565
rect 215782 53513 215834 53565
rect 217174 53513 217226 53565
rect 217462 53513 217514 53565
rect 228502 53513 228554 53565
rect 398326 53513 398378 53565
rect 423574 53513 423626 53565
rect 443350 53513 443402 53565
rect 460822 53513 460874 53565
rect 490966 53587 491018 53639
rect 209206 53439 209258 53491
rect 216358 53439 216410 53491
rect 209398 53365 209450 53417
rect 219670 53439 219722 53491
rect 256246 53439 256298 53491
rect 443446 53439 443498 53491
rect 209782 53291 209834 53343
rect 213430 53291 213482 53343
rect 209686 53217 209738 53269
rect 213718 53217 213770 53269
rect 207286 53143 207338 53195
rect 255958 53365 256010 53417
rect 256150 53365 256202 53417
rect 443350 53365 443402 53417
rect 460822 53365 460874 53417
rect 293686 53291 293738 53343
rect 403414 53291 403466 53343
rect 423382 53291 423434 53343
rect 443638 53291 443690 53343
rect 490966 53291 491018 53343
rect 512278 53291 512330 53343
rect 273622 53217 273674 53269
rect 210742 53069 210794 53121
rect 207094 52995 207146 53047
rect 220342 52995 220394 53047
rect 221398 52995 221450 53047
rect 276406 53069 276458 53121
rect 276598 53069 276650 53121
rect 321046 53217 321098 53269
rect 383062 53217 383114 53269
rect 443734 53217 443786 53269
rect 331126 53143 331178 53195
rect 362710 53143 362762 53195
rect 362998 53143 363050 53195
rect 403126 53143 403178 53195
rect 403318 53143 403370 53195
rect 440662 53143 440714 53195
rect 525910 53217 525962 53269
rect 321046 52995 321098 53047
rect 331126 52995 331178 53047
rect 208150 52921 208202 52973
rect 220054 52921 220106 52973
rect 210166 52847 210218 52899
rect 218902 52847 218954 52899
rect 151414 52699 151466 52751
rect 217270 52699 217322 52751
rect 443350 52551 443402 52603
rect 460726 52551 460778 52603
rect 211894 52477 211946 52529
rect 220918 52477 220970 52529
rect 212182 52329 212234 52381
rect 226966 52329 227018 52381
rect 137494 52255 137546 52307
rect 239062 52255 239114 52307
rect 151318 52181 151370 52233
rect 219862 52181 219914 52233
rect 146710 52107 146762 52159
rect 212182 52107 212234 52159
rect 144406 52033 144458 52085
rect 211894 52033 211946 52085
rect 144598 51959 144650 52011
rect 225718 52107 225770 52159
rect 212374 52033 212426 52085
rect 213430 52033 213482 52085
rect 146422 51885 146474 51937
rect 331126 51959 331178 52011
rect 342550 51959 342602 52011
rect 460822 51959 460874 52011
rect 470806 51959 470858 52011
rect 625942 51959 625994 52011
rect 639670 51959 639722 52011
rect 227542 51885 227594 51937
rect 213430 51811 213482 51863
rect 237430 51811 237482 51863
rect 239062 51811 239114 51863
rect 244150 51811 244202 51863
rect 254422 51811 254474 51863
rect 211222 51737 211274 51789
rect 322582 51811 322634 51863
rect 331126 51811 331178 51863
rect 342742 51811 342794 51863
rect 368470 51811 368522 51863
rect 368566 51811 368618 51863
rect 408886 51811 408938 51863
rect 408982 51811 409034 51863
rect 449206 51811 449258 51863
rect 449302 51811 449354 51863
rect 460822 51811 460874 51863
rect 509782 51811 509834 51863
rect 541366 51885 541418 51937
rect 209878 51663 209930 51715
rect 214102 51663 214154 51715
rect 308086 51737 308138 51789
rect 308182 51737 308234 51789
rect 322486 51737 322538 51789
rect 541462 51811 541514 51863
rect 558742 51885 558794 51937
rect 558838 51737 558890 51789
rect 590326 51811 590378 51863
rect 590422 51811 590474 51863
rect 645526 51737 645578 51789
rect 251926 51663 251978 51715
rect 209590 51589 209642 51641
rect 214486 51589 214538 51641
rect 253558 51589 253610 51641
rect 308086 51589 308138 51641
rect 308182 51589 308234 51641
rect 322390 51663 322442 51715
rect 145366 51515 145418 51567
rect 236758 51515 236810 51567
rect 237430 51515 237482 51567
rect 145942 51441 145994 51493
rect 237142 51441 237194 51493
rect 144790 51367 144842 51419
rect 233590 51367 233642 51419
rect 322390 51515 322442 51567
rect 342742 51589 342794 51641
rect 342646 51515 342698 51567
rect 362998 51589 363050 51641
rect 374422 51589 374474 51641
rect 394486 51589 394538 51641
rect 414646 51663 414698 51715
rect 470806 51663 470858 51715
rect 509686 51663 509738 51715
rect 518326 51663 518378 51715
rect 362806 51515 362858 51567
rect 417526 51515 417578 51567
rect 423286 51589 423338 51641
rect 423382 51589 423434 51641
rect 457942 51589 457994 51641
rect 480886 51589 480938 51641
rect 498262 51589 498314 51641
rect 604726 51663 604778 51715
rect 538582 51589 538634 51641
rect 541462 51589 541514 51641
rect 584662 51589 584714 51641
rect 625942 51589 625994 51641
rect 251926 51441 251978 51493
rect 253462 51441 253514 51493
rect 478006 51441 478058 51493
rect 480886 51441 480938 51493
rect 254422 51367 254474 51419
rect 414646 51367 414698 51419
rect 417526 51367 417578 51419
rect 144982 51293 145034 51345
rect 234550 51293 234602 51345
rect 145654 51219 145706 51271
rect 235318 51219 235370 51271
rect 145846 51145 145898 51197
rect 234934 51145 234986 51197
rect 146230 51071 146282 51123
rect 232342 51071 232394 51123
rect 146806 50997 146858 51049
rect 231958 50997 232010 51049
rect 146614 50923 146666 50975
rect 230998 50923 231050 50975
rect 145558 50849 145610 50901
rect 231382 50849 231434 50901
rect 146038 50775 146090 50827
rect 230518 50775 230570 50827
rect 145078 50701 145130 50753
rect 228310 50701 228362 50753
rect 145462 50627 145514 50679
rect 228694 50627 228746 50679
rect 145270 50553 145322 50605
rect 229750 50553 229802 50605
rect 145174 50479 145226 50531
rect 228790 50479 228842 50531
rect 144502 50405 144554 50457
rect 208054 50405 208106 50457
rect 144118 50331 144170 50383
rect 207958 50331 208010 50383
rect 208246 50331 208298 50383
rect 216118 50331 216170 50383
rect 146134 50257 146186 50309
rect 207862 50257 207914 50309
rect 208438 50257 208490 50309
rect 216886 50257 216938 50309
rect 144310 50183 144362 50235
rect 208342 50183 208394 50235
rect 208534 50183 208586 50235
rect 217654 50183 217706 50235
rect 144214 50109 144266 50161
rect 235798 50109 235850 50161
rect 146518 50035 146570 50087
rect 235414 50035 235466 50087
rect 144694 49961 144746 50013
rect 232726 49961 232778 50013
rect 208054 49887 208106 49939
rect 224950 49887 225002 49939
rect 208342 49813 208394 49865
rect 224278 49813 224330 49865
rect 207958 49739 208010 49791
rect 225334 49739 225386 49791
rect 145750 49665 145802 49717
rect 211606 49665 211658 49717
rect 645814 49739 645866 49791
rect 207862 49591 207914 49643
rect 226582 49591 226634 49643
rect 215830 49443 215882 49495
rect 215926 49443 215978 49495
rect 218806 49443 218858 49495
rect 218806 49295 218858 49347
rect 241174 49295 241226 49347
rect 443446 48999 443498 49051
rect 210070 48925 210122 48977
rect 220726 48925 220778 48977
rect 223702 48925 223754 48977
rect 229654 48925 229706 48977
rect 282358 48925 282410 48977
rect 302422 48925 302474 48977
rect 471382 48925 471434 48977
rect 222262 48851 222314 48903
rect 645142 48851 645194 48903
rect 209014 48777 209066 48829
rect 222070 48777 222122 48829
rect 222934 48777 222986 48829
rect 645238 48777 645290 48829
rect 208630 48703 208682 48755
rect 221686 48703 221738 48755
rect 224086 48703 224138 48755
rect 645334 48703 645386 48755
rect 148246 48629 148298 48681
rect 236374 48629 236426 48681
rect 148822 48555 148874 48607
rect 234166 48555 234218 48607
rect 185686 48481 185738 48533
rect 240214 48481 240266 48533
rect 197206 48407 197258 48459
rect 239830 48407 239882 48459
rect 194326 48333 194378 48385
rect 239734 48333 239786 48385
rect 202966 48259 203018 48311
rect 241558 48259 241610 48311
rect 149302 48185 149354 48237
rect 208534 48185 208586 48237
rect 208918 48185 208970 48237
rect 222454 48185 222506 48237
rect 149398 48111 149450 48163
rect 208630 48111 208682 48163
rect 208822 48111 208874 48163
rect 222742 48111 222794 48163
rect 148054 48037 148106 48089
rect 219478 48037 219530 48089
rect 148150 47963 148202 48015
rect 219094 47963 219146 48015
rect 149494 47889 149546 47941
rect 221302 47889 221354 47941
rect 149590 47815 149642 47867
rect 220534 47815 220586 47867
rect 149686 47741 149738 47793
rect 220246 47741 220298 47793
rect 147670 47667 147722 47719
rect 216502 47667 216554 47719
rect 147766 47593 147818 47645
rect 218038 47593 218090 47645
rect 218518 47593 218570 47645
rect 645622 47593 645674 47645
rect 147958 47519 148010 47571
rect 218710 47519 218762 47571
rect 147862 47445 147914 47497
rect 218326 47445 218378 47497
rect 177046 47371 177098 47423
rect 238006 47371 238058 47423
rect 179926 47297 179978 47349
rect 238582 47297 238634 47349
rect 200086 47223 200138 47275
rect 238966 47223 239018 47275
rect 148918 47149 148970 47201
rect 233302 47149 233354 47201
rect 188566 47075 188618 47127
rect 239350 47075 239402 47127
rect 148534 47001 148586 47053
rect 230902 47001 230954 47053
rect 191446 46927 191498 46979
rect 240790 46927 240842 46979
rect 148726 46853 148778 46905
rect 227926 46853 227978 46905
rect 148438 46779 148490 46831
rect 233110 46779 233162 46831
rect 149206 46705 149258 46757
rect 208438 46705 208490 46757
rect 208726 46705 208778 46757
rect 223510 46705 223562 46757
rect 149014 46631 149066 46683
rect 230134 46631 230186 46683
rect 207766 46557 207818 46609
rect 223894 46557 223946 46609
rect 149110 46483 149162 46535
rect 208342 46483 208394 46535
rect 208630 46483 208682 46535
rect 223126 46483 223178 46535
rect 148630 46409 148682 46461
rect 229174 46409 229226 46461
rect 208534 46335 208586 46387
rect 224662 46335 224714 46387
rect 208438 46261 208490 46313
rect 226102 46261 226154 46313
rect 208342 46187 208394 46239
rect 226486 46187 226538 46239
rect 398326 46113 398378 46165
rect 408886 46039 408938 46091
rect 211414 45299 211466 45351
rect 361750 45299 361802 45351
rect 213238 45225 213290 45277
rect 406102 45225 406154 45277
rect 212854 45151 212906 45203
rect 411574 45151 411626 45203
rect 213910 45077 213962 45129
rect 443926 45077 443978 45129
rect 215062 45003 215114 45055
rect 509686 45003 509738 45055
rect 214678 44929 214730 44981
rect 508246 44929 508298 44981
rect 508246 43227 508298 43279
rect 406102 43153 406154 43205
rect 410998 43153 411050 43205
rect 521494 43153 521546 43205
rect 133654 42783 133706 42835
rect 136534 42783 136586 42835
rect 212470 42339 212522 42391
rect 310102 42339 310154 42391
rect 206902 42117 206954 42169
rect 405238 42117 405290 42169
rect 213622 42043 213674 42095
rect 460054 42043 460106 42095
rect 214294 41969 214346 42021
rect 514870 41969 514922 42021
rect 459190 41525 459242 41577
rect 443926 37381 443978 37433
rect 459190 37381 459242 37433
<< metal2 >>
rect 148532 1015974 148588 1015983
rect 148532 1015909 148588 1015918
rect 251348 1015974 251404 1015983
rect 251348 1015909 251404 1015918
rect 353396 1015974 353452 1015983
rect 353396 1015909 353452 1015918
rect 148546 1007991 148574 1015909
rect 145364 1007982 145420 1007991
rect 145364 1007917 145420 1007926
rect 148532 1007982 148588 1007991
rect 148532 1007917 148588 1007926
rect 143926 1002615 143978 1002621
rect 143926 1002557 143978 1002563
rect 143734 1002541 143786 1002547
rect 143734 1002483 143786 1002489
rect 143746 999532 143774 1002483
rect 143830 1002393 143882 1002399
rect 143830 1002335 143882 1002341
rect 143650 999504 143774 999532
rect 92662 999433 92714 999439
rect 92662 999375 92714 999381
rect 126646 999433 126698 999439
rect 126646 999375 126698 999381
rect 81044 995846 81100 995855
rect 80784 995804 81044 995832
rect 85728 995813 85982 995832
rect 91248 995813 91550 995832
rect 85728 995807 85994 995813
rect 85728 995804 85942 995807
rect 81044 995781 81100 995790
rect 91248 995807 91562 995813
rect 91248 995804 91510 995807
rect 85942 995749 85994 995755
rect 91510 995749 91562 995755
rect 81620 995698 81676 995707
rect 81408 995656 81620 995684
rect 81620 995633 81676 995642
rect 85364 995550 85420 995559
rect 77088 995508 77342 995536
rect 69142 995141 69194 995147
rect 69142 995083 69194 995089
rect 61846 993587 61898 993593
rect 61846 993529 61898 993535
rect 47638 988333 47690 988339
rect 47638 988275 47690 988281
rect 44758 988259 44810 988265
rect 44758 988201 44810 988207
rect 43126 987889 43178 987895
rect 43126 987831 43178 987837
rect 42178 968771 42206 969252
rect 42164 968762 42220 968771
rect 42164 968697 42220 968706
rect 41794 967143 41822 967402
rect 43138 967323 43166 987831
rect 42166 967317 42218 967323
rect 42166 967259 42218 967265
rect 43126 967317 43178 967323
rect 43126 967259 43178 967265
rect 41780 967134 41836 967143
rect 41780 967069 41836 967078
rect 42178 966736 42206 967259
rect 41794 965071 41822 965552
rect 41780 965062 41836 965071
rect 41780 964997 41836 965006
rect 42178 964035 42206 964368
rect 42164 964026 42220 964035
rect 42164 963961 42220 963970
rect 41794 963443 41822 963702
rect 41780 963434 41836 963443
rect 41780 963369 41836 963378
rect 41794 962703 41822 963081
rect 41780 962694 41836 962703
rect 41780 962629 41836 962638
rect 41890 962259 41918 962518
rect 42164 962398 42220 962407
rect 42220 962356 42302 962384
rect 42164 962333 42220 962342
rect 41876 962250 41932 962259
rect 41876 962185 41932 962194
rect 42178 961200 42206 961260
rect 42274 961200 42302 962356
rect 42452 962102 42508 962111
rect 42452 962037 42508 962046
rect 42178 961172 42302 961200
rect 42466 961033 42494 962037
rect 42166 961027 42218 961033
rect 42166 960969 42218 960975
rect 42454 961027 42506 961033
rect 42454 960969 42506 960975
rect 42178 960594 42206 960969
rect 41794 959743 41822 960045
rect 41780 959734 41836 959743
rect 41780 959669 41836 959678
rect 41890 959151 41918 959410
rect 41876 959142 41932 959151
rect 41876 959077 41932 959086
rect 41794 958559 41822 958744
rect 41780 958550 41836 958559
rect 41780 958485 41836 958494
rect 42178 957819 42206 958226
rect 42164 957810 42220 957819
rect 42164 957745 42220 957754
rect 42082 956191 42110 956376
rect 42068 956182 42124 956191
rect 42068 956117 42124 956126
rect 42082 955261 42110 955710
rect 42070 955255 42122 955261
rect 42070 955197 42122 955203
rect 42838 955255 42890 955261
rect 42838 955197 42890 955203
rect 41794 954669 41822 955077
rect 41782 954663 41834 954669
rect 41782 954605 41834 954611
rect 41782 954441 41834 954447
rect 41782 954383 41834 954389
rect 40436 943010 40492 943019
rect 40436 942945 40492 942954
rect 40342 942379 40394 942385
rect 40342 942321 40394 942327
rect 40052 941974 40108 941983
rect 40052 941909 40108 941918
rect 39956 941826 40012 941835
rect 39956 941761 40012 941770
rect 39970 939171 39998 941761
rect 40066 940355 40094 941909
rect 40052 940346 40108 940355
rect 40052 940281 40108 940290
rect 39956 939162 40012 939171
rect 39956 939097 40012 939106
rect 35252 932650 35308 932659
rect 35252 932585 35308 932594
rect 35266 932215 35294 932585
rect 35252 932206 35308 932215
rect 35252 932141 35308 932150
rect 40354 816775 40382 942321
rect 40450 817219 40478 942945
rect 41794 941983 41822 954383
rect 42550 944673 42602 944679
rect 42548 944638 42550 944647
rect 42602 944638 42604 944647
rect 42548 944573 42604 944582
rect 42550 944229 42602 944235
rect 42548 944194 42550 944203
rect 42602 944194 42604 944203
rect 42548 944129 42604 944138
rect 42550 944081 42602 944087
rect 42548 944046 42550 944055
rect 42602 944046 42604 944055
rect 42548 943981 42604 943990
rect 42550 943045 42602 943051
rect 42548 943010 42550 943019
rect 42602 943010 42604 943019
rect 42548 942945 42604 942954
rect 42550 942897 42602 942903
rect 42550 942839 42602 942845
rect 42562 942427 42590 942839
rect 42548 942418 42604 942427
rect 42548 942353 42550 942362
rect 42602 942353 42604 942362
rect 42550 942321 42602 942327
rect 42562 942293 42590 942321
rect 41780 941974 41836 941983
rect 41780 941909 41836 941918
rect 42850 937839 42878 955197
rect 42836 937830 42892 937839
rect 42836 937765 42892 937774
rect 42548 933242 42604 933251
rect 42548 933177 42604 933186
rect 42562 932215 42590 933177
rect 42548 932206 42604 932215
rect 42548 932141 42550 932150
rect 42602 932141 42604 932150
rect 42550 932109 42602 932115
rect 42550 819317 42602 819323
rect 42548 819282 42550 819291
rect 42602 819282 42604 819291
rect 42548 819217 42604 819226
rect 42838 818577 42890 818583
rect 42836 818542 42838 818551
rect 42890 818542 42892 818551
rect 42836 818477 42892 818486
rect 42550 818281 42602 818287
rect 42548 818246 42550 818255
rect 42602 818246 42604 818255
rect 42548 818181 42604 818190
rect 43220 817506 43276 817515
rect 43220 817441 43276 817450
rect 40436 817210 40492 817219
rect 40436 817145 40492 817154
rect 40340 816766 40396 816775
rect 40340 816701 40396 816710
rect 41684 814990 41740 814999
rect 41684 814925 41740 814934
rect 40244 813954 40300 813963
rect 40244 813889 40300 813898
rect 40148 811734 40204 811743
rect 40148 811669 40204 811678
rect 35156 806850 35212 806859
rect 35156 806785 35212 806794
rect 35170 806415 35198 806785
rect 35156 806406 35212 806415
rect 35156 806341 35212 806350
rect 40162 801975 40190 811669
rect 40258 802123 40286 813889
rect 41492 810550 41548 810559
rect 41492 810485 41548 810494
rect 40244 802114 40300 802123
rect 40244 802049 40300 802058
rect 40148 801966 40204 801975
rect 40148 801901 40204 801910
rect 41506 800791 41534 810485
rect 41588 808922 41644 808931
rect 41588 808857 41644 808866
rect 41492 800782 41548 800791
rect 41492 800717 41548 800726
rect 41602 800643 41630 808857
rect 41588 800634 41644 800643
rect 41588 800569 41644 800578
rect 41698 800495 41726 814925
rect 42548 814398 42604 814407
rect 42548 814333 42604 814342
rect 41972 813362 42028 813371
rect 41972 813297 42028 813306
rect 41876 812326 41932 812335
rect 41876 812261 41932 812270
rect 41780 808478 41836 808487
rect 41780 808413 41836 808422
rect 41684 800486 41740 800495
rect 41684 800421 41740 800430
rect 41794 800347 41822 808413
rect 41780 800338 41836 800347
rect 41780 800273 41836 800282
rect 41890 800231 41918 812261
rect 41986 802081 42014 813297
rect 42068 812770 42124 812779
rect 42068 812705 42124 812714
rect 42082 802451 42110 812705
rect 42164 809514 42220 809523
rect 42164 809449 42220 809458
rect 42070 802445 42122 802451
rect 42070 802387 42122 802393
rect 41974 802075 42026 802081
rect 41974 802017 42026 802023
rect 42178 800347 42206 809449
rect 42562 807483 42590 814333
rect 43124 811438 43180 811447
rect 43124 811373 43180 811382
rect 42932 810402 42988 810411
rect 42932 810337 42988 810346
rect 42550 807477 42602 807483
rect 42550 807419 42602 807425
rect 42838 807477 42890 807483
rect 42838 807419 42890 807425
rect 42454 802075 42506 802081
rect 42454 802017 42506 802023
rect 42466 801952 42494 802017
rect 42466 801924 42590 801952
rect 42164 800338 42220 800347
rect 42164 800273 42220 800282
rect 41878 800225 41930 800231
rect 41878 800167 41930 800173
rect 41878 800003 41930 800009
rect 41878 799945 41930 799951
rect 41890 799422 41918 799945
rect 42166 798153 42218 798159
rect 42166 798095 42218 798101
rect 42178 797605 42206 798095
rect 42070 797339 42122 797345
rect 42070 797281 42122 797287
rect 42082 796980 42110 797281
rect 42166 796303 42218 796309
rect 42166 796245 42218 796251
rect 42178 795765 42206 796245
rect 42166 795045 42218 795051
rect 42166 794987 42218 794993
rect 42178 794569 42206 794987
rect 42068 794270 42124 794279
rect 42068 794205 42124 794214
rect 42082 793946 42110 794205
rect 41780 793826 41836 793835
rect 41780 793761 41836 793770
rect 41794 793280 41822 793761
rect 42166 793195 42218 793201
rect 42166 793137 42218 793143
rect 42178 792729 42206 793137
rect 42452 792198 42508 792207
rect 42562 792184 42590 801924
rect 42850 798381 42878 807419
rect 42946 798381 42974 810337
rect 43028 808182 43084 808191
rect 43028 808117 43084 808126
rect 42838 798375 42890 798381
rect 42838 798317 42890 798323
rect 42934 798375 42986 798381
rect 42934 798317 42986 798323
rect 42742 798079 42794 798085
rect 42742 798021 42794 798027
rect 42754 796309 42782 798021
rect 42742 796303 42794 796309
rect 42742 796245 42794 796251
rect 42740 796194 42796 796203
rect 42740 796129 42796 796138
rect 42508 792156 42590 792184
rect 42452 792133 42508 792142
rect 42452 791902 42508 791911
rect 42452 791837 42508 791846
rect 42082 791171 42110 791430
rect 42068 791162 42124 791171
rect 42068 791097 42124 791106
rect 41794 790579 41822 790797
rect 42166 790679 42218 790685
rect 42166 790621 42218 790627
rect 41780 790570 41836 790579
rect 41780 790505 41836 790514
rect 42178 790246 42206 790621
rect 42166 789939 42218 789945
rect 42166 789881 42218 789887
rect 42178 789580 42206 789881
rect 42166 789495 42218 789501
rect 42166 789437 42218 789443
rect 42178 788957 42206 789437
rect 42466 788835 42494 791837
rect 42754 790685 42782 796129
rect 43042 795051 43070 808117
rect 43138 802599 43166 811373
rect 43126 802593 43178 802599
rect 43126 802535 43178 802541
rect 43126 802445 43178 802451
rect 43126 802387 43178 802393
rect 43030 795045 43082 795051
rect 43030 794987 43082 794993
rect 43138 793201 43166 802387
rect 43126 793195 43178 793201
rect 43126 793137 43178 793143
rect 42836 791902 42892 791911
rect 42836 791837 42892 791846
rect 42742 790679 42794 790685
rect 42742 790621 42794 790627
rect 42850 789945 42878 791837
rect 42932 791754 42988 791763
rect 42932 791689 42988 791698
rect 42838 789939 42890 789945
rect 42838 789881 42890 789887
rect 42836 789386 42892 789395
rect 42836 789321 42892 789330
rect 42740 789238 42796 789247
rect 42740 789173 42796 789182
rect 42166 788829 42218 788835
rect 42166 788771 42218 788777
rect 42454 788829 42506 788835
rect 42454 788771 42506 788777
rect 42178 788396 42206 788771
rect 42166 787053 42218 787059
rect 42166 786995 42218 787001
rect 42178 786546 42206 786995
rect 42754 786467 42782 789173
rect 42166 786461 42218 786467
rect 42166 786403 42218 786409
rect 42742 786461 42794 786467
rect 42742 786403 42794 786409
rect 42178 785921 42206 786403
rect 42850 785653 42878 789321
rect 42946 787059 42974 791689
rect 42934 787053 42986 787059
rect 42934 786995 42986 787001
rect 42070 785647 42122 785653
rect 42070 785589 42122 785595
rect 42838 785647 42890 785653
rect 42838 785589 42890 785595
rect 42082 785288 42110 785589
rect 42742 775953 42794 775959
rect 42740 775918 42742 775927
rect 42794 775918 42796 775927
rect 42740 775853 42796 775862
rect 42742 775361 42794 775367
rect 42740 775326 42742 775335
rect 42794 775326 42796 775335
rect 42740 775261 42796 775270
rect 42742 774843 42794 774849
rect 42740 774808 42742 774817
rect 42794 774808 42796 774817
rect 42740 774743 42796 774752
rect 43234 774424 43262 817441
rect 44660 806554 44716 806563
rect 44660 806489 44716 806498
rect 43414 802593 43466 802599
rect 43414 802535 43466 802541
rect 43318 800669 43370 800675
rect 43318 800611 43370 800617
rect 43330 797345 43358 800611
rect 43318 797339 43370 797345
rect 43318 797281 43370 797287
rect 43426 789501 43454 802535
rect 43414 789495 43466 789501
rect 43414 789437 43466 789443
rect 43234 774396 43454 774424
rect 43220 774290 43276 774299
rect 43220 774225 43276 774234
rect 42932 772070 42988 772079
rect 42932 772005 42988 772014
rect 41972 771182 42028 771191
rect 41972 771117 42028 771126
rect 40244 770738 40300 770747
rect 40244 770673 40300 770682
rect 35156 763634 35212 763643
rect 35156 763569 35212 763578
rect 35170 763199 35198 763569
rect 35156 763190 35212 763199
rect 35156 763125 35212 763134
rect 40258 757723 40286 770673
rect 41492 770146 41548 770155
rect 41492 770081 41548 770090
rect 40244 757714 40300 757723
rect 40244 757649 40300 757658
rect 41506 757427 41534 770081
rect 41780 769554 41836 769563
rect 41780 769489 41836 769498
rect 41588 767482 41644 767491
rect 41588 767417 41644 767426
rect 41492 757418 41548 757427
rect 41602 757385 41630 767417
rect 41684 766298 41740 766307
rect 41684 766233 41740 766242
rect 41492 757353 41548 757362
rect 41590 757379 41642 757385
rect 41590 757321 41642 757327
rect 41698 757311 41726 766233
rect 41686 757305 41738 757311
rect 41794 757279 41822 769489
rect 41876 769110 41932 769119
rect 41876 769045 41932 769054
rect 41686 757247 41738 757253
rect 41780 757270 41836 757279
rect 41780 757205 41836 757214
rect 41890 757015 41918 769045
rect 41986 757131 42014 771117
rect 42068 766298 42124 766307
rect 42068 766233 42124 766242
rect 41972 757122 42028 757131
rect 41972 757057 42028 757066
rect 42082 757015 42110 766233
rect 42838 758637 42890 758643
rect 42838 758579 42890 758585
rect 41878 757009 41930 757015
rect 41878 756951 41930 756957
rect 42070 757009 42122 757015
rect 42070 756951 42122 756957
rect 41878 756787 41930 756793
rect 41878 756729 41930 756735
rect 41890 756245 41918 756729
rect 42850 756719 42878 758579
rect 42838 756713 42890 756719
rect 42838 756655 42890 756661
rect 41876 754902 41932 754911
rect 41876 754837 41932 754846
rect 41890 754430 41918 754837
rect 42166 754123 42218 754129
rect 42166 754065 42218 754071
rect 42178 753764 42206 754065
rect 42070 753087 42122 753093
rect 42070 753029 42122 753035
rect 42082 752580 42110 753029
rect 42946 751951 42974 772005
rect 43124 767186 43180 767195
rect 43124 767121 43180 767130
rect 43028 765558 43084 765567
rect 43028 765493 43084 765502
rect 43042 758643 43070 765493
rect 43030 758637 43082 758643
rect 43030 758579 43082 758585
rect 43138 758144 43166 767121
rect 43234 761844 43262 774225
rect 43426 773707 43454 774396
rect 43412 773698 43468 773707
rect 43412 773633 43468 773642
rect 43234 761816 43742 761844
rect 43138 758116 43358 758144
rect 43330 757700 43358 758116
rect 43030 757675 43082 757681
rect 43030 757617 43082 757623
rect 43138 757672 43358 757700
rect 43042 754277 43070 757617
rect 43030 754271 43082 754277
rect 43030 754213 43082 754219
rect 43030 754123 43082 754129
rect 43030 754065 43082 754071
rect 42932 751942 42988 751951
rect 42932 751877 42988 751886
rect 42068 751794 42124 751803
rect 42068 751729 42124 751738
rect 42934 751755 42986 751761
rect 42082 751396 42110 751729
rect 42934 751697 42986 751703
rect 42946 751169 42974 751697
rect 42070 751163 42122 751169
rect 42070 751105 42122 751111
rect 42934 751163 42986 751169
rect 42934 751105 42986 751111
rect 42082 750730 42110 751105
rect 42932 751054 42988 751063
rect 42932 750989 42988 750998
rect 42166 750423 42218 750429
rect 42166 750365 42218 750371
rect 42178 750064 42206 750365
rect 42068 749870 42124 749879
rect 42068 749805 42124 749814
rect 42082 749546 42110 749805
rect 42452 749278 42508 749287
rect 42452 749213 42508 749222
rect 41986 747807 42014 748214
rect 41972 747798 42028 747807
rect 41972 747733 42028 747742
rect 41794 747215 41822 747622
rect 42166 747315 42218 747321
rect 42166 747257 42218 747263
rect 41780 747206 41836 747215
rect 41780 747141 41836 747150
rect 42178 747030 42206 747257
rect 42166 746945 42218 746951
rect 42166 746887 42218 746893
rect 42178 746401 42206 746887
rect 42068 746318 42124 746327
rect 42068 746253 42124 746262
rect 42082 745772 42110 746253
rect 42166 745687 42218 745693
rect 42166 745629 42218 745635
rect 42178 745180 42206 745629
rect 42466 745545 42494 749213
rect 42946 745693 42974 750989
rect 43042 750429 43070 754065
rect 43138 753093 43166 757672
rect 43510 757379 43562 757385
rect 43510 757321 43562 757327
rect 43414 757305 43466 757311
rect 43414 757247 43466 757253
rect 43318 757009 43370 757015
rect 43318 756951 43370 756957
rect 43222 756713 43274 756719
rect 43222 756655 43274 756661
rect 43234 754129 43262 756655
rect 43222 754123 43274 754129
rect 43222 754065 43274 754071
rect 43330 753112 43358 756951
rect 43126 753087 43178 753093
rect 43126 753029 43178 753035
rect 43234 753084 43358 753112
rect 43234 752964 43262 753084
rect 43138 752936 43262 752964
rect 43138 751835 43166 752936
rect 43426 752594 43454 757247
rect 43330 752566 43454 752594
rect 43126 751829 43178 751835
rect 43126 751771 43178 751777
rect 43330 751632 43358 752566
rect 43138 751604 43358 751632
rect 43414 751681 43466 751687
rect 43414 751623 43466 751629
rect 43030 750423 43082 750429
rect 43030 750365 43082 750371
rect 43030 750275 43082 750281
rect 43030 750217 43082 750223
rect 43042 747025 43070 750217
rect 43138 747321 43166 751604
rect 43126 747315 43178 747321
rect 43126 747257 43178 747263
rect 43124 747058 43180 747067
rect 43030 747019 43082 747025
rect 43124 746993 43180 747002
rect 43030 746961 43082 746967
rect 43028 746910 43084 746919
rect 43028 746845 43084 746854
rect 42934 745687 42986 745693
rect 42934 745629 42986 745635
rect 42454 745539 42506 745545
rect 42454 745481 42506 745487
rect 42934 745539 42986 745545
rect 42934 745481 42986 745487
rect 42946 743843 42974 745481
rect 42166 743837 42218 743843
rect 42166 743779 42218 743785
rect 42934 743837 42986 743843
rect 42934 743779 42986 743785
rect 42178 743365 42206 743779
rect 42070 743245 42122 743251
rect 42070 743187 42122 743193
rect 42082 742738 42110 743187
rect 43042 742659 43070 746845
rect 43138 743251 43166 746993
rect 43126 743245 43178 743251
rect 43126 743187 43178 743193
rect 42166 742653 42218 742659
rect 42166 742595 42218 742601
rect 43030 742653 43082 742659
rect 43030 742595 43082 742601
rect 42178 742072 42206 742595
rect 42838 732737 42890 732743
rect 42836 732702 42838 732711
rect 42890 732702 42892 732711
rect 42836 732637 42892 732646
rect 42838 732145 42890 732151
rect 42836 732110 42838 732119
rect 42890 732110 42892 732119
rect 42836 732045 42892 732054
rect 42838 731849 42890 731855
rect 42836 731814 42838 731823
rect 42890 731814 42892 731823
rect 42836 731749 42892 731758
rect 43426 730491 43454 751623
rect 43522 750281 43550 757321
rect 43714 751687 43742 761816
rect 43702 751681 43754 751687
rect 43702 751623 43754 751629
rect 43510 750275 43562 750281
rect 43510 750217 43562 750223
rect 43700 731074 43756 731083
rect 43700 731009 43756 731018
rect 43412 730482 43468 730491
rect 43412 730417 43468 730426
rect 41492 728706 41548 728715
rect 41492 728641 41548 728650
rect 35156 720418 35212 720427
rect 35156 720353 35212 720362
rect 35170 719983 35198 720353
rect 35156 719974 35212 719983
rect 35156 719909 35212 719918
rect 41506 714243 41534 728641
rect 42452 727966 42508 727975
rect 42508 727924 42590 727952
rect 42452 727901 42508 727910
rect 41588 726930 41644 726939
rect 41588 726865 41644 726874
rect 41494 714237 41546 714243
rect 41494 714179 41546 714185
rect 41602 714169 41630 726865
rect 41876 725894 41932 725903
rect 41876 725829 41932 725838
rect 41684 724710 41740 724719
rect 41684 724645 41740 724654
rect 41590 714163 41642 714169
rect 41590 714105 41642 714111
rect 41698 714095 41726 724645
rect 41780 724266 41836 724275
rect 41780 724201 41836 724210
rect 41686 714089 41738 714095
rect 41686 714031 41738 714037
rect 41794 713915 41822 724201
rect 41780 713906 41836 713915
rect 41890 713873 41918 725829
rect 41972 723674 42028 723683
rect 41972 723609 42028 723618
rect 41986 713873 42014 723609
rect 42068 722638 42124 722647
rect 42068 722573 42124 722582
rect 42082 714063 42110 722573
rect 42164 722046 42220 722055
rect 42164 721981 42220 721990
rect 42452 722046 42508 722055
rect 42562 722032 42590 727924
rect 43124 726338 43180 726347
rect 43124 726273 43180 726282
rect 42508 722004 42590 722032
rect 42452 721981 42508 721990
rect 42068 714054 42124 714063
rect 42068 713989 42124 713998
rect 42178 713915 42206 721981
rect 42452 721602 42508 721611
rect 42452 721537 42508 721546
rect 42164 713906 42220 713915
rect 41780 713841 41836 713850
rect 41878 713867 41930 713873
rect 41878 713809 41930 713815
rect 41974 713867 42026 713873
rect 42164 713841 42220 713850
rect 41974 713809 42026 713815
rect 41878 713571 41930 713577
rect 41878 713513 41930 713519
rect 41890 713064 41918 713513
rect 42466 713323 42494 721537
rect 43138 717277 43166 726273
rect 43316 722046 43372 722055
rect 43316 721981 43372 721990
rect 43126 717271 43178 717277
rect 43126 717213 43178 717219
rect 43126 717123 43178 717129
rect 43126 717065 43178 717071
rect 42452 713314 42508 713323
rect 42452 713249 42508 713258
rect 42070 711721 42122 711727
rect 42070 711663 42122 711669
rect 42082 711214 42110 711663
rect 43138 711524 43166 717065
rect 43222 713867 43274 713873
rect 43222 713809 43274 713815
rect 43234 711653 43262 713809
rect 43330 711727 43358 721981
rect 43510 714237 43562 714243
rect 43510 714179 43562 714185
rect 43414 714089 43466 714095
rect 43414 714031 43466 714037
rect 43318 711721 43370 711727
rect 43318 711663 43370 711669
rect 43426 711653 43454 714031
rect 43222 711647 43274 711653
rect 43222 711589 43274 711595
rect 43414 711647 43466 711653
rect 43414 711589 43466 711595
rect 43138 711496 43454 711524
rect 43126 711425 43178 711431
rect 43318 711425 43370 711431
rect 43126 711367 43178 711373
rect 43220 711390 43276 711399
rect 43028 711094 43084 711103
rect 43028 711029 43084 711038
rect 42166 710907 42218 710913
rect 42166 710849 42218 710855
rect 42178 710548 42206 710849
rect 42166 709945 42218 709951
rect 42166 709887 42218 709893
rect 42178 709364 42206 709887
rect 42068 708578 42124 708587
rect 42068 708513 42124 708522
rect 42082 708180 42110 708513
rect 41780 707986 41836 707995
rect 41780 707921 41836 707930
rect 41794 707514 41822 707921
rect 42740 707838 42796 707847
rect 42740 707773 42796 707782
rect 42164 707394 42220 707403
rect 42164 707329 42220 707338
rect 42178 706881 42206 707329
rect 42166 706763 42218 706769
rect 42166 706705 42218 706711
rect 42178 706330 42206 706705
rect 42452 705470 42508 705479
rect 42452 705405 42508 705414
rect 41890 704739 41918 705041
rect 41876 704730 41932 704739
rect 41876 704665 41932 704674
rect 41794 704147 41822 704406
rect 42166 704321 42218 704327
rect 42166 704263 42218 704269
rect 41780 704138 41836 704147
rect 41780 704073 41836 704082
rect 42178 703845 42206 704263
rect 42070 703729 42122 703735
rect 42070 703671 42122 703677
rect 42082 703222 42110 703671
rect 42166 702915 42218 702921
rect 42166 702857 42218 702863
rect 42178 702556 42206 702857
rect 42166 702323 42218 702329
rect 42166 702265 42218 702271
rect 42178 702005 42206 702265
rect 42070 700473 42122 700479
rect 42070 700415 42122 700421
rect 42082 700188 42110 700415
rect 42466 700109 42494 705405
rect 42754 704327 42782 707773
rect 42742 704321 42794 704327
rect 42742 704263 42794 704269
rect 42742 704173 42794 704179
rect 42742 704115 42794 704121
rect 42754 702329 42782 704115
rect 43042 703735 43070 711029
rect 43138 709951 43166 711367
rect 43318 711367 43370 711373
rect 43220 711325 43276 711334
rect 43126 709945 43178 709951
rect 43126 709887 43178 709893
rect 43234 706621 43262 711325
rect 43222 706615 43274 706621
rect 43222 706557 43274 706563
rect 43330 706492 43358 711367
rect 43426 710913 43454 711496
rect 43414 710907 43466 710913
rect 43414 710849 43466 710855
rect 43138 706464 43358 706492
rect 43030 703729 43082 703735
rect 43030 703671 43082 703677
rect 43028 703546 43084 703555
rect 43028 703481 43084 703490
rect 42742 702323 42794 702329
rect 42742 702265 42794 702271
rect 42166 700103 42218 700109
rect 42166 700045 42218 700051
rect 42454 700103 42506 700109
rect 42454 700045 42506 700051
rect 42178 699522 42206 700045
rect 42454 699881 42506 699887
rect 42454 699823 42506 699829
rect 42166 699215 42218 699221
rect 42166 699157 42218 699163
rect 42178 698856 42206 699157
rect 42466 689199 42494 699823
rect 43042 699221 43070 703481
rect 43138 702921 43166 706464
rect 43222 706393 43274 706399
rect 43222 706335 43274 706341
rect 43126 702915 43178 702921
rect 43126 702857 43178 702863
rect 43126 702767 43178 702773
rect 43126 702709 43178 702715
rect 43138 700479 43166 702709
rect 43126 700473 43178 700479
rect 43126 700415 43178 700421
rect 43030 699215 43082 699221
rect 43030 699157 43082 699163
rect 42838 689521 42890 689527
rect 42836 689486 42838 689495
rect 42890 689486 42892 689495
rect 42836 689421 42892 689430
rect 42452 689190 42508 689199
rect 42452 689125 42508 689134
rect 42454 688633 42506 688639
rect 42452 688598 42454 688607
rect 42506 688598 42508 688607
rect 42452 688533 42508 688542
rect 43234 687719 43262 706335
rect 43522 702773 43550 714179
rect 43606 714163 43658 714169
rect 43606 714105 43658 714111
rect 43618 704179 43646 714105
rect 43714 711399 43742 731009
rect 43798 717271 43850 717277
rect 43798 717213 43850 717219
rect 43700 711390 43756 711399
rect 43700 711325 43756 711334
rect 43810 706769 43838 717213
rect 43798 706763 43850 706769
rect 43798 706705 43850 706711
rect 43606 704173 43658 704179
rect 43606 704115 43658 704121
rect 43510 702767 43562 702773
rect 43510 702709 43562 702715
rect 43220 687710 43276 687719
rect 43220 687645 43276 687654
rect 43220 687562 43276 687571
rect 43220 687497 43276 687506
rect 41876 685490 41932 685499
rect 41876 685425 41932 685434
rect 40244 684306 40300 684315
rect 40244 684241 40300 684250
rect 35252 677202 35308 677211
rect 35252 677137 35308 677146
rect 35266 676767 35294 677137
rect 35252 676758 35308 676767
rect 35252 676693 35308 676702
rect 40258 673363 40286 684241
rect 41684 683714 41740 683723
rect 41684 683649 41740 683658
rect 41588 683122 41644 683131
rect 41588 683057 41644 683066
rect 40532 681050 40588 681059
rect 40532 680985 40588 680994
rect 40244 673354 40300 673363
rect 40244 673289 40300 673298
rect 40546 671143 40574 680985
rect 40628 679866 40684 679875
rect 40628 679801 40684 679810
rect 41492 679866 41548 679875
rect 41492 679801 41548 679810
rect 40532 671134 40588 671143
rect 40532 671069 40588 671078
rect 40642 670995 40670 679801
rect 40628 670986 40684 670995
rect 40628 670921 40684 670930
rect 41506 670879 41534 679801
rect 41602 670995 41630 683057
rect 41698 671027 41726 683649
rect 41686 671021 41738 671027
rect 41588 670986 41644 670995
rect 41686 670963 41738 670969
rect 41588 670921 41644 670930
rect 41494 670873 41546 670879
rect 41890 670824 41918 685425
rect 42452 684898 42508 684907
rect 42452 684833 42508 684842
rect 41972 682678 42028 682687
rect 41972 682613 42028 682622
rect 41494 670815 41546 670821
rect 41794 670796 41918 670824
rect 41794 670699 41822 670796
rect 41780 670690 41836 670699
rect 41986 670657 42014 682613
rect 42164 681494 42220 681503
rect 42164 681429 42220 681438
rect 42068 678386 42124 678395
rect 42068 678321 42124 678330
rect 42082 670657 42110 678321
rect 42178 671027 42206 681429
rect 42166 671021 42218 671027
rect 42166 670963 42218 670969
rect 41780 670625 41836 670634
rect 41974 670651 42026 670657
rect 41974 670593 42026 670599
rect 42070 670651 42122 670657
rect 42070 670593 42122 670599
rect 41974 670355 42026 670361
rect 41974 670297 42026 670303
rect 41986 669848 42014 670297
rect 42466 670139 42494 684833
rect 43028 680754 43084 680763
rect 43028 680689 43084 680698
rect 43042 670287 43070 680689
rect 43124 679126 43180 679135
rect 43124 679061 43180 679070
rect 43138 670847 43166 679061
rect 43124 670838 43180 670847
rect 43124 670773 43180 670782
rect 43126 670651 43178 670657
rect 43126 670593 43178 670599
rect 43030 670281 43082 670287
rect 43030 670223 43082 670229
rect 42454 670133 42506 670139
rect 42454 670075 42506 670081
rect 43030 670133 43082 670139
rect 43030 670075 43082 670081
rect 43042 668955 43070 670075
rect 43030 668949 43082 668955
rect 43030 668891 43082 668897
rect 42740 668618 42796 668627
rect 42166 668579 42218 668585
rect 42740 668553 42796 668562
rect 42166 668521 42218 668527
rect 42178 667998 42206 668521
rect 42166 667913 42218 667919
rect 42166 667855 42218 667861
rect 42178 667361 42206 667855
rect 42166 666729 42218 666735
rect 42166 666671 42218 666677
rect 42178 666148 42206 666671
rect 42166 665397 42218 665403
rect 42166 665339 42218 665345
rect 42178 664964 42206 665339
rect 41780 664622 41836 664631
rect 41780 664557 41836 664566
rect 41794 664298 41822 664557
rect 42164 664178 42220 664187
rect 42164 664113 42220 664122
rect 42178 664016 42206 664113
rect 42082 663988 42206 664016
rect 42082 663706 42110 663988
rect 42754 663553 42782 668553
rect 42838 668505 42890 668511
rect 42838 668447 42890 668453
rect 42850 666735 42878 668447
rect 42838 666729 42890 666735
rect 42838 666671 42890 666677
rect 42838 666581 42890 666587
rect 42838 666523 42890 666529
rect 42742 663547 42794 663553
rect 42742 663489 42794 663495
rect 42166 663399 42218 663405
rect 42166 663341 42218 663347
rect 42742 663399 42794 663405
rect 42742 663341 42794 663347
rect 42178 663114 42206 663341
rect 42452 662846 42508 662855
rect 42452 662781 42508 662790
rect 41780 661514 41836 661523
rect 41780 661449 41836 661458
rect 41794 661190 41822 661449
rect 41890 661375 41918 661856
rect 41876 661366 41932 661375
rect 41876 661301 41932 661310
rect 42070 661105 42122 661111
rect 42070 661047 42122 661053
rect 42082 660672 42110 661047
rect 41780 660330 41836 660339
rect 41780 660265 41836 660274
rect 41794 660006 41822 660265
rect 42166 659921 42218 659927
rect 42166 659863 42218 659869
rect 42178 659340 42206 659863
rect 42166 659255 42218 659261
rect 42166 659197 42218 659203
rect 42178 659132 42206 659197
rect 42082 659104 42206 659132
rect 42082 658822 42110 659104
rect 42466 657411 42494 662781
rect 42754 659927 42782 663341
rect 42850 661111 42878 666523
rect 43138 665403 43166 670593
rect 43126 665397 43178 665403
rect 43126 665339 43178 665345
rect 43126 665249 43178 665255
rect 43126 665191 43178 665197
rect 42838 661105 42890 661111
rect 42838 661047 42890 661053
rect 42742 659921 42794 659927
rect 42742 659863 42794 659869
rect 43138 659261 43166 665191
rect 43126 659255 43178 659261
rect 43126 659197 43178 659203
rect 43124 659146 43180 659155
rect 43124 659081 43180 659090
rect 42070 657405 42122 657411
rect 42070 657347 42122 657353
rect 42454 657405 42506 657411
rect 42454 657347 42506 657353
rect 42082 656972 42110 657347
rect 42934 656739 42986 656745
rect 42934 656681 42986 656687
rect 42166 656665 42218 656671
rect 42166 656607 42218 656613
rect 42178 656306 42206 656607
rect 42164 656186 42220 656195
rect 42164 656121 42220 656130
rect 42178 655677 42206 656121
rect 42946 646279 42974 656681
rect 43138 656671 43166 659081
rect 43126 656665 43178 656671
rect 43126 656607 43178 656613
rect 42932 646270 42988 646279
rect 42932 646205 42988 646214
rect 42452 645530 42508 645539
rect 42452 645465 42508 645474
rect 42466 645127 42494 645465
rect 42934 645269 42986 645275
rect 42932 645234 42934 645243
rect 42986 645234 42988 645243
rect 42932 645169 42988 645178
rect 42454 645121 42506 645127
rect 42454 645063 42506 645069
rect 43234 644503 43262 687497
rect 43414 673907 43466 673913
rect 43414 673849 43466 673855
rect 43426 670972 43454 673849
rect 43702 671021 43754 671027
rect 43426 670944 43646 670972
rect 43702 670963 43754 670969
rect 43414 670873 43466 670879
rect 43414 670815 43466 670821
rect 43318 670281 43370 670287
rect 43318 670223 43370 670229
rect 43330 668511 43358 670223
rect 43318 668505 43370 668511
rect 43318 668447 43370 668453
rect 43426 666587 43454 670815
rect 43510 670799 43562 670805
rect 43510 670741 43562 670747
rect 43414 666581 43466 666587
rect 43414 666523 43466 666529
rect 43522 665255 43550 670741
rect 43618 667919 43646 670944
rect 43606 667913 43658 667919
rect 43606 667855 43658 667861
rect 43510 665249 43562 665255
rect 43510 665191 43562 665197
rect 43714 663405 43742 670963
rect 43702 663399 43754 663405
rect 43702 663341 43754 663347
rect 43796 647158 43852 647167
rect 43796 647093 43852 647102
rect 43604 647010 43660 647019
rect 43604 646945 43660 646954
rect 43412 644642 43468 644651
rect 43412 644577 43468 644586
rect 43220 644494 43276 644503
rect 43220 644429 43276 644438
rect 41492 642274 41548 642283
rect 41492 642209 41548 642218
rect 39860 641090 39916 641099
rect 39860 641025 39916 641034
rect 35156 633986 35212 633995
rect 35156 633921 35212 633930
rect 35170 633551 35198 633921
rect 35156 633542 35212 633551
rect 35156 633477 35212 633486
rect 39874 627927 39902 641025
rect 40244 638870 40300 638879
rect 40244 638805 40300 638814
rect 40258 628075 40286 638805
rect 41300 638426 41356 638435
rect 41300 638361 41356 638370
rect 40244 628066 40300 628075
rect 40244 628001 40300 628010
rect 39860 627918 39916 627927
rect 39860 627853 39916 627862
rect 41314 627779 41342 638361
rect 41506 627927 41534 642209
rect 42932 641978 42988 641987
rect 42932 641913 42988 641922
rect 41588 640498 41644 640507
rect 41588 640433 41644 640442
rect 41492 627918 41548 627927
rect 41492 627853 41548 627862
rect 41602 627779 41630 640433
rect 41684 640054 41740 640063
rect 41684 639989 41740 639998
rect 41300 627770 41356 627779
rect 41300 627705 41356 627714
rect 41588 627770 41644 627779
rect 41698 627737 41726 639989
rect 41876 639462 41932 639471
rect 41876 639397 41932 639406
rect 41588 627705 41644 627714
rect 41686 627731 41738 627737
rect 41686 627673 41738 627679
rect 41890 627441 41918 639397
rect 42068 636798 42124 636807
rect 42068 636733 42124 636742
rect 41972 636206 42028 636215
rect 41972 636141 42028 636150
rect 41986 627483 42014 636141
rect 41972 627474 42028 627483
rect 41878 627435 41930 627441
rect 42082 627441 42110 636733
rect 42164 635614 42220 635623
rect 42164 635549 42220 635558
rect 42178 627663 42206 635549
rect 42166 627657 42218 627663
rect 42166 627599 42218 627605
rect 41972 627409 42028 627418
rect 42070 627435 42122 627441
rect 41878 627377 41930 627383
rect 42070 627377 42122 627383
rect 41878 627213 41930 627219
rect 41878 627155 41930 627161
rect 41890 626632 41918 627155
rect 42946 625369 42974 641913
rect 43124 638130 43180 638139
rect 43124 638065 43180 638074
rect 43028 635614 43084 635623
rect 43028 635549 43084 635558
rect 43042 627885 43070 635549
rect 43138 628033 43166 638065
rect 43426 630716 43454 644577
rect 43618 643023 43646 646945
rect 43810 643615 43838 647093
rect 43796 643606 43852 643615
rect 43796 643541 43852 643550
rect 43604 643014 43660 643023
rect 43604 642949 43660 642958
rect 43330 630688 43454 630716
rect 43126 628027 43178 628033
rect 43126 627969 43178 627975
rect 43030 627879 43082 627885
rect 43030 627821 43082 627827
rect 43030 627731 43082 627737
rect 43030 627673 43082 627679
rect 42166 625363 42218 625369
rect 42166 625305 42218 625311
rect 42934 625363 42986 625369
rect 42934 625305 42986 625311
rect 42178 624782 42206 625305
rect 42934 625215 42986 625221
rect 42934 625157 42986 625163
rect 42166 624697 42218 624703
rect 42166 624639 42218 624645
rect 42178 624161 42206 624639
rect 42164 623478 42220 623487
rect 42164 623413 42220 623422
rect 42178 622965 42206 623413
rect 42166 622255 42218 622261
rect 42166 622197 42218 622203
rect 42178 621748 42206 622197
rect 42166 621663 42218 621669
rect 42166 621605 42218 621611
rect 42178 621125 42206 621605
rect 42946 620929 42974 625157
rect 42070 620923 42122 620929
rect 42070 620865 42122 620871
rect 42934 620923 42986 620929
rect 42934 620865 42986 620871
rect 42082 620490 42110 620865
rect 43042 620411 43070 627673
rect 43126 627657 43178 627663
rect 43178 627605 43262 627608
rect 43126 627599 43262 627605
rect 43138 627580 43262 627599
rect 43126 627435 43178 627441
rect 43126 627377 43178 627383
rect 43138 621669 43166 627377
rect 43234 625221 43262 627580
rect 43222 625215 43274 625221
rect 43222 625157 43274 625163
rect 43126 621663 43178 621669
rect 43126 621605 43178 621611
rect 43124 621554 43180 621563
rect 43124 621489 43180 621498
rect 42166 620405 42218 620411
rect 42166 620347 42218 620353
rect 43030 620405 43082 620411
rect 43030 620347 43082 620353
rect 42178 619929 42206 620347
rect 42452 619630 42508 619639
rect 42452 619565 42508 619574
rect 41794 618455 41822 618640
rect 41780 618446 41836 618455
rect 41780 618381 41836 618390
rect 41780 618298 41836 618307
rect 41780 618233 41836 618242
rect 41794 617974 41822 618233
rect 41972 617854 42028 617863
rect 41972 617789 42028 617798
rect 41986 617456 42014 617789
rect 42166 617223 42218 617229
rect 42166 617165 42218 617171
rect 42178 616790 42206 617165
rect 41780 616670 41836 616679
rect 41780 616605 41836 616614
rect 41794 616157 41822 616605
rect 42466 616045 42494 619565
rect 42166 616039 42218 616045
rect 42166 615981 42218 615987
rect 42454 616039 42506 616045
rect 42454 615981 42506 615987
rect 42178 615606 42206 615981
rect 43138 614195 43166 621489
rect 42166 614189 42218 614195
rect 42166 614131 42218 614137
rect 43126 614189 43178 614195
rect 43126 614131 43178 614137
rect 42178 613756 42206 614131
rect 42164 613562 42220 613571
rect 42164 613497 42220 613506
rect 42838 613523 42890 613529
rect 42178 613121 42206 613497
rect 42838 613465 42890 613471
rect 41780 612822 41836 612831
rect 41780 612757 41836 612766
rect 41794 612498 41822 612757
rect 42850 603169 42878 613465
rect 42166 603163 42218 603169
rect 42166 603105 42218 603111
rect 42838 603163 42890 603169
rect 42838 603105 42890 603111
rect 42178 602175 42206 603105
rect 42836 603054 42892 603063
rect 42836 602989 42892 602998
rect 42740 602314 42796 602323
rect 42740 602249 42742 602258
rect 42794 602249 42796 602258
rect 42742 602217 42794 602223
rect 42164 602166 42220 602175
rect 42164 602101 42220 602110
rect 42850 601911 42878 602989
rect 42838 601905 42890 601911
rect 42838 601847 42890 601853
rect 43330 601287 43358 630688
rect 43510 627953 43562 627959
rect 43510 627895 43562 627901
rect 43414 627879 43466 627885
rect 43414 627821 43466 627827
rect 43426 622261 43454 627821
rect 43522 624703 43550 627895
rect 43510 624697 43562 624703
rect 43510 624639 43562 624645
rect 43414 622255 43466 622261
rect 43414 622197 43466 622203
rect 43316 601278 43372 601287
rect 43316 601213 43372 601222
rect 43618 599807 43646 642949
rect 43702 628027 43754 628033
rect 43702 627969 43754 627975
rect 43714 617229 43742 627969
rect 43702 617223 43754 617229
rect 43702 617165 43754 617171
rect 43810 600399 43838 643541
rect 43988 601426 44044 601435
rect 43988 601361 44044 601370
rect 43796 600390 43852 600399
rect 43796 600325 43852 600334
rect 43604 599798 43660 599807
rect 43604 599733 43660 599742
rect 43124 599206 43180 599215
rect 43124 599141 43180 599150
rect 41972 598466 42028 598475
rect 41972 598401 42028 598410
rect 41588 597282 41644 597291
rect 41588 597217 41644 597226
rect 41492 596838 41548 596847
rect 41492 596773 41548 596782
rect 41506 584521 41534 596773
rect 41602 584711 41630 597217
rect 41876 596246 41932 596255
rect 41876 596181 41932 596190
rect 41780 595210 41836 595219
rect 41780 595145 41836 595154
rect 41684 594618 41740 594627
rect 41684 594553 41740 594562
rect 41588 584702 41644 584711
rect 41588 584637 41644 584646
rect 41698 584563 41726 594553
rect 41684 584554 41740 584563
rect 41494 584515 41546 584521
rect 41684 584489 41740 584498
rect 41494 584457 41546 584463
rect 41794 584299 41822 595145
rect 41782 584293 41834 584299
rect 41782 584235 41834 584241
rect 41890 584225 41918 596181
rect 41986 584267 42014 598401
rect 42164 593582 42220 593591
rect 42164 593517 42220 593526
rect 42068 592990 42124 592999
rect 42068 592925 42124 592934
rect 42082 584415 42110 592925
rect 42068 584406 42124 584415
rect 42068 584341 42124 584350
rect 42178 584267 42206 593517
rect 42836 592768 42892 592777
rect 42836 592703 42892 592712
rect 42740 588402 42796 588411
rect 42740 588337 42796 588346
rect 42754 584392 42782 588337
rect 42850 584563 42878 592703
rect 43138 584836 43166 599141
rect 43138 584808 43550 584836
rect 43126 584737 43178 584743
rect 43126 584679 43178 584685
rect 42836 584554 42892 584563
rect 42836 584489 42892 584498
rect 42754 584364 42878 584392
rect 41972 584258 42028 584267
rect 41878 584219 41930 584225
rect 41972 584193 42028 584202
rect 42164 584258 42220 584267
rect 42164 584193 42220 584202
rect 41878 584161 41930 584167
rect 41878 583997 41930 584003
rect 41878 583939 41930 583945
rect 41890 583445 41918 583939
rect 42850 583855 42878 584364
rect 42838 583849 42890 583855
rect 42838 583791 42890 583797
rect 41876 582038 41932 582047
rect 41876 581973 41932 581982
rect 41890 581605 41918 581973
rect 43030 581555 43082 581561
rect 43030 581497 43082 581503
rect 42070 581481 42122 581487
rect 42070 581423 42122 581429
rect 42082 580974 42110 581423
rect 41780 580262 41836 580271
rect 41780 580197 41836 580206
rect 41794 579790 41822 580197
rect 43042 579045 43070 581497
rect 43138 581487 43166 584679
rect 43222 584515 43274 584521
rect 43222 584457 43274 584463
rect 43126 581481 43178 581487
rect 43126 581423 43178 581429
rect 43234 581284 43262 584457
rect 43414 584293 43466 584299
rect 43414 584235 43466 584241
rect 43318 583849 43370 583855
rect 43318 583791 43370 583797
rect 43330 581561 43358 583791
rect 43318 581555 43370 581561
rect 43318 581497 43370 581503
rect 43138 581256 43262 581284
rect 43138 579064 43166 581256
rect 42166 579039 42218 579045
rect 42166 578981 42218 578987
rect 43030 579039 43082 579045
rect 43138 579036 43262 579064
rect 43030 578981 43082 578987
rect 42178 578569 42206 578981
rect 43030 578891 43082 578897
rect 43030 578833 43082 578839
rect 42068 578486 42124 578495
rect 42068 578421 42124 578430
rect 42082 577940 42110 578421
rect 42932 578338 42988 578347
rect 42932 578273 42988 578282
rect 42164 577598 42220 577607
rect 42164 577533 42220 577542
rect 42178 577274 42206 577533
rect 42166 577189 42218 577195
rect 42166 577131 42218 577137
rect 42178 576992 42206 577131
rect 42082 576964 42206 576992
rect 42082 576756 42110 576964
rect 42082 574943 42110 575424
rect 42068 574934 42124 574943
rect 42068 574869 42124 574878
rect 41794 574499 41822 574797
rect 42068 574638 42124 574647
rect 42068 574573 42124 574582
rect 41780 574490 41836 574499
rect 41780 574425 41836 574434
rect 42082 574240 42110 574573
rect 41780 574046 41836 574055
rect 41780 573981 41836 573990
rect 41794 573574 41822 573981
rect 42166 573489 42218 573495
rect 42166 573431 42218 573437
rect 42178 573292 42206 573431
rect 42082 573264 42206 573292
rect 42082 572982 42110 573264
rect 42946 572681 42974 578273
rect 43042 573495 43070 578833
rect 43234 578768 43262 579036
rect 43426 578897 43454 584235
rect 43414 578891 43466 578897
rect 43414 578833 43466 578839
rect 43138 578740 43262 578768
rect 43138 577195 43166 578740
rect 43522 577732 43550 584808
rect 43234 577704 43550 577732
rect 43126 577189 43178 577195
rect 43126 577131 43178 577137
rect 43234 576992 43262 577704
rect 43618 577584 43646 599733
rect 43138 576964 43262 576992
rect 43522 577556 43646 577584
rect 43030 573489 43082 573495
rect 43030 573431 43082 573437
rect 42166 572675 42218 572681
rect 42166 572617 42218 572623
rect 42934 572675 42986 572681
rect 42934 572617 42986 572623
rect 42178 572390 42206 572617
rect 43138 571053 43166 576964
rect 43220 573158 43276 573167
rect 43220 573093 43276 573102
rect 42166 571047 42218 571053
rect 42166 570989 42218 570995
rect 43126 571047 43178 571053
rect 43126 570989 43178 570995
rect 42178 570540 42206 570989
rect 43234 570924 43262 573093
rect 43138 570896 43262 570924
rect 41780 570494 41836 570503
rect 41780 570429 41836 570438
rect 41794 569948 41822 570429
rect 42934 570307 42986 570313
rect 42934 570249 42986 570255
rect 42070 569715 42122 569721
rect 42070 569657 42122 569663
rect 42082 569282 42110 569657
rect 42836 559690 42892 559699
rect 42836 559625 42892 559634
rect 42850 558917 42878 559625
rect 42838 558911 42890 558917
rect 42838 558853 42890 558859
rect 42946 558811 42974 570249
rect 43138 569721 43166 570896
rect 43126 569715 43178 569721
rect 43126 569657 43178 569663
rect 43028 559394 43084 559403
rect 43028 559329 43030 559338
rect 43082 559329 43084 559338
rect 43030 559297 43082 559303
rect 43522 559107 43550 577556
rect 43508 559098 43564 559107
rect 43508 559033 43564 559042
rect 42932 558802 42988 558811
rect 42932 558737 42988 558746
rect 43412 557174 43468 557183
rect 43412 557109 43468 557118
rect 41588 555842 41644 555851
rect 41588 555777 41644 555786
rect 41492 554066 41548 554075
rect 41492 554001 41548 554010
rect 41396 549774 41452 549783
rect 41396 549709 41452 549718
rect 35156 547554 35212 547563
rect 35156 547489 35212 547498
rect 35170 547119 35198 547489
rect 35156 547110 35212 547119
rect 35156 547045 35212 547054
rect 41410 541347 41438 549709
rect 41506 541495 41534 554001
rect 41492 541486 41548 541495
rect 41492 541421 41548 541430
rect 41396 541338 41452 541347
rect 41602 541305 41630 555777
rect 41876 555250 41932 555259
rect 41876 555185 41932 555194
rect 41780 551402 41836 551411
rect 41780 551337 41836 551346
rect 41684 549182 41740 549191
rect 41684 549117 41740 549126
rect 41698 541347 41726 549117
rect 41684 541338 41740 541347
rect 41396 541273 41452 541282
rect 41590 541299 41642 541305
rect 41684 541273 41740 541282
rect 41590 541241 41642 541247
rect 41794 541051 41822 551337
rect 41890 544265 41918 555185
rect 42164 553622 42220 553631
rect 42164 553557 42220 553566
rect 41972 551994 42028 552003
rect 41972 551929 42028 551938
rect 41878 544259 41930 544265
rect 41878 544201 41930 544207
rect 41780 541042 41836 541051
rect 41986 541009 42014 551929
rect 42068 550366 42124 550375
rect 42068 550301 42124 550310
rect 42082 541231 42110 550301
rect 42070 541225 42122 541231
rect 42178 541199 42206 553557
rect 42452 553030 42508 553039
rect 42452 552965 42508 552974
rect 42070 541167 42122 541173
rect 42164 541190 42220 541199
rect 42466 541157 42494 552965
rect 43124 550810 43180 550819
rect 43124 550745 43180 550754
rect 43138 549168 43166 550745
rect 43042 549140 43166 549168
rect 42934 544259 42986 544265
rect 42934 544201 42986 544207
rect 42164 541125 42220 541134
rect 42454 541151 42506 541157
rect 42454 541093 42506 541099
rect 41780 540977 41836 540986
rect 41974 541003 42026 541009
rect 41974 540945 42026 540951
rect 42454 541003 42506 541009
rect 42454 540945 42506 540951
rect 42466 540880 42494 540945
rect 42466 540852 42590 540880
rect 42166 540781 42218 540787
rect 42166 540723 42218 540729
rect 42178 540245 42206 540723
rect 42070 538931 42122 538937
rect 42070 538873 42122 538879
rect 42082 538424 42110 538873
rect 42166 538191 42218 538197
rect 42166 538133 42218 538139
rect 42178 537758 42206 538133
rect 42068 537046 42124 537055
rect 42068 536981 42124 536990
rect 42082 536574 42110 536981
rect 42070 535823 42122 535829
rect 42070 535765 42122 535771
rect 42082 535390 42110 535765
rect 42166 535083 42218 535089
rect 42166 535025 42218 535031
rect 42178 534724 42206 535025
rect 41780 534382 41836 534391
rect 41780 534317 41836 534326
rect 41794 534058 41822 534317
rect 41972 533790 42028 533799
rect 41972 533725 42028 533734
rect 41986 533540 42014 533725
rect 42562 533332 42590 540852
rect 42946 538937 42974 544201
rect 43042 541643 43070 549140
rect 43124 549034 43180 549043
rect 43124 548969 43180 548978
rect 43028 541634 43084 541643
rect 43028 541569 43084 541578
rect 43030 541521 43082 541527
rect 43030 541463 43082 541469
rect 42934 538931 42986 538937
rect 42934 538873 42986 538879
rect 42934 538783 42986 538789
rect 42934 538725 42986 538731
rect 42946 535089 42974 538725
rect 43042 538197 43070 541463
rect 43030 538191 43082 538197
rect 43030 538133 43082 538139
rect 43028 538082 43084 538091
rect 43028 538017 43084 538026
rect 42934 535083 42986 535089
rect 42934 535025 42986 535031
rect 42466 533304 42590 533332
rect 42068 532754 42124 532763
rect 42068 532689 42124 532698
rect 42082 532241 42110 532689
rect 41780 531866 41836 531875
rect 41780 531801 41836 531810
rect 41794 531616 41822 531801
rect 41780 531274 41836 531283
rect 41780 531209 41836 531218
rect 41794 531024 41822 531209
rect 42166 530939 42218 530945
rect 42166 530881 42218 530887
rect 42178 530401 42206 530881
rect 42466 530279 42494 533304
rect 42932 532606 42988 532615
rect 42932 532541 42988 532550
rect 42070 530273 42122 530279
rect 42070 530215 42122 530221
rect 42454 530273 42506 530279
rect 42454 530215 42506 530221
rect 42082 529766 42110 530215
rect 42454 530125 42506 530131
rect 42454 530067 42506 530073
rect 42164 529498 42220 529507
rect 42164 529433 42220 529442
rect 42178 529205 42206 529433
rect 42466 529243 42494 530067
rect 42946 529391 42974 532541
rect 43042 530945 43070 538017
rect 43138 535829 43166 548969
rect 43222 541225 43274 541231
rect 43222 541167 43274 541173
rect 43234 538789 43262 541167
rect 43222 538783 43274 538789
rect 43222 538725 43274 538731
rect 43126 535823 43178 535829
rect 43126 535765 43178 535771
rect 43126 535675 43178 535681
rect 43126 535617 43178 535623
rect 43030 530939 43082 530945
rect 43030 530881 43082 530887
rect 43138 530205 43166 535617
rect 43126 530199 43178 530205
rect 43126 530141 43178 530147
rect 43028 530090 43084 530099
rect 43084 530048 43166 530076
rect 43028 530025 43084 530034
rect 43030 529977 43082 529983
rect 43030 529919 43082 529925
rect 42934 529385 42986 529391
rect 42934 529327 42986 529333
rect 42454 529237 42506 529243
rect 42454 529179 42506 529185
rect 42934 529237 42986 529243
rect 42934 529179 42986 529185
rect 42838 528941 42890 528947
rect 42838 528883 42890 528889
rect 42166 527683 42218 527689
rect 42166 527625 42218 527631
rect 42178 527365 42206 527625
rect 42070 527091 42122 527097
rect 42070 527033 42122 527039
rect 42082 526732 42110 527033
rect 42850 526505 42878 528883
rect 42946 527689 42974 529179
rect 42934 527683 42986 527689
rect 42934 527625 42986 527631
rect 42166 526499 42218 526505
rect 42166 526441 42218 526447
rect 42838 526499 42890 526505
rect 42838 526441 42890 526447
rect 42178 526066 42206 526441
rect 43042 519845 43070 529919
rect 43138 529539 43166 530048
rect 43318 530051 43370 530057
rect 43318 529993 43370 529999
rect 43126 529533 43178 529539
rect 43126 529475 43178 529481
rect 43126 529385 43178 529391
rect 43126 529327 43178 529333
rect 43138 527097 43166 529327
rect 43126 527091 43178 527097
rect 43126 527033 43178 527039
rect 43330 524179 43358 529993
rect 43124 524170 43180 524179
rect 43124 524105 43180 524114
rect 43316 524170 43372 524179
rect 43316 524105 43372 524114
rect 41878 519839 41930 519845
rect 41878 519781 41930 519787
rect 43030 519839 43082 519845
rect 43030 519781 43082 519787
rect 41890 431383 41918 519781
rect 42164 509962 42220 509971
rect 42164 509897 42220 509906
rect 42178 504051 42206 509897
rect 43138 509781 43166 524105
rect 43126 509775 43178 509781
rect 43126 509717 43178 509723
rect 43318 509775 43370 509781
rect 43318 509717 43370 509723
rect 42164 504042 42220 504051
rect 42164 503977 42220 503986
rect 42068 483766 42124 483775
rect 42068 483701 42124 483710
rect 42082 463943 42110 483701
rect 43330 469451 43358 509717
rect 43318 469445 43370 469451
rect 43318 469387 43370 469393
rect 42068 463934 42124 463943
rect 42068 463869 42124 463878
rect 43222 449317 43274 449323
rect 43222 449259 43274 449265
rect 42838 432297 42890 432303
rect 42836 432262 42838 432271
rect 42890 432262 42892 432271
rect 42836 432197 42892 432206
rect 42550 432001 42602 432007
rect 42548 431966 42550 431975
rect 42602 431966 42604 431975
rect 42548 431901 42604 431910
rect 41876 431374 41932 431383
rect 41876 431309 41932 431318
rect 42932 430634 42988 430643
rect 42932 430569 42988 430578
rect 42548 427674 42604 427683
rect 42604 427632 42686 427660
rect 42548 427609 42604 427618
rect 40244 425454 40300 425463
rect 40244 425389 40300 425398
rect 39956 422790 40012 422799
rect 39956 422725 40012 422734
rect 35156 419978 35212 419987
rect 35156 419913 35212 419922
rect 35170 419543 35198 419913
rect 35156 419534 35212 419543
rect 35156 419469 35212 419478
rect 39970 415949 39998 422725
rect 40148 422198 40204 422207
rect 40148 422133 40204 422142
rect 40052 421606 40108 421615
rect 40052 421541 40108 421550
rect 39958 415943 40010 415949
rect 39958 415885 40010 415891
rect 40066 415431 40094 421541
rect 40054 415425 40106 415431
rect 40054 415367 40106 415373
rect 40162 414765 40190 422133
rect 40258 420537 40286 425389
rect 42356 423382 42412 423391
rect 42356 423317 42412 423326
rect 40246 420531 40298 420537
rect 40246 420473 40298 420479
rect 41782 420531 41834 420537
rect 41782 420473 41834 420479
rect 40150 414759 40202 414765
rect 40150 414701 40202 414707
rect 41794 413433 41822 420473
rect 41782 413427 41834 413433
rect 41782 413369 41834 413375
rect 41782 413205 41834 413211
rect 41782 413147 41834 413153
rect 41794 412624 41822 413147
rect 42166 410985 42218 410991
rect 42166 410927 42218 410933
rect 42178 410805 42206 410927
rect 42178 409733 42206 410182
rect 42166 409727 42218 409733
rect 42166 409669 42218 409675
rect 42370 409511 42398 423317
rect 42452 419534 42508 419543
rect 42452 419469 42508 419478
rect 42466 417651 42494 419469
rect 42454 417645 42506 417651
rect 42454 417587 42506 417593
rect 42454 415943 42506 415949
rect 42454 415885 42506 415891
rect 42466 411435 42494 415885
rect 42454 411429 42506 411435
rect 42454 411371 42506 411377
rect 42658 411232 42686 427632
rect 42946 423423 42974 430569
rect 43234 430199 43262 449259
rect 43220 430190 43276 430199
rect 43220 430125 43276 430134
rect 43124 429746 43180 429755
rect 43426 429732 43454 557109
rect 43180 429704 43454 429732
rect 43124 429681 43180 429690
rect 43522 429015 43550 559033
rect 43700 558506 43756 558515
rect 43700 558441 43756 558450
rect 43606 541299 43658 541305
rect 43606 541241 43658 541247
rect 43618 535681 43646 541241
rect 43606 535675 43658 535681
rect 43606 535617 43658 535623
rect 43714 530057 43742 558441
rect 43810 557183 43838 600325
rect 44002 558071 44030 601361
rect 43988 558062 44044 558071
rect 43988 557997 44044 558006
rect 43796 557174 43852 557183
rect 43796 557109 43852 557118
rect 44564 547406 44620 547415
rect 44564 547341 44620 547350
rect 43702 530051 43754 530057
rect 43702 529993 43754 529999
rect 43606 469445 43658 469451
rect 43606 469387 43658 469393
rect 43618 449323 43646 469387
rect 43606 449317 43658 449323
rect 43606 449259 43658 449265
rect 43508 429006 43564 429015
rect 43508 428941 43564 428950
rect 43124 424122 43180 424131
rect 43124 424057 43180 424066
rect 42934 423417 42986 423423
rect 42934 423359 42986 423365
rect 42932 421458 42988 421467
rect 42932 421393 42988 421402
rect 42562 411204 42686 411232
rect 42562 410991 42590 411204
rect 42550 410985 42602 410991
rect 42550 410927 42602 410933
rect 42550 409727 42602 409733
rect 42550 409669 42602 409675
rect 42166 409505 42218 409511
rect 42166 409447 42218 409453
rect 42358 409505 42410 409511
rect 42358 409447 42410 409453
rect 42178 408965 42206 409447
rect 42358 409357 42410 409363
rect 42358 409299 42410 409305
rect 42370 408253 42398 409299
rect 42166 408247 42218 408253
rect 42166 408189 42218 408195
rect 42358 408247 42410 408253
rect 42358 408189 42410 408195
rect 42178 407769 42206 408189
rect 42356 408138 42412 408147
rect 42356 408073 42412 408082
rect 42070 407507 42122 407513
rect 42070 407449 42122 407455
rect 42082 407148 42110 407449
rect 42166 407063 42218 407069
rect 42166 407005 42218 407011
rect 42178 406482 42206 407005
rect 42068 406066 42124 406075
rect 42068 406001 42124 406010
rect 42082 405929 42110 406001
rect 42082 404299 42110 404632
rect 42068 404290 42124 404299
rect 42068 404225 42124 404234
rect 41794 403855 41822 403997
rect 41780 403846 41836 403855
rect 41780 403781 41836 403790
rect 42370 403462 42398 408073
rect 42562 406107 42590 409669
rect 42946 409363 42974 421393
rect 43138 415524 43166 424057
rect 43702 423417 43754 423423
rect 43702 423359 43754 423365
rect 43138 415496 43358 415524
rect 43126 415425 43178 415431
rect 43126 415367 43178 415373
rect 43030 414759 43082 414765
rect 43030 414701 43082 414707
rect 42934 409357 42986 409363
rect 43042 409331 43070 414701
rect 42934 409299 42986 409305
rect 43028 409322 43084 409331
rect 43028 409257 43084 409266
rect 43138 409160 43166 415367
rect 43222 411429 43274 411435
rect 43222 411371 43274 411377
rect 42946 409132 43166 409160
rect 42946 407069 42974 409132
rect 43030 409061 43082 409067
rect 43234 409012 43262 411371
rect 43330 409141 43358 415496
rect 43318 409135 43370 409141
rect 43318 409077 43370 409083
rect 43030 409003 43082 409009
rect 42934 407063 42986 407069
rect 42934 407005 42986 407011
rect 42550 406101 42602 406107
rect 42550 406043 42602 406049
rect 42192 403434 42398 403462
rect 43042 403221 43070 409003
rect 43138 408984 43262 409012
rect 43138 407513 43166 408984
rect 43714 408979 43742 423359
rect 43330 408951 43742 408979
rect 43126 407507 43178 407513
rect 43126 407449 43178 407455
rect 43330 403221 43358 408951
rect 42166 403215 42218 403221
rect 42166 403157 42218 403163
rect 43030 403215 43082 403221
rect 43030 403157 43082 403163
rect 43318 403215 43370 403221
rect 43318 403157 43370 403163
rect 42178 402782 42206 403157
rect 42934 403141 42986 403147
rect 42934 403083 42986 403089
rect 41780 402662 41836 402671
rect 41780 402597 41836 402606
rect 41794 402157 41822 402597
rect 41780 401922 41836 401931
rect 41780 401857 41836 401866
rect 41794 401598 41822 401857
rect 41780 400146 41836 400155
rect 41780 400081 41836 400090
rect 41794 399748 41822 400081
rect 41780 399554 41836 399563
rect 41780 399489 41836 399498
rect 41794 399121 41822 399489
rect 41780 398814 41836 398823
rect 41780 398749 41836 398758
rect 41794 398490 41822 398749
rect 42358 389377 42410 389383
rect 42356 389342 42358 389351
rect 42410 389342 42412 389351
rect 42356 389277 42412 389286
rect 42646 388785 42698 388791
rect 42644 388750 42646 388759
rect 42698 388750 42700 388759
rect 42644 388685 42700 388694
rect 42646 388045 42698 388051
rect 42644 388010 42646 388019
rect 42698 388010 42700 388019
rect 42644 387945 42700 387954
rect 42946 387131 42974 403083
rect 43412 387270 43468 387279
rect 43412 387205 43468 387214
rect 42932 387122 42988 387131
rect 42932 387057 42988 387066
rect 42740 384754 42796 384763
rect 42740 384689 42796 384698
rect 42356 382238 42412 382247
rect 42356 382173 42412 382182
rect 39956 380610 40012 380619
rect 39956 380545 40012 380554
rect 35156 376762 35212 376771
rect 35156 376697 35212 376706
rect 35170 376327 35198 376697
rect 35156 376318 35212 376327
rect 35156 376253 35212 376262
rect 39970 371623 39998 380545
rect 40052 380166 40108 380175
rect 40052 380101 40108 380110
rect 40066 374361 40094 380101
rect 40244 378390 40300 378399
rect 40244 378325 40300 378334
rect 40054 374355 40106 374361
rect 40054 374297 40106 374303
rect 40258 373695 40286 378325
rect 40246 373689 40298 373695
rect 40246 373631 40298 373637
rect 39958 371617 40010 371623
rect 39958 371559 40010 371565
rect 42370 369995 42398 382173
rect 42644 377650 42700 377659
rect 42644 377585 42700 377594
rect 42658 376623 42686 377585
rect 42644 376614 42700 376623
rect 42644 376549 42646 376558
rect 42698 376549 42700 376558
rect 42646 376517 42698 376523
rect 42754 370513 42782 384689
rect 43028 379870 43084 379879
rect 43028 379805 43084 379814
rect 42932 378242 42988 378251
rect 42932 378177 42988 378186
rect 42838 373689 42890 373695
rect 42838 373631 42890 373637
rect 42742 370507 42794 370513
rect 42742 370449 42794 370455
rect 42166 369989 42218 369995
rect 42166 369931 42218 369937
rect 42358 369989 42410 369995
rect 42358 369931 42410 369937
rect 42178 369445 42206 369931
rect 42850 369847 42878 373631
rect 42358 369841 42410 369847
rect 42358 369783 42410 369789
rect 42838 369841 42890 369847
rect 42838 369783 42890 369789
rect 42070 368139 42122 368145
rect 42070 368081 42122 368087
rect 42082 367632 42110 368081
rect 42070 367399 42122 367405
rect 42070 367341 42122 367347
rect 42082 366966 42110 367341
rect 42070 366289 42122 366295
rect 42070 366231 42122 366237
rect 42082 365782 42110 366231
rect 42166 365031 42218 365037
rect 42166 364973 42218 364979
rect 42178 364569 42206 364973
rect 42070 364291 42122 364297
rect 42070 364233 42122 364239
rect 42082 363932 42110 364233
rect 42370 363853 42398 369783
rect 42946 369644 42974 378177
rect 42850 369616 42974 369644
rect 42850 365037 42878 369616
rect 42934 369545 42986 369551
rect 42934 369487 42986 369493
rect 42946 366295 42974 369487
rect 42934 366289 42986 366295
rect 42934 366231 42986 366237
rect 42838 365031 42890 365037
rect 42838 364973 42890 364979
rect 43042 364297 43070 379805
rect 43126 374355 43178 374361
rect 43126 374297 43178 374303
rect 43138 369551 43166 374297
rect 43318 371617 43370 371623
rect 43318 371559 43370 371565
rect 43222 370507 43274 370513
rect 43222 370449 43274 370455
rect 43126 369545 43178 369551
rect 43126 369487 43178 369493
rect 43234 369348 43262 370449
rect 43138 369320 43262 369348
rect 43138 368145 43166 369320
rect 43222 369249 43274 369255
rect 43222 369191 43274 369197
rect 43234 368145 43262 369191
rect 43126 368139 43178 368145
rect 43126 368081 43178 368087
rect 43222 368139 43274 368145
rect 43222 368081 43274 368087
rect 43330 368016 43358 371559
rect 43426 369255 43454 387205
rect 43414 369249 43466 369255
rect 43414 369191 43466 369197
rect 43138 367988 43358 368016
rect 43030 364291 43082 364297
rect 43030 364233 43082 364239
rect 42166 363847 42218 363853
rect 42166 363789 42218 363795
rect 42358 363847 42410 363853
rect 42358 363789 42410 363795
rect 42178 363266 42206 363789
rect 41780 362850 41836 362859
rect 41780 362785 41836 362794
rect 41794 362748 41822 362785
rect 42164 361962 42220 361971
rect 42164 361897 42220 361906
rect 42178 361416 42206 361897
rect 42260 361222 42316 361231
rect 42260 361157 42316 361166
rect 42178 360639 42206 360824
rect 42164 360630 42220 360639
rect 42164 360565 42220 360574
rect 42274 360246 42302 361157
rect 42192 360218 42302 360246
rect 43138 360153 43166 367988
rect 43222 367917 43274 367923
rect 43222 367859 43274 367865
rect 42166 360147 42218 360153
rect 42166 360089 42218 360095
rect 43126 360147 43178 360153
rect 43126 360089 43178 360095
rect 42178 359601 42206 360089
rect 42068 359446 42124 359455
rect 42068 359381 42124 359390
rect 42082 358974 42110 359381
rect 41780 358706 41836 358715
rect 41780 358641 41836 358650
rect 41794 358382 41822 358641
rect 41780 356930 41836 356939
rect 41780 356865 41836 356874
rect 41794 356565 41822 356865
rect 41780 356486 41836 356495
rect 41780 356421 41836 356430
rect 41794 355940 41822 356421
rect 41780 355598 41836 355607
rect 41780 355533 41836 355542
rect 41794 355274 41822 355533
rect 42838 345939 42890 345945
rect 42836 345904 42838 345913
rect 42890 345904 42892 345913
rect 42836 345839 42892 345848
rect 42838 345421 42890 345427
rect 42836 345386 42838 345395
rect 42890 345386 42892 345395
rect 42836 345321 42892 345330
rect 42838 344829 42890 344835
rect 42836 344794 42838 344803
rect 42890 344794 42892 344803
rect 42836 344729 42892 344738
rect 43234 343767 43262 367859
rect 43412 344202 43468 344211
rect 43412 344137 43468 344146
rect 43220 343758 43276 343767
rect 43220 343693 43276 343702
rect 42836 341538 42892 341547
rect 42836 341473 42892 341482
rect 41780 339022 41836 339031
rect 41780 338957 41836 338966
rect 40052 336950 40108 336959
rect 40052 336885 40108 336894
rect 35156 333546 35212 333555
rect 35156 333481 35212 333490
rect 35170 333111 35198 333481
rect 35156 333102 35212 333111
rect 35156 333037 35212 333046
rect 40066 329369 40094 336885
rect 40148 336358 40204 336367
rect 40148 336293 40204 336302
rect 40162 329591 40190 336293
rect 40150 329585 40202 329591
rect 40150 329527 40202 329533
rect 40054 329363 40106 329369
rect 40054 329305 40106 329311
rect 41794 327075 41822 338957
rect 42260 337542 42316 337551
rect 42260 337477 42316 337486
rect 41782 327069 41834 327075
rect 41782 327011 41834 327017
rect 42274 327001 42302 337477
rect 42548 334730 42604 334739
rect 42548 334665 42604 334674
rect 42262 326995 42314 327001
rect 42262 326937 42314 326943
rect 41782 326773 41834 326779
rect 41782 326715 41834 326721
rect 41794 326266 41822 326715
rect 42070 324923 42122 324929
rect 42070 324865 42122 324871
rect 42082 324416 42110 324865
rect 42166 324183 42218 324189
rect 42166 324125 42218 324131
rect 42178 323750 42206 324125
rect 42166 323147 42218 323153
rect 42166 323089 42218 323095
rect 42178 322566 42206 323089
rect 42562 321821 42590 334665
rect 42850 324929 42878 341473
rect 43220 333398 43276 333407
rect 43220 333333 43276 333342
rect 43234 332255 43262 333333
rect 43222 332249 43274 332255
rect 43222 332191 43274 332197
rect 43030 329585 43082 329591
rect 43030 329527 43082 329533
rect 42934 326995 42986 327001
rect 42934 326937 42986 326943
rect 42838 324923 42890 324929
rect 42838 324865 42890 324871
rect 42836 324814 42892 324823
rect 42836 324749 42892 324758
rect 42070 321815 42122 321821
rect 42070 321757 42122 321763
rect 42550 321815 42602 321821
rect 42550 321757 42602 321763
rect 42082 321382 42110 321757
rect 42166 321075 42218 321081
rect 42166 321017 42218 321023
rect 42178 320716 42206 321017
rect 41780 320522 41836 320531
rect 41780 320457 41836 320466
rect 41794 320081 41822 320457
rect 42068 319782 42124 319791
rect 42068 319717 42124 319726
rect 42082 319532 42110 319717
rect 42850 318787 42878 324749
rect 42262 318781 42314 318787
rect 42262 318723 42314 318729
rect 42838 318781 42890 318787
rect 42838 318723 42890 318729
rect 42164 318450 42220 318459
rect 42164 318385 42220 318394
rect 42178 318241 42206 318385
rect 42068 318006 42124 318015
rect 42068 317941 42124 317950
rect 42082 317608 42110 317941
rect 42274 317059 42302 318723
rect 42192 317031 42302 317059
rect 42946 316937 42974 326937
rect 43042 321081 43070 329527
rect 43126 329363 43178 329369
rect 43126 329305 43178 329311
rect 43138 323153 43166 329305
rect 43426 328352 43454 344137
rect 43234 328324 43454 328352
rect 43126 323147 43178 323153
rect 43126 323089 43178 323095
rect 43030 321075 43082 321081
rect 43030 321017 43082 321023
rect 42070 316931 42122 316937
rect 42070 316873 42122 316879
rect 42934 316931 42986 316937
rect 42934 316873 42986 316879
rect 42082 316424 42110 316873
rect 41780 316230 41836 316239
rect 41780 316165 41836 316174
rect 41794 315758 41822 316165
rect 41780 315490 41836 315499
rect 41780 315425 41836 315434
rect 41794 315205 41822 315425
rect 41876 313714 41932 313723
rect 41876 313649 41932 313658
rect 41890 313390 41918 313649
rect 41780 313270 41836 313279
rect 41780 313205 41836 313214
rect 41794 312724 41822 313205
rect 41780 312382 41836 312391
rect 41780 312317 41836 312326
rect 41794 312058 41822 312317
rect 42838 302723 42890 302729
rect 42836 302688 42838 302697
rect 42890 302688 42892 302697
rect 42836 302623 42892 302632
rect 42454 302353 42506 302359
rect 42452 302318 42454 302327
rect 42506 302318 42508 302327
rect 42452 302253 42508 302262
rect 42838 301687 42890 301693
rect 42838 301629 42890 301635
rect 42850 301587 42878 301629
rect 42836 301578 42892 301587
rect 42836 301513 42892 301522
rect 43124 300986 43180 300995
rect 43124 300921 43180 300930
rect 43138 300380 43166 300921
rect 43234 300551 43262 328324
rect 43220 300542 43276 300551
rect 43220 300477 43276 300486
rect 43138 300352 43262 300380
rect 41780 298026 41836 298035
rect 41780 297961 41836 297970
rect 40244 293734 40300 293743
rect 40244 293669 40300 293678
rect 40052 293142 40108 293151
rect 40052 293077 40108 293086
rect 39956 292550 40012 292559
rect 39956 292485 40012 292494
rect 35156 290478 35212 290487
rect 35156 290413 35212 290422
rect 35170 289895 35198 290413
rect 35156 289886 35212 289895
rect 35156 289821 35212 289830
rect 39970 285413 39998 292485
rect 39958 285407 40010 285413
rect 39958 285349 40010 285355
rect 40066 285339 40094 293077
rect 40148 292106 40204 292115
rect 40148 292041 40204 292050
rect 40054 285333 40106 285339
rect 40054 285275 40106 285281
rect 40162 285265 40190 292041
rect 40150 285259 40202 285265
rect 40150 285201 40202 285207
rect 40258 285191 40286 293669
rect 40246 285185 40298 285191
rect 40246 285127 40298 285133
rect 41794 284544 41822 297961
rect 42260 295806 42316 295815
rect 42260 295741 42316 295750
rect 42274 284692 42302 295741
rect 42356 294326 42412 294335
rect 42356 294261 42412 294270
rect 42370 284863 42398 294261
rect 42836 290182 42892 290191
rect 42836 290117 42838 290126
rect 42890 290117 42892 290126
rect 42838 290085 42890 290091
rect 43126 285333 43178 285339
rect 43126 285275 43178 285281
rect 43030 285259 43082 285265
rect 43030 285201 43082 285207
rect 42934 285185 42986 285191
rect 42934 285127 42986 285133
rect 42356 284854 42412 284863
rect 42356 284789 42412 284798
rect 42274 284664 42494 284692
rect 41794 284516 42398 284544
rect 42178 282971 42206 283050
rect 42166 282965 42218 282971
rect 42166 282907 42218 282913
rect 42370 281787 42398 284516
rect 42466 282971 42494 284664
rect 42454 282965 42506 282971
rect 42454 282907 42506 282913
rect 42166 281781 42218 281787
rect 42166 281723 42218 281729
rect 42358 281781 42410 281787
rect 42358 281723 42410 281729
rect 42178 281200 42206 281723
rect 42356 281598 42412 281607
rect 42356 281533 42412 281542
rect 42166 281115 42218 281121
rect 42166 281057 42218 281063
rect 42178 280534 42206 281057
rect 42166 279931 42218 279937
rect 42166 279873 42218 279879
rect 42178 279350 42206 279873
rect 42164 278638 42220 278647
rect 42164 278573 42220 278582
rect 42178 278166 42206 278573
rect 42166 277859 42218 277865
rect 42166 277801 42218 277807
rect 42178 277500 42206 277801
rect 42070 277415 42122 277421
rect 42070 277357 42122 277363
rect 42082 276908 42110 277357
rect 42068 276566 42124 276575
rect 42068 276501 42124 276510
rect 42082 276316 42110 276501
rect 42262 275491 42314 275497
rect 42262 275433 42314 275439
rect 41972 274790 42028 274799
rect 41972 274725 42028 274734
rect 41986 274392 42014 274725
rect 42178 274651 42206 275058
rect 42164 274642 42220 274651
rect 42164 274577 42220 274586
rect 42274 273859 42302 275433
rect 42192 273831 42302 273859
rect 42370 273222 42398 281533
rect 42946 279937 42974 285127
rect 42934 279931 42986 279937
rect 42934 279873 42986 279879
rect 42934 279783 42986 279789
rect 42934 279725 42986 279731
rect 42946 275497 42974 279725
rect 43042 277421 43070 285201
rect 43138 277865 43166 285275
rect 43126 277859 43178 277865
rect 43126 277801 43178 277807
rect 43030 277415 43082 277421
rect 43030 277357 43082 277363
rect 42934 275491 42986 275497
rect 42934 275433 42986 275439
rect 42192 273194 42398 273222
rect 41780 273014 41836 273023
rect 41780 272949 41836 272958
rect 41794 272542 41822 272949
rect 41780 272274 41836 272283
rect 41780 272209 41836 272218
rect 41794 272024 41822 272209
rect 41780 270646 41836 270655
rect 41780 270581 41836 270590
rect 43124 270646 43180 270655
rect 43124 270581 43180 270590
rect 41794 270174 41822 270581
rect 41780 270054 41836 270063
rect 41780 269989 41836 269998
rect 41794 269508 41822 269989
rect 41780 269166 41836 269175
rect 41780 269101 41836 269110
rect 41794 268877 41822 269101
rect 42550 259729 42602 259735
rect 42548 259694 42550 259703
rect 42602 259694 42604 259703
rect 42548 259629 42604 259638
rect 42646 258989 42698 258995
rect 42644 258954 42646 258963
rect 42698 258954 42700 258963
rect 42644 258889 42700 258898
rect 42550 258249 42602 258255
rect 42548 258214 42550 258223
rect 42602 258214 42604 258223
rect 42548 258149 42604 258158
rect 43138 257811 43166 270581
rect 42262 257805 42314 257811
rect 42262 257747 42314 257753
rect 43126 257805 43178 257811
rect 43126 257747 43178 257753
rect 41780 252590 41836 252599
rect 41780 252525 41836 252534
rect 40244 250518 40300 250527
rect 40244 250453 40300 250462
rect 39956 249926 40012 249935
rect 39956 249861 40012 249870
rect 35252 247262 35308 247271
rect 35252 247197 35308 247206
rect 35266 246827 35294 247197
rect 35252 246818 35308 246827
rect 35252 246753 35308 246762
rect 39970 242123 39998 249861
rect 40052 249334 40108 249343
rect 40052 249269 40108 249278
rect 40066 242197 40094 249269
rect 40148 248890 40204 248899
rect 40148 248825 40204 248834
rect 40054 242191 40106 242197
rect 40054 242133 40106 242139
rect 39958 242117 40010 242123
rect 39958 242059 40010 242065
rect 40162 242049 40190 248825
rect 40150 242043 40202 242049
rect 40150 241985 40202 241991
rect 40258 241975 40286 250453
rect 40246 241969 40298 241975
rect 40246 241911 40298 241917
rect 41794 240643 41822 252525
rect 42274 243867 42302 257747
rect 42548 257622 42604 257631
rect 42548 257557 42604 257566
rect 42562 257219 42590 257557
rect 43234 257335 43262 300352
rect 43318 285407 43370 285413
rect 43318 285349 43370 285355
rect 43330 279789 43358 285349
rect 43318 279783 43370 279789
rect 43318 279725 43370 279731
rect 43220 257326 43276 257335
rect 43220 257261 43276 257270
rect 42550 257213 42602 257219
rect 42550 257155 42602 257161
rect 43222 257213 43274 257219
rect 43222 257155 43274 257161
rect 43028 255106 43084 255115
rect 43028 255041 43084 255050
rect 42548 247854 42604 247863
rect 42548 247789 42604 247798
rect 42562 247271 42590 247789
rect 42548 247262 42604 247271
rect 42548 247197 42604 247206
rect 42562 244935 42590 247197
rect 42550 244929 42602 244935
rect 42550 244871 42602 244877
rect 42260 243858 42316 243867
rect 42260 243793 42316 243802
rect 42262 242191 42314 242197
rect 42262 242133 42314 242139
rect 42274 240759 42302 242133
rect 42934 242117 42986 242123
rect 42934 242059 42986 242065
rect 42550 242043 42602 242049
rect 42550 241985 42602 241991
rect 42358 241969 42410 241975
rect 42358 241911 42410 241917
rect 42260 240750 42316 240759
rect 42260 240685 42316 240694
rect 41782 240637 41834 240643
rect 41782 240579 41834 240585
rect 41782 240415 41834 240421
rect 41782 240357 41834 240363
rect 41794 239834 41822 240357
rect 42166 238565 42218 238571
rect 42166 238507 42218 238513
rect 42178 237984 42206 238507
rect 42166 237899 42218 237905
rect 42166 237841 42218 237847
rect 42178 237361 42206 237841
rect 42370 236721 42398 241911
rect 42562 239237 42590 241985
rect 42550 239231 42602 239237
rect 42550 239173 42602 239179
rect 42454 238935 42506 238941
rect 42454 238877 42506 238883
rect 42166 236715 42218 236721
rect 42166 236657 42218 236663
rect 42358 236715 42410 236721
rect 42358 236657 42410 236663
rect 42178 236165 42206 236657
rect 42356 236606 42412 236615
rect 42356 236541 42412 236550
rect 42166 235457 42218 235463
rect 42166 235399 42218 235405
rect 42178 234950 42206 235399
rect 42166 234865 42218 234871
rect 42166 234807 42218 234813
rect 42178 234325 42206 234807
rect 42070 234199 42122 234205
rect 42070 234141 42122 234147
rect 42082 233692 42110 234141
rect 41780 233350 41836 233359
rect 41780 233285 41836 233294
rect 41794 233129 41822 233285
rect 41986 231731 42014 231842
rect 41972 231722 42028 231731
rect 41972 231657 42028 231666
rect 41794 231139 41822 231176
rect 41780 231130 41836 231139
rect 41780 231065 41836 231074
rect 42370 230672 42398 236541
rect 42466 234205 42494 238877
rect 42946 234871 42974 242059
rect 43042 238571 43070 255041
rect 43124 248594 43180 248603
rect 43124 248529 43180 248538
rect 43030 238565 43082 238571
rect 43030 238507 43082 238513
rect 43138 235463 43166 248529
rect 43126 235457 43178 235463
rect 43126 235399 43178 235405
rect 42934 234865 42986 234871
rect 42934 234807 42986 234813
rect 42454 234199 42506 234205
rect 42454 234141 42506 234147
rect 42192 230644 42398 230672
rect 41780 230390 41836 230399
rect 41780 230325 41836 230334
rect 41794 229992 41822 230325
rect 41780 229650 41836 229659
rect 41780 229585 41836 229594
rect 41794 229357 41822 229585
rect 41780 229058 41836 229067
rect 41780 228993 41836 229002
rect 41794 228808 41822 228993
rect 41780 227430 41836 227439
rect 41780 227365 41836 227374
rect 41794 226958 41822 227365
rect 41780 226838 41836 226847
rect 41780 226773 41836 226782
rect 41794 226321 41822 226773
rect 41780 225950 41836 225959
rect 41780 225885 41836 225894
rect 41794 225700 41822 225885
rect 42742 216365 42794 216371
rect 42740 216330 42742 216339
rect 42794 216330 42796 216339
rect 42740 216265 42796 216274
rect 42742 215773 42794 215779
rect 42740 215738 42742 215747
rect 42794 215738 42796 215747
rect 42740 215673 42796 215682
rect 42742 215255 42794 215261
rect 42740 215220 42742 215229
rect 42794 215220 42796 215229
rect 42740 215155 42796 215164
rect 43234 214119 43262 257155
rect 43412 256734 43468 256743
rect 43412 256669 43468 256678
rect 43316 255846 43372 255855
rect 43316 255781 43372 255790
rect 43330 242831 43358 255781
rect 43426 246119 43454 256669
rect 44578 246267 44606 547341
rect 44566 246261 44618 246267
rect 44674 246235 44702 806489
rect 44770 627959 44798 988201
rect 44854 988185 44906 988191
rect 44854 988127 44906 988133
rect 44866 673913 44894 988127
rect 44950 988111 45002 988117
rect 44950 988053 45002 988059
rect 44962 717129 44990 988053
rect 45046 988037 45098 988043
rect 45046 987979 45098 987985
rect 45058 757681 45086 987979
rect 45142 987963 45194 987969
rect 45142 987905 45194 987911
rect 45154 800675 45182 987905
rect 47542 986705 47594 986711
rect 47542 986647 47594 986653
rect 47446 986557 47498 986563
rect 47446 986499 47498 986505
rect 46102 959103 46154 959109
rect 46102 959045 46154 959051
rect 46114 944087 46142 959045
rect 46102 944081 46154 944087
rect 46102 944023 46154 944029
rect 47458 941687 47486 986499
rect 47554 943051 47582 986647
rect 47542 943045 47594 943051
rect 47542 942987 47594 942993
rect 47444 941678 47500 941687
rect 47444 941613 47500 941622
rect 47542 872671 47594 872677
rect 47542 872613 47594 872619
rect 47446 858315 47498 858321
rect 47446 858257 47498 858263
rect 45142 800669 45194 800675
rect 45142 800611 45194 800617
rect 45046 757675 45098 757681
rect 45046 757617 45098 757623
rect 44950 717123 45002 717129
rect 44950 717065 45002 717071
rect 44854 673907 44906 673913
rect 44854 673849 44906 673855
rect 44758 627953 44810 627959
rect 44758 627895 44810 627901
rect 44758 486761 44810 486767
rect 44758 486703 44810 486709
rect 44770 388051 44798 486703
rect 44854 472405 44906 472411
rect 44854 472347 44906 472353
rect 44866 389383 44894 472347
rect 45046 414759 45098 414765
rect 45046 414701 45098 414707
rect 44854 389377 44906 389383
rect 44854 389319 44906 389325
rect 44758 388045 44810 388051
rect 44758 387987 44810 387993
rect 44950 385973 45002 385979
rect 44950 385915 45002 385921
rect 44758 376575 44810 376581
rect 44758 376517 44810 376523
rect 44770 246341 44798 376517
rect 44854 313971 44906 313977
rect 44854 313913 44906 313919
rect 44758 246335 44810 246341
rect 44758 246277 44810 246283
rect 44566 246203 44618 246209
rect 44660 246226 44716 246235
rect 44660 246161 44716 246170
rect 43414 246113 43466 246119
rect 43414 246055 43466 246061
rect 43316 242822 43372 242831
rect 43316 242757 43372 242766
rect 43220 214110 43276 214119
rect 43220 214045 43276 214054
rect 43330 213083 43358 242757
rect 43426 213675 43454 246055
rect 44866 215261 44894 313913
rect 44962 302729 44990 385915
rect 45058 345427 45086 414701
rect 47458 367405 47486 858257
rect 47554 818583 47582 872613
rect 47542 818577 47594 818583
rect 47542 818519 47594 818525
rect 47542 786313 47594 786319
rect 47542 786255 47594 786261
rect 47554 731855 47582 786255
rect 47542 731849 47594 731855
rect 47542 731791 47594 731797
rect 47542 728667 47594 728673
rect 47542 728609 47594 728615
rect 47554 688639 47582 728609
rect 47542 688633 47594 688639
rect 47542 688575 47594 688581
rect 47542 685525 47594 685531
rect 47542 685467 47594 685473
rect 47446 367399 47498 367405
rect 47446 367341 47498 367347
rect 47446 357187 47498 357193
rect 47446 357129 47498 357135
rect 45046 345421 45098 345427
rect 45046 345363 45098 345369
rect 45046 332249 45098 332255
rect 45046 332191 45098 332197
rect 44950 302723 45002 302729
rect 44950 302665 45002 302671
rect 44950 299615 45002 299621
rect 44950 299557 45002 299563
rect 44962 216371 44990 299557
rect 45058 249153 45086 332191
rect 45142 285185 45194 285191
rect 45142 285127 45194 285133
rect 45046 249147 45098 249153
rect 45046 249089 45098 249095
rect 44950 216365 45002 216371
rect 44950 216307 45002 216313
rect 45154 215779 45182 285127
rect 47458 258255 47486 357129
rect 47446 258249 47498 258255
rect 47446 258191 47498 258197
rect 47554 237905 47582 685467
rect 47650 584743 47678 988275
rect 47734 986631 47786 986637
rect 47734 986573 47786 986579
rect 47746 942903 47774 986573
rect 59444 975422 59500 975431
rect 59444 975357 59500 975366
rect 59458 973539 59486 975357
rect 50518 973533 50570 973539
rect 50518 973475 50570 973481
rect 59446 973533 59498 973539
rect 59446 973475 59498 973481
rect 47734 942897 47786 942903
rect 47734 942839 47786 942845
rect 50326 901531 50378 901537
rect 50326 901473 50378 901479
rect 47734 829529 47786 829535
rect 47734 829471 47786 829477
rect 47746 775959 47774 829471
rect 50338 818287 50366 901473
rect 50326 818281 50378 818287
rect 50326 818223 50378 818229
rect 50422 815099 50474 815105
rect 50422 815041 50474 815047
rect 50326 800669 50378 800675
rect 50326 800611 50378 800617
rect 47734 775953 47786 775959
rect 47734 775895 47786 775901
rect 47638 584737 47690 584743
rect 47638 584679 47690 584685
rect 48886 559355 48938 559361
rect 48886 559297 48938 559303
rect 48898 544709 48926 559297
rect 48886 544703 48938 544709
rect 48886 544645 48938 544651
rect 47734 501191 47786 501197
rect 47734 501133 47786 501139
rect 47746 432007 47774 501133
rect 47734 432001 47786 432007
rect 47734 431943 47786 431949
rect 47638 429189 47690 429195
rect 47638 429131 47690 429137
rect 47650 345945 47678 429131
rect 47734 371617 47786 371623
rect 47734 371559 47786 371565
rect 47638 345939 47690 345945
rect 47638 345881 47690 345887
rect 47746 302359 47774 371559
rect 50338 324189 50366 800611
rect 50434 775367 50462 815041
rect 50422 775361 50474 775367
rect 50422 775303 50474 775309
rect 50422 714311 50474 714317
rect 50422 714253 50474 714259
rect 50434 689527 50462 714253
rect 50422 689521 50474 689527
rect 50422 689463 50474 689469
rect 50422 671095 50474 671101
rect 50422 671037 50474 671043
rect 50434 645275 50462 671037
rect 50422 645269 50474 645275
rect 50422 645211 50474 645217
rect 50422 627879 50474 627885
rect 50422 627821 50474 627827
rect 50326 324183 50378 324189
rect 50326 324125 50378 324131
rect 47734 302353 47786 302359
rect 47734 302295 47786 302301
rect 47638 290143 47690 290149
rect 47638 290085 47690 290091
rect 47650 246711 47678 290085
rect 47638 246705 47690 246711
rect 47638 246647 47690 246653
rect 50326 241969 50378 241975
rect 50326 241911 50378 241917
rect 47542 237899 47594 237905
rect 47542 237841 47594 237847
rect 45142 215773 45194 215779
rect 45142 215715 45194 215721
rect 44854 215255 44906 215261
rect 44854 215197 44906 215203
rect 43412 213666 43468 213675
rect 43412 213601 43468 213610
rect 43316 213074 43372 213083
rect 43316 213009 43372 213018
rect 41972 211594 42028 211603
rect 41972 211529 42028 211538
rect 40244 209522 40300 209531
rect 40244 209457 40300 209466
rect 40258 206825 40286 209457
rect 40246 206819 40298 206825
rect 40246 206761 40298 206767
rect 41782 206819 41834 206825
rect 41782 206761 41834 206767
rect 40148 206710 40204 206719
rect 40148 206645 40204 206654
rect 40052 206118 40108 206127
rect 40052 206053 40108 206062
rect 35156 204046 35212 204055
rect 35156 203981 35212 203990
rect 35170 203611 35198 203981
rect 35156 203602 35212 203611
rect 35156 203537 35212 203546
rect 40066 198907 40094 206053
rect 40162 199055 40190 206645
rect 40244 205674 40300 205683
rect 40244 205609 40300 205618
rect 40150 199049 40202 199055
rect 40150 198991 40202 198997
rect 40054 198901 40106 198907
rect 40054 198843 40106 198849
rect 40258 198759 40286 205609
rect 40246 198753 40298 198759
rect 40246 198695 40298 198701
rect 41794 197427 41822 206761
rect 41986 201127 42014 211529
rect 42356 209966 42412 209975
rect 42356 209901 42412 209910
rect 42370 201243 42398 209901
rect 42740 207746 42796 207755
rect 42740 207681 42796 207690
rect 42754 205068 42782 207681
rect 42932 207302 42988 207311
rect 42932 207237 42988 207246
rect 42754 205040 42878 205068
rect 42740 204860 42796 204869
rect 42740 204795 42796 204804
rect 42754 204457 42782 204795
rect 42742 204451 42794 204457
rect 42742 204393 42794 204399
rect 42754 203759 42782 204393
rect 42740 203750 42796 203759
rect 42740 203685 42796 203694
rect 42356 201234 42412 201243
rect 42356 201169 42412 201178
rect 41974 201121 42026 201127
rect 41974 201063 42026 201069
rect 42358 201121 42410 201127
rect 42358 201063 42410 201069
rect 42166 199049 42218 199055
rect 42166 198991 42218 198997
rect 42178 197543 42206 198991
rect 42164 197534 42220 197543
rect 42164 197469 42220 197478
rect 41782 197421 41834 197427
rect 41782 197363 41834 197369
rect 41782 197199 41834 197205
rect 41782 197141 41834 197147
rect 41794 196618 41822 197141
rect 42370 195355 42398 201063
rect 42166 195349 42218 195355
rect 42166 195291 42218 195297
rect 42358 195349 42410 195355
rect 42358 195291 42410 195297
rect 42178 194805 42206 195291
rect 42356 195166 42412 195175
rect 42356 195101 42412 195110
rect 42070 194535 42122 194541
rect 42070 194477 42122 194483
rect 42082 194176 42110 194477
rect 42070 193499 42122 193505
rect 42070 193441 42122 193447
rect 42082 192992 42110 193441
rect 42166 192241 42218 192247
rect 42166 192183 42218 192189
rect 42178 191769 42206 192183
rect 42370 191507 42398 195101
rect 42070 191501 42122 191507
rect 42070 191443 42122 191449
rect 42358 191501 42410 191507
rect 42358 191443 42410 191449
rect 42082 191142 42110 191443
rect 42166 191057 42218 191063
rect 42166 190999 42218 191005
rect 42178 190476 42206 190999
rect 42068 190282 42124 190291
rect 42068 190217 42124 190226
rect 42082 189929 42110 190217
rect 41972 189098 42028 189107
rect 41972 189033 42028 189042
rect 41986 188626 42014 189033
rect 41780 188358 41836 188367
rect 41780 188293 41836 188302
rect 41794 188011 41822 188293
rect 41794 187997 42398 188011
rect 41808 187983 42398 187997
rect 42262 187949 42314 187955
rect 42262 187891 42314 187897
rect 42274 187456 42302 187891
rect 42192 187428 42302 187456
rect 42166 187135 42218 187141
rect 42166 187077 42218 187083
rect 42178 186776 42206 187077
rect 41780 186730 41836 186739
rect 41780 186665 41836 186674
rect 41794 186184 41822 186665
rect 41780 185842 41836 185851
rect 41780 185777 41836 185786
rect 41794 185592 41822 185777
rect 42370 184792 42398 187983
rect 42850 187141 42878 205040
rect 42946 193505 42974 207237
rect 43028 205378 43084 205387
rect 43028 205313 43084 205322
rect 42934 193499 42986 193505
rect 42934 193441 42986 193447
rect 42934 193351 42986 193357
rect 42934 193293 42986 193299
rect 42946 187955 42974 193293
rect 43042 192247 43070 205313
rect 50338 204457 50366 241911
rect 50326 204451 50378 204457
rect 50326 204393 50378 204399
rect 43126 198901 43178 198907
rect 43178 198849 43262 198852
rect 43126 198843 43262 198849
rect 43138 198824 43262 198843
rect 43126 198753 43178 198759
rect 43126 198695 43178 198701
rect 43030 192241 43082 192247
rect 43030 192183 43082 192189
rect 43138 191063 43166 198695
rect 43234 193357 43262 198824
rect 50434 194541 50462 627821
rect 50530 541527 50558 973475
rect 61858 962111 61886 993529
rect 62036 992146 62092 992155
rect 62036 992081 62092 992090
rect 62050 962407 62078 992081
rect 69154 987988 69182 995083
rect 77314 993667 77342 995508
rect 77698 993815 77726 995522
rect 77686 993809 77738 993815
rect 78370 993783 78398 995522
rect 77686 993751 77738 993757
rect 78356 993774 78412 993783
rect 80194 993741 80222 995522
rect 82032 995517 82334 995536
rect 82032 995511 82346 995517
rect 82032 995508 82294 995511
rect 82294 995453 82346 995459
rect 78356 993709 78412 993718
rect 80182 993735 80234 993741
rect 80182 993677 80234 993683
rect 77302 993661 77354 993667
rect 77302 993603 77354 993609
rect 82594 993593 82622 995522
rect 83232 995508 83486 995536
rect 84528 995508 84830 995536
rect 85104 995508 85364 995536
rect 83458 993635 83486 995508
rect 84802 995411 84830 995508
rect 85364 995485 85420 995494
rect 84788 995402 84844 995411
rect 86338 995369 86366 995522
rect 87552 995508 87806 995536
rect 84788 995337 84844 995346
rect 86326 995363 86378 995369
rect 86326 995305 86378 995311
rect 87778 995263 87806 995508
rect 87764 995254 87820 995263
rect 87764 995189 87820 995198
rect 88738 993931 88766 995522
rect 89410 994967 89438 995522
rect 89396 994958 89452 994967
rect 89396 994893 89452 994902
rect 88724 993922 88780 993931
rect 88724 993857 88780 993866
rect 92674 993635 92702 999375
rect 104660 996586 104716 996595
rect 97942 996547 97994 996553
rect 104660 996521 104662 996530
rect 97942 996489 97994 996495
rect 104714 996521 104716 996530
rect 104662 996489 104714 996495
rect 94966 995955 95018 995961
rect 94966 995897 95018 995903
rect 94978 995855 95006 995897
rect 94964 995846 95020 995855
rect 94964 995781 95020 995790
rect 94966 995733 95018 995739
rect 94964 995698 94966 995707
rect 95018 995698 95020 995707
rect 94964 995633 95020 995642
rect 95062 995659 95114 995665
rect 95062 995601 95114 995607
rect 93526 995585 93578 995591
rect 93526 995527 93578 995533
rect 83444 993626 83500 993635
rect 82582 993587 82634 993593
rect 83444 993561 83500 993570
rect 92660 993626 92716 993635
rect 92660 993561 92716 993570
rect 82582 993529 82634 993535
rect 83458 992155 83486 993561
rect 83444 992146 83500 992155
rect 73366 992107 73418 992113
rect 83444 992081 83500 992090
rect 73366 992049 73418 992055
rect 69058 987960 69182 987988
rect 65110 986779 65162 986785
rect 65110 986721 65162 986727
rect 63286 986483 63338 986489
rect 63286 986425 63338 986431
rect 62036 962398 62092 962407
rect 62036 962333 62092 962342
rect 61844 962102 61900 962111
rect 61844 962037 61900 962046
rect 59540 960918 59596 960927
rect 59540 960853 59596 960862
rect 59554 959109 59582 960853
rect 59542 959103 59594 959109
rect 59542 959045 59594 959051
rect 59540 946710 59596 946719
rect 59540 946645 59596 946654
rect 59554 944679 59582 946645
rect 59542 944673 59594 944679
rect 59542 944615 59594 944621
rect 51862 944229 51914 944235
rect 51862 944171 51914 944177
rect 51874 930545 51902 944171
rect 59540 932206 59596 932215
rect 53206 932167 53258 932173
rect 59540 932141 59596 932150
rect 53206 932109 53258 932115
rect 51862 930539 51914 930545
rect 51862 930481 51914 930487
rect 51862 602275 51914 602281
rect 51862 602217 51914 602223
rect 51874 586001 51902 602217
rect 51862 585995 51914 586001
rect 51862 585937 51914 585943
rect 50518 541521 50570 541527
rect 50518 541463 50570 541469
rect 50518 457975 50570 457981
rect 50518 457917 50570 457923
rect 50530 388791 50558 457917
rect 50518 388785 50570 388791
rect 50518 388727 50570 388733
rect 50518 342831 50570 342837
rect 50518 342773 50570 342779
rect 50530 259735 50558 342773
rect 50518 259729 50570 259735
rect 50518 259671 50570 259677
rect 53218 246489 53246 932109
rect 59554 930545 59582 932141
rect 59542 930539 59594 930545
rect 59542 930481 59594 930487
rect 59540 917850 59596 917859
rect 59540 917785 59596 917794
rect 59554 915893 59582 917785
rect 53398 915887 53450 915893
rect 53398 915829 53450 915835
rect 59542 915887 59594 915893
rect 59542 915829 59594 915835
rect 53302 843885 53354 843891
rect 53302 843827 53354 843833
rect 53314 774849 53342 843827
rect 53302 774843 53354 774849
rect 53302 774785 53354 774791
rect 53300 763338 53356 763347
rect 53300 763273 53356 763282
rect 53206 246483 53258 246489
rect 53206 246425 53258 246431
rect 53314 246383 53342 763273
rect 53410 406107 53438 915829
rect 59540 903494 59596 903503
rect 59540 903429 59596 903438
rect 59554 901537 59582 903429
rect 59542 901531 59594 901537
rect 59542 901473 59594 901479
rect 59540 889138 59596 889147
rect 59540 889073 59596 889082
rect 59554 887181 59582 889073
rect 53494 887175 53546 887181
rect 53494 887117 53546 887123
rect 59542 887175 59594 887181
rect 59542 887117 59594 887123
rect 53506 819323 53534 887117
rect 59540 874782 59596 874791
rect 59540 874717 59596 874726
rect 59554 872677 59582 874717
rect 59542 872671 59594 872677
rect 59542 872613 59594 872619
rect 58580 860426 58636 860435
rect 58580 860361 58636 860370
rect 58594 858321 58622 860361
rect 58582 858315 58634 858321
rect 58582 858257 58634 858263
rect 59540 846070 59596 846079
rect 59540 846005 59596 846014
rect 59554 843891 59582 846005
rect 59542 843885 59594 843891
rect 59542 843827 59594 843833
rect 59540 831714 59596 831723
rect 59540 831649 59596 831658
rect 59554 829535 59582 831649
rect 59542 829529 59594 829535
rect 59542 829471 59594 829477
rect 53494 819317 53546 819323
rect 53494 819259 53546 819265
rect 59540 817358 59596 817367
rect 59540 817293 59596 817302
rect 59554 815105 59582 817293
rect 59542 815099 59594 815105
rect 59542 815041 59594 815047
rect 59540 802854 59596 802863
rect 59540 802789 59596 802798
rect 59554 800675 59582 802789
rect 59542 800669 59594 800675
rect 59542 800611 59594 800617
rect 59540 788646 59596 788655
rect 59540 788581 59596 788590
rect 59554 786319 59582 788581
rect 59542 786313 59594 786319
rect 59542 786255 59594 786261
rect 59540 774142 59596 774151
rect 59540 774077 59596 774086
rect 59554 771889 59582 774077
rect 53494 771883 53546 771889
rect 53494 771825 53546 771831
rect 59542 771883 59594 771889
rect 59542 771825 59594 771831
rect 53506 732743 53534 771825
rect 59540 759786 59596 759795
rect 59540 759721 59596 759730
rect 59554 757533 59582 759721
rect 53686 757527 53738 757533
rect 53686 757469 53738 757475
rect 59542 757527 59594 757533
rect 59542 757469 59594 757475
rect 53590 743097 53642 743103
rect 53590 743039 53642 743045
rect 53494 732737 53546 732743
rect 53494 732679 53546 732685
rect 53492 720122 53548 720131
rect 53492 720057 53548 720066
rect 53398 406101 53450 406107
rect 53398 406043 53450 406049
rect 53398 328401 53450 328407
rect 53398 328343 53450 328349
rect 53410 258995 53438 328343
rect 53398 258989 53450 258995
rect 53398 258931 53450 258937
rect 53506 246563 53534 720057
rect 53602 281121 53630 743039
rect 53698 732151 53726 757469
rect 59540 745578 59596 745587
rect 59540 745513 59596 745522
rect 59554 743103 59582 745513
rect 59542 743097 59594 743103
rect 59542 743039 59594 743045
rect 53686 732145 53738 732151
rect 53686 732087 53738 732093
rect 59540 731074 59596 731083
rect 59540 731009 59596 731018
rect 59554 728673 59582 731009
rect 59542 728667 59594 728673
rect 59542 728609 59594 728615
rect 59540 716718 59596 716727
rect 59540 716653 59596 716662
rect 59554 714317 59582 716653
rect 59542 714311 59594 714317
rect 59542 714253 59594 714259
rect 59540 702362 59596 702371
rect 59540 702297 59596 702306
rect 59554 699887 59582 702297
rect 59542 699881 59594 699887
rect 59542 699823 59594 699829
rect 59540 688006 59596 688015
rect 59540 687941 59596 687950
rect 59554 685531 59582 687941
rect 59542 685525 59594 685531
rect 59542 685467 59594 685473
rect 53684 676906 53740 676915
rect 53684 676841 53740 676850
rect 53590 281115 53642 281121
rect 53590 281057 53642 281063
rect 53494 246557 53546 246563
rect 53698 246531 53726 676841
rect 59540 673650 59596 673659
rect 59540 673585 59596 673594
rect 59554 671101 59582 673585
rect 59542 671095 59594 671101
rect 59542 671037 59594 671043
rect 59540 659294 59596 659303
rect 59540 659229 59596 659238
rect 59554 656745 59582 659229
rect 59542 656739 59594 656745
rect 59542 656681 59594 656687
rect 59542 645121 59594 645127
rect 59542 645063 59594 645069
rect 59554 644947 59582 645063
rect 59540 644938 59596 644947
rect 59540 644873 59596 644882
rect 56084 633986 56140 633995
rect 56084 633921 56140 633930
rect 53780 590622 53836 590631
rect 53780 590557 53836 590566
rect 53794 249227 53822 590557
rect 53974 515547 54026 515553
rect 53974 515489 54026 515495
rect 53878 443619 53930 443625
rect 53878 443561 53930 443567
rect 53890 344835 53918 443561
rect 53986 432303 54014 515489
rect 53974 432297 54026 432303
rect 53974 432239 54026 432245
rect 53878 344829 53930 344835
rect 53878 344771 53930 344777
rect 53782 249221 53834 249227
rect 53782 249163 53834 249169
rect 56098 246637 56126 633921
rect 59540 630582 59596 630591
rect 59540 630517 59596 630526
rect 59554 627885 59582 630517
rect 59542 627879 59594 627885
rect 59542 627821 59594 627827
rect 59540 616226 59596 616235
rect 59540 616161 59596 616170
rect 59554 613529 59582 616161
rect 59542 613523 59594 613529
rect 59542 613465 59594 613471
rect 59542 601905 59594 601911
rect 59540 601870 59542 601879
rect 59594 601870 59596 601879
rect 59540 601805 59596 601814
rect 59540 587514 59596 587523
rect 59540 587449 59596 587458
rect 59554 586001 59582 587449
rect 59542 585995 59594 586001
rect 59542 585937 59594 585943
rect 59540 573010 59596 573019
rect 59540 572945 59596 572954
rect 59554 570313 59582 572945
rect 59542 570307 59594 570313
rect 59542 570249 59594 570255
rect 59540 558950 59596 558959
rect 59540 558885 59542 558894
rect 59594 558885 59596 558894
rect 59542 558853 59594 558859
rect 59542 544703 59594 544709
rect 59542 544645 59594 544651
rect 59554 544455 59582 544645
rect 59540 544446 59596 544455
rect 59540 544381 59596 544390
rect 59540 530090 59596 530099
rect 59540 530025 59596 530034
rect 59554 529983 59582 530025
rect 59542 529977 59594 529983
rect 59542 529919 59594 529925
rect 59540 515734 59596 515743
rect 59540 515669 59596 515678
rect 59554 515553 59582 515669
rect 59542 515547 59594 515553
rect 59542 515489 59594 515495
rect 59540 501230 59596 501239
rect 59540 501165 59542 501174
rect 59594 501165 59596 501174
rect 59542 501133 59594 501139
rect 58580 486874 58636 486883
rect 58580 486809 58636 486818
rect 58594 486767 58622 486809
rect 58582 486761 58634 486767
rect 58582 486703 58634 486709
rect 59540 472518 59596 472527
rect 59540 472453 59596 472462
rect 59554 472411 59582 472453
rect 59542 472405 59594 472411
rect 59542 472347 59594 472353
rect 59540 458162 59596 458171
rect 59540 458097 59596 458106
rect 59554 457981 59582 458097
rect 59542 457975 59594 457981
rect 59542 457917 59594 457923
rect 59540 443806 59596 443815
rect 59540 443741 59596 443750
rect 59554 443625 59582 443741
rect 59542 443619 59594 443625
rect 59542 443561 59594 443567
rect 59540 429450 59596 429459
rect 59540 429385 59596 429394
rect 59554 429195 59582 429385
rect 59542 429189 59594 429195
rect 59542 429131 59594 429137
rect 56182 417645 56234 417651
rect 56182 417587 56234 417593
rect 56194 249301 56222 417587
rect 58388 415094 58444 415103
rect 58388 415029 58444 415038
rect 58402 414765 58430 415029
rect 58390 414759 58442 414765
rect 58390 414701 58442 414707
rect 57620 400738 57676 400747
rect 57620 400673 57676 400682
rect 57634 400409 57662 400673
rect 56278 400403 56330 400409
rect 56278 400345 56330 400351
rect 57622 400403 57674 400409
rect 57622 400345 57674 400351
rect 56290 301693 56318 400345
rect 59252 386382 59308 386391
rect 59252 386317 59308 386326
rect 59266 385979 59294 386317
rect 59254 385973 59306 385979
rect 59254 385915 59306 385921
rect 59540 371878 59596 371887
rect 59540 371813 59596 371822
rect 59554 371623 59582 371813
rect 59542 371617 59594 371623
rect 59542 371559 59594 371565
rect 59540 357670 59596 357679
rect 59540 357605 59596 357614
rect 59554 357193 59582 357605
rect 59542 357187 59594 357193
rect 59542 357129 59594 357135
rect 58388 343166 58444 343175
rect 58388 343101 58444 343110
rect 58402 342837 58430 343101
rect 58390 342831 58442 342837
rect 58390 342773 58442 342779
rect 57812 328810 57868 328819
rect 57812 328745 57868 328754
rect 57826 328407 57854 328745
rect 57814 328401 57866 328407
rect 57814 328343 57866 328349
rect 58004 314602 58060 314611
rect 58004 314537 58060 314546
rect 58018 313977 58046 314537
rect 58006 313971 58058 313977
rect 58006 313913 58058 313919
rect 56278 301687 56330 301693
rect 56278 301629 56330 301635
rect 59444 300098 59500 300107
rect 59444 300033 59500 300042
rect 59458 299621 59486 300033
rect 59446 299615 59498 299621
rect 59446 299557 59498 299563
rect 58100 285890 58156 285899
rect 58100 285825 58156 285834
rect 58114 285191 58142 285825
rect 58102 285185 58154 285191
rect 58102 285127 58154 285133
rect 56182 249295 56234 249301
rect 56182 249237 56234 249243
rect 63298 246785 63326 986425
rect 64918 986187 64970 986193
rect 64918 986129 64970 986135
rect 64822 983597 64874 983603
rect 64822 983539 64874 983545
rect 64834 278605 64862 983539
rect 64822 278599 64874 278605
rect 64822 278541 64874 278547
rect 64930 277939 64958 986129
rect 65014 983523 65066 983529
rect 65014 983465 65066 983471
rect 64918 277933 64970 277939
rect 64918 277875 64970 277881
rect 65026 267875 65054 983465
rect 65014 267869 65066 267875
rect 65014 267811 65066 267817
rect 63286 246779 63338 246785
rect 63286 246721 63338 246727
rect 65014 246705 65066 246711
rect 65014 246647 65066 246653
rect 56086 246631 56138 246637
rect 56086 246573 56138 246579
rect 53494 246499 53546 246505
rect 53684 246522 53740 246531
rect 53684 246457 53740 246466
rect 53300 246374 53356 246383
rect 53300 246309 53356 246318
rect 65026 246193 65054 246647
rect 65014 246187 65066 246193
rect 65014 246129 65066 246135
rect 65122 246087 65150 986721
rect 65206 986409 65258 986415
rect 65206 986351 65258 986357
rect 65218 246711 65246 986351
rect 69058 986193 69086 987960
rect 69046 986187 69098 986193
rect 69046 986129 69098 986135
rect 73378 983548 73406 992049
rect 89590 989295 89642 989301
rect 89590 989237 89642 989243
rect 73378 983520 73488 983548
rect 89602 983534 89630 989237
rect 93538 986785 93566 995527
rect 95074 993815 95102 995601
rect 97954 995115 97982 996489
rect 107542 996325 107594 996331
rect 107542 996267 107594 996273
rect 99764 995994 99820 996003
rect 99764 995929 99820 995938
rect 102836 995994 102892 996003
rect 102836 995929 102838 995938
rect 98036 995846 98092 995855
rect 98036 995781 98092 995790
rect 98050 995591 98078 995781
rect 98038 995585 98090 995591
rect 98038 995527 98090 995533
rect 99778 995369 99806 995929
rect 102890 995929 102892 995938
rect 102838 995897 102890 995903
rect 101206 995881 101258 995887
rect 100724 995846 100780 995855
rect 100724 995781 100780 995790
rect 101204 995846 101206 995855
rect 101258 995846 101260 995855
rect 101204 995781 101260 995790
rect 102452 995846 102508 995855
rect 102452 995781 102508 995790
rect 103988 995846 104044 995855
rect 103988 995781 103990 995790
rect 100738 995517 100766 995781
rect 102466 995739 102494 995781
rect 104042 995781 104044 995790
rect 103990 995749 104042 995755
rect 102454 995733 102506 995739
rect 102356 995698 102412 995707
rect 107554 995707 107582 996267
rect 107926 996103 107978 996109
rect 107926 996045 107978 996051
rect 107938 995855 107966 996045
rect 108982 996029 109034 996035
rect 108980 995994 108982 996003
rect 109034 995994 109036 996003
rect 108980 995929 109036 995938
rect 109556 995994 109612 996003
rect 109556 995929 109612 995938
rect 107924 995846 107980 995855
rect 107924 995781 107980 995790
rect 102454 995675 102506 995681
rect 105332 995698 105388 995707
rect 102356 995633 102358 995642
rect 102410 995633 102412 995642
rect 105332 995633 105388 995642
rect 105908 995698 105964 995707
rect 105908 995633 105964 995642
rect 107540 995698 107596 995707
rect 107540 995633 107596 995642
rect 102358 995601 102410 995607
rect 100726 995511 100778 995517
rect 100726 995453 100778 995459
rect 99766 995363 99818 995369
rect 99766 995305 99818 995311
rect 97940 995106 97996 995115
rect 97940 995041 97996 995050
rect 95062 993809 95114 993815
rect 95062 993751 95114 993757
rect 105346 993741 105374 995633
rect 105334 993735 105386 993741
rect 105334 993677 105386 993683
rect 105922 993667 105950 995633
rect 106772 995254 106828 995263
rect 106772 995189 106828 995198
rect 106786 993783 106814 995189
rect 106772 993774 106828 993783
rect 106772 993709 106828 993718
rect 105910 993661 105962 993667
rect 105910 993603 105962 993609
rect 105814 990553 105866 990559
rect 105814 990495 105866 990501
rect 93526 986779 93578 986785
rect 93526 986721 93578 986727
rect 105826 983534 105854 990495
rect 107554 986563 107582 995633
rect 107938 986637 107966 995781
rect 109172 995698 109228 995707
rect 109172 995633 109228 995642
rect 109186 986711 109214 995633
rect 109364 995550 109420 995559
rect 109364 995485 109420 995494
rect 109378 989301 109406 995485
rect 109570 990559 109598 995929
rect 110132 995698 110188 995707
rect 110132 995633 110188 995642
rect 110146 992113 110174 995633
rect 126658 993635 126686 999375
rect 126742 996325 126794 996331
rect 126742 996267 126794 996273
rect 126754 995591 126782 996267
rect 136464 995813 136862 995832
rect 138960 995813 139358 995832
rect 142656 995813 143006 995832
rect 136464 995807 136874 995813
rect 136464 995804 136822 995807
rect 138960 995807 139370 995813
rect 138960 995804 139318 995807
rect 136822 995749 136874 995755
rect 142656 995807 143018 995813
rect 142656 995804 142966 995807
rect 139318 995749 139370 995755
rect 142966 995749 143018 995755
rect 137974 995733 138026 995739
rect 137136 995665 137438 995684
rect 137760 995681 137974 995684
rect 137760 995675 138026 995681
rect 137136 995659 137450 995665
rect 137136 995656 137398 995659
rect 137760 995656 138014 995675
rect 143650 995665 143678 999504
rect 143734 999433 143786 999439
rect 143734 999375 143786 999381
rect 143746 995813 143774 999375
rect 143734 995807 143786 995813
rect 143734 995749 143786 995755
rect 143842 995739 143870 1002335
rect 143938 995887 143966 1002557
rect 144022 1002467 144074 1002473
rect 144022 1002409 144074 1002415
rect 144034 995961 144062 1002409
rect 144118 1002319 144170 1002325
rect 144118 1002261 144170 1002267
rect 144022 995955 144074 995961
rect 144022 995897 144074 995903
rect 143926 995881 143978 995887
rect 143926 995823 143978 995829
rect 143830 995733 143882 995739
rect 143830 995675 143882 995681
rect 143638 995659 143690 995665
rect 137398 995601 137450 995607
rect 143638 995601 143690 995607
rect 144130 995591 144158 1002261
rect 144214 996325 144266 996331
rect 144214 996267 144266 996273
rect 144226 995665 144254 996267
rect 144214 995659 144266 995665
rect 144214 995601 144266 995607
rect 126742 995585 126794 995591
rect 143830 995585 143882 995591
rect 133652 995550 133708 995559
rect 126742 995527 126794 995533
rect 128482 993667 128510 995522
rect 129120 995508 129374 995536
rect 129346 993815 129374 995508
rect 129730 994079 129758 995522
rect 131616 995508 131870 995536
rect 129716 994070 129772 994079
rect 129716 994005 129772 994014
rect 129334 993809 129386 993815
rect 129334 993751 129386 993757
rect 131842 993741 131870 995508
rect 132130 995295 132158 995522
rect 132118 995289 132170 995295
rect 132118 995231 132170 995237
rect 132802 994523 132830 995522
rect 133440 995508 133652 995536
rect 133652 995485 133708 995494
rect 133954 995508 134016 995536
rect 134338 995508 134640 995536
rect 135936 995508 136190 995536
rect 140160 995508 140414 995536
rect 143830 995527 143882 995533
rect 144118 995585 144170 995591
rect 144118 995527 144170 995533
rect 132788 994514 132844 994523
rect 132788 994449 132844 994458
rect 131830 993735 131882 993741
rect 131830 993677 131882 993683
rect 128470 993661 128522 993667
rect 126644 993626 126700 993635
rect 128470 993603 128522 993609
rect 133954 993593 133982 995508
rect 134338 993783 134366 995508
rect 136162 994227 136190 995508
rect 136148 994218 136204 994227
rect 136148 994153 136204 994162
rect 140386 993783 140414 995508
rect 140770 994375 140798 995522
rect 140756 994366 140812 994375
rect 140756 994301 140812 994310
rect 134324 993774 134380 993783
rect 134324 993709 134380 993718
rect 140372 993774 140428 993783
rect 140372 993709 140428 993718
rect 143842 993593 143870 995527
rect 126644 993561 126700 993570
rect 133942 993587 133994 993593
rect 133942 993529 133994 993535
rect 143830 993587 143882 993593
rect 143830 993529 143882 993535
rect 110134 992107 110186 992113
rect 110134 992049 110186 992055
rect 109558 990553 109610 990559
rect 109558 990495 109610 990501
rect 109366 989295 109418 989301
rect 109366 989237 109418 989243
rect 138262 989295 138314 989301
rect 138262 989237 138314 989243
rect 122038 988333 122090 988339
rect 122038 988275 122090 988281
rect 109174 986705 109226 986711
rect 109174 986647 109226 986653
rect 107926 986631 107978 986637
rect 107926 986573 107978 986579
rect 107542 986557 107594 986563
rect 107542 986499 107594 986505
rect 122050 983534 122078 988275
rect 138274 983534 138302 989237
rect 145378 986489 145406 1007917
rect 164278 1005279 164330 1005285
rect 164278 1005221 164330 1005227
rect 172822 1005279 172874 1005285
rect 172822 1005221 172874 1005227
rect 160436 1003246 160492 1003255
rect 160436 1003181 160438 1003190
rect 160490 1003181 160492 1003190
rect 161492 1003209 161548 1003218
rect 164290 1003213 164318 1005221
rect 160438 1003149 160490 1003155
rect 161492 1003144 161548 1003153
rect 164278 1003207 164330 1003213
rect 164278 1003149 164330 1003155
rect 161506 1002991 161534 1003144
rect 161494 1002985 161546 1002991
rect 161494 1002927 161546 1002933
rect 169942 1002985 169994 1002991
rect 169942 1002927 169994 1002933
rect 153332 1002654 153388 1002663
rect 153332 1002589 153334 1002598
rect 153386 1002589 153388 1002598
rect 153334 1002557 153386 1002563
rect 152662 1002541 152714 1002547
rect 151604 1002506 151660 1002515
rect 151604 1002441 151606 1002450
rect 151658 1002441 151660 1002450
rect 152660 1002506 152662 1002515
rect 152714 1002506 152716 1002515
rect 152660 1002441 152716 1002450
rect 151606 1002409 151658 1002415
rect 151030 1002393 151082 1002399
rect 151028 1002358 151030 1002367
rect 151082 1002358 151084 1002367
rect 151028 1002293 151084 1002302
rect 155542 999433 155594 999439
rect 155540 999398 155542 999407
rect 155594 999398 155596 999407
rect 155540 999333 155596 999342
rect 159188 996290 159244 996299
rect 159188 996225 159190 996234
rect 159242 996225 159244 996234
rect 159190 996193 159242 996199
rect 159764 996142 159820 996151
rect 159764 996077 159766 996086
rect 159818 996077 159820 996086
rect 159766 996045 159818 996051
rect 160438 996029 160490 996035
rect 156596 995994 156652 996003
rect 156596 995929 156652 995938
rect 160436 995994 160438 996003
rect 160490 995994 160492 996003
rect 160436 995929 160492 995938
rect 154868 995846 154924 995855
rect 149590 995807 149642 995813
rect 154868 995781 154870 995790
rect 149590 995749 149642 995755
rect 154922 995781 154924 995790
rect 154870 995749 154922 995755
rect 146806 995289 146858 995295
rect 146804 995254 146806 995263
rect 146858 995254 146860 995263
rect 146804 995189 146860 995198
rect 149602 993815 149630 995749
rect 149684 995402 149740 995411
rect 149684 995337 149740 995346
rect 149698 994523 149726 995337
rect 156404 995254 156460 995263
rect 156130 995212 156404 995240
rect 149684 994514 149740 994523
rect 149684 994449 149740 994458
rect 156130 994375 156158 995212
rect 156404 995189 156460 995198
rect 156116 994366 156172 994375
rect 156116 994301 156172 994310
rect 149590 993809 149642 993815
rect 149590 993751 149642 993757
rect 156610 993741 156638 995929
rect 161492 995846 161548 995855
rect 161492 995781 161548 995790
rect 157268 995402 157324 995411
rect 157268 995337 157324 995346
rect 156598 993735 156650 993741
rect 156598 993677 156650 993683
rect 157282 993667 157310 995337
rect 157270 993661 157322 993667
rect 157270 993603 157322 993609
rect 154486 989369 154538 989375
rect 154486 989311 154538 989317
rect 145366 986483 145418 986489
rect 145366 986425 145418 986431
rect 154498 983534 154526 989311
rect 161506 989301 161534 995781
rect 161684 995254 161740 995263
rect 161684 995189 161740 995198
rect 161698 989375 161726 995189
rect 161686 989369 161738 989375
rect 161686 989311 161738 989317
rect 161494 989295 161546 989301
rect 161494 989237 161546 989243
rect 169954 983548 169982 1002927
rect 172834 995961 172862 1005221
rect 218806 1005205 218858 1005211
rect 213812 1005170 213868 1005179
rect 213812 1005105 213868 1005114
rect 218804 1005170 218806 1005179
rect 222646 1005205 222698 1005211
rect 218858 1005170 218860 1005179
rect 222646 1005147 222698 1005153
rect 218804 1005105 218860 1005114
rect 195286 1003281 195338 1003287
rect 195286 1003223 195338 1003229
rect 209108 1003246 209164 1003255
rect 175702 1002319 175754 1002325
rect 175702 1002261 175754 1002267
rect 172822 995955 172874 995961
rect 172822 995897 172874 995903
rect 175714 995813 175742 1002261
rect 195190 999507 195242 999513
rect 195190 999449 195242 999455
rect 195094 999433 195146 999439
rect 195094 999375 195146 999381
rect 183764 995846 183820 995855
rect 175702 995807 175754 995813
rect 183552 995804 183764 995832
rect 192500 995846 192556 995855
rect 185218 995818 185424 995832
rect 185218 995813 185438 995818
rect 183764 995781 183820 995790
rect 185206 995807 185438 995813
rect 175702 995749 175754 995755
rect 185258 995804 185438 995807
rect 188544 995813 188894 995832
rect 190368 995813 190622 995832
rect 188544 995807 188906 995813
rect 188544 995804 188854 995807
rect 185206 995749 185258 995755
rect 179842 993741 179870 995522
rect 180514 993889 180542 995522
rect 181152 995508 181406 995536
rect 180502 993883 180554 993889
rect 180502 993825 180554 993831
rect 181378 993815 181406 995508
rect 183010 995221 183038 995522
rect 184162 995295 184190 995522
rect 184848 995508 185150 995536
rect 185122 995443 185150 995508
rect 185110 995437 185162 995443
rect 185110 995379 185162 995385
rect 184150 995289 184202 995295
rect 184150 995231 184202 995237
rect 182998 995215 183050 995221
rect 182998 995157 183050 995163
rect 181366 993809 181418 993815
rect 181366 993751 181418 993757
rect 179830 993735 179882 993741
rect 179830 993677 179882 993683
rect 185410 993667 185438 995804
rect 190368 995807 190634 995813
rect 190368 995804 190582 995807
rect 188854 995749 188906 995755
rect 192192 995804 192500 995832
rect 192500 995781 192556 995790
rect 190582 995749 190634 995755
rect 188086 995733 188138 995739
rect 186048 995656 186206 995684
rect 187872 995681 188086 995684
rect 187872 995675 188138 995681
rect 187872 995656 188126 995675
rect 194064 995665 194462 995684
rect 195106 995665 195134 999375
rect 194064 995659 194474 995665
rect 194064 995656 194422 995659
rect 185398 993661 185450 993667
rect 186178 993635 186206 995656
rect 194422 995601 194474 995607
rect 195094 995659 195146 995665
rect 195094 995601 195146 995607
rect 195202 995591 195230 999449
rect 195298 995855 195326 1003223
rect 209108 1003181 209110 1003190
rect 209162 1003181 209164 1003190
rect 211796 1003246 211852 1003255
rect 213826 1003213 213854 1005105
rect 211796 1003181 211798 1003190
rect 209110 1003149 209162 1003155
rect 211850 1003181 211852 1003190
rect 213814 1003207 213866 1003213
rect 211798 1003149 211850 1003155
rect 213814 1003149 213866 1003155
rect 195478 999655 195530 999661
rect 195478 999597 195530 999603
rect 195284 995846 195340 995855
rect 195284 995781 195340 995790
rect 191926 995585 191978 995591
rect 189428 995550 189484 995559
rect 187330 994079 187358 995522
rect 189168 995508 189428 995536
rect 191568 995533 191926 995536
rect 191568 995527 191978 995533
rect 195190 995585 195242 995591
rect 195190 995527 195242 995533
rect 191568 995508 191966 995527
rect 189428 995485 189484 995494
rect 187316 994070 187372 994079
rect 187316 994005 187372 994014
rect 195490 993635 195518 999597
rect 206902 999433 206954 999439
rect 206900 999398 206902 999407
rect 206954 999398 206956 999407
rect 206900 999333 206956 999342
rect 196822 996695 196874 996701
rect 196822 996637 196874 996643
rect 195766 996547 195818 996553
rect 195766 996489 195818 996495
rect 195778 995295 195806 996489
rect 195766 995289 195818 995295
rect 195766 995231 195818 995237
rect 196834 995221 196862 996637
rect 205172 996586 205228 996595
rect 205172 996521 205174 996530
rect 205226 996521 205228 996530
rect 207956 996586 208012 996595
rect 207956 996521 207958 996530
rect 205174 996489 205226 996495
rect 208010 996521 208012 996530
rect 207958 996489 208010 996495
rect 210164 996142 210220 996151
rect 210164 996077 210166 996086
rect 210218 996077 210220 996086
rect 210166 996045 210218 996051
rect 222658 996035 222686 1005147
rect 226006 999507 226058 999513
rect 226006 999449 226058 999455
rect 222934 999433 222986 999439
rect 222934 999375 222986 999381
rect 210646 996029 210698 996035
rect 204020 995994 204076 996003
rect 204020 995929 204076 995938
rect 210644 995994 210646 996003
rect 222646 996029 222698 996035
rect 210698 995994 210700 996003
rect 210644 995929 210700 995938
rect 211796 995994 211852 996003
rect 211796 995929 211798 995938
rect 204034 995887 204062 995929
rect 211850 995929 211852 995938
rect 219092 995994 219148 996003
rect 222646 995971 222698 995977
rect 219092 995929 219148 995938
rect 211798 995897 211850 995903
rect 204022 995881 204074 995887
rect 203060 995846 203116 995855
rect 203060 995781 203116 995790
rect 203636 995846 203692 995855
rect 204022 995823 204074 995829
rect 204692 995846 204748 995855
rect 203636 995781 203692 995790
rect 204692 995781 204694 995790
rect 203074 995739 203102 995781
rect 203062 995733 203114 995739
rect 197204 995698 197260 995707
rect 203062 995675 203114 995681
rect 197204 995633 197260 995642
rect 196822 995215 196874 995221
rect 196822 995157 196874 995163
rect 185398 993603 185450 993609
rect 186164 993626 186220 993635
rect 186164 993561 186220 993570
rect 195476 993626 195532 993635
rect 195476 993561 195532 993570
rect 186934 988259 186986 988265
rect 186934 988201 186986 988207
rect 169954 983520 170736 983548
rect 186946 983534 186974 988201
rect 197218 986415 197246 995633
rect 203650 995443 203678 995781
rect 204746 995781 204748 995790
rect 213332 995846 213388 995855
rect 213332 995781 213388 995790
rect 204694 995749 204746 995755
rect 203638 995437 203690 995443
rect 203638 995379 203690 995385
rect 208724 995402 208780 995411
rect 208724 995337 208780 995346
rect 198644 995254 198700 995263
rect 198644 995189 198700 995198
rect 198658 993889 198686 995189
rect 198646 993883 198698 993889
rect 198646 993825 198698 993831
rect 208738 993741 208766 995337
rect 209780 995254 209836 995263
rect 209780 995189 209836 995198
rect 209794 993815 209822 995189
rect 209782 993809 209834 993815
rect 209782 993751 209834 993757
rect 208726 993735 208778 993741
rect 208726 993677 208778 993683
rect 213346 989375 213374 995781
rect 216020 995698 216076 995707
rect 216020 995633 216076 995642
rect 203158 989369 203210 989375
rect 203158 989311 203210 989317
rect 213334 989369 213386 989375
rect 213334 989311 213386 989317
rect 197206 986409 197258 986415
rect 197206 986351 197258 986357
rect 203170 983534 203198 989311
rect 216034 989301 216062 995633
rect 216022 989295 216074 989301
rect 216022 989237 216074 989243
rect 219106 983548 219134 995929
rect 222946 995073 222974 999375
rect 225238 996399 225290 996405
rect 225238 996341 225290 996347
rect 225250 996109 225278 996341
rect 225238 996103 225290 996109
rect 225238 996045 225290 996051
rect 226018 995813 226046 999449
rect 246550 999433 246602 999439
rect 246550 999375 246602 999381
rect 239540 995846 239596 995855
rect 236256 995813 236510 995832
rect 226006 995807 226058 995813
rect 236256 995807 236522 995813
rect 236256 995804 236470 995807
rect 226006 995749 226058 995755
rect 239280 995804 239540 995832
rect 239540 995781 239596 995790
rect 236470 995749 236522 995755
rect 246562 995739 246590 999375
rect 247510 996103 247562 996109
rect 247510 996045 247562 996051
rect 245686 995733 245738 995739
rect 240788 995698 240844 995707
rect 237238 995659 237290 995665
rect 240576 995656 240788 995684
rect 245424 995681 245686 995684
rect 245424 995675 245738 995681
rect 246550 995733 246602 995739
rect 246550 995675 246602 995681
rect 245424 995656 245726 995675
rect 240788 995633 240844 995642
rect 237238 995601 237290 995607
rect 237250 995536 237278 995601
rect 243860 995550 243916 995559
rect 231264 995508 231518 995536
rect 231936 995508 232190 995536
rect 222934 995067 222986 995073
rect 222934 995009 222986 995015
rect 231490 993815 231518 995508
rect 232162 994523 232190 995508
rect 232148 994514 232204 994523
rect 232148 994449 232204 994458
rect 231478 993809 231530 993815
rect 231478 993751 231530 993757
rect 232546 993741 232574 995522
rect 234370 994227 234398 995522
rect 234356 994218 234412 994227
rect 234356 994153 234412 994162
rect 234946 993963 234974 995522
rect 235584 995508 235838 995536
rect 237250 995522 237456 995536
rect 235810 994671 235838 995508
rect 235796 994662 235852 994671
rect 235796 994597 235852 994606
rect 234934 993957 234986 993963
rect 234934 993899 234986 993905
rect 232534 993735 232586 993741
rect 232534 993677 232586 993683
rect 236770 993667 236798 995522
rect 237250 995508 237470 995522
rect 237442 994999 237470 995508
rect 237430 994993 237482 994999
rect 237430 994935 237482 994941
rect 238690 993889 238718 995522
rect 239952 995508 240254 995536
rect 240226 995411 240254 995508
rect 240212 995402 240268 995411
rect 240212 995337 240268 995346
rect 241762 995263 241790 995522
rect 242976 995508 243230 995536
rect 243600 995508 243860 995536
rect 241748 995254 241804 995263
rect 241748 995189 241804 995198
rect 239446 994105 239498 994111
rect 243202 994079 243230 995508
rect 243860 995485 243916 995494
rect 247522 994523 247550 996045
rect 250486 995955 250538 995961
rect 250486 995897 250538 995903
rect 250498 995855 250526 995897
rect 250484 995846 250540 995855
rect 250484 995781 250540 995790
rect 250390 995733 250442 995739
rect 250390 995675 250442 995681
rect 247606 995659 247658 995665
rect 247606 995601 247658 995607
rect 247618 994671 247646 995601
rect 250100 995550 250156 995559
rect 250100 995485 250156 995494
rect 250114 995115 250142 995485
rect 250100 995106 250156 995115
rect 250100 995041 250156 995050
rect 247604 994662 247660 994671
rect 247604 994597 247660 994606
rect 247508 994514 247564 994523
rect 247508 994449 247564 994458
rect 239446 994047 239498 994053
rect 243188 994070 243244 994079
rect 238678 993883 238730 993889
rect 238678 993825 238730 993831
rect 239458 993667 239486 994047
rect 243188 994005 243244 994014
rect 250402 993963 250430 995675
rect 250486 994993 250538 994999
rect 250486 994935 250538 994941
rect 250390 993957 250442 993963
rect 250390 993899 250442 993905
rect 250498 993667 250526 994935
rect 236758 993661 236810 993667
rect 236758 993603 236810 993609
rect 239446 993661 239498 993667
rect 239446 993603 239498 993609
rect 250486 993661 250538 993667
rect 250486 993603 250538 993609
rect 251362 993593 251390 1015909
rect 348884 1007834 348940 1007843
rect 348884 1007769 348940 1007778
rect 353300 1007834 353356 1007843
rect 353410 1007820 353438 1015909
rect 452182 1008165 452234 1008171
rect 452182 1008107 452234 1008113
rect 472150 1008165 472202 1008171
rect 472150 1008107 472202 1008113
rect 434998 1008091 435050 1008097
rect 434998 1008033 435050 1008039
rect 434710 1008017 434762 1008023
rect 434710 1007959 434762 1007965
rect 353356 1007792 353438 1007820
rect 353300 1007769 353356 1007778
rect 316822 1005205 316874 1005211
rect 316822 1005147 316874 1005153
rect 331222 1005205 331274 1005211
rect 331222 1005147 331274 1005153
rect 316436 1003246 316492 1003255
rect 316834 1003232 316862 1005147
rect 316492 1003204 316862 1003232
rect 316436 1003181 316492 1003190
rect 298294 1002985 298346 1002991
rect 312118 1002985 312170 1002991
rect 298294 1002927 298346 1002933
rect 308852 1002950 308908 1002959
rect 258358 999433 258410 999439
rect 258356 999398 258358 999407
rect 298198 999433 298250 999439
rect 258410 999398 258412 999407
rect 298198 999375 298250 999381
rect 258356 999333 258412 999342
rect 270644 997178 270700 997187
rect 270644 997113 270700 997122
rect 298100 997178 298156 997187
rect 298100 997113 298102 997122
rect 262484 996438 262540 996447
rect 270658 996405 270686 997113
rect 298154 997113 298156 997122
rect 298102 997081 298154 997087
rect 262484 996373 262486 996382
rect 262538 996373 262540 996382
rect 270646 996399 270698 996405
rect 262486 996341 262538 996347
rect 270646 996341 270698 996347
rect 263062 996177 263114 996183
rect 257780 996142 257836 996151
rect 257780 996077 257782 996086
rect 257834 996077 257836 996086
rect 262004 996142 262060 996151
rect 262004 996077 262006 996086
rect 257782 996045 257834 996051
rect 262058 996077 262060 996086
rect 263060 996142 263062 996151
rect 263114 996142 263116 996151
rect 263060 996077 263116 996086
rect 262006 996045 262058 996051
rect 263254 996029 263306 996035
rect 254516 995994 254572 996003
rect 254516 995929 254518 995938
rect 254570 995929 254572 995938
rect 254900 995994 254956 996003
rect 254900 995929 254956 995938
rect 261044 995994 261100 996003
rect 261044 995929 261100 995938
rect 263252 995994 263254 996003
rect 263306 995994 263308 996003
rect 263252 995929 263308 995938
rect 254518 995897 254570 995903
rect 254914 995813 254942 995929
rect 256148 995846 256204 995855
rect 254902 995807 254954 995813
rect 256148 995781 256204 995790
rect 257108 995846 257164 995855
rect 257108 995781 257164 995790
rect 259220 995846 259276 995855
rect 259220 995781 259276 995790
rect 254902 995749 254954 995755
rect 255956 995698 256012 995707
rect 255956 995633 255958 995642
rect 256010 995633 256012 995642
rect 255958 995601 256010 995607
rect 256162 995263 256190 995781
rect 257122 995739 257150 995781
rect 257110 995733 257162 995739
rect 257110 995675 257162 995681
rect 259028 995550 259084 995559
rect 259028 995485 259084 995494
rect 256148 995254 256204 995263
rect 256148 995189 256204 995198
rect 259042 993889 259070 995485
rect 259234 994227 259262 995781
rect 260084 995254 260140 995263
rect 260084 995189 260140 995198
rect 259220 994218 259276 994227
rect 259220 994153 259276 994162
rect 259030 993883 259082 993889
rect 259030 993825 259082 993831
rect 260098 993815 260126 995189
rect 260086 993809 260138 993815
rect 260086 993751 260138 993757
rect 261058 993741 261086 995929
rect 270740 995846 270796 995855
rect 287924 995846 287980 995855
rect 283536 995813 283742 995832
rect 283536 995807 283754 995813
rect 283536 995804 283702 995807
rect 270740 995781 270796 995790
rect 267860 995698 267916 995707
rect 267860 995633 267916 995642
rect 261046 993735 261098 993741
rect 261046 993677 261098 993683
rect 237430 993587 237482 993593
rect 237430 993529 237482 993535
rect 251350 993587 251402 993593
rect 251350 993529 251402 993535
rect 235606 989295 235658 989301
rect 235606 989237 235658 989243
rect 219106 983520 219408 983548
rect 235618 983534 235646 989237
rect 237442 983603 237470 993529
rect 251830 988185 251882 988191
rect 251830 988127 251882 988133
rect 237430 983597 237482 983603
rect 237430 983539 237482 983545
rect 251842 983534 251870 988127
rect 267874 983548 267902 995633
rect 267956 995550 268012 995559
rect 267956 995485 268012 995494
rect 267970 989301 267998 995485
rect 270754 989375 270782 995781
rect 287856 995804 287924 995832
rect 290352 995813 290654 995832
rect 292176 995813 292574 995832
rect 290352 995807 290666 995813
rect 290352 995804 290614 995807
rect 287924 995781 287980 995790
rect 283702 995749 283754 995755
rect 292176 995807 292586 995813
rect 292176 995804 292534 995807
rect 290614 995749 290666 995755
rect 292534 995749 292586 995755
rect 291190 995733 291242 995739
rect 286772 995698 286828 995707
rect 286560 995656 286772 995684
rect 290880 995681 291190 995684
rect 290880 995675 291242 995681
rect 290880 995656 291230 995675
rect 297072 995665 297374 995684
rect 298210 995665 298238 999375
rect 297072 995659 297386 995665
rect 297072 995656 297334 995659
rect 286772 995633 286828 995642
rect 297334 995601 297386 995607
rect 298198 995659 298250 995665
rect 298198 995601 298250 995607
rect 298306 995591 298334 1002927
rect 299350 1002911 299402 1002917
rect 308852 1002885 308854 1002894
rect 299350 1002853 299402 1002859
rect 308906 1002885 308908 1002894
rect 312116 1002950 312118 1002959
rect 312170 1002950 312172 1002959
rect 312116 1002885 312172 1002894
rect 308854 1002853 308906 1002859
rect 299254 1002763 299306 1002769
rect 299254 1002705 299306 1002711
rect 298390 997953 298442 997959
rect 298390 997895 298442 997901
rect 295414 995585 295466 995591
rect 287444 995550 287500 995559
rect 279286 994105 279338 994111
rect 279286 994047 279338 994053
rect 279298 993593 279326 994047
rect 282850 993815 282878 995522
rect 284160 995508 284414 995536
rect 282838 993809 282890 993815
rect 282838 993751 282890 993757
rect 284386 993741 284414 995508
rect 286018 994523 286046 995522
rect 287184 995508 287444 995536
rect 287444 995485 287500 995494
rect 288130 995508 288384 995536
rect 289056 995508 289310 995536
rect 286004 994514 286060 994523
rect 286004 994449 286060 994458
rect 284374 993735 284426 993741
rect 284374 993677 284426 993683
rect 288130 993593 288158 995508
rect 289282 994851 289310 995508
rect 291490 995263 291518 995522
rect 293376 995517 293726 995536
rect 295200 995533 295414 995536
rect 295200 995527 295466 995533
rect 298294 995585 298346 995591
rect 298294 995527 298346 995533
rect 293376 995511 293738 995517
rect 293376 995508 293686 995511
rect 293686 995453 293738 995459
rect 291476 995254 291532 995263
rect 291476 995189 291532 995198
rect 289270 994845 289322 994851
rect 289270 994787 289322 994793
rect 289282 993667 289310 994787
rect 294562 994227 294590 995522
rect 295200 995508 295454 995527
rect 298402 995147 298430 997895
rect 298964 995698 299020 995707
rect 298964 995633 299020 995642
rect 298390 995141 298442 995147
rect 298390 995083 298442 995089
rect 296662 994845 296714 994851
rect 296662 994787 296714 994793
rect 296674 994375 296702 994787
rect 296660 994366 296716 994375
rect 296660 994301 296716 994310
rect 294548 994218 294604 994227
rect 294548 994153 294604 994162
rect 289270 993661 289322 993667
rect 289270 993603 289322 993609
rect 279286 993587 279338 993593
rect 279286 993529 279338 993535
rect 288118 993587 288170 993593
rect 288118 993529 288170 993535
rect 298978 991817 299006 995633
rect 299266 995559 299294 1002705
rect 299362 995855 299390 1002853
rect 299446 1002837 299498 1002843
rect 309334 1002837 309386 1002843
rect 299446 1002779 299498 1002785
rect 308276 1002802 308332 1002811
rect 299458 995961 299486 1002779
rect 308276 1002737 308278 1002746
rect 308330 1002737 308332 1002746
rect 309332 1002802 309334 1002811
rect 309386 1002802 309388 1002811
rect 309332 1002737 309388 1002746
rect 308278 1002705 308330 1002711
rect 309910 999433 309962 999439
rect 309908 999398 309910 999407
rect 309962 999398 309964 999407
rect 309908 999333 309964 999342
rect 313750 999359 313802 999365
rect 313750 999301 313802 999307
rect 328342 999359 328394 999365
rect 328342 999301 328394 999307
rect 313762 997187 313790 999301
rect 314804 997918 314860 997927
rect 314804 997853 314806 997862
rect 314858 997853 314860 997862
rect 314806 997821 314858 997827
rect 328354 997811 328382 999301
rect 328342 997805 328394 997811
rect 328342 997747 328394 997753
rect 313748 997178 313804 997187
rect 313748 997113 313750 997122
rect 313802 997113 313804 997122
rect 313750 997081 313802 997087
rect 311540 996586 311596 996595
rect 309910 996547 309962 996553
rect 311540 996521 311542 996530
rect 309910 996489 309962 996495
rect 311594 996521 311596 996530
rect 311542 996489 311594 996495
rect 299540 996142 299596 996151
rect 299540 996077 299596 996086
rect 299446 995955 299498 995961
rect 299446 995897 299498 995903
rect 299348 995846 299404 995855
rect 299348 995781 299404 995790
rect 299554 995559 299582 996077
rect 303956 995994 304012 996003
rect 304340 995994 304396 996003
rect 304012 995952 304340 995980
rect 303956 995929 304012 995938
rect 304340 995929 304396 995938
rect 305492 995994 305548 996003
rect 305492 995929 305548 995938
rect 305506 995813 305534 995929
rect 305972 995846 306028 995855
rect 305494 995807 305546 995813
rect 305972 995781 306028 995790
rect 307604 995846 307660 995855
rect 307604 995781 307660 995790
rect 305494 995749 305546 995755
rect 305986 995739 306014 995781
rect 305974 995733 306026 995739
rect 305974 995675 306026 995681
rect 299252 995550 299308 995559
rect 299252 995485 299308 995494
rect 299540 995550 299596 995559
rect 307618 995517 307646 995781
rect 299540 995485 299596 995494
rect 307606 995511 307658 995517
rect 307606 995453 307658 995459
rect 309922 993815 309950 996489
rect 313174 996473 313226 996479
rect 313174 996415 313226 996421
rect 313186 996151 313214 996415
rect 314806 996177 314858 996183
rect 313172 996142 313228 996151
rect 313172 996077 313174 996086
rect 313226 996077 313228 996086
rect 314804 996142 314806 996151
rect 314858 996142 314860 996151
rect 314804 996077 314860 996086
rect 313174 996045 313226 996051
rect 310292 995994 310348 996003
rect 310292 995929 310348 995938
rect 319604 995994 319660 996003
rect 319604 995929 319660 995938
rect 310306 995887 310334 995929
rect 310294 995881 310346 995887
rect 310294 995823 310346 995829
rect 312788 995402 312844 995411
rect 312788 995337 312844 995346
rect 309910 993809 309962 993815
rect 309910 993751 309962 993757
rect 312802 993741 312830 995337
rect 312790 993735 312842 993741
rect 312790 993677 312842 993683
rect 290902 991811 290954 991817
rect 290902 991753 290954 991759
rect 298966 991811 299018 991817
rect 298966 991753 299018 991759
rect 270742 989369 270794 989375
rect 270742 989311 270794 989317
rect 284278 989369 284330 989375
rect 284278 989311 284330 989317
rect 267958 989295 268010 989301
rect 267958 989237 268010 989243
rect 267874 983520 268080 983548
rect 284290 983534 284318 989311
rect 290914 985028 290942 991753
rect 319618 989375 319646 995929
rect 319700 995698 319756 995707
rect 319700 995633 319756 995642
rect 319606 989369 319658 989375
rect 319606 989311 319658 989317
rect 319714 989301 319742 995633
rect 331234 992631 331262 1005147
rect 348898 997959 348926 1007769
rect 367222 1005501 367274 1005507
rect 367222 1005443 367274 1005449
rect 383638 1005501 383690 1005507
rect 383638 1005443 383690 1005449
rect 434614 1005501 434666 1005507
rect 434614 1005443 434666 1005449
rect 357428 1003246 357484 1003255
rect 357428 1003181 357430 1003190
rect 357482 1003181 357484 1003190
rect 362516 1003246 362572 1003255
rect 367234 1003213 367262 1005443
rect 377302 1003281 377354 1003287
rect 377302 1003223 377354 1003229
rect 362516 1003181 362518 1003190
rect 357430 1003149 357482 1003155
rect 362570 1003181 362572 1003190
rect 367222 1003207 367274 1003213
rect 362518 1003149 362570 1003155
rect 367222 1003149 367274 1003155
rect 358580 1002802 358636 1002811
rect 358580 1002737 358582 1002746
rect 358634 1002737 358636 1002746
rect 373366 1002763 373418 1002769
rect 358582 1002705 358634 1002711
rect 373366 1002705 373418 1002711
rect 358006 1002689 358058 1002695
rect 358004 1002654 358006 1002663
rect 372502 1002689 372554 1002695
rect 358058 1002654 358060 1002663
rect 372502 1002631 372554 1002637
rect 358004 1002589 358060 1002598
rect 361846 1002541 361898 1002547
rect 361844 1002506 361846 1002515
rect 371542 1002541 371594 1002547
rect 361898 1002506 361900 1002515
rect 371542 1002483 371594 1002489
rect 361844 1002441 361900 1002450
rect 362902 1002393 362954 1002399
rect 359060 1002358 359116 1002367
rect 359060 1002293 359062 1002302
rect 359114 1002293 359116 1002302
rect 362900 1002358 362902 1002367
rect 362954 1002358 362956 1002367
rect 362900 1002293 362956 1002302
rect 365782 1002319 365834 1002325
rect 359062 1002261 359114 1002267
rect 365782 1002261 365834 1002267
rect 361366 1002245 361418 1002251
rect 361364 1002210 361366 1002219
rect 361418 1002210 361420 1002219
rect 361364 1002145 361420 1002154
rect 356372 1001322 356428 1001331
rect 356372 1001257 356374 1001266
rect 356426 1001257 356428 1001266
rect 356374 1001225 356426 1001231
rect 357044 1001174 357100 1001183
rect 357100 1001141 357182 1001160
rect 357100 1001135 357194 1001141
rect 357100 1001132 357142 1001135
rect 357044 1001109 357100 1001118
rect 357142 1001077 357194 1001083
rect 365794 1000993 365822 1002261
rect 365782 1000987 365834 1000993
rect 365782 1000929 365834 1000935
rect 360214 1000913 360266 1000919
rect 359636 1000878 359692 1000887
rect 359636 1000813 359638 1000822
rect 359690 1000813 359692 1000822
rect 360212 1000878 360214 1000887
rect 360266 1000878 360268 1000887
rect 360212 1000813 360268 1000822
rect 359638 1000781 359690 1000787
rect 371554 999513 371582 1002483
rect 371638 1002393 371690 1002399
rect 371638 1002335 371690 1002341
rect 371542 999507 371594 999513
rect 371542 999449 371594 999455
rect 371650 999439 371678 1002335
rect 371638 999433 371690 999439
rect 364532 999398 364588 999407
rect 371638 999375 371690 999381
rect 364532 999333 364534 999342
rect 364586 999333 364588 999342
rect 364534 999301 364586 999307
rect 348886 997953 348938 997959
rect 348886 997895 348938 997901
rect 364546 997811 364574 999301
rect 365204 997918 365260 997927
rect 365204 997853 365206 997862
rect 365258 997853 365260 997862
rect 365206 997821 365258 997827
rect 364534 997805 364586 997811
rect 364534 997747 364586 997753
rect 363958 996473 364010 996479
rect 363958 996415 364010 996421
rect 363970 996035 363998 996415
rect 368662 996177 368714 996183
rect 368662 996119 368714 996125
rect 363958 996029 364010 996035
rect 363956 995994 363958 996003
rect 364010 995994 364012 996003
rect 363956 995929 364012 995938
rect 360884 995846 360940 995855
rect 366164 995846 366220 995855
rect 360884 995781 360886 995790
rect 360938 995781 360940 995790
rect 365782 995807 365834 995813
rect 360886 995749 360938 995755
rect 366164 995781 366220 995790
rect 366740 995846 366796 995855
rect 366740 995781 366742 995790
rect 365782 995749 365834 995755
rect 365794 993667 365822 995749
rect 366178 995739 366206 995781
rect 366794 995781 366796 995790
rect 366742 995749 366794 995755
rect 366166 995733 366218 995739
rect 368674 995707 368702 996119
rect 371540 995846 371596 995855
rect 371540 995781 371596 995790
rect 371638 995807 371690 995813
rect 366166 995675 366218 995681
rect 368660 995698 368716 995707
rect 368660 995633 368716 995642
rect 365782 993661 365834 993667
rect 365782 993603 365834 993609
rect 331222 992625 331274 992631
rect 331222 992567 331274 992573
rect 332566 992625 332618 992631
rect 332566 992567 332618 992573
rect 300502 989295 300554 989301
rect 300502 989237 300554 989243
rect 319702 989295 319754 989301
rect 319702 989237 319754 989243
rect 290818 985000 290942 985028
rect 290818 983529 290846 985000
rect 300514 983534 300542 989237
rect 316726 988111 316778 988117
rect 316726 988053 316778 988059
rect 316738 983534 316766 988053
rect 332578 983548 332606 992567
rect 371554 989375 371582 995781
rect 371638 995749 371690 995755
rect 371650 989449 371678 995749
rect 371734 995733 371786 995739
rect 371734 995675 371786 995681
rect 371638 989443 371690 989449
rect 371638 989385 371690 989391
rect 348502 989369 348554 989375
rect 348502 989311 348554 989317
rect 371542 989369 371594 989375
rect 371542 989311 371594 989317
rect 348514 983696 348542 989311
rect 371746 989301 371774 995675
rect 372514 993741 372542 1002631
rect 373378 994523 373406 1002705
rect 377314 999883 377342 1003223
rect 379990 1002245 380042 1002251
rect 379990 1002187 380042 1002193
rect 379798 1001283 379850 1001289
rect 379798 1001225 379850 1001231
rect 377302 999877 377354 999883
rect 377302 999819 377354 999825
rect 379810 995443 379838 1001225
rect 379894 999433 379946 999439
rect 379894 999375 379946 999381
rect 379906 996553 379934 999375
rect 380002 998921 380030 1002187
rect 380086 1001135 380138 1001141
rect 380086 1001077 380138 1001083
rect 379990 998915 380042 998921
rect 379990 998857 380042 998863
rect 379894 996547 379946 996553
rect 379894 996489 379946 996495
rect 380098 995517 380126 1001077
rect 383158 1000987 383210 1000993
rect 383158 1000929 383210 1000935
rect 380374 999359 380426 999365
rect 380374 999301 380426 999307
rect 380386 996109 380414 999301
rect 383062 998915 383114 998921
rect 383062 998857 383114 998863
rect 382966 996547 383018 996553
rect 382966 996489 383018 996495
rect 380374 996103 380426 996109
rect 380374 996045 380426 996051
rect 382978 995961 383006 996489
rect 382966 995955 383018 995961
rect 382966 995897 383018 995903
rect 383074 995707 383102 998857
rect 383060 995698 383116 995707
rect 383060 995633 383116 995642
rect 383170 995591 383198 1000929
rect 383446 1000913 383498 1000919
rect 383446 1000855 383498 1000861
rect 383254 1000839 383306 1000845
rect 383254 1000781 383306 1000787
rect 383266 995665 383294 1000781
rect 383350 999877 383402 999883
rect 383350 999819 383402 999825
rect 383362 995887 383390 999819
rect 383350 995881 383402 995887
rect 383350 995823 383402 995829
rect 383458 995739 383486 1000855
rect 383542 999359 383594 999365
rect 383542 999301 383594 999307
rect 383554 995855 383582 999301
rect 383540 995846 383596 995855
rect 383650 995813 383678 1005443
rect 434626 1003287 434654 1005443
rect 434614 1003281 434666 1003287
rect 428660 1003246 428716 1003255
rect 434614 1003223 434666 1003229
rect 428660 1003181 428662 1003190
rect 428714 1003181 428716 1003190
rect 429526 1003207 429578 1003213
rect 428662 1003149 428714 1003155
rect 429526 1003149 429578 1003155
rect 425398 1003133 425450 1003139
rect 425396 1003098 425398 1003107
rect 425450 1003098 425452 1003107
rect 425396 1003033 425452 1003042
rect 428276 1003098 428332 1003107
rect 428276 1003033 428278 1003042
rect 428330 1003033 428332 1003042
rect 429142 1003059 429194 1003065
rect 428278 1003001 428330 1003007
rect 429142 1003001 429194 1003007
rect 426070 1002985 426122 1002991
rect 423860 1002950 423916 1002959
rect 423860 1002885 423862 1002894
rect 423914 1002885 423916 1002894
rect 426068 1002950 426070 1002959
rect 426122 1002950 426124 1002959
rect 426068 1002885 426124 1002894
rect 423862 1002853 423914 1002859
rect 424342 1002837 424394 1002843
rect 424340 1002802 424342 1002811
rect 424394 1002802 424396 1002811
rect 424340 1002737 424396 1002746
rect 424820 1002802 424876 1002811
rect 424820 1002737 424822 1002746
rect 424874 1002737 424876 1002746
rect 424822 1002705 424874 1002711
rect 427606 1002689 427658 1002695
rect 427604 1002654 427606 1002663
rect 427658 1002654 427660 1002663
rect 427604 1002589 427660 1002598
rect 426646 1002541 426698 1002547
rect 426644 1002506 426646 1002515
rect 426698 1002506 426700 1002515
rect 426644 1002441 426700 1002450
rect 427124 1002506 427180 1002515
rect 427124 1002441 427126 1002450
rect 427178 1002441 427180 1002450
rect 427126 1002409 427178 1002415
rect 429154 1002399 429182 1003001
rect 429538 1002843 429566 1003149
rect 430292 1003098 430348 1003107
rect 430292 1003033 430294 1003042
rect 430346 1003033 430348 1003042
rect 430294 1003001 430346 1003007
rect 429526 1002837 429578 1002843
rect 432022 1002837 432074 1002843
rect 429526 1002779 429578 1002785
rect 432020 1002802 432022 1002811
rect 432074 1002802 432076 1002811
rect 432020 1002737 432076 1002746
rect 429236 1002654 429292 1002663
rect 434722 1002621 434750 1007959
rect 434902 1005353 434954 1005359
rect 434902 1005295 434954 1005301
rect 434914 1003065 434942 1005295
rect 434902 1003059 434954 1003065
rect 434902 1003001 434954 1003007
rect 435010 1002843 435038 1008033
rect 452194 1008023 452222 1008107
rect 471574 1008091 471626 1008097
rect 471574 1008033 471626 1008039
rect 452182 1008017 452234 1008023
rect 452182 1007959 452234 1007965
rect 435284 1006354 435340 1006363
rect 435284 1006289 435340 1006298
rect 465620 1006354 465676 1006363
rect 465620 1006289 465676 1006298
rect 435188 1006058 435244 1006067
rect 435188 1005993 435244 1006002
rect 435092 1005910 435148 1005919
rect 435092 1005845 435148 1005854
rect 434998 1002837 435050 1002843
rect 434998 1002779 435050 1002785
rect 429236 1002589 429238 1002598
rect 429290 1002589 429292 1002598
rect 434710 1002615 434762 1002621
rect 429238 1002557 429290 1002563
rect 434710 1002557 434762 1002563
rect 429142 1002393 429194 1002399
rect 429142 1002335 429194 1002341
rect 430966 1000913 431018 1000919
rect 429908 1000878 429964 1000887
rect 429908 1000813 429910 1000822
rect 429962 1000813 429964 1000822
rect 430964 1000878 430966 1000887
rect 431018 1000878 431020 1000887
rect 430964 1000813 431020 1000822
rect 429910 1000781 429962 1000787
rect 432500 996290 432556 996299
rect 432418 996248 432500 996276
rect 432418 996183 432446 996248
rect 432500 996225 432556 996234
rect 432406 996177 432458 996183
rect 432502 996177 432554 996183
rect 432406 996119 432458 996125
rect 432500 996142 432502 996151
rect 432554 996142 432556 996151
rect 435010 996109 435038 1002779
rect 435106 1002695 435134 1005845
rect 435094 1002689 435146 1002695
rect 435094 1002631 435146 1002637
rect 435202 1002547 435230 1005993
rect 435190 1002541 435242 1002547
rect 435190 1002483 435242 1002489
rect 435298 1002473 435326 1006289
rect 465236 1005910 465292 1005919
rect 465236 1005845 465292 1005854
rect 437494 1005279 437546 1005285
rect 437494 1005221 437546 1005227
rect 435382 1003059 435434 1003065
rect 435382 1003001 435434 1003007
rect 435394 1002917 435422 1003001
rect 435382 1002911 435434 1002917
rect 435382 1002853 435434 1002859
rect 435286 1002467 435338 1002473
rect 435286 1002409 435338 1002415
rect 432500 996077 432556 996086
rect 434998 996103 435050 996109
rect 434998 996045 435050 996051
rect 437506 996035 437534 1005221
rect 439126 1003281 439178 1003287
rect 439126 1003223 439178 1003229
rect 439138 1002769 439166 1003223
rect 439222 1002985 439274 1002991
rect 439222 1002927 439274 1002933
rect 439234 1002843 439262 1002927
rect 439222 1002837 439274 1002843
rect 439222 1002779 439274 1002785
rect 439126 1002763 439178 1002769
rect 439126 1002705 439178 1002711
rect 443542 1002393 443594 1002399
rect 443542 1002335 443594 1002341
rect 430966 996029 431018 996035
rect 421556 995994 421612 996003
rect 421556 995929 421612 995938
rect 430964 995994 430966 996003
rect 437494 996029 437546 996035
rect 431018 995994 431020 996003
rect 437494 995971 437546 995977
rect 437876 995994 437932 996003
rect 430964 995929 431020 995938
rect 437876 995929 437932 995938
rect 421570 995887 421598 995929
rect 417526 995881 417578 995887
rect 387476 995846 387532 995855
rect 384418 995813 384672 995832
rect 383540 995781 383596 995790
rect 383638 995807 383690 995813
rect 383638 995749 383690 995755
rect 384406 995807 384672 995813
rect 384458 995804 384672 995807
rect 387532 995804 387792 995832
rect 389410 995813 389664 995832
rect 396706 995813 397008 995832
rect 417526 995823 417578 995829
rect 421558 995881 421610 995887
rect 421558 995823 421610 995829
rect 389398 995807 389664 995813
rect 387476 995781 387532 995790
rect 384406 995749 384458 995755
rect 389450 995804 389664 995807
rect 396694 995807 397008 995813
rect 389398 995749 389450 995755
rect 396746 995804 397008 995807
rect 396694 995749 396746 995755
rect 383446 995733 383498 995739
rect 383446 995675 383498 995681
rect 384982 995733 385034 995739
rect 391796 995698 391852 995707
rect 385034 995681 385296 995684
rect 384982 995675 385296 995681
rect 383254 995659 383306 995665
rect 384994 995656 385296 995675
rect 388066 995665 388368 995684
rect 388054 995659 388368 995665
rect 383254 995601 383306 995607
rect 388106 995656 388368 995659
rect 391852 995656 392112 995684
rect 391796 995633 391852 995642
rect 388054 995601 388106 995607
rect 383158 995585 383210 995591
rect 383158 995527 383210 995533
rect 388822 995585 388874 995591
rect 388874 995533 388992 995536
rect 388822 995527 388992 995533
rect 380086 995511 380138 995517
rect 380086 995453 380138 995459
rect 379798 995437 379850 995443
rect 379798 995379 379850 995385
rect 385954 995263 385982 995522
rect 388834 995508 388992 995527
rect 385940 995254 385996 995263
rect 385940 995189 385996 995198
rect 377300 994810 377356 994819
rect 377300 994745 377356 994754
rect 373364 994514 373420 994523
rect 373364 994449 373420 994458
rect 377314 994375 377342 994745
rect 377300 994366 377356 994375
rect 377300 994301 377356 994310
rect 372502 993735 372554 993741
rect 372502 993677 372554 993683
rect 390178 993593 390206 995522
rect 390850 994819 390878 995522
rect 392386 995517 392688 995536
rect 392374 995511 392688 995517
rect 392426 995508 392688 995511
rect 393058 995508 393312 995536
rect 393730 995508 393984 995536
rect 392374 995453 392426 995459
rect 390836 994810 390892 994819
rect 390836 994745 390892 994754
rect 393058 993741 393086 995508
rect 393730 995443 393758 995508
rect 393718 995437 393770 995443
rect 393718 995379 393770 995385
rect 395170 994523 395198 995522
rect 396322 995263 396350 995522
rect 396308 995254 396364 995263
rect 396308 995189 396364 995198
rect 395156 994514 395212 994523
rect 395156 994449 395212 994458
rect 393046 993735 393098 993741
rect 393046 993677 393098 993683
rect 398818 993667 398846 995522
rect 398806 993661 398858 993667
rect 398806 993603 398858 993609
rect 403124 993626 403180 993635
rect 390166 993587 390218 993593
rect 403124 993561 403126 993570
rect 390166 993529 390218 993535
rect 403178 993561 403180 993570
rect 403126 993529 403178 993535
rect 397846 989443 397898 989449
rect 397846 989385 397898 989391
rect 365398 989295 365450 989301
rect 365398 989237 365450 989243
rect 371734 989295 371786 989301
rect 371734 989237 371786 989243
rect 348514 983668 348830 983696
rect 348802 983548 348830 983668
rect 290806 983523 290858 983529
rect 332578 983520 332976 983548
rect 348802 983520 349200 983548
rect 365410 983534 365438 989237
rect 381622 988037 381674 988043
rect 381622 987979 381674 987985
rect 381634 983534 381662 987979
rect 397858 983534 397886 989385
rect 414070 989369 414122 989375
rect 414070 989311 414122 989317
rect 414082 983534 414110 989311
rect 417538 983529 417566 995823
rect 437780 995698 437836 995707
rect 437780 995633 437836 995642
rect 437794 989449 437822 995633
rect 437782 989443 437834 989449
rect 437782 989385 437834 989391
rect 437890 989375 437918 995929
rect 437972 995550 438028 995559
rect 437972 995485 438028 995494
rect 437878 989369 437930 989375
rect 437878 989311 437930 989317
rect 437986 989301 438014 995485
rect 443554 993667 443582 1002335
rect 465250 1001067 465278 1005845
rect 465526 1002985 465578 1002991
rect 465526 1002927 465578 1002933
rect 465238 1001061 465290 1001067
rect 465238 1001003 465290 1001009
rect 465538 998995 465566 1002927
rect 465526 998989 465578 998995
rect 465526 998931 465578 998937
rect 465634 995559 465662 1006289
rect 466100 1006058 466156 1006067
rect 466100 1005993 466156 1006002
rect 465620 995550 465676 995559
rect 465620 995485 465676 995494
rect 466114 995411 466142 1005993
rect 469366 1005353 469418 1005359
rect 469366 1005295 469418 1005301
rect 466486 1003281 466538 1003287
rect 466486 1003223 466538 1003229
rect 466390 1003207 466442 1003213
rect 466390 1003149 466442 1003155
rect 466294 1003133 466346 1003139
rect 466294 1003075 466346 1003081
rect 466198 1003059 466250 1003065
rect 466198 1003001 466250 1003007
rect 466210 995517 466238 1003001
rect 466306 999291 466334 1003075
rect 466294 999285 466346 999291
rect 466294 999227 466346 999233
rect 466402 995961 466430 1003149
rect 466498 999069 466526 1003223
rect 469378 999384 469406 1005295
rect 470134 1005279 470186 1005285
rect 470134 1005221 470186 1005227
rect 469378 999356 469502 999384
rect 466486 999063 466538 999069
rect 466486 999005 466538 999011
rect 466390 995955 466442 995961
rect 466390 995897 466442 995903
rect 466198 995511 466250 995517
rect 466198 995453 466250 995459
rect 466100 995402 466156 995411
rect 466100 995337 466156 995346
rect 469474 995221 469502 999356
rect 470146 996035 470174 1005221
rect 471586 996109 471614 1008033
rect 471862 1005501 471914 1005507
rect 471862 1005443 471914 1005449
rect 471574 996103 471626 996109
rect 471574 996045 471626 996051
rect 470134 996029 470186 996035
rect 470134 995971 470186 995977
rect 471874 995443 471902 1005443
rect 472054 999285 472106 999291
rect 472054 999227 472106 999233
rect 471958 998989 472010 998995
rect 471958 998931 472010 998937
rect 471970 995961 471998 998931
rect 471958 995955 472010 995961
rect 471958 995897 472010 995903
rect 472066 995707 472094 999227
rect 472052 995698 472108 995707
rect 472052 995633 472108 995642
rect 472162 995591 472190 1008107
rect 519670 1003281 519722 1003287
rect 502388 1003246 502444 1003255
rect 519670 1003223 519722 1003229
rect 502388 1003181 502390 1003190
rect 502442 1003181 502444 1003190
rect 502390 1003149 502442 1003155
rect 501332 1003098 501388 1003107
rect 501332 1003033 501334 1003042
rect 501386 1003033 501388 1003042
rect 502964 1003098 503020 1003107
rect 502964 1003033 502966 1003042
rect 501334 1003001 501386 1003007
rect 503018 1003033 503020 1003042
rect 502966 1003001 503018 1003007
rect 489142 1002319 489194 1002325
rect 489142 1002261 489194 1002267
rect 519094 1002319 519146 1002325
rect 519094 1002261 519146 1002267
rect 472534 1001061 472586 1001067
rect 472534 1001003 472586 1001009
rect 472438 1000913 472490 1000919
rect 472438 1000855 472490 1000861
rect 472246 999063 472298 999069
rect 472246 999005 472298 999011
rect 472258 995855 472286 999005
rect 472244 995846 472300 995855
rect 472244 995781 472300 995790
rect 472450 995665 472478 1000855
rect 472546 995739 472574 1001003
rect 472630 1000839 472682 1000845
rect 472630 1000781 472682 1000787
rect 472642 995813 472670 1000781
rect 488950 999433 489002 999439
rect 488950 999375 489002 999381
rect 478388 995846 478444 995855
rect 473314 995813 473664 995832
rect 472630 995807 472682 995813
rect 472630 995749 472682 995755
rect 473302 995807 473664 995813
rect 473354 995804 473664 995807
rect 478444 995804 478656 995832
rect 481378 995813 481680 995832
rect 483874 995813 484176 995832
rect 481366 995807 481680 995813
rect 478388 995781 478444 995790
rect 473302 995749 473354 995755
rect 481418 995804 481680 995807
rect 483862 995807 484176 995813
rect 481366 995749 481418 995755
rect 483914 995804 484176 995807
rect 485376 995813 485726 995832
rect 488962 995813 488990 999375
rect 485376 995807 485738 995813
rect 485376 995804 485686 995807
rect 483862 995749 483914 995755
rect 485686 995749 485738 995755
rect 488950 995807 489002 995813
rect 488950 995749 489002 995755
rect 472534 995733 472586 995739
rect 472534 995675 472586 995681
rect 474070 995733 474122 995739
rect 482036 995698 482092 995707
rect 474122 995681 474336 995684
rect 474070 995675 474336 995681
rect 472438 995659 472490 995665
rect 474082 995656 474336 995675
rect 474658 995665 474960 995684
rect 474646 995659 474960 995665
rect 472438 995601 472490 995607
rect 474698 995656 474960 995659
rect 482092 995656 482352 995684
rect 482036 995633 482092 995642
rect 474646 995601 474698 995607
rect 472150 995585 472202 995591
rect 472150 995527 472202 995533
rect 476374 995585 476426 995591
rect 477044 995550 477100 995559
rect 476426 995533 476784 995536
rect 476374 995527 476784 995533
rect 476386 995508 476784 995527
rect 477100 995508 477360 995536
rect 477730 995508 477984 995536
rect 477044 995485 477100 995494
rect 471862 995437 471914 995443
rect 477730 995411 477758 995508
rect 471862 995379 471914 995385
rect 477716 995402 477772 995411
rect 477716 995337 477772 995346
rect 469462 995215 469514 995221
rect 469462 995157 469514 995163
rect 443542 993661 443594 993667
rect 479170 993635 479198 995522
rect 479842 994523 479870 995522
rect 480994 995508 481104 995536
rect 482722 995517 482976 995536
rect 482710 995511 482976 995517
rect 480994 995443 481022 995508
rect 482762 995508 482976 995511
rect 482710 995453 482762 995459
rect 480982 995437 481034 995443
rect 480982 995379 481034 995385
rect 485986 995221 486014 995522
rect 485974 995215 486026 995221
rect 485974 995157 486026 995163
rect 479828 994514 479884 994523
rect 479828 994449 479884 994458
rect 487810 993667 487838 995522
rect 487798 993661 487850 993667
rect 443542 993603 443594 993609
rect 479156 993626 479212 993635
rect 489154 993635 489182 1002261
rect 506324 1001026 506380 1001035
rect 506324 1000961 506326 1000970
rect 506378 1000961 506380 1000970
rect 515542 1000987 515594 1000993
rect 506326 1000929 506378 1000935
rect 515542 1000929 515594 1000935
rect 507860 1000878 507916 1000887
rect 507860 1000813 507862 1000822
rect 507914 1000813 507916 1000822
rect 512662 1000839 512714 1000845
rect 507862 1000781 507914 1000787
rect 512662 1000781 512714 1000787
rect 506900 1000730 506956 1000739
rect 506900 1000665 506902 1000674
rect 506954 1000665 506956 1000674
rect 512182 1000691 512234 1000697
rect 506902 1000633 506954 1000639
rect 512182 1000633 512234 1000639
rect 504694 999877 504746 999883
rect 504692 999842 504694 999851
rect 512086 999877 512138 999883
rect 504746 999842 504748 999851
rect 512084 999842 512086 999851
rect 512138 999842 512140 999851
rect 504692 999777 504748 999786
rect 509686 999803 509738 999809
rect 512084 999777 512140 999786
rect 509686 999745 509738 999751
rect 503638 999729 503690 999735
rect 500756 999694 500812 999703
rect 500756 999629 500758 999638
rect 500810 999629 500812 999638
rect 503636 999694 503638 999703
rect 503690 999694 503692 999703
rect 503636 999629 503692 999638
rect 500758 999597 500810 999603
rect 503638 999581 503690 999587
rect 502004 999546 502060 999555
rect 502004 999481 502006 999490
rect 502058 999481 502060 999490
rect 503636 999546 503638 999555
rect 503690 999546 503692 999555
rect 503636 999481 503692 999490
rect 502006 999449 502058 999455
rect 509698 999439 509726 999745
rect 512084 999694 512140 999703
rect 511990 999655 512042 999661
rect 512084 999629 512086 999638
rect 511990 999597 512042 999603
rect 512138 999629 512140 999638
rect 512086 999597 512138 999603
rect 509686 999433 509738 999439
rect 509686 999375 509738 999381
rect 512002 996775 512030 999597
rect 512194 999555 512222 1000633
rect 512674 1000147 512702 1000781
rect 515554 1000295 515582 1000929
rect 515540 1000286 515596 1000295
rect 515540 1000221 515596 1000230
rect 512660 1000138 512716 1000147
rect 512660 1000073 512716 1000082
rect 512276 999990 512332 999999
rect 512276 999925 512332 999934
rect 512290 999735 512318 999925
rect 512278 999729 512330 999735
rect 512278 999671 512330 999677
rect 512180 999546 512236 999555
rect 512086 999507 512138 999513
rect 512180 999481 512236 999490
rect 512086 999449 512138 999455
rect 512098 999407 512126 999449
rect 512084 999398 512140 999407
rect 512084 999333 512140 999342
rect 511990 996769 512042 996775
rect 511990 996711 512042 996717
rect 518326 996769 518378 996775
rect 518326 996711 518378 996717
rect 507478 996621 507530 996627
rect 505748 996586 505804 996595
rect 505748 996521 505750 996530
rect 505802 996521 505804 996530
rect 507476 996586 507478 996595
rect 507530 996586 507532 996595
rect 507476 996521 507532 996530
rect 505750 996489 505802 996495
rect 509590 996177 509642 996183
rect 508916 996142 508972 996151
rect 508916 996077 508918 996086
rect 508970 996077 508972 996086
rect 509588 996142 509590 996151
rect 509974 996177 510026 996183
rect 509642 996142 509644 996151
rect 509974 996119 510026 996125
rect 509588 996077 509644 996086
rect 508918 996045 508970 996051
rect 508342 996029 508394 996035
rect 508340 995994 508342 996003
rect 508394 995994 508396 996003
rect 508340 995929 508396 995938
rect 499316 995846 499372 995855
rect 499316 995781 499372 995790
rect 499330 995559 499358 995781
rect 509986 995707 510014 996119
rect 515540 995994 515596 996003
rect 515540 995929 515596 995938
rect 509972 995698 510028 995707
rect 509972 995633 510028 995642
rect 510262 995585 510314 995591
rect 499316 995550 499372 995559
rect 499316 995485 499372 995494
rect 501812 995550 501868 995559
rect 501812 995485 501868 995494
rect 510260 995550 510262 995559
rect 510314 995550 510316 995559
rect 510260 995485 510316 995494
rect 501826 995221 501854 995485
rect 501814 995215 501866 995221
rect 501814 995157 501866 995163
rect 487798 993603 487850 993609
rect 489140 993626 489196 993635
rect 479156 993561 479212 993570
rect 489140 993561 489196 993570
rect 462742 989443 462794 989449
rect 462742 989385 462794 989391
rect 430294 989295 430346 989301
rect 430294 989237 430346 989243
rect 437974 989295 438026 989301
rect 437974 989237 438026 989243
rect 430306 983534 430334 989237
rect 446518 987963 446570 987969
rect 446518 987905 446570 987911
rect 446530 983534 446558 987905
rect 462754 983534 462782 989385
rect 515554 989375 515582 995929
rect 515636 995698 515692 995707
rect 515636 995633 515692 995642
rect 515650 989449 515678 995633
rect 515732 995550 515788 995559
rect 515732 995485 515788 995494
rect 515638 989443 515690 989449
rect 515638 989385 515690 989391
rect 478966 989369 479018 989375
rect 478966 989311 479018 989317
rect 515542 989369 515594 989375
rect 515542 989311 515594 989317
rect 478978 983534 479006 989311
rect 515746 989301 515774 995485
rect 518338 994671 518366 996711
rect 519106 995295 519134 1002261
rect 519190 996547 519242 996553
rect 519190 996489 519242 996495
rect 519202 995443 519230 996489
rect 519682 995559 519710 1003223
rect 519766 1003207 519818 1003213
rect 519766 1003149 519818 1003155
rect 519778 996003 519806 1003149
rect 555380 1003098 555436 1003107
rect 519862 1003059 519914 1003065
rect 555380 1003033 555382 1003042
rect 519862 1003001 519914 1003007
rect 555434 1003033 555436 1003042
rect 572758 1003059 572810 1003065
rect 555382 1003001 555434 1003007
rect 572758 1003001 572810 1003007
rect 519874 996151 519902 1003001
rect 554326 1002985 554378 1002991
rect 553748 1002950 553804 1002959
rect 553748 1002885 553750 1002894
rect 553802 1002885 553804 1002894
rect 554324 1002950 554326 1002959
rect 554378 1002950 554380 1002959
rect 554324 1002885 554380 1002894
rect 570742 1002911 570794 1002917
rect 553750 1002853 553802 1002859
rect 570742 1002853 570794 1002859
rect 554900 1002802 554956 1002811
rect 554900 1002737 554902 1002746
rect 554954 1002737 554956 1002746
rect 554902 1002705 554954 1002711
rect 553268 1002654 553324 1002663
rect 553268 1002589 553270 1002598
rect 553322 1002589 553324 1002598
rect 553270 1002557 553322 1002563
rect 552308 1000878 552364 1000887
rect 552308 1000813 552310 1000822
rect 552362 1000813 552364 1000822
rect 552310 1000781 552362 1000787
rect 523508 1000286 523564 1000295
rect 523508 1000221 523564 1000230
rect 519958 999803 520010 999809
rect 519958 999745 520010 999751
rect 519860 996142 519916 996151
rect 519860 996077 519916 996086
rect 519764 995994 519820 996003
rect 519764 995929 519820 995938
rect 519668 995550 519724 995559
rect 519668 995485 519724 995494
rect 519190 995437 519242 995443
rect 519190 995379 519242 995385
rect 519094 995289 519146 995295
rect 519094 995231 519146 995237
rect 519970 995147 519998 999745
rect 521302 996621 521354 996627
rect 521302 996563 521354 996569
rect 521314 995369 521342 996563
rect 523522 995707 523550 1000221
rect 523604 1000138 523660 1000147
rect 523604 1000073 523660 1000082
rect 523508 995698 523564 995707
rect 523508 995633 523564 995642
rect 521398 995585 521450 995591
rect 521398 995527 521450 995533
rect 521302 995363 521354 995369
rect 521302 995305 521354 995311
rect 519958 995141 520010 995147
rect 519958 995083 520010 995089
rect 518324 994662 518380 994671
rect 518324 994597 518380 994606
rect 521410 993667 521438 995527
rect 523618 995517 523646 1000073
rect 523700 999990 523756 999999
rect 523700 999925 523756 999934
rect 523714 995855 523742 999925
rect 523988 999842 524044 999851
rect 523988 999777 524044 999786
rect 523796 999694 523852 999703
rect 523796 999629 523852 999638
rect 523700 995846 523756 995855
rect 523700 995781 523756 995790
rect 523810 995591 523838 999629
rect 523892 999546 523948 999555
rect 523892 999481 523948 999490
rect 523906 995665 523934 999481
rect 524002 995739 524030 999777
rect 552982 999433 553034 999439
rect 524084 999398 524140 999407
rect 524084 999333 524140 999342
rect 552884 999398 552940 999407
rect 552940 999381 552982 999384
rect 552940 999375 553034 999381
rect 552940 999356 553022 999375
rect 567382 999359 567434 999365
rect 552884 999333 552940 999342
rect 524098 995813 524126 999333
rect 567382 999301 567434 999307
rect 558838 999285 558890 999291
rect 558836 999250 558838 999259
rect 558890 999250 558892 999259
rect 558836 999185 558892 999194
rect 557206 998841 557258 998847
rect 557204 998806 557206 998815
rect 557258 998806 557260 998815
rect 557204 998741 557260 998750
rect 555956 997918 556012 997927
rect 555956 997853 555958 997862
rect 556010 997853 556012 997862
rect 555958 997821 556010 997827
rect 558166 997805 558218 997811
rect 558164 997770 558166 997779
rect 558218 997770 558220 997779
rect 558164 997705 558220 997714
rect 557782 997657 557834 997663
rect 557780 997622 557782 997631
rect 557834 997622 557836 997631
rect 557780 997557 557836 997566
rect 559412 997622 559468 997631
rect 559412 997557 559414 997566
rect 559466 997557 559468 997566
rect 559414 997525 559466 997531
rect 561046 996177 561098 996183
rect 561044 996142 561046 996151
rect 561098 996142 561100 996151
rect 560182 996103 560234 996109
rect 561044 996077 561100 996086
rect 560182 996045 560234 996051
rect 559606 996029 559658 996035
rect 559606 995971 559658 995977
rect 528404 995846 528460 995855
rect 524086 995807 524138 995813
rect 532820 995846 532876 995855
rect 528460 995804 528768 995832
rect 529846 995807 529898 995813
rect 528404 995781 528460 995790
rect 524086 995749 524138 995755
rect 550484 995846 550540 995855
rect 532876 995804 533088 995832
rect 532820 995781 532876 995790
rect 550484 995781 550540 995790
rect 556532 995846 556588 995855
rect 556532 995781 556534 995790
rect 529846 995749 529898 995755
rect 523990 995733 524042 995739
rect 525334 995733 525386 995739
rect 523990 995675 524042 995681
rect 524770 995665 525072 995684
rect 527828 995698 527884 995707
rect 525386 995681 525744 995684
rect 525334 995675 525744 995681
rect 523894 995659 523946 995665
rect 523894 995601 523946 995607
rect 524758 995659 525072 995665
rect 524810 995656 525072 995659
rect 525346 995656 525744 995675
rect 529858 995684 529886 995749
rect 533396 995698 533452 995707
rect 527884 995656 528192 995684
rect 529858 995656 530064 995684
rect 527828 995633 527884 995642
rect 533452 995656 533712 995684
rect 533396 995633 533452 995642
rect 524758 995601 524810 995607
rect 523798 995585 523850 995591
rect 528982 995585 529034 995591
rect 523798 995527 523850 995533
rect 526114 995517 526368 995536
rect 550498 995559 550526 995781
rect 556586 995781 556588 995790
rect 556534 995749 556586 995755
rect 559618 995707 559646 995971
rect 560194 995707 560222 996045
rect 563254 995807 563306 995813
rect 563254 995749 563306 995755
rect 558932 995698 558988 995707
rect 558932 995633 558988 995642
rect 559604 995698 559660 995707
rect 559604 995633 559606 995642
rect 535316 995550 535372 995559
rect 529034 995533 529392 995536
rect 528982 995527 529392 995533
rect 523606 995511 523658 995517
rect 523606 995453 523658 995459
rect 526102 995511 526368 995517
rect 526154 995508 526368 995511
rect 528994 995508 529392 995527
rect 526102 995453 526154 995459
rect 530578 995295 530606 995522
rect 530566 995289 530618 995295
rect 530566 995231 530618 995237
rect 528214 995215 528266 995221
rect 528214 995157 528266 995163
rect 521398 993661 521450 993667
rect 521398 993603 521450 993609
rect 527638 989443 527690 989449
rect 527638 989385 527690 989391
rect 495190 989295 495242 989301
rect 495190 989237 495242 989243
rect 515734 989295 515786 989301
rect 515734 989237 515786 989243
rect 495202 983534 495230 989237
rect 511414 987889 511466 987895
rect 511414 987831 511466 987837
rect 511426 983534 511454 987831
rect 527650 983534 527678 989385
rect 528226 983603 528254 995157
rect 531202 994523 531230 995522
rect 532258 995517 532512 995536
rect 532246 995511 532512 995517
rect 532298 995508 532512 995511
rect 532246 995453 532298 995459
rect 534370 994671 534398 995522
rect 550484 995550 550540 995559
rect 535372 995508 535584 995536
rect 535316 995485 535372 995494
rect 534356 994662 534412 994671
rect 534356 994597 534412 994606
rect 531188 994514 531244 994523
rect 531188 994449 531244 994458
rect 536770 993931 536798 995522
rect 537394 995369 537422 995522
rect 538978 995508 539232 995536
rect 537382 995363 537434 995369
rect 537382 995305 537434 995311
rect 533684 993922 533740 993931
rect 533684 993857 533740 993866
rect 536756 993922 536812 993931
rect 536756 993857 536812 993866
rect 533698 989449 533726 993857
rect 538978 993667 539006 995508
rect 550484 995485 550540 995494
rect 558946 995221 558974 995633
rect 559658 995633 559660 995642
rect 560180 995698 560236 995707
rect 560180 995633 560236 995642
rect 559606 995601 559658 995607
rect 560194 995591 560222 995633
rect 560182 995585 560234 995591
rect 560182 995527 560234 995533
rect 558934 995215 558986 995221
rect 558934 995157 558986 995163
rect 563266 993889 563294 995749
rect 564598 995659 564650 995665
rect 564598 995601 564650 995607
rect 564502 995585 564554 995591
rect 564502 995527 564554 995533
rect 563254 993883 563306 993889
rect 563254 993825 563306 993831
rect 538966 993661 539018 993667
rect 538966 993603 539018 993609
rect 533686 989443 533738 989449
rect 533686 989385 533738 989391
rect 543766 989369 543818 989375
rect 543766 989311 543818 989317
rect 528214 983597 528266 983603
rect 528214 983539 528266 983545
rect 543778 983534 543806 989311
rect 560086 989295 560138 989301
rect 560086 989237 560138 989243
rect 560098 983534 560126 989237
rect 564514 986489 564542 995527
rect 564502 986483 564554 986489
rect 564502 986425 564554 986431
rect 564610 986415 564638 995601
rect 567284 995402 567340 995411
rect 567284 995337 567340 995346
rect 567298 989301 567326 995337
rect 567394 993815 567422 999301
rect 569972 995846 570028 995855
rect 569972 995781 570028 995790
rect 569876 995698 569932 995707
rect 569876 995633 569932 995642
rect 569780 995550 569836 995559
rect 569780 995485 569836 995494
rect 567382 993809 567434 993815
rect 567382 993751 567434 993757
rect 569794 989375 569822 995485
rect 569890 989597 569918 995633
rect 569878 989591 569930 989597
rect 569878 989533 569930 989539
rect 569986 989523 570014 995781
rect 570754 993963 570782 1002853
rect 571222 1002763 571274 1002769
rect 571222 1002705 571274 1002711
rect 571234 997737 571262 1002705
rect 572770 997959 572798 1003001
rect 573046 1002985 573098 1002991
rect 573046 1002927 573098 1002933
rect 572950 1002615 573002 1002621
rect 572950 1002557 573002 1002563
rect 572758 997953 572810 997959
rect 572758 997895 572810 997901
rect 571222 997731 571274 997737
rect 571222 997673 571274 997679
rect 572962 997441 572990 1002557
rect 572950 997435 573002 997441
rect 572950 997377 573002 997383
rect 570742 993957 570794 993963
rect 570742 993899 570794 993905
rect 573058 993741 573086 1002927
rect 573142 1000839 573194 1000845
rect 573142 1000781 573194 1000787
rect 573154 997515 573182 1000781
rect 613462 999803 613514 999809
rect 613462 999745 613514 999751
rect 625846 999803 625898 999809
rect 625846 999745 625898 999751
rect 610582 999729 610634 999735
rect 610582 999671 610634 999677
rect 604246 999655 604298 999661
rect 604246 999597 604298 999603
rect 596182 999507 596234 999513
rect 596182 999449 596234 999455
rect 593302 999433 593354 999439
rect 593302 999375 593354 999381
rect 573718 999285 573770 999291
rect 573718 999227 573770 999233
rect 573142 997509 573194 997515
rect 573142 997451 573194 997457
rect 573730 994671 573758 999227
rect 573910 998841 573962 998847
rect 573910 998783 573962 998789
rect 573922 994819 573950 998783
rect 593314 997885 593342 999375
rect 593302 997879 593354 997885
rect 593302 997821 593354 997827
rect 596194 997811 596222 999449
rect 604258 997959 604286 999597
rect 609046 999581 609098 999587
rect 609046 999523 609098 999529
rect 604246 997953 604298 997959
rect 604246 997895 604298 997901
rect 596182 997805 596234 997811
rect 596182 997747 596234 997753
rect 609058 997515 609086 999523
rect 610594 997737 610622 999671
rect 610582 997731 610634 997737
rect 610582 997673 610634 997679
rect 613474 997663 613502 999745
rect 625558 999729 625610 999735
rect 625558 999671 625610 999677
rect 625858 999680 625886 999745
rect 625462 999581 625514 999587
rect 625462 999523 625514 999529
rect 613462 997657 613514 997663
rect 613462 997599 613514 997605
rect 622006 997583 622058 997589
rect 622006 997525 622058 997531
rect 609046 997509 609098 997515
rect 609046 997451 609098 997457
rect 621910 997435 621962 997441
rect 621910 997377 621962 997383
rect 621922 995887 621950 997377
rect 621910 995881 621962 995887
rect 621910 995823 621962 995829
rect 622018 995813 622046 997525
rect 625474 995961 625502 999523
rect 625462 995955 625514 995961
rect 625462 995897 625514 995903
rect 622006 995807 622058 995813
rect 622006 995749 622058 995755
rect 625570 995517 625598 999671
rect 625654 999655 625706 999661
rect 625858 999652 625982 999680
rect 625654 999597 625706 999603
rect 625666 995591 625694 999597
rect 625846 999507 625898 999513
rect 625846 999449 625898 999455
rect 625750 999433 625802 999439
rect 625750 999375 625802 999381
rect 625762 995665 625790 999375
rect 625858 995739 625886 999449
rect 625954 995855 625982 999652
rect 625940 995846 625996 995855
rect 629588 995846 629644 995855
rect 627874 995813 628176 995832
rect 625940 995781 625996 995790
rect 627862 995807 628176 995813
rect 627914 995804 628176 995807
rect 629644 995804 630000 995832
rect 631522 995813 631824 995832
rect 635842 995813 636144 995832
rect 631510 995807 631824 995813
rect 629588 995781 629644 995790
rect 627862 995749 627914 995755
rect 631562 995804 631824 995807
rect 635830 995807 636144 995813
rect 631510 995749 631562 995755
rect 635882 995804 636144 995807
rect 638544 995813 638846 995832
rect 638544 995807 638858 995813
rect 638544 995804 638806 995807
rect 635830 995749 635882 995755
rect 638806 995749 638858 995755
rect 649942 995807 649994 995813
rect 649942 995749 649994 995755
rect 625846 995733 625898 995739
rect 625846 995675 625898 995681
rect 626518 995733 626570 995739
rect 626570 995681 626880 995684
rect 626518 995675 626880 995681
rect 625750 995659 625802 995665
rect 626530 995656 626880 995675
rect 627106 995665 627504 995684
rect 627094 995659 627504 995665
rect 625750 995601 625802 995607
rect 627146 995656 627504 995659
rect 627094 995601 627146 995607
rect 625654 995585 625706 995591
rect 625654 995527 625706 995533
rect 630166 995585 630218 995591
rect 630218 995533 630576 995536
rect 630166 995527 630576 995533
rect 625558 995511 625610 995517
rect 630178 995508 630576 995527
rect 630946 995517 631200 995536
rect 630934 995511 631200 995517
rect 625558 995453 625610 995459
rect 630986 995508 631200 995511
rect 630934 995453 630986 995459
rect 632386 995295 632414 995522
rect 633024 995508 633086 995536
rect 632374 995289 632426 995295
rect 627668 995254 627724 995263
rect 632374 995231 632426 995237
rect 627668 995189 627724 995198
rect 573908 994810 573964 994819
rect 573908 994745 573964 994754
rect 573716 994662 573772 994671
rect 573716 994597 573772 994606
rect 573046 993735 573098 993741
rect 573046 993677 573098 993683
rect 627682 992113 627710 995189
rect 627670 992107 627722 992113
rect 627670 992049 627722 992055
rect 592438 989591 592490 989597
rect 592438 989533 592490 989539
rect 569974 989517 570026 989523
rect 569974 989459 570026 989465
rect 576310 989443 576362 989449
rect 576310 989385 576362 989391
rect 569782 989369 569834 989375
rect 569782 989311 569834 989317
rect 567286 989295 567338 989301
rect 567286 989237 567338 989243
rect 564598 986409 564650 986415
rect 564598 986351 564650 986357
rect 576322 983534 576350 989385
rect 592450 983534 592478 989533
rect 608758 989517 608810 989523
rect 608758 989459 608810 989465
rect 608770 983534 608798 989459
rect 624982 989369 625034 989375
rect 624982 989311 625034 989317
rect 624994 983534 625022 989311
rect 632386 983751 632414 995231
rect 633058 994523 633086 995508
rect 634306 994819 634334 995522
rect 634292 994810 634348 994819
rect 634292 994745 634348 994754
rect 633044 994514 633100 994523
rect 633044 994449 633100 994458
rect 632374 983745 632426 983751
rect 632374 983687 632426 983693
rect 633058 983677 633086 994449
rect 634882 993815 634910 995522
rect 635266 995508 635520 995536
rect 635266 993963 635294 995508
rect 635254 993957 635306 993963
rect 635254 993899 635306 993905
rect 634870 993809 634922 993815
rect 634870 993751 634922 993757
rect 637378 993741 637406 995522
rect 639202 994671 639230 995522
rect 639188 994662 639244 994671
rect 639188 994597 639244 994606
rect 640532 993922 640588 993931
rect 641026 993889 641054 995522
rect 649366 995215 649418 995221
rect 649366 995157 649418 995163
rect 643316 994218 643372 994227
rect 643316 994153 643372 994162
rect 640532 993857 640588 993866
rect 641014 993883 641066 993889
rect 637366 993735 637418 993741
rect 637366 993677 637418 993683
rect 640546 989967 640574 993857
rect 641014 993825 641066 993831
rect 641108 993774 641164 993783
rect 641108 993709 641164 993718
rect 640534 989961 640586 989967
rect 640534 989903 640586 989909
rect 633046 983671 633098 983677
rect 633046 983613 633098 983619
rect 641122 983534 641150 993709
rect 643330 989375 643358 994153
rect 643318 989369 643370 989375
rect 643318 989311 643370 989317
rect 417526 983523 417578 983529
rect 290806 983465 290858 983471
rect 417526 983465 417578 983471
rect 368564 278638 368620 278647
rect 293794 278605 294014 278624
rect 67222 278599 67274 278605
rect 67222 278541 67274 278547
rect 268150 278599 268202 278605
rect 268150 278541 268202 278547
rect 293782 278599 294014 278605
rect 293834 278596 294014 278599
rect 293782 278541 293834 278547
rect 65890 272907 65918 277870
rect 65878 272901 65930 272907
rect 65878 272843 65930 272849
rect 67042 272167 67070 277870
rect 67234 273573 67262 278541
rect 255190 278525 255242 278531
rect 233520 278457 233822 278476
rect 254928 278473 255190 278476
rect 257588 278490 257644 278499
rect 254928 278467 255242 278473
rect 233520 278451 233834 278457
rect 233520 278448 233782 278451
rect 254928 278448 255230 278467
rect 257506 278448 257588 278476
rect 233782 278393 233834 278399
rect 240720 278161 241022 278180
rect 240720 278155 241034 278161
rect 240720 278152 240982 278155
rect 240982 278097 241034 278103
rect 222864 278013 223166 278032
rect 222864 278007 223178 278013
rect 222864 278004 223126 278007
rect 223126 277949 223178 277955
rect 184342 277933 184394 277939
rect 67222 273567 67274 273573
rect 67222 273509 67274 273515
rect 67030 272161 67082 272167
rect 67030 272103 67082 272109
rect 68194 270761 68222 277870
rect 69442 272135 69470 277870
rect 70594 272579 70622 277870
rect 70580 272570 70636 272579
rect 70580 272505 70636 272514
rect 71746 272431 71774 277870
rect 71732 272422 71788 272431
rect 71732 272357 71788 272366
rect 69428 272126 69484 272135
rect 69428 272061 69484 272070
rect 72994 271395 73022 277870
rect 74146 272283 74174 277870
rect 74132 272274 74188 272283
rect 74132 272209 74188 272218
rect 72980 271386 73036 271395
rect 72980 271321 73036 271330
rect 75394 270761 75422 277870
rect 76546 272727 76574 277870
rect 76532 272718 76588 272727
rect 76532 272653 76588 272662
rect 77794 270951 77822 277870
rect 78946 272875 78974 277870
rect 80208 277856 80606 277884
rect 79030 273567 79082 273573
rect 79030 273509 79082 273515
rect 78932 272866 78988 272875
rect 78932 272801 78988 272810
rect 77780 270942 77836 270951
rect 77780 270877 77836 270886
rect 68182 270755 68234 270761
rect 68182 270697 68234 270703
rect 69046 270755 69098 270761
rect 69046 270697 69098 270703
rect 75382 270755 75434 270761
rect 75382 270697 75434 270703
rect 77686 270755 77738 270761
rect 77686 270697 77738 270703
rect 67606 267869 67658 267875
rect 67606 267811 67658 267817
rect 67618 253445 67646 267811
rect 67606 253439 67658 253445
rect 67606 253381 67658 253387
rect 65206 246705 65258 246711
rect 65206 246647 65258 246653
rect 65108 246078 65164 246087
rect 65108 246013 65164 246022
rect 69058 243381 69086 270697
rect 74902 253439 74954 253445
rect 74902 253381 74954 253387
rect 74914 249375 74942 253381
rect 74902 249369 74954 249375
rect 74902 249311 74954 249317
rect 77698 243455 77726 270697
rect 79042 269947 79070 273509
rect 79030 269941 79082 269947
rect 79030 269883 79082 269889
rect 80470 246853 80522 246859
rect 80470 246795 80522 246801
rect 80482 246679 80510 246795
rect 80468 246670 80524 246679
rect 80468 246605 80524 246614
rect 80470 246409 80522 246415
rect 80470 246351 80522 246357
rect 80482 246193 80510 246351
rect 80470 246187 80522 246193
rect 80470 246129 80522 246135
rect 80578 243529 80606 277856
rect 81346 273023 81374 277870
rect 81332 273014 81388 273023
rect 81332 272949 81388 272958
rect 82594 271247 82622 277870
rect 83650 273467 83678 277870
rect 83636 273458 83692 273467
rect 83636 273393 83692 273402
rect 84898 272389 84926 277870
rect 86050 273171 86078 277870
rect 86036 273162 86092 273171
rect 86036 273097 86092 273106
rect 84886 272383 84938 272389
rect 84886 272325 84938 272331
rect 86326 272383 86378 272389
rect 86326 272325 86378 272331
rect 82580 271238 82636 271247
rect 82580 271173 82636 271182
rect 83446 269941 83498 269947
rect 83446 269883 83498 269889
rect 83458 264860 83486 269883
rect 83458 264832 83582 264860
rect 83554 259365 83582 264832
rect 83542 259359 83594 259365
rect 83542 259301 83594 259307
rect 86338 243603 86366 272325
rect 87202 271099 87230 277870
rect 88450 273615 88478 277870
rect 88436 273606 88492 273615
rect 88436 273541 88492 273550
rect 89602 272093 89630 277870
rect 89590 272087 89642 272093
rect 89590 272029 89642 272035
rect 90850 271987 90878 277870
rect 92002 273499 92030 277870
rect 91990 273493 92042 273499
rect 91990 273435 92042 273441
rect 92086 272087 92138 272093
rect 92086 272029 92138 272035
rect 90836 271978 90892 271987
rect 90836 271913 90892 271922
rect 87188 271090 87244 271099
rect 87188 271025 87244 271034
rect 90646 249369 90698 249375
rect 90646 249311 90698 249317
rect 86518 246853 86570 246859
rect 86518 246795 86570 246801
rect 86530 246679 86558 246795
rect 86516 246670 86572 246679
rect 86516 246605 86572 246614
rect 90658 244713 90686 249311
rect 90646 244707 90698 244713
rect 90646 244649 90698 244655
rect 92098 243677 92126 272029
rect 93250 271839 93278 277870
rect 94416 277856 95006 277884
rect 93236 271830 93292 271839
rect 93236 271765 93292 271774
rect 94978 243751 95006 277856
rect 95650 273129 95678 277870
rect 95638 273123 95690 273129
rect 95638 273065 95690 273071
rect 96802 271691 96830 277870
rect 96788 271682 96844 271691
rect 96788 271617 96844 271626
rect 98050 270021 98078 277870
rect 99202 272019 99230 277870
rect 99190 272013 99242 272019
rect 99190 271955 99242 271961
rect 100354 271543 100382 277870
rect 100726 273123 100778 273129
rect 100726 273065 100778 273071
rect 100738 271649 100766 273065
rect 101506 272833 101534 277870
rect 101494 272827 101546 272833
rect 101494 272769 101546 272775
rect 100726 271643 100778 271649
rect 100726 271585 100778 271591
rect 100340 271534 100396 271543
rect 100340 271469 100396 271478
rect 102658 271427 102686 277870
rect 103606 272827 103658 272833
rect 103606 272769 103658 272775
rect 102646 271421 102698 271427
rect 102646 271363 102698 271369
rect 98038 270015 98090 270021
rect 98038 269957 98090 269963
rect 100726 270015 100778 270021
rect 100726 269957 100778 269963
rect 95062 259211 95114 259217
rect 95062 259153 95114 259159
rect 95074 244787 95102 259153
rect 95062 244781 95114 244787
rect 95062 244723 95114 244729
rect 100738 243825 100766 269957
rect 103618 243899 103646 272769
rect 103906 272241 103934 277870
rect 105058 272833 105086 277870
rect 105046 272827 105098 272833
rect 105046 272769 105098 272775
rect 103894 272235 103946 272241
rect 103894 272177 103946 272183
rect 106306 271057 106334 277870
rect 106486 272827 106538 272833
rect 106486 272769 106538 272775
rect 106294 271051 106346 271057
rect 106294 270993 106346 270999
rect 106498 243973 106526 272769
rect 107458 272315 107486 277870
rect 108720 277856 109406 277884
rect 107446 272309 107498 272315
rect 107446 272251 107498 272257
rect 109378 244047 109406 277856
rect 109858 271131 109886 277870
rect 111106 272389 111134 277870
rect 111094 272383 111146 272389
rect 111094 272325 111146 272331
rect 109846 271125 109898 271131
rect 109846 271067 109898 271073
rect 112258 244121 112286 277870
rect 113506 271353 113534 277870
rect 114658 276533 114686 277870
rect 114646 276527 114698 276533
rect 114646 276469 114698 276475
rect 115810 272833 115838 277870
rect 115798 272827 115850 272833
rect 115798 272769 115850 272775
rect 113494 271347 113546 271353
rect 113494 271289 113546 271295
rect 116962 271279 116990 277870
rect 118006 272827 118058 272833
rect 118006 272769 118058 272775
rect 116950 271273 117002 271279
rect 116950 271215 117002 271221
rect 118018 244195 118046 272769
rect 118114 272463 118142 277870
rect 119362 272833 119390 277870
rect 119350 272827 119402 272833
rect 119350 272769 119402 272775
rect 118102 272457 118154 272463
rect 118102 272399 118154 272405
rect 120514 271205 120542 277870
rect 120886 272827 120938 272833
rect 120886 272769 120938 272775
rect 120502 271199 120554 271205
rect 120502 271141 120554 271147
rect 120898 244269 120926 272769
rect 121762 272537 121790 277870
rect 122914 272833 122942 277870
rect 124162 272833 124190 277870
rect 122902 272827 122954 272833
rect 122902 272769 122954 272775
rect 123766 272827 123818 272833
rect 123766 272769 123818 272775
rect 124150 272827 124202 272833
rect 124150 272769 124202 272775
rect 121750 272531 121802 272537
rect 121750 272473 121802 272479
rect 121174 271643 121226 271649
rect 121174 271585 121226 271591
rect 121186 271520 121214 271585
rect 120994 271501 121214 271520
rect 120982 271495 121214 271501
rect 121034 271492 121214 271495
rect 120982 271437 121034 271443
rect 123778 244343 123806 272769
rect 125314 272611 125342 277870
rect 126576 277856 126686 277884
rect 126550 272827 126602 272833
rect 126550 272769 126602 272775
rect 125302 272605 125354 272611
rect 125302 272547 125354 272553
rect 126562 247377 126590 272769
rect 126550 247371 126602 247377
rect 126550 247313 126602 247319
rect 126658 244417 126686 277856
rect 127714 272833 127742 277870
rect 128962 273203 128990 277870
rect 128950 273197 129002 273203
rect 128950 273139 129002 273145
rect 130114 272981 130142 277870
rect 130102 272975 130154 272981
rect 130102 272917 130154 272923
rect 131266 272833 131294 277870
rect 132514 273129 132542 277870
rect 132502 273123 132554 273129
rect 132502 273065 132554 273071
rect 133570 272981 133598 277870
rect 134832 277856 135230 277884
rect 132406 272975 132458 272981
rect 132406 272917 132458 272923
rect 133558 272975 133610 272981
rect 133558 272917 133610 272923
rect 127702 272827 127754 272833
rect 127702 272769 127754 272775
rect 129526 272827 129578 272833
rect 129526 272769 129578 272775
rect 131254 272827 131306 272833
rect 131254 272769 131306 272775
rect 132310 272827 132362 272833
rect 132310 272769 132362 272775
rect 129538 247303 129566 272769
rect 129526 247297 129578 247303
rect 129526 247239 129578 247245
rect 132322 247229 132350 272769
rect 132310 247223 132362 247229
rect 132310 247165 132362 247171
rect 132418 244491 132446 272917
rect 135202 247155 135230 277856
rect 135286 272975 135338 272981
rect 135286 272917 135338 272923
rect 135190 247149 135242 247155
rect 135190 247091 135242 247097
rect 135298 244565 135326 272917
rect 135970 272759 135998 277870
rect 137218 272833 137246 277870
rect 137206 272827 137258 272833
rect 137206 272769 137258 272775
rect 138166 272827 138218 272833
rect 138166 272769 138218 272775
rect 135958 272753 136010 272759
rect 135958 272695 136010 272701
rect 138178 244639 138206 272769
rect 138370 267505 138398 277870
rect 139618 272981 139646 277870
rect 139606 272975 139658 272981
rect 139606 272917 139658 272923
rect 140770 270021 140798 277870
rect 142018 272833 142046 277870
rect 143170 273055 143198 277870
rect 144418 273351 144446 277870
rect 144406 273345 144458 273351
rect 144406 273287 144458 273293
rect 143158 273049 143210 273055
rect 143158 272991 143210 272997
rect 142006 272827 142058 272833
rect 142006 272769 142058 272775
rect 143926 272827 143978 272833
rect 143926 272769 143978 272775
rect 140758 270015 140810 270021
rect 140758 269957 140810 269963
rect 141046 270015 141098 270021
rect 141046 269957 141098 269963
rect 138358 267499 138410 267505
rect 138358 267441 138410 267447
rect 140950 267499 141002 267505
rect 140950 267441 141002 267447
rect 140962 247081 140990 267441
rect 140950 247075 141002 247081
rect 140950 247017 141002 247023
rect 139990 244781 140042 244787
rect 139990 244723 140042 244729
rect 138166 244633 138218 244639
rect 138166 244575 138218 244581
rect 135286 244559 135338 244565
rect 135286 244501 135338 244507
rect 132406 244485 132458 244491
rect 132406 244427 132458 244433
rect 126646 244411 126698 244417
rect 126646 244353 126698 244359
rect 123766 244337 123818 244343
rect 123766 244279 123818 244285
rect 120886 244263 120938 244269
rect 120886 244205 120938 244211
rect 118006 244189 118058 244195
rect 118006 244131 118058 244137
rect 112246 244115 112298 244121
rect 112246 244057 112298 244063
rect 109366 244041 109418 244047
rect 109366 243983 109418 243989
rect 106486 243967 106538 243973
rect 106486 243909 106538 243915
rect 103606 243893 103658 243899
rect 103606 243835 103658 243841
rect 100726 243819 100778 243825
rect 100726 243761 100778 243767
rect 94966 243745 95018 243751
rect 94966 243687 95018 243693
rect 92086 243671 92138 243677
rect 92086 243613 92138 243619
rect 86326 243597 86378 243603
rect 86326 243539 86378 243545
rect 80566 243523 80618 243529
rect 80566 243465 80618 243471
rect 77686 243449 77738 243455
rect 77686 243391 77738 243397
rect 69046 243375 69098 243381
rect 69046 243317 69098 243323
rect 54754 242928 54878 242956
rect 54754 242831 54782 242928
rect 54740 242822 54796 242831
rect 54740 242757 54796 242766
rect 54850 242535 54878 242928
rect 106580 242674 106636 242683
rect 106580 242609 106636 242618
rect 126644 242674 126700 242683
rect 126836 242674 126892 242683
rect 126700 242632 126836 242660
rect 126644 242609 126700 242618
rect 126836 242609 126892 242618
rect 138260 242674 138316 242683
rect 138260 242609 138316 242618
rect 54836 242526 54892 242535
rect 54836 242461 54892 242470
rect 95060 242526 95116 242535
rect 106594 242493 106622 242609
rect 138274 242493 138302 242609
rect 95060 242461 95062 242470
rect 95114 242461 95116 242470
rect 106582 242487 106634 242493
rect 95062 242429 95114 242435
rect 106582 242429 106634 242435
rect 138262 242487 138314 242493
rect 138262 242429 138314 242435
rect 140002 239237 140030 244723
rect 139990 239231 140042 239237
rect 139990 239173 140042 239179
rect 141058 224659 141086 269957
rect 143938 247007 143966 272769
rect 145570 272093 145598 277870
rect 146518 273419 146570 273425
rect 146518 273361 146570 273367
rect 146530 273203 146558 273361
rect 146518 273197 146570 273203
rect 146518 273139 146570 273145
rect 146722 273129 146750 277870
rect 146806 273345 146858 273351
rect 146806 273287 146858 273293
rect 146710 273123 146762 273129
rect 146710 273065 146762 273071
rect 146710 272827 146762 272833
rect 146626 272787 146710 272815
rect 146626 272759 146654 272787
rect 146710 272769 146762 272775
rect 146614 272753 146666 272759
rect 146614 272695 146666 272701
rect 145558 272087 145610 272093
rect 145558 272029 145610 272035
rect 146710 272087 146762 272093
rect 146710 272029 146762 272035
rect 143926 247001 143978 247007
rect 143926 246943 143978 246949
rect 146722 246933 146750 272029
rect 146710 246927 146762 246933
rect 146710 246869 146762 246875
rect 145846 246409 145898 246415
rect 145846 246351 145898 246357
rect 145858 246193 145886 246351
rect 145846 246187 145898 246193
rect 145846 246129 145898 246135
rect 142486 244707 142538 244713
rect 142486 244649 142538 244655
rect 142498 237651 142526 244649
rect 144020 242378 144076 242387
rect 144020 242313 144076 242322
rect 144034 242049 144062 242313
rect 144022 242043 144074 242049
rect 144022 241985 144074 241991
rect 146036 240602 146092 240611
rect 146036 240537 146092 240546
rect 144116 238678 144172 238687
rect 144116 238613 144172 238622
rect 142484 237642 142540 237651
rect 142484 237577 142540 237586
rect 144020 236310 144076 236319
rect 144020 236245 144022 236254
rect 144074 236245 144076 236254
rect 144022 236213 144074 236219
rect 144130 236203 144158 238613
rect 144118 236197 144170 236203
rect 144118 236139 144170 236145
rect 144020 233646 144076 233655
rect 144020 233581 144076 233590
rect 144034 233317 144062 233581
rect 144022 233311 144074 233317
rect 144022 233253 144074 233259
rect 144116 232166 144172 232175
rect 144116 232101 144172 232110
rect 144020 231426 144076 231435
rect 144020 231361 144076 231370
rect 144034 230579 144062 231361
rect 144022 230573 144074 230579
rect 144022 230515 144074 230521
rect 144130 230505 144158 232101
rect 144118 230499 144170 230505
rect 144118 230441 144170 230447
rect 144212 230242 144268 230251
rect 144212 230177 144268 230186
rect 144116 228466 144172 228475
rect 144116 228401 144172 228410
rect 144020 227874 144076 227883
rect 144020 227809 144076 227818
rect 144034 227767 144062 227809
rect 144022 227761 144074 227767
rect 144022 227703 144074 227709
rect 144130 227693 144158 228401
rect 144118 227687 144170 227693
rect 144118 227629 144170 227635
rect 144226 227619 144254 230177
rect 144214 227613 144266 227619
rect 144214 227555 144266 227561
rect 141046 224653 141098 224659
rect 141046 224595 141098 224601
rect 144404 223730 144460 223739
rect 144404 223665 144460 223674
rect 144418 221847 144446 223665
rect 144406 221841 144458 221847
rect 144406 221783 144458 221789
rect 144404 220178 144460 220187
rect 144404 220113 144460 220122
rect 144418 218961 144446 220113
rect 144406 218955 144458 218961
rect 144406 218897 144458 218903
rect 146050 216020 146078 240537
rect 146818 237628 146846 273287
rect 147970 273203 147998 277870
rect 149136 277856 149630 277884
rect 147862 273197 147914 273203
rect 147862 273139 147914 273145
rect 147958 273197 148010 273203
rect 147958 273139 148010 273145
rect 147874 272759 147902 273139
rect 147862 272753 147914 272759
rect 147862 272695 147914 272701
rect 149602 245791 149630 277856
rect 149686 273197 149738 273203
rect 149686 273139 149738 273145
rect 149588 245782 149644 245791
rect 149588 245717 149644 245726
rect 146434 237600 146846 237628
rect 148342 237603 148394 237609
rect 146228 236902 146284 236911
rect 146228 236837 146284 236846
rect 146132 225062 146188 225071
rect 146132 224997 146188 225006
rect 146146 224733 146174 224997
rect 146134 224727 146186 224733
rect 146134 224669 146186 224675
rect 146242 216149 146270 236837
rect 146434 224585 146462 237600
rect 148342 237545 148394 237551
rect 146516 235126 146572 235135
rect 146516 235061 146572 235070
rect 146422 224579 146474 224585
rect 146422 224521 146474 224527
rect 146230 216143 146282 216149
rect 146230 216085 146282 216091
rect 146326 216069 146378 216075
rect 146050 215992 146270 216020
rect 146326 216011 146378 216017
rect 144404 215294 144460 215303
rect 144404 215229 144460 215238
rect 144418 213189 144446 215229
rect 145364 214554 145420 214563
rect 145364 214489 145420 214498
rect 144406 213183 144458 213189
rect 144406 213125 144458 213131
rect 145268 211742 145324 211751
rect 145268 211677 145324 211686
rect 145282 210303 145310 211677
rect 145270 210297 145322 210303
rect 145270 210239 145322 210245
rect 144020 203306 144076 203315
rect 144020 203241 144076 203250
rect 144034 201645 144062 203241
rect 144022 201639 144074 201645
rect 144022 201581 144074 201587
rect 144500 199606 144556 199615
rect 144500 199541 144556 199550
rect 144020 199014 144076 199023
rect 144020 198949 144022 198958
rect 144074 198949 144076 198958
rect 144022 198917 144074 198923
rect 144514 198759 144542 199541
rect 144502 198753 144554 198759
rect 144502 198695 144554 198701
rect 144692 197830 144748 197839
rect 144692 197765 144748 197774
rect 144596 196646 144652 196655
rect 144596 196581 144652 196590
rect 144404 194870 144460 194879
rect 144404 194805 144460 194814
rect 50422 194535 50474 194541
rect 50422 194477 50474 194483
rect 43222 193351 43274 193357
rect 43222 193293 43274 193299
rect 144308 192946 144364 192955
rect 144308 192881 144364 192890
rect 144020 191762 144076 191771
rect 144020 191697 144076 191706
rect 43126 191057 43178 191063
rect 43126 190999 43178 191005
rect 144034 190175 144062 191697
rect 144322 190249 144350 192881
rect 144310 190243 144362 190249
rect 144310 190185 144362 190191
rect 144022 190169 144074 190175
rect 144022 190111 144074 190117
rect 144020 188210 144076 188219
rect 144020 188145 144076 188154
rect 42934 187949 42986 187955
rect 42934 187891 42986 187897
rect 144034 187289 144062 188145
rect 144022 187283 144074 187289
rect 144022 187225 144074 187231
rect 42838 187135 42890 187141
rect 42838 187077 42890 187083
rect 42370 184764 42494 184792
rect 41780 184214 41836 184223
rect 41780 184149 41836 184158
rect 41794 183742 41822 184149
rect 41780 183622 41836 183631
rect 41780 183557 41836 183566
rect 41794 183121 41822 183557
rect 41780 182882 41836 182891
rect 41780 182817 41836 182826
rect 41794 182484 41822 182817
rect 42466 125351 42494 184764
rect 144020 184510 144076 184519
rect 144020 184445 144076 184454
rect 144034 184403 144062 184445
rect 144022 184397 144074 184403
rect 144022 184339 144074 184345
rect 144212 183326 144268 183335
rect 144212 183261 144268 183270
rect 144020 181846 144076 181855
rect 144020 181781 144076 181790
rect 144034 181517 144062 181781
rect 144226 181591 144254 183261
rect 144214 181585 144266 181591
rect 144214 181527 144266 181533
rect 144022 181511 144074 181517
rect 144022 181453 144074 181459
rect 144116 180514 144172 180523
rect 144116 180449 144172 180458
rect 144130 178705 144158 180449
rect 144118 178699 144170 178705
rect 144118 178641 144170 178647
rect 144022 178625 144074 178631
rect 144020 178590 144022 178599
rect 144074 178590 144076 178599
rect 144020 178525 144076 178534
rect 144020 176814 144076 176823
rect 144020 176749 144076 176758
rect 144034 175745 144062 176749
rect 144022 175739 144074 175745
rect 144022 175681 144074 175687
rect 144116 174446 144172 174455
rect 144116 174381 144172 174390
rect 144020 173410 144076 173419
rect 144020 173345 144076 173354
rect 144034 172859 144062 173345
rect 144130 172933 144158 174381
rect 144118 172927 144170 172933
rect 144118 172869 144170 172875
rect 144022 172853 144074 172859
rect 144022 172795 144074 172801
rect 144118 172779 144170 172785
rect 144118 172721 144170 172727
rect 144020 171338 144076 171347
rect 144020 171273 144076 171282
rect 144034 170269 144062 171273
rect 144022 170263 144074 170269
rect 144022 170205 144074 170211
rect 144020 167638 144076 167647
rect 144020 167573 144076 167582
rect 144034 167309 144062 167573
rect 144022 167303 144074 167309
rect 144022 167245 144074 167251
rect 144020 157574 144076 157583
rect 143938 157532 144020 157560
rect 143938 155488 143966 157532
rect 144020 157509 144076 157518
rect 144130 155765 144158 172721
rect 144212 163642 144268 163651
rect 144212 163577 144268 163586
rect 144118 155759 144170 155765
rect 144118 155701 144170 155707
rect 143938 155460 144062 155488
rect 144034 146164 144062 155460
rect 144116 146918 144172 146927
rect 144116 146853 144172 146862
rect 144130 146293 144158 146853
rect 144118 146287 144170 146293
rect 144118 146229 144170 146235
rect 144034 146136 144158 146164
rect 144020 146030 144076 146039
rect 144020 145965 144076 145974
rect 144034 144073 144062 145965
rect 144022 144067 144074 144073
rect 144022 144009 144074 144015
rect 144020 143218 144076 143227
rect 144020 143153 144076 143162
rect 144034 142593 144062 143153
rect 144022 142587 144074 142593
rect 144022 142529 144074 142535
rect 144020 142478 144076 142487
rect 144020 142413 144076 142422
rect 144034 141187 144062 142413
rect 144022 141181 144074 141187
rect 144022 141123 144074 141129
rect 144020 140998 144076 141007
rect 144020 140933 144076 140942
rect 143734 139775 143786 139781
rect 143734 139717 143786 139723
rect 143746 126683 143774 139717
rect 144034 138764 144062 140933
rect 143938 138736 144062 138764
rect 143938 132455 143966 138736
rect 144020 138630 144076 138639
rect 144020 138565 144076 138574
rect 144034 138301 144062 138565
rect 144022 138295 144074 138301
rect 144022 138237 144074 138243
rect 144020 134782 144076 134791
rect 144020 134717 144076 134726
rect 144034 132973 144062 134717
rect 144022 132967 144074 132973
rect 144022 132909 144074 132915
rect 144020 132858 144076 132867
rect 144020 132793 144076 132802
rect 144034 132529 144062 132793
rect 144022 132523 144074 132529
rect 144022 132465 144074 132471
rect 143926 132449 143978 132455
rect 144130 132400 144158 146136
rect 143926 132391 143978 132397
rect 144034 132372 144158 132400
rect 144034 130328 144062 132372
rect 144116 131082 144172 131091
rect 144116 131017 144172 131026
rect 143938 130300 144062 130328
rect 143938 129440 143966 130300
rect 144020 130194 144076 130203
rect 144020 130129 144076 130138
rect 144034 129643 144062 130129
rect 144130 129717 144158 131017
rect 144118 129711 144170 129717
rect 144118 129653 144170 129659
rect 144022 129637 144074 129643
rect 144022 129579 144074 129585
rect 143938 129412 144158 129440
rect 144020 129306 144076 129315
rect 144020 129241 144076 129250
rect 144034 127053 144062 129241
rect 144022 127047 144074 127053
rect 144022 126989 144074 126995
rect 143926 126899 143978 126905
rect 143926 126841 143978 126847
rect 143938 126776 143966 126841
rect 143938 126748 144062 126776
rect 143734 126677 143786 126683
rect 143734 126619 143786 126625
rect 143926 126677 143978 126683
rect 143926 126619 143978 126625
rect 39862 125345 39914 125351
rect 39860 125310 39862 125319
rect 42454 125345 42506 125351
rect 39914 125310 39916 125319
rect 42454 125287 42506 125293
rect 39860 125245 39916 125254
rect 143938 120930 143966 126619
rect 144034 124537 144062 126748
rect 144130 125277 144158 129412
rect 144118 125271 144170 125277
rect 144118 125213 144170 125219
rect 144116 125162 144172 125171
rect 144116 125097 144172 125106
rect 144022 124531 144074 124537
rect 144022 124473 144074 124479
rect 144020 124422 144076 124431
rect 144020 124357 144076 124366
rect 144034 124019 144062 124357
rect 144022 124013 144074 124019
rect 144022 123955 144074 123961
rect 144130 123945 144158 125097
rect 144118 123939 144170 123945
rect 144118 123881 144170 123887
rect 144116 122794 144172 122803
rect 144116 122729 144172 122738
rect 144020 121610 144076 121619
rect 144130 121577 144158 122729
rect 144020 121545 144076 121554
rect 144118 121571 144170 121577
rect 144034 121059 144062 121545
rect 144118 121513 144170 121519
rect 144022 121053 144074 121059
rect 144022 120995 144074 121001
rect 143938 120902 144062 120930
rect 141044 118650 141100 118659
rect 141044 118585 141100 118594
rect 141058 118363 141086 118585
rect 144034 118488 144062 120902
rect 144116 120870 144172 120879
rect 144116 120805 144172 120814
rect 143938 118460 144062 118488
rect 141044 118354 141100 118363
rect 141044 118289 141100 118298
rect 143938 118025 143966 118460
rect 144020 118354 144076 118363
rect 144020 118289 144022 118298
rect 144074 118289 144076 118298
rect 144022 118257 144074 118263
rect 144130 118173 144158 120805
rect 144022 118167 144074 118173
rect 144022 118109 144074 118115
rect 144118 118167 144170 118173
rect 144118 118109 144170 118115
rect 143926 118019 143978 118025
rect 143926 117961 143978 117967
rect 144034 114344 144062 118109
rect 144118 118019 144170 118025
rect 144118 117961 144170 117967
rect 143938 114316 144062 114344
rect 143830 113283 143882 113289
rect 143830 113225 143882 113231
rect 143638 107215 143690 107221
rect 143638 107157 143690 107163
rect 143650 103373 143678 107157
rect 143734 107141 143786 107147
rect 143734 107083 143786 107089
rect 143746 106555 143774 107083
rect 143842 107073 143870 113225
rect 143938 112272 143966 114316
rect 144020 114210 144076 114219
rect 144020 114145 144076 114154
rect 144034 112697 144062 114145
rect 144130 113289 144158 117961
rect 144118 113283 144170 113289
rect 144118 113225 144170 113231
rect 144116 113174 144172 113183
rect 144116 113109 144172 113118
rect 144022 112691 144074 112697
rect 144022 112633 144074 112639
rect 144130 112475 144158 113109
rect 144118 112469 144170 112475
rect 144020 112434 144076 112443
rect 144118 112411 144170 112417
rect 144020 112369 144022 112378
rect 144074 112369 144076 112378
rect 144022 112337 144074 112343
rect 143938 112244 144062 112272
rect 144034 109904 144062 112244
rect 144116 111250 144172 111259
rect 144116 111185 144172 111194
rect 143938 109876 144062 109904
rect 143938 109312 143966 109876
rect 144020 109770 144076 109779
rect 144020 109705 144076 109714
rect 144034 109515 144062 109705
rect 144130 109589 144158 111185
rect 144118 109583 144170 109589
rect 144118 109525 144170 109531
rect 144022 109509 144074 109515
rect 144022 109451 144074 109457
rect 144118 109435 144170 109441
rect 144118 109377 144170 109383
rect 143938 109284 144062 109312
rect 144034 107684 144062 109284
rect 143938 107656 144062 107684
rect 143830 107067 143882 107073
rect 143830 107009 143882 107015
rect 143938 106967 143966 107656
rect 144020 107550 144076 107559
rect 144020 107485 144076 107494
rect 143924 106958 143980 106967
rect 143830 106919 143882 106925
rect 143924 106893 143980 106902
rect 143830 106861 143882 106867
rect 143842 106648 143870 106861
rect 144034 106777 144062 107485
rect 144130 107221 144158 109377
rect 144118 107215 144170 107221
rect 144118 107157 144170 107163
rect 144118 107067 144170 107073
rect 144118 107009 144170 107015
rect 144022 106771 144074 106777
rect 144022 106713 144074 106719
rect 143842 106620 143966 106648
rect 143734 106549 143786 106555
rect 143734 106491 143786 106497
rect 143938 103984 143966 106620
rect 144022 106623 144074 106629
rect 144022 106565 144074 106571
rect 144034 106037 144062 106565
rect 144022 106031 144074 106037
rect 144022 105973 144074 105979
rect 144020 105922 144076 105931
rect 144020 105857 144076 105866
rect 144034 104409 144062 105857
rect 144130 104927 144158 107009
rect 144226 106185 144254 163577
rect 144308 159942 144364 159951
rect 144308 159877 144364 159886
rect 144322 139633 144350 159877
rect 144310 139627 144362 139633
rect 144310 139569 144362 139575
rect 144308 139518 144364 139527
rect 144308 139453 144364 139462
rect 144322 138449 144350 139453
rect 144310 138443 144362 138449
rect 144310 138385 144362 138391
rect 144308 134042 144364 134051
rect 144308 133977 144364 133986
rect 144322 132603 144350 133977
rect 144310 132597 144362 132603
rect 144310 132539 144362 132545
rect 144310 132449 144362 132455
rect 144310 132391 144362 132397
rect 144214 106179 144266 106185
rect 144214 106121 144266 106127
rect 144214 106031 144266 106037
rect 144214 105973 144266 105979
rect 144118 104921 144170 104927
rect 144118 104863 144170 104869
rect 144116 104738 144172 104747
rect 144116 104673 144172 104682
rect 144022 104403 144074 104409
rect 144022 104345 144074 104351
rect 144020 104294 144076 104303
rect 144020 104229 144022 104238
rect 144074 104229 144076 104238
rect 144022 104197 144074 104203
rect 143938 103956 144062 103984
rect 143638 103367 143690 103373
rect 143638 103309 143690 103315
rect 144034 101764 144062 103956
rect 144130 103743 144158 104673
rect 144118 103737 144170 103743
rect 144118 103679 144170 103685
rect 144116 102814 144172 102823
rect 144116 102749 144172 102758
rect 143938 101736 144062 101764
rect 143938 101468 143966 101736
rect 144020 101630 144076 101639
rect 144020 101565 144022 101574
rect 144074 101565 144076 101574
rect 144022 101533 144074 101539
rect 143938 101440 144062 101468
rect 144034 100709 144062 101440
rect 144130 100857 144158 102749
rect 144118 100851 144170 100857
rect 144118 100793 144170 100799
rect 144226 100783 144254 105973
rect 144214 100777 144266 100783
rect 144214 100719 144266 100725
rect 144022 100703 144074 100709
rect 144022 100645 144074 100651
rect 144212 99854 144268 99863
rect 144212 99789 144268 99798
rect 144116 99114 144172 99123
rect 144116 99049 144172 99058
rect 144022 98113 144074 98119
rect 144020 98078 144022 98087
rect 144074 98078 144076 98087
rect 144130 98045 144158 99049
rect 144020 98013 144076 98022
rect 144118 98039 144170 98045
rect 144118 97981 144170 97987
rect 144226 97971 144254 99789
rect 144214 97965 144266 97971
rect 144214 97907 144266 97913
rect 144116 96302 144172 96311
rect 144116 96237 144172 96246
rect 144020 95562 144076 95571
rect 144020 95497 144076 95506
rect 144034 95159 144062 95497
rect 144022 95153 144074 95159
rect 144022 95095 144074 95101
rect 144130 95085 144158 96237
rect 144118 95079 144170 95085
rect 144118 95021 144170 95027
rect 144116 94378 144172 94387
rect 144116 94313 144172 94322
rect 144020 92898 144076 92907
rect 144020 92833 144076 92842
rect 144034 92199 144062 92833
rect 144130 92273 144158 94313
rect 144118 92267 144170 92273
rect 144118 92209 144170 92215
rect 144022 92193 144074 92199
rect 144022 92135 144074 92141
rect 144212 91418 144268 91427
rect 144212 91353 144268 91362
rect 144116 90826 144172 90835
rect 144116 90761 144172 90770
rect 144020 89642 144076 89651
rect 144020 89577 144076 89586
rect 144034 89461 144062 89577
rect 144022 89455 144074 89461
rect 144022 89397 144074 89403
rect 144130 89387 144158 90761
rect 144118 89381 144170 89387
rect 144118 89323 144170 89329
rect 144226 89313 144254 91353
rect 144214 89307 144266 89313
rect 144214 89249 144266 89255
rect 144116 87126 144172 87135
rect 144116 87061 144172 87070
rect 144020 85942 144076 85951
rect 144020 85877 144076 85886
rect 144034 85021 144062 85877
rect 144022 85015 144074 85021
rect 144022 84957 144074 84963
rect 144020 82390 144076 82399
rect 144020 82325 144076 82334
rect 144034 82135 144062 82325
rect 144022 82129 144074 82135
rect 144022 82071 144074 82077
rect 144022 80871 144074 80877
rect 144022 80813 144074 80819
rect 144034 79712 144062 80813
rect 143842 79684 144062 79712
rect 143842 72663 143870 79684
rect 144130 79564 144158 87061
rect 144034 79536 144158 79564
rect 144034 78824 144062 79536
rect 144116 79430 144172 79439
rect 144116 79365 144172 79374
rect 143938 78796 144062 78824
rect 143938 77640 143966 78796
rect 144020 78690 144076 78699
rect 144020 78625 144076 78634
rect 144034 77843 144062 78625
rect 144130 77917 144158 79365
rect 144118 77911 144170 77917
rect 144118 77853 144170 77859
rect 144022 77837 144074 77843
rect 144022 77779 144074 77785
rect 143938 77612 144062 77640
rect 144034 75864 144062 77612
rect 144116 77506 144172 77515
rect 144116 77441 144172 77450
rect 143938 75836 144062 75864
rect 143938 75013 143966 75836
rect 144020 75730 144076 75739
rect 144020 75665 144076 75674
rect 144034 75105 144062 75665
rect 144022 75099 144074 75105
rect 144022 75041 144074 75047
rect 143938 74985 144062 75013
rect 144034 74088 144062 74985
rect 144130 74957 144158 77441
rect 144214 76431 144266 76437
rect 144214 76373 144266 76379
rect 144118 74951 144170 74957
rect 144118 74893 144170 74899
rect 144118 74285 144170 74291
rect 144118 74227 144170 74233
rect 143938 74060 144062 74088
rect 143830 72657 143882 72663
rect 143830 72599 143882 72605
rect 143938 70684 143966 74060
rect 144020 73954 144076 73963
rect 144020 73889 144076 73898
rect 144034 72071 144062 73889
rect 144130 72779 144158 74227
rect 144116 72770 144172 72779
rect 144116 72705 144172 72714
rect 144118 72657 144170 72663
rect 144118 72599 144170 72605
rect 144022 72065 144074 72071
rect 144022 72007 144074 72013
rect 144020 71290 144076 71299
rect 144020 71225 144076 71234
rect 144034 70887 144062 71225
rect 144022 70881 144074 70887
rect 144022 70823 144074 70829
rect 143938 70656 144062 70684
rect 144034 69944 144062 70656
rect 143938 69916 144062 69944
rect 143938 69056 143966 69916
rect 144020 69810 144076 69819
rect 144020 69745 144076 69754
rect 144034 69185 144062 69745
rect 144022 69179 144074 69185
rect 144022 69121 144074 69127
rect 143938 69028 144062 69056
rect 144034 67872 144062 69028
rect 143938 67844 144062 67872
rect 143938 67280 143966 67844
rect 144020 67738 144076 67747
rect 144020 67673 144076 67682
rect 144034 67409 144062 67673
rect 144022 67403 144074 67409
rect 144022 67345 144074 67351
rect 143938 67252 144062 67280
rect 144034 66743 144062 67252
rect 144022 66737 144074 66743
rect 144022 66679 144074 66685
rect 144022 66293 144074 66299
rect 144022 66235 144074 66241
rect 144034 65633 144062 66235
rect 144022 65627 144074 65633
rect 144022 65569 144074 65575
rect 144020 65518 144076 65527
rect 144020 65453 144076 65462
rect 144034 64893 144062 65453
rect 144022 64887 144074 64893
rect 144022 64829 144074 64835
rect 144020 62706 144076 62715
rect 144020 62641 144076 62650
rect 144034 62229 144062 62641
rect 144022 62223 144074 62229
rect 144022 62165 144074 62171
rect 144022 59633 144074 59639
rect 144020 59598 144022 59607
rect 144074 59598 144076 59607
rect 144020 59533 144076 59542
rect 144022 59041 144074 59047
rect 144022 58983 144074 58989
rect 144034 58719 144062 58983
rect 144020 58710 144076 58719
rect 144020 58645 144076 58654
rect 144022 57117 144074 57123
rect 144020 57082 144022 57091
rect 144074 57082 144076 57091
rect 144020 57017 144076 57026
rect 144022 56525 144074 56531
rect 144022 56467 144074 56473
rect 144034 56203 144062 56467
rect 144020 56194 144076 56203
rect 144020 56129 144076 56138
rect 144020 54714 144076 54723
rect 144020 54649 144022 54658
rect 144074 54649 144076 54658
rect 144022 54617 144074 54623
rect 144022 54157 144074 54163
rect 144022 54099 144074 54105
rect 144034 53835 144062 54099
rect 144020 53826 144076 53835
rect 144020 53761 144076 53770
rect 137494 52307 137546 52313
rect 137494 52249 137546 52255
rect 137506 51888 137534 52249
rect 137280 51860 137534 51888
rect 144130 50389 144158 72599
rect 144226 66521 144254 76373
rect 144214 66515 144266 66521
rect 144214 66457 144266 66463
rect 144212 66406 144268 66415
rect 144212 66341 144268 66350
rect 144226 66299 144254 66341
rect 144214 66293 144266 66299
rect 144214 66235 144266 66241
rect 144214 65627 144266 65633
rect 144214 65569 144266 65575
rect 144118 50383 144170 50389
rect 144118 50325 144170 50331
rect 144226 50167 144254 65569
rect 144322 50241 144350 132391
rect 144418 124685 144446 194805
rect 144502 175665 144554 175671
rect 144502 175607 144554 175613
rect 144514 155691 144542 175607
rect 144502 155685 144554 155691
rect 144502 155627 144554 155633
rect 144500 154466 144556 154475
rect 144500 154401 144556 154410
rect 144514 152731 144542 154401
rect 144502 152725 144554 152731
rect 144502 152667 144554 152673
rect 144500 151654 144556 151663
rect 144500 151589 144556 151598
rect 144514 149919 144542 151589
rect 144502 149913 144554 149919
rect 144502 149855 144554 149861
rect 144500 149730 144556 149739
rect 144500 149665 144556 149674
rect 144514 147033 144542 149665
rect 144502 147027 144554 147033
rect 144502 146969 144554 146975
rect 144502 146435 144554 146441
rect 144502 146377 144554 146383
rect 144514 139781 144542 146377
rect 144502 139775 144554 139781
rect 144502 139717 144554 139723
rect 144502 139627 144554 139633
rect 144502 139569 144554 139575
rect 144514 126905 144542 139569
rect 144502 126899 144554 126905
rect 144502 126841 144554 126847
rect 144500 126790 144556 126799
rect 144500 126725 144556 126734
rect 144406 124679 144458 124685
rect 144406 124621 144458 124627
rect 144406 124531 144458 124537
rect 144406 124473 144458 124479
rect 144418 107147 144446 124473
rect 144406 107141 144458 107147
rect 144406 107083 144458 107089
rect 144406 106993 144458 106999
rect 144406 106935 144458 106941
rect 144418 103521 144446 106935
rect 144406 103515 144458 103521
rect 144406 103457 144458 103463
rect 144406 103367 144458 103373
rect 144406 103309 144458 103315
rect 144418 92125 144446 103309
rect 144406 92119 144458 92125
rect 144406 92061 144458 92067
rect 144406 86421 144458 86427
rect 144406 86363 144458 86369
rect 144418 80877 144446 86363
rect 144406 80871 144458 80877
rect 144406 80813 144458 80819
rect 144404 80762 144460 80771
rect 144404 80697 144460 80706
rect 144418 52091 144446 80697
rect 144406 52085 144458 52091
rect 144406 52027 144458 52033
rect 144514 50463 144542 126725
rect 144610 125425 144638 196581
rect 144706 195873 144734 197765
rect 145078 197273 145130 197279
rect 145078 197215 145130 197221
rect 144694 195867 144746 195873
rect 144694 195809 144746 195815
rect 144884 179774 144940 179783
rect 144884 179709 144940 179718
rect 144692 166602 144748 166611
rect 144692 166537 144748 166546
rect 144706 164201 144734 166537
rect 144898 165607 144926 179709
rect 145090 172637 145118 197215
rect 145268 176074 145324 176083
rect 145268 176009 145324 176018
rect 145078 172631 145130 172637
rect 145078 172573 145130 172579
rect 145172 172078 145228 172087
rect 145172 172013 145228 172022
rect 144980 170154 145036 170163
rect 144980 170089 145036 170098
rect 144886 165601 144938 165607
rect 144886 165543 144938 165549
rect 144884 164826 144940 164835
rect 144884 164761 144940 164770
rect 144694 164195 144746 164201
rect 144694 164137 144746 164143
rect 144692 162902 144748 162911
rect 144692 162837 144748 162846
rect 144706 161315 144734 162837
rect 144788 161422 144844 161431
rect 144788 161357 144844 161366
rect 144694 161309 144746 161315
rect 144694 161251 144746 161257
rect 144692 159350 144748 159359
rect 144692 159285 144748 159294
rect 144706 158503 144734 159285
rect 144694 158497 144746 158503
rect 144694 158439 144746 158445
rect 144692 156390 144748 156399
rect 144692 156325 144748 156334
rect 144706 155617 144734 156325
rect 144694 155611 144746 155617
rect 144694 155553 144746 155559
rect 144694 153169 144746 153175
rect 144694 153111 144746 153117
rect 144706 146441 144734 153111
rect 144694 146435 144746 146441
rect 144694 146377 144746 146383
rect 144694 146287 144746 146293
rect 144694 146229 144746 146235
rect 144706 126683 144734 146229
rect 144694 126677 144746 126683
rect 144694 126619 144746 126625
rect 144598 125419 144650 125425
rect 144598 125361 144650 125367
rect 144598 125271 144650 125277
rect 144598 125213 144650 125219
rect 144610 109441 144638 125213
rect 144694 124679 144746 124685
rect 144694 124621 144746 124627
rect 144598 109435 144650 109441
rect 144598 109377 144650 109383
rect 144706 108424 144734 124621
rect 144610 108396 144734 108424
rect 144610 106851 144638 108396
rect 144692 108290 144748 108299
rect 144692 108225 144748 108234
rect 144598 106845 144650 106851
rect 144598 106787 144650 106793
rect 144596 106662 144652 106671
rect 144706 106629 144734 108225
rect 144596 106597 144652 106606
rect 144694 106623 144746 106629
rect 144610 105020 144638 106597
rect 144694 106565 144746 106571
rect 144610 104992 144734 105020
rect 144598 104921 144650 104927
rect 144598 104863 144650 104869
rect 144610 86427 144638 104863
rect 144706 103595 144734 104992
rect 144694 103589 144746 103595
rect 144694 103531 144746 103537
rect 144598 86421 144650 86427
rect 144598 86363 144650 86369
rect 144692 83574 144748 83583
rect 144692 83509 144748 83518
rect 144598 72509 144650 72515
rect 144598 72451 144650 72457
rect 144610 67261 144638 72451
rect 144598 67255 144650 67261
rect 144598 67197 144650 67203
rect 144706 67132 144734 83509
rect 144610 67104 144734 67132
rect 144610 52017 144638 67104
rect 144694 67033 144746 67039
rect 144694 66975 144746 66981
rect 144598 52011 144650 52017
rect 144598 51953 144650 51959
rect 144502 50457 144554 50463
rect 144502 50399 144554 50405
rect 144310 50235 144362 50241
rect 144310 50177 144362 50183
rect 144214 50161 144266 50167
rect 144214 50103 144266 50109
rect 144706 50019 144734 66975
rect 144802 51425 144830 161357
rect 144898 64912 144926 164761
rect 144994 65041 145022 170089
rect 145076 168378 145132 168387
rect 145076 168313 145132 168322
rect 144982 65035 145034 65041
rect 144982 64977 145034 64983
rect 144898 64884 145022 64912
rect 144886 64813 144938 64819
rect 144884 64778 144886 64787
rect 144938 64778 144940 64787
rect 144884 64713 144940 64722
rect 144790 51419 144842 51425
rect 144790 51361 144842 51367
rect 144994 51351 145022 64884
rect 144982 51345 145034 51351
rect 144982 51287 145034 51293
rect 145090 50759 145118 168313
rect 145078 50753 145130 50759
rect 145078 50695 145130 50701
rect 145186 50537 145214 172013
rect 145282 50611 145310 176009
rect 145378 51573 145406 214489
rect 145460 210558 145516 210567
rect 145460 210493 145516 210502
rect 145474 76437 145502 210493
rect 145556 208042 145612 208051
rect 145556 207977 145612 207986
rect 145462 76431 145514 76437
rect 145462 76373 145514 76379
rect 145570 76308 145598 207977
rect 145652 205674 145708 205683
rect 145652 205609 145708 205618
rect 145474 76280 145598 76308
rect 145474 65189 145502 76280
rect 145558 76209 145610 76215
rect 145558 76151 145610 76157
rect 145462 65183 145514 65189
rect 145462 65125 145514 65131
rect 145462 65035 145514 65041
rect 145462 64977 145514 64983
rect 145366 51567 145418 51573
rect 145366 51509 145418 51515
rect 145474 50685 145502 64977
rect 145570 50907 145598 76151
rect 145666 51277 145694 205609
rect 145748 205082 145804 205091
rect 145748 205017 145804 205026
rect 145762 201516 145790 205017
rect 145844 202122 145900 202131
rect 145844 202057 145900 202066
rect 145858 201719 145886 202057
rect 145846 201713 145898 201719
rect 145846 201655 145898 201661
rect 145762 201488 145886 201516
rect 145748 201382 145804 201391
rect 145748 201317 145804 201326
rect 145654 51271 145706 51277
rect 145654 51213 145706 51219
rect 145558 50901 145610 50907
rect 145558 50843 145610 50849
rect 145462 50679 145514 50685
rect 145462 50621 145514 50627
rect 145270 50605 145322 50611
rect 145270 50547 145322 50553
rect 145174 50531 145226 50537
rect 145174 50473 145226 50479
rect 144694 50013 144746 50019
rect 144694 49955 144746 49961
rect 145762 49723 145790 201317
rect 145858 51203 145886 201488
rect 146242 197279 146270 215992
rect 146230 197273 146282 197279
rect 146230 197215 146282 197221
rect 145940 193686 145996 193695
rect 145940 193621 145996 193630
rect 145954 51499 145982 193621
rect 146036 190134 146092 190143
rect 146036 190069 146092 190078
rect 146050 76479 146078 190069
rect 146228 189394 146284 189403
rect 146228 189329 146284 189338
rect 146132 186434 146188 186443
rect 146132 186369 146188 186378
rect 146146 175912 146174 186369
rect 146242 176041 146270 189329
rect 146338 184625 146366 216011
rect 146420 185250 146476 185259
rect 146420 185185 146476 185194
rect 146326 184619 146378 184625
rect 146326 184561 146378 184567
rect 146434 182128 146462 185185
rect 146338 182100 146462 182128
rect 146338 176060 146366 182100
rect 146530 176189 146558 235061
rect 146804 226690 146860 226699
rect 146804 226625 146860 226634
rect 146818 226435 146846 226625
rect 146806 226429 146858 226435
rect 146806 226371 146858 226377
rect 146804 222990 146860 222999
rect 146804 222925 146860 222934
rect 146710 221989 146762 221995
rect 146710 221931 146762 221937
rect 146722 221815 146750 221931
rect 146818 221921 146846 222925
rect 146806 221915 146858 221921
rect 146806 221857 146858 221863
rect 146708 221806 146764 221815
rect 146708 221741 146764 221750
rect 146804 218254 146860 218263
rect 146804 218189 146860 218198
rect 146818 216593 146846 218189
rect 146806 216587 146858 216593
rect 146806 216529 146858 216535
rect 146804 213370 146860 213379
rect 146804 213305 146860 213314
rect 146818 213263 146846 213305
rect 146806 213257 146858 213263
rect 146806 213199 146858 213205
rect 148246 210297 148298 210303
rect 148246 210239 148298 210245
rect 146612 209818 146668 209827
rect 146612 209753 146668 209762
rect 146626 207491 146654 209753
rect 146614 207485 146666 207491
rect 146614 207427 146666 207433
rect 146804 207450 146860 207459
rect 146804 207385 146806 207394
rect 146858 207385 146860 207394
rect 146806 207353 146858 207359
rect 146806 184619 146858 184625
rect 146806 184561 146858 184567
rect 146818 181980 146846 184561
rect 146818 181952 146942 181980
rect 146614 181585 146666 181591
rect 146614 181527 146666 181533
rect 146518 176183 146570 176189
rect 146518 176125 146570 176131
rect 146230 176035 146282 176041
rect 146338 176032 146558 176060
rect 146230 175977 146282 175983
rect 146146 175884 146366 175912
rect 146230 175813 146282 175819
rect 146230 175755 146282 175761
rect 146134 155833 146186 155839
rect 146134 155775 146186 155781
rect 146146 135341 146174 155775
rect 146134 135335 146186 135341
rect 146134 135277 146186 135283
rect 146132 135226 146188 135235
rect 146132 135161 146188 135170
rect 146146 126799 146174 135161
rect 146132 126790 146188 126799
rect 146132 126725 146188 126734
rect 146134 126677 146186 126683
rect 146134 126619 146186 126625
rect 146146 107073 146174 126619
rect 146134 107067 146186 107073
rect 146134 107009 146186 107015
rect 146242 106819 146270 175755
rect 146228 106810 146284 106819
rect 146228 106745 146284 106754
rect 146228 106514 146284 106523
rect 146228 106449 146284 106458
rect 146134 101443 146186 101449
rect 146134 101385 146186 101391
rect 146146 86501 146174 101385
rect 146134 86495 146186 86501
rect 146134 86437 146186 86443
rect 146036 76470 146092 76479
rect 146036 76405 146092 76414
rect 146038 76357 146090 76363
rect 146038 76299 146090 76305
rect 145942 51493 145994 51499
rect 145942 51435 145994 51441
rect 145846 51197 145898 51203
rect 145846 51139 145898 51145
rect 146050 50833 146078 76299
rect 146134 66885 146186 66891
rect 146134 66827 146186 66833
rect 146038 50827 146090 50833
rect 146038 50769 146090 50775
rect 146146 50315 146174 66827
rect 146242 51129 146270 106449
rect 146338 101449 146366 175884
rect 146422 155759 146474 155765
rect 146422 155701 146474 155707
rect 146434 125795 146462 155701
rect 146422 125789 146474 125795
rect 146422 125731 146474 125737
rect 146422 125419 146474 125425
rect 146422 125361 146474 125367
rect 146434 106925 146462 125361
rect 146422 106919 146474 106925
rect 146422 106861 146474 106867
rect 146422 106179 146474 106185
rect 146422 106121 146474 106127
rect 146326 101443 146378 101449
rect 146326 101385 146378 101391
rect 146434 94641 146462 106121
rect 146422 94635 146474 94641
rect 146422 94577 146474 94583
rect 146420 87866 146476 87875
rect 146420 87801 146476 87810
rect 146326 86495 146378 86501
rect 146326 86437 146378 86443
rect 146338 66225 146366 86437
rect 146326 66219 146378 66225
rect 146326 66161 146378 66167
rect 146434 51943 146462 87801
rect 146530 76215 146558 176032
rect 146518 76209 146570 76215
rect 146518 76151 146570 76157
rect 146516 76026 146572 76035
rect 146516 75961 146572 75970
rect 146530 72515 146558 75961
rect 146518 72509 146570 72515
rect 146518 72451 146570 72457
rect 146516 69070 146572 69079
rect 146516 69005 146572 69014
rect 146530 66373 146558 69005
rect 146518 66367 146570 66373
rect 146518 66309 146570 66315
rect 146518 65183 146570 65189
rect 146518 65125 146570 65131
rect 146422 51937 146474 51943
rect 146422 51879 146474 51885
rect 146230 51123 146282 51129
rect 146230 51065 146282 51071
rect 146134 50309 146186 50315
rect 146134 50251 146186 50257
rect 146530 50093 146558 65125
rect 146626 50981 146654 181527
rect 146914 181388 146942 181952
rect 146818 181360 146942 181388
rect 146818 178724 146846 181360
rect 146818 178696 146942 178724
rect 146914 178428 146942 178696
rect 146722 178400 146942 178428
rect 146722 172785 146750 178400
rect 146998 176183 147050 176189
rect 146998 176125 147050 176131
rect 146806 175665 146858 175671
rect 147010 175653 147038 176125
rect 146858 175625 147038 175653
rect 146806 175607 146858 175613
rect 146710 172779 146762 172785
rect 146710 172721 146762 172727
rect 146710 172631 146762 172637
rect 146710 172573 146762 172579
rect 146722 155839 146750 172573
rect 146806 165601 146858 165607
rect 146806 165543 146858 165549
rect 146710 155833 146762 155839
rect 146710 155775 146762 155781
rect 146710 155685 146762 155691
rect 146710 155627 146762 155633
rect 146722 153175 146750 155627
rect 146710 153169 146762 153175
rect 146710 153111 146762 153117
rect 146818 153120 146846 165543
rect 146902 155685 146954 155691
rect 146900 155650 146902 155659
rect 146954 155650 146956 155659
rect 146900 155585 146956 155594
rect 146818 153092 146942 153120
rect 146804 152986 146860 152995
rect 146804 152921 146860 152930
rect 146818 152805 146846 152921
rect 146806 152799 146858 152805
rect 146806 152741 146858 152747
rect 146914 152676 146942 153092
rect 146818 152648 146942 152676
rect 146818 151048 146846 152648
rect 146818 151020 146942 151048
rect 146804 150914 146860 150923
rect 146804 150849 146860 150858
rect 146818 149845 146846 150849
rect 146806 149839 146858 149845
rect 146806 149781 146858 149787
rect 146914 149728 146942 151020
rect 146818 149700 146942 149728
rect 146818 148088 146846 149700
rect 146818 148060 146942 148088
rect 146804 147954 146860 147963
rect 146804 147889 146860 147898
rect 146818 146959 146846 147889
rect 146806 146953 146858 146959
rect 146806 146895 146858 146901
rect 146708 144254 146764 144263
rect 146708 144189 146764 144198
rect 146722 135679 146750 144189
rect 146708 135670 146764 135679
rect 146708 135605 146764 135614
rect 146914 135415 146942 148060
rect 146996 136114 147052 136123
rect 146996 136049 146998 136058
rect 147050 136049 147052 136058
rect 146998 136017 147050 136023
rect 146710 135409 146762 135415
rect 146710 135351 146762 135357
rect 146902 135409 146954 135415
rect 146902 135351 146954 135357
rect 146722 131068 146750 135351
rect 146998 135261 147050 135267
rect 146998 135203 147050 135209
rect 146722 131040 146846 131068
rect 146708 127530 146764 127539
rect 146708 127465 146764 127474
rect 146722 126757 146750 127465
rect 146710 126751 146762 126757
rect 146710 126693 146762 126699
rect 146710 125789 146762 125795
rect 146710 125731 146762 125737
rect 146722 118247 146750 125731
rect 146818 118340 146846 131040
rect 146900 119094 146956 119103
rect 146900 119029 146902 119038
rect 146954 119029 146956 119038
rect 146902 118997 146954 119003
rect 146818 118312 146942 118340
rect 146710 118241 146762 118247
rect 146710 118183 146762 118189
rect 146914 117896 146942 118312
rect 146818 117868 146942 117896
rect 146710 106549 146762 106555
rect 146710 106491 146762 106497
rect 146722 94937 146750 106491
rect 146710 94931 146762 94937
rect 146710 94873 146762 94879
rect 146708 84166 146764 84175
rect 146708 84101 146764 84110
rect 146722 66891 146750 84101
rect 146818 76363 146846 117868
rect 146900 116726 146956 116735
rect 146900 116661 146902 116670
rect 146954 116661 146956 116670
rect 146902 116629 146954 116635
rect 146900 115986 146956 115995
rect 146900 115921 146902 115930
rect 146954 115921 146956 115930
rect 146902 115889 146954 115895
rect 147010 103669 147038 135203
rect 147092 126938 147148 126947
rect 147092 126873 147094 126882
rect 147146 126873 147148 126882
rect 147094 126841 147146 126847
rect 148054 116687 148106 116693
rect 148054 116629 148106 116635
rect 147958 112469 148010 112475
rect 147958 112411 148010 112417
rect 147862 112395 147914 112401
rect 147862 112337 147914 112343
rect 147766 109583 147818 109589
rect 147766 109525 147818 109531
rect 146998 103663 147050 103669
rect 146998 103605 147050 103611
rect 147670 100851 147722 100857
rect 147670 100793 147722 100799
rect 146806 76357 146858 76363
rect 146806 76299 146858 76305
rect 146900 75138 146956 75147
rect 146900 75073 146956 75082
rect 146914 75031 146942 75073
rect 146902 75025 146954 75031
rect 146902 74967 146954 74973
rect 146710 66885 146762 66891
rect 146710 66827 146762 66833
rect 146710 66737 146762 66743
rect 146710 66679 146762 66685
rect 146722 52165 146750 66679
rect 146806 66219 146858 66225
rect 146806 66161 146858 66167
rect 146710 52159 146762 52165
rect 146710 52101 146762 52107
rect 146818 51055 146846 66161
rect 146902 63407 146954 63413
rect 146902 63349 146954 63355
rect 146914 62419 146942 63349
rect 146900 62410 146956 62419
rect 146900 62345 146956 62354
rect 146900 60782 146956 60791
rect 146900 60717 146956 60726
rect 146914 60453 146942 60717
rect 146902 60447 146954 60453
rect 146902 60389 146954 60395
rect 146806 51049 146858 51055
rect 146806 50991 146858 50997
rect 146614 50975 146666 50981
rect 146614 50917 146666 50923
rect 146518 50087 146570 50093
rect 146518 50029 146570 50035
rect 145750 49717 145802 49723
rect 145750 49659 145802 49665
rect 147682 47725 147710 100793
rect 147670 47719 147722 47725
rect 147670 47661 147722 47667
rect 147778 47651 147806 109525
rect 147766 47645 147818 47651
rect 147766 47587 147818 47593
rect 147874 47503 147902 112337
rect 147970 47577 147998 112411
rect 148066 48095 148094 116629
rect 148150 115947 148202 115953
rect 148150 115889 148202 115895
rect 148054 48089 148106 48095
rect 148054 48031 148106 48037
rect 148162 48021 148190 115889
rect 148258 48687 148286 210239
rect 148354 74291 148382 237545
rect 149698 224511 149726 273139
rect 150274 272093 150302 277870
rect 151126 273419 151178 273425
rect 151126 273361 151178 273367
rect 151138 272685 151166 273361
rect 151426 273203 151454 277870
rect 152674 273203 152702 277870
rect 153826 273573 153854 277870
rect 155088 277856 155486 277884
rect 153814 273567 153866 273573
rect 153814 273509 153866 273515
rect 151414 273197 151466 273203
rect 151414 273139 151466 273145
rect 152566 273197 152618 273203
rect 152566 273139 152618 273145
rect 152662 273197 152714 273203
rect 152662 273139 152714 273145
rect 155350 273197 155402 273203
rect 155350 273139 155402 273145
rect 151126 272679 151178 272685
rect 151126 272621 151178 272627
rect 150262 272087 150314 272093
rect 150262 272029 150314 272035
rect 152470 239231 152522 239237
rect 152470 239173 152522 239179
rect 152482 237799 152510 239173
rect 152468 237790 152524 237799
rect 152468 237725 152524 237734
rect 151126 230573 151178 230579
rect 151126 230515 151178 230521
rect 149686 224505 149738 224511
rect 149686 224447 149738 224453
rect 148438 190169 148490 190175
rect 148438 190111 148490 190117
rect 148342 74285 148394 74291
rect 148342 74227 148394 74233
rect 148342 60521 148394 60527
rect 148342 60463 148394 60469
rect 148354 54163 148382 60463
rect 148342 54157 148394 54163
rect 148342 54099 148394 54105
rect 148246 48681 148298 48687
rect 148246 48623 148298 48629
rect 148150 48015 148202 48021
rect 148150 47957 148202 47963
rect 147958 47571 148010 47577
rect 147958 47513 148010 47519
rect 147862 47497 147914 47503
rect 147862 47439 147914 47445
rect 133618 46708 133646 46990
rect 148450 46837 148478 190111
rect 148534 178699 148586 178705
rect 148534 178641 148586 178647
rect 148546 47059 148574 178641
rect 148630 172927 148682 172933
rect 148630 172869 148682 172875
rect 148534 47053 148586 47059
rect 148534 46995 148586 47001
rect 148438 46831 148490 46837
rect 148438 46773 148490 46779
rect 133618 46680 133694 46708
rect 133666 42841 133694 46680
rect 148642 46467 148670 172869
rect 148726 164195 148778 164201
rect 148726 164137 148778 164143
rect 148738 46911 148766 164137
rect 148822 161309 148874 161315
rect 148822 161251 148874 161257
rect 148834 48613 148862 161251
rect 148918 158497 148970 158503
rect 148918 158439 148970 158445
rect 148822 48607 148874 48613
rect 148822 48549 148874 48555
rect 148930 47207 148958 158439
rect 149014 155685 149066 155691
rect 149014 155627 149066 155633
rect 148918 47201 148970 47207
rect 148918 47143 148970 47149
rect 148726 46905 148778 46911
rect 148726 46847 148778 46853
rect 149026 46689 149054 155627
rect 149110 149913 149162 149919
rect 149110 149855 149162 149861
rect 149014 46683 149066 46689
rect 149014 46625 149066 46631
rect 149122 46541 149150 149855
rect 149206 147027 149258 147033
rect 149206 146969 149258 146975
rect 149218 46763 149246 146969
rect 149302 142587 149354 142593
rect 149302 142529 149354 142535
rect 149314 48243 149342 142529
rect 149398 136075 149450 136081
rect 149398 136017 149450 136023
rect 149302 48237 149354 48243
rect 149302 48179 149354 48185
rect 149410 48169 149438 136017
rect 149494 126899 149546 126905
rect 149494 126841 149546 126847
rect 149398 48163 149450 48169
rect 149398 48105 149450 48111
rect 149506 47947 149534 126841
rect 149590 121571 149642 121577
rect 149590 121513 149642 121519
rect 149494 47941 149546 47947
rect 149494 47883 149546 47889
rect 149602 47873 149630 121513
rect 149686 121053 149738 121059
rect 149686 120995 149738 121001
rect 149590 47867 149642 47873
rect 149590 47809 149642 47815
rect 149698 47799 149726 120995
rect 151138 100635 151166 230515
rect 152578 224437 152606 273139
rect 155362 245495 155390 273139
rect 155348 245486 155404 245495
rect 155348 245421 155404 245430
rect 152566 224431 152618 224437
rect 152566 224373 152618 224379
rect 155458 221773 155486 277856
rect 156226 273203 156254 277870
rect 157474 273351 157502 277870
rect 157462 273345 157514 273351
rect 157462 273287 157514 273293
rect 158626 273277 158654 277870
rect 158614 273271 158666 273277
rect 158614 273213 158666 273219
rect 159874 273203 159902 277870
rect 161026 273425 161054 277870
rect 161014 273419 161066 273425
rect 161014 273361 161066 273367
rect 161206 273271 161258 273277
rect 161206 273213 161258 273219
rect 156214 273197 156266 273203
rect 156214 273139 156266 273145
rect 158326 273197 158378 273203
rect 158326 273139 158378 273145
rect 159862 273197 159914 273203
rect 159862 273139 159914 273145
rect 161110 273197 161162 273203
rect 161110 273139 161162 273145
rect 156886 271643 156938 271649
rect 156886 271585 156938 271591
rect 156898 271427 156926 271585
rect 156886 271421 156938 271427
rect 156886 271363 156938 271369
rect 155542 246039 155594 246045
rect 155542 245981 155594 245987
rect 155554 245823 155582 245981
rect 155542 245817 155594 245823
rect 155542 245759 155594 245765
rect 158338 245199 158366 273139
rect 160918 246335 160970 246341
rect 160918 246277 160970 246283
rect 160930 245897 160958 246277
rect 161014 246261 161066 246267
rect 161014 246203 161066 246209
rect 161026 245971 161054 246203
rect 161014 245965 161066 245971
rect 161014 245907 161066 245913
rect 160918 245891 160970 245897
rect 160918 245833 160970 245839
rect 158324 245190 158380 245199
rect 158324 245125 158380 245134
rect 161122 245051 161150 273139
rect 161108 245042 161164 245051
rect 161108 244977 161164 244986
rect 156886 226429 156938 226435
rect 156886 226371 156938 226377
rect 155446 221767 155498 221773
rect 155446 221709 155498 221715
rect 154006 216587 154058 216593
rect 154006 216529 154058 216535
rect 151222 190243 151274 190249
rect 151222 190185 151274 190191
rect 151126 100629 151178 100635
rect 151126 100571 151178 100577
rect 151234 94863 151262 190185
rect 151510 129711 151562 129717
rect 151510 129653 151562 129659
rect 151318 119055 151370 119061
rect 151318 118997 151370 119003
rect 151222 94857 151274 94863
rect 151222 94799 151274 94805
rect 151126 89455 151178 89461
rect 151126 89397 151178 89403
rect 151138 71997 151166 89397
rect 151126 71991 151178 71997
rect 151126 71933 151178 71939
rect 149782 70881 149834 70887
rect 149782 70823 149834 70829
rect 149794 69037 149822 70823
rect 149782 69031 149834 69037
rect 149782 68973 149834 68979
rect 149782 62223 149834 62229
rect 149782 62165 149834 62171
rect 149794 60379 149822 62165
rect 151126 60595 151178 60601
rect 151126 60537 151178 60543
rect 149782 60373 149834 60379
rect 149782 60315 149834 60321
rect 151138 54681 151166 60537
rect 151126 54675 151178 54681
rect 151126 54617 151178 54623
rect 151330 52239 151358 118997
rect 151414 104403 151466 104409
rect 151414 104345 151466 104351
rect 151426 52757 151454 104345
rect 151522 83541 151550 129653
rect 154018 97897 154046 216529
rect 154102 144067 154154 144073
rect 154102 144009 154154 144015
rect 154006 97891 154058 97897
rect 154006 97833 154058 97839
rect 154006 92267 154058 92273
rect 154006 92209 154058 92215
rect 151510 83535 151562 83541
rect 151510 83477 151562 83483
rect 154018 74883 154046 92209
rect 154114 86427 154142 144009
rect 156898 97823 156926 226371
rect 161218 221699 161246 273213
rect 162178 273203 162206 277870
rect 163440 277856 164030 277884
rect 163126 273567 163178 273573
rect 163126 273509 163178 273515
rect 163138 273277 163166 273509
rect 163126 273271 163178 273277
rect 163126 273213 163178 273219
rect 162166 273197 162218 273203
rect 162166 273139 162218 273145
rect 164002 247715 164030 277856
rect 164086 273197 164138 273203
rect 164086 273139 164138 273145
rect 164182 273197 164234 273203
rect 164182 273139 164234 273145
rect 163988 247706 164044 247715
rect 163988 247641 164044 247650
rect 161302 246409 161354 246415
rect 161302 246351 161354 246357
rect 161314 246119 161342 246351
rect 163702 246261 163754 246267
rect 163702 246203 163754 246209
rect 161302 246113 161354 246119
rect 161302 246055 161354 246061
rect 161494 246113 161546 246119
rect 161494 246055 161546 246061
rect 161506 245823 161534 246055
rect 163714 245971 163742 246203
rect 163702 245965 163754 245971
rect 163702 245907 163754 245913
rect 161494 245817 161546 245823
rect 161494 245759 161546 245765
rect 161206 221693 161258 221699
rect 161206 221635 161258 221641
rect 164098 221625 164126 273139
rect 164194 272093 164222 273139
rect 164578 272093 164606 277870
rect 165826 273573 165854 277870
rect 165814 273567 165866 273573
rect 165814 273509 165866 273515
rect 164182 272087 164234 272093
rect 164182 272029 164234 272035
rect 164566 272087 164618 272093
rect 164566 272029 164618 272035
rect 166882 246975 166910 277870
rect 166966 273567 167018 273573
rect 166966 273509 167018 273515
rect 166868 246966 166924 246975
rect 166868 246901 166924 246910
rect 165526 246335 165578 246341
rect 165526 246277 165578 246283
rect 165538 245897 165566 246277
rect 165526 245891 165578 245897
rect 165526 245833 165578 245839
rect 165526 230499 165578 230505
rect 165526 230441 165578 230447
rect 164086 221619 164138 221625
rect 164086 221561 164138 221567
rect 162646 201713 162698 201719
rect 162646 201655 162698 201661
rect 159766 198975 159818 198981
rect 159766 198917 159818 198923
rect 156982 167303 157034 167309
rect 156982 167245 157034 167251
rect 156886 97817 156938 97823
rect 156886 97759 156938 97765
rect 156994 89239 157022 167245
rect 157078 101591 157130 101597
rect 157078 101533 157130 101539
rect 156982 89233 157034 89239
rect 156982 89175 157034 89181
rect 154102 86421 154154 86427
rect 154102 86363 154154 86369
rect 157090 77769 157118 101533
rect 159778 100561 159806 198917
rect 159862 170263 159914 170269
rect 159862 170205 159914 170211
rect 159766 100555 159818 100561
rect 159766 100497 159818 100503
rect 159874 89165 159902 170205
rect 161108 137594 161164 137603
rect 161108 137529 161164 137538
rect 161122 135508 161150 137529
rect 161206 135631 161258 135637
rect 161206 135573 161258 135579
rect 161218 135508 161246 135573
rect 161122 135480 161246 135508
rect 159958 104255 160010 104261
rect 159958 104197 160010 104203
rect 159862 89159 159914 89165
rect 159862 89101 159914 89107
rect 157078 77763 157130 77769
rect 157078 77705 157130 77711
rect 159970 77695 159998 104197
rect 162658 100487 162686 201655
rect 162742 172853 162794 172859
rect 162742 172795 162794 172801
rect 162646 100481 162698 100487
rect 162646 100423 162698 100429
rect 162754 89091 162782 172795
rect 162838 106771 162890 106777
rect 162838 106713 162890 106719
rect 162742 89085 162794 89091
rect 162742 89027 162794 89033
rect 159958 77689 160010 77695
rect 159958 77631 160010 77637
rect 162850 77621 162878 106713
rect 162838 77615 162890 77621
rect 162838 77557 162890 77563
rect 160534 75099 160586 75105
rect 160534 75041 160586 75047
rect 156886 75025 156938 75031
rect 156886 74967 156938 74973
rect 154006 74877 154058 74883
rect 154006 74819 154058 74825
rect 154582 72065 154634 72071
rect 154582 72007 154634 72013
rect 154594 68963 154622 72007
rect 154582 68957 154634 68963
rect 154582 68899 154634 68905
rect 156898 68889 156926 74967
rect 156886 68883 156938 68889
rect 156886 68825 156938 68831
rect 160546 68815 160574 75041
rect 161590 74951 161642 74957
rect 161590 74893 161642 74899
rect 161602 71923 161630 74893
rect 161590 71917 161642 71923
rect 161590 71859 161642 71865
rect 160534 68809 160586 68815
rect 160534 68751 160586 68757
rect 152662 67403 152714 67409
rect 152662 67345 152714 67351
rect 152674 66151 152702 67345
rect 157654 66367 157706 66373
rect 157654 66309 157706 66315
rect 152662 66145 152714 66151
rect 152662 66087 152714 66093
rect 157666 66077 157694 66309
rect 157654 66071 157706 66077
rect 157654 66013 157706 66019
rect 160534 60817 160586 60823
rect 160534 60759 160586 60765
rect 156310 60743 156362 60749
rect 156310 60685 156362 60691
rect 152662 60669 152714 60675
rect 152662 60611 152714 60617
rect 152674 56531 152702 60611
rect 156322 57123 156350 60685
rect 160546 59639 160574 60759
rect 160534 59633 160586 59639
rect 160534 59575 160586 59581
rect 156310 57117 156362 57123
rect 156310 57059 156362 57065
rect 152662 56525 152714 56531
rect 152662 56467 152714 56473
rect 151414 52751 151466 52757
rect 151414 52693 151466 52699
rect 151318 52233 151370 52239
rect 151318 52175 151370 52181
rect 165538 48211 165566 230441
rect 166978 221551 167006 273509
rect 168130 270909 168158 277870
rect 169296 277856 169886 277884
rect 168118 270903 168170 270909
rect 168118 270845 168170 270851
rect 168406 236271 168458 236277
rect 168406 236213 168458 236219
rect 166966 221545 167018 221551
rect 166966 221487 167018 221493
rect 165622 207485 165674 207491
rect 165622 207427 165674 207433
rect 165634 94789 165662 207427
rect 166978 135637 167102 135656
rect 166966 135631 167114 135637
rect 167018 135628 167062 135631
rect 166966 135573 167018 135579
rect 167062 135573 167114 135579
rect 165718 132967 165770 132973
rect 165718 132909 165770 132915
rect 165622 94783 165674 94789
rect 165622 94725 165674 94731
rect 165622 89381 165674 89387
rect 165622 89323 165674 89329
rect 165634 71849 165662 89323
rect 165730 83467 165758 132909
rect 167158 118389 167210 118395
rect 166978 118337 167158 118340
rect 166978 118331 167210 118337
rect 166978 118321 167198 118331
rect 166966 118315 167198 118321
rect 167018 118312 167198 118315
rect 166966 118257 167018 118263
rect 165718 83461 165770 83467
rect 165718 83403 165770 83409
rect 165622 71843 165674 71849
rect 165622 71785 165674 71791
rect 168418 48803 168446 236213
rect 169858 221477 169886 277856
rect 170530 273573 170558 277870
rect 170518 273567 170570 273573
rect 170518 273509 170570 273515
rect 171682 271797 171710 277870
rect 172726 273567 172778 273573
rect 172726 273509 172778 273515
rect 171670 271791 171722 271797
rect 171670 271733 171722 271739
rect 171286 246853 171338 246859
rect 171286 246795 171338 246801
rect 171298 246711 171326 246795
rect 171286 246705 171338 246711
rect 172738 246679 172766 273509
rect 172930 271945 172958 277870
rect 174082 273573 174110 277870
rect 174070 273567 174122 273573
rect 174070 273509 174122 273515
rect 172918 271939 172970 271945
rect 172918 271881 172970 271887
rect 175330 271723 175358 277870
rect 175510 273567 175562 273573
rect 175510 273509 175562 273515
rect 175318 271717 175370 271723
rect 175318 271659 175370 271665
rect 175522 247567 175550 273509
rect 176482 271945 176510 277870
rect 177634 273573 177662 277870
rect 177622 273567 177674 273573
rect 177622 273509 177674 273515
rect 178390 273567 178442 273573
rect 178390 273509 178442 273515
rect 175606 271939 175658 271945
rect 175606 271881 175658 271887
rect 176470 271939 176522 271945
rect 176470 271881 176522 271887
rect 175508 247558 175564 247567
rect 175508 247493 175564 247502
rect 171286 246647 171338 246653
rect 172724 246670 172780 246679
rect 172724 246605 172780 246614
rect 171380 242674 171436 242683
rect 171380 242609 171436 242618
rect 171394 242493 171422 242609
rect 171382 242487 171434 242493
rect 171382 242429 171434 242435
rect 174166 236197 174218 236203
rect 174166 236139 174218 236145
rect 171286 233311 171338 233317
rect 171286 233253 171338 233259
rect 169846 221471 169898 221477
rect 169846 221413 169898 221419
rect 168502 213257 168554 213263
rect 168502 213199 168554 213205
rect 168514 94715 168542 213199
rect 168598 138443 168650 138449
rect 168598 138385 168650 138391
rect 168502 94709 168554 94715
rect 168502 94651 168554 94657
rect 168502 89307 168554 89313
rect 168502 89249 168554 89255
rect 168514 71775 168542 89249
rect 168610 83393 168638 138385
rect 168598 83387 168650 83393
rect 168598 83329 168650 83335
rect 168502 71769 168554 71775
rect 168502 71711 168554 71717
rect 168404 48794 168460 48803
rect 168404 48729 168460 48738
rect 171298 48655 171326 233253
rect 171382 213183 171434 213189
rect 171382 213125 171434 213131
rect 171394 97749 171422 213125
rect 171478 141181 171530 141187
rect 171478 141123 171530 141129
rect 171382 97743 171434 97749
rect 171382 97685 171434 97691
rect 171382 92193 171434 92199
rect 171382 92135 171434 92141
rect 171394 71701 171422 92135
rect 171490 83319 171518 141123
rect 171478 83313 171530 83319
rect 171478 83255 171530 83261
rect 171382 71695 171434 71701
rect 171382 71637 171434 71643
rect 171284 48646 171340 48655
rect 171284 48581 171340 48590
rect 174178 48507 174206 236139
rect 174262 218955 174314 218961
rect 174262 218897 174314 218903
rect 174274 97675 174302 218897
rect 175618 218887 175646 271881
rect 177046 271495 177098 271501
rect 177046 271437 177098 271443
rect 177058 270835 177086 271437
rect 177046 270829 177098 270835
rect 177046 270771 177098 270777
rect 178402 243571 178430 273509
rect 178486 271939 178538 271945
rect 178486 271881 178538 271887
rect 178388 243562 178444 243571
rect 178388 243497 178444 243506
rect 175702 242413 175754 242419
rect 175700 242378 175702 242387
rect 175754 242378 175756 242387
rect 175700 242313 175756 242322
rect 177046 221989 177098 221995
rect 177046 221931 177098 221937
rect 175606 218881 175658 218887
rect 175606 218823 175658 218829
rect 174358 146953 174410 146959
rect 174358 146895 174410 146901
rect 174262 97669 174314 97675
rect 174262 97611 174314 97617
rect 174370 86353 174398 146895
rect 174454 95153 174506 95159
rect 174454 95095 174506 95101
rect 174358 86347 174410 86353
rect 174358 86289 174410 86295
rect 174466 74809 174494 95095
rect 174454 74803 174506 74809
rect 174454 74745 174506 74751
rect 174164 48498 174220 48507
rect 174164 48433 174220 48442
rect 165524 48202 165580 48211
rect 165524 48137 165580 48146
rect 149686 47793 149738 47799
rect 149686 47735 149738 47741
rect 177058 47429 177086 221931
rect 178498 218813 178526 271881
rect 178882 271649 178910 277870
rect 180034 273573 180062 277870
rect 180022 273567 180074 273573
rect 180022 273509 180074 273515
rect 178870 271643 178922 271649
rect 178870 271585 178922 271591
rect 181282 247419 181310 277870
rect 181366 273567 181418 273573
rect 181366 273509 181418 273515
rect 181268 247410 181324 247419
rect 181268 247345 181324 247354
rect 181378 247123 181406 273509
rect 182434 271723 182462 277870
rect 183600 277856 184286 277884
rect 184342 277875 184394 277881
rect 182422 271717 182474 271723
rect 182422 271659 182474 271665
rect 181364 247114 181420 247123
rect 181364 247049 181420 247058
rect 181366 246853 181418 246859
rect 181366 246795 181418 246801
rect 181378 246711 181406 246795
rect 181366 246705 181418 246711
rect 181366 246647 181418 246653
rect 180982 246631 181034 246637
rect 180982 246573 181034 246579
rect 181270 246631 181322 246637
rect 181270 246573 181322 246579
rect 180994 246508 181022 246573
rect 181282 246508 181310 246573
rect 180994 246480 181310 246508
rect 181364 245930 181420 245939
rect 181364 245865 181420 245874
rect 179926 221915 179978 221921
rect 179926 221857 179978 221863
rect 178486 218807 178538 218813
rect 178486 218749 178538 218755
rect 177142 149839 177194 149845
rect 177142 149781 177194 149787
rect 177154 86279 177182 149781
rect 177238 95079 177290 95085
rect 177238 95021 177290 95027
rect 177142 86273 177194 86279
rect 177142 86215 177194 86221
rect 177250 74735 177278 95021
rect 177238 74729 177290 74735
rect 177238 74671 177290 74677
rect 177046 47423 177098 47429
rect 177046 47365 177098 47371
rect 179938 47355 179966 221857
rect 181378 218739 181406 245865
rect 182806 242043 182858 242049
rect 182806 241985 182858 241991
rect 181366 218733 181418 218739
rect 181366 218675 181418 218681
rect 180022 152799 180074 152805
rect 180022 152741 180074 152747
rect 180034 86205 180062 152741
rect 181462 118537 181514 118543
rect 181462 118479 181514 118485
rect 181474 118395 181502 118479
rect 181462 118389 181514 118395
rect 181462 118331 181514 118337
rect 180118 98113 180170 98119
rect 180118 98055 180170 98061
rect 180022 86199 180074 86205
rect 180022 86141 180074 86147
rect 180130 74661 180158 98055
rect 180118 74655 180170 74661
rect 180118 74597 180170 74603
rect 182818 48359 182846 241985
rect 182902 221841 182954 221847
rect 182902 221783 182954 221789
rect 182914 97601 182942 221783
rect 184258 218665 184286 277856
rect 184354 274239 184382 277875
rect 184342 274233 184394 274239
rect 184342 274175 184394 274181
rect 184738 273573 184766 277870
rect 184726 273567 184778 273573
rect 184726 273509 184778 273515
rect 185986 271649 186014 277870
rect 187030 273567 187082 273573
rect 187030 273509 187082 273515
rect 185974 271643 186026 271649
rect 185974 271585 186026 271591
rect 187042 247271 187070 273509
rect 187028 247262 187084 247271
rect 187028 247197 187084 247206
rect 184246 218659 184298 218665
rect 184246 218601 184298 218607
rect 187138 216001 187166 277870
rect 188386 270761 188414 277870
rect 189538 271575 189566 277870
rect 189526 271569 189578 271575
rect 189526 271511 189578 271517
rect 190786 270761 190814 277870
rect 191446 271051 191498 271057
rect 191446 270993 191498 270999
rect 188374 270755 188426 270761
rect 188374 270697 188426 270703
rect 190006 270755 190058 270761
rect 190006 270697 190058 270703
rect 190774 270755 190826 270761
rect 190774 270697 190826 270703
rect 187220 247706 187276 247715
rect 187220 247641 187276 247650
rect 187234 247123 187262 247641
rect 187220 247114 187276 247123
rect 187220 247049 187276 247058
rect 190018 245939 190046 270697
rect 190004 245930 190060 245939
rect 190004 245865 190060 245874
rect 191458 238835 191486 270993
rect 191938 270983 191966 277870
rect 193090 271057 193118 277870
rect 193078 271051 193130 271057
rect 193078 270993 193130 270999
rect 191926 270977 191978 270983
rect 191926 270919 191978 270925
rect 192886 270755 192938 270761
rect 192886 270697 192938 270703
rect 191444 238826 191500 238835
rect 191444 238761 191500 238770
rect 188566 227761 188618 227767
rect 188566 227703 188618 227709
rect 187126 215995 187178 216001
rect 187126 215937 187178 215943
rect 185686 195867 185738 195873
rect 185686 195809 185738 195815
rect 182998 152725 183050 152731
rect 182998 152667 183050 152673
rect 182902 97595 182954 97601
rect 182902 97537 182954 97543
rect 183010 86131 183038 152667
rect 183094 98039 183146 98045
rect 183094 97981 183146 97987
rect 182998 86125 183050 86131
rect 182998 86067 183050 86073
rect 183106 74587 183134 97981
rect 183094 74581 183146 74587
rect 183094 74523 183146 74529
rect 185698 48539 185726 195809
rect 185782 175739 185834 175745
rect 185782 175681 185834 175687
rect 185794 89017 185822 175681
rect 185878 109509 185930 109515
rect 185878 109451 185930 109457
rect 185782 89011 185834 89017
rect 185782 88953 185834 88959
rect 185890 77547 185918 109451
rect 187222 77911 187274 77917
rect 187222 77853 187274 77859
rect 185878 77541 185930 77547
rect 185878 77483 185930 77489
rect 187234 77473 187262 77853
rect 187222 77467 187274 77473
rect 187222 77409 187274 77415
rect 185686 48533 185738 48539
rect 185686 48475 185738 48481
rect 182804 48350 182860 48359
rect 182804 48285 182860 48294
rect 179926 47349 179978 47355
rect 179926 47291 179978 47297
rect 188578 47133 188606 227703
rect 192898 215927 192926 270697
rect 194338 270021 194366 277870
rect 195490 270835 195518 277870
rect 196738 275497 196766 277870
rect 197890 276607 197918 277870
rect 197878 276601 197930 276607
rect 197878 276543 197930 276549
rect 196726 275491 196778 275497
rect 196726 275433 196778 275439
rect 198646 273567 198698 273573
rect 198646 273509 198698 273515
rect 198658 272907 198686 273509
rect 198646 272901 198698 272907
rect 198646 272843 198698 272849
rect 198742 272901 198794 272907
rect 198742 272843 198794 272849
rect 198754 272019 198782 272843
rect 198742 272013 198794 272019
rect 198742 271955 198794 271961
rect 198838 272013 198890 272019
rect 198838 271955 198890 271961
rect 195766 271495 195818 271501
rect 195766 271437 195818 271443
rect 195478 270829 195530 270835
rect 195478 270771 195530 270777
rect 195778 270761 195806 271437
rect 198850 271427 198878 271955
rect 198838 271421 198890 271427
rect 198838 271363 198890 271369
rect 199138 271279 199166 277870
rect 200194 275275 200222 277870
rect 200182 275269 200234 275275
rect 200182 275211 200234 275217
rect 200086 274233 200138 274239
rect 200086 274175 200138 274181
rect 199126 271273 199178 271279
rect 199126 271215 199178 271221
rect 195766 270755 195818 270761
rect 195766 270697 195818 270703
rect 194326 270015 194378 270021
rect 194326 269957 194378 269963
rect 200098 247747 200126 274175
rect 201442 265063 201470 277870
rect 202594 271131 202622 277870
rect 201526 271125 201578 271131
rect 201526 271067 201578 271073
rect 202582 271125 202634 271131
rect 202582 271067 202634 271073
rect 201538 270655 201566 271067
rect 201524 270646 201580 270655
rect 201524 270581 201580 270590
rect 203842 270539 203870 277870
rect 203830 270533 203882 270539
rect 203830 270475 203882 270481
rect 204994 267801 205022 277870
rect 206036 277010 206092 277019
rect 206036 276945 206092 276954
rect 206050 273499 206078 276945
rect 206038 273493 206090 273499
rect 206038 273435 206090 273441
rect 206242 270761 206270 277870
rect 207394 274239 207422 277870
rect 208546 276681 208574 277870
rect 208534 276675 208586 276681
rect 208534 276617 208586 276623
rect 207382 274233 207434 274239
rect 207382 274175 207434 274181
rect 209794 271501 209822 277870
rect 206614 271495 206666 271501
rect 206614 271437 206666 271443
rect 209782 271495 209834 271501
rect 209782 271437 209834 271443
rect 206230 270755 206282 270761
rect 206230 270697 206282 270703
rect 204982 267795 205034 267801
rect 204982 267737 205034 267743
rect 201430 265057 201482 265063
rect 201430 264999 201482 265005
rect 205558 249295 205610 249301
rect 205558 249237 205610 249243
rect 200086 247741 200138 247747
rect 196916 247706 196972 247715
rect 200086 247683 200138 247689
rect 196916 247641 196972 247650
rect 205270 247667 205322 247673
rect 196930 247419 196958 247641
rect 205270 247609 205322 247615
rect 197396 247558 197452 247567
rect 197026 247516 197396 247544
rect 196916 247410 196972 247419
rect 196916 247345 196972 247354
rect 196916 247262 196972 247271
rect 196916 247197 196972 247206
rect 196930 246383 196958 247197
rect 197026 247123 197054 247516
rect 197396 247493 197452 247502
rect 197012 247114 197068 247123
rect 197012 247049 197068 247058
rect 204598 246779 204650 246785
rect 204598 246721 204650 246727
rect 204502 246557 204554 246563
rect 197300 246522 197356 246531
rect 204502 246499 204554 246505
rect 197300 246457 197356 246466
rect 196724 246374 196780 246383
rect 196724 246309 196780 246318
rect 196916 246374 196972 246383
rect 196916 246309 196972 246318
rect 196738 244903 196766 246309
rect 197204 246226 197260 246235
rect 197204 246161 197260 246170
rect 197218 245643 197246 246161
rect 197204 245634 197260 245643
rect 197204 245569 197260 245578
rect 197314 245347 197342 246457
rect 197588 246374 197644 246383
rect 197588 246309 197644 246318
rect 199606 246335 199658 246341
rect 197602 245939 197630 246309
rect 199606 246277 199658 246283
rect 198742 246261 198794 246267
rect 198794 246209 198878 246212
rect 198742 246203 198878 246209
rect 198754 246184 198878 246203
rect 197588 245930 197644 245939
rect 197588 245865 197644 245874
rect 198850 245453 198878 246184
rect 198838 245447 198890 245453
rect 198838 245389 198890 245395
rect 197300 245338 197356 245347
rect 197300 245273 197356 245282
rect 196724 244894 196780 244903
rect 196724 244829 196780 244838
rect 199618 243307 199646 246277
rect 199606 243301 199658 243307
rect 199606 243243 199658 243249
rect 195764 242526 195820 242535
rect 195764 242461 195820 242470
rect 195778 242419 195806 242461
rect 195766 242413 195818 242419
rect 195766 242355 195818 242361
rect 204514 231583 204542 246499
rect 204610 232619 204638 246721
rect 204790 246631 204842 246637
rect 204790 246573 204842 246579
rect 204694 246483 204746 246489
rect 204694 246425 204746 246431
rect 204596 232610 204652 232619
rect 204596 232545 204652 232554
rect 204706 232175 204734 246425
rect 204692 232166 204748 232175
rect 204692 232101 204748 232110
rect 204500 231574 204556 231583
rect 204500 231509 204556 231518
rect 204802 230991 204830 246573
rect 205174 244485 205226 244491
rect 205174 244427 205226 244433
rect 204982 244189 205034 244195
rect 204982 244131 205034 244137
rect 204788 230982 204844 230991
rect 204788 230917 204844 230926
rect 204994 227735 205022 244131
rect 204980 227726 205036 227735
rect 194326 227687 194378 227693
rect 204980 227661 205036 227670
rect 194326 227629 194378 227635
rect 192886 215921 192938 215927
rect 192886 215863 192938 215869
rect 191446 198753 191498 198759
rect 191446 198695 191498 198701
rect 188662 181511 188714 181517
rect 188662 181453 188714 181459
rect 188674 92051 188702 181453
rect 188758 118537 188810 118543
rect 188758 118479 188810 118485
rect 188662 92045 188714 92051
rect 188662 91987 188714 91993
rect 188770 80655 188798 118479
rect 188758 80649 188810 80655
rect 188758 80591 188810 80597
rect 188566 47127 188618 47133
rect 188566 47069 188618 47075
rect 191458 46985 191486 198695
rect 191542 178625 191594 178631
rect 191542 178567 191594 178573
rect 191554 88943 191582 178567
rect 191638 112691 191690 112697
rect 191638 112633 191690 112639
rect 191542 88937 191594 88943
rect 191542 88879 191594 88885
rect 191650 77399 191678 112633
rect 191638 77393 191690 77399
rect 191638 77335 191690 77341
rect 194338 48391 194366 227629
rect 197206 227613 197258 227619
rect 197206 227555 197258 227561
rect 194422 184397 194474 184403
rect 194422 184339 194474 184345
rect 194434 91977 194462 184339
rect 194518 118167 194570 118173
rect 194518 118109 194570 118115
rect 194422 91971 194474 91977
rect 194422 91913 194474 91919
rect 194530 80581 194558 118109
rect 194518 80575 194570 80581
rect 194518 80517 194570 80523
rect 197218 48465 197246 227555
rect 205186 225663 205214 244427
rect 205282 243011 205310 247609
rect 205570 244584 205598 249237
rect 206626 244607 206654 271437
rect 210946 268689 210974 277870
rect 212208 277856 212510 277884
rect 212374 273567 212426 273573
rect 212374 273509 212426 273515
rect 211606 272901 211658 272907
rect 211606 272843 211658 272849
rect 210934 268683 210986 268689
rect 210934 268625 210986 268631
rect 211508 268278 211564 268287
rect 211508 268213 211564 268222
rect 210646 264909 210698 264915
rect 210646 264851 210698 264857
rect 207188 261322 207244 261331
rect 207188 261257 207244 261266
rect 207092 249334 207148 249343
rect 207092 249269 207148 249278
rect 206902 249147 206954 249153
rect 206902 249089 206954 249095
rect 206914 245749 206942 249089
rect 206902 245743 206954 245749
rect 206902 245685 206954 245691
rect 207106 244732 207134 249269
rect 206818 244704 207134 244732
rect 205474 244556 205598 244584
rect 206612 244598 206668 244607
rect 205366 244337 205418 244343
rect 205366 244279 205418 244285
rect 205270 243005 205322 243011
rect 205270 242947 205322 242953
rect 205268 232610 205324 232619
rect 205268 232545 205324 232554
rect 205282 227915 205310 232545
rect 205270 227909 205322 227915
rect 205270 227851 205322 227857
rect 205378 226699 205406 244279
rect 205474 230547 205502 244556
rect 206612 244533 206668 244542
rect 205558 244411 205610 244417
rect 205558 244353 205610 244359
rect 205460 230538 205516 230547
rect 205460 230473 205516 230482
rect 205364 226690 205420 226699
rect 205364 226625 205420 226634
rect 205570 226107 205598 244353
rect 205654 244263 205706 244269
rect 205654 244205 205706 244211
rect 205666 228008 205694 244205
rect 206614 244115 206666 244121
rect 206614 244057 206666 244063
rect 205750 244041 205802 244047
rect 205750 243983 205802 243989
rect 205762 228211 205790 243983
rect 206518 243967 206570 243973
rect 206518 243909 206570 243915
rect 206326 243893 206378 243899
rect 206326 243835 206378 243841
rect 206230 243745 206282 243751
rect 206230 243687 206282 243693
rect 206038 243671 206090 243677
rect 206038 243613 206090 243619
rect 205942 243449 205994 243455
rect 205942 243391 205994 243397
rect 205846 241969 205898 241975
rect 205846 241911 205898 241917
rect 205750 228205 205802 228211
rect 205750 228147 205802 228153
rect 205666 227980 205790 228008
rect 205654 227909 205706 227915
rect 205654 227851 205706 227857
rect 205556 226098 205612 226107
rect 205556 226033 205612 226042
rect 205172 225654 205228 225663
rect 205172 225589 205228 225598
rect 200086 224727 200138 224733
rect 200086 224669 200138 224675
rect 197302 187283 197354 187289
rect 197302 187225 197354 187231
rect 197314 91829 197342 187225
rect 197398 124013 197450 124019
rect 197398 123955 197450 123961
rect 197302 91823 197354 91829
rect 197302 91765 197354 91771
rect 197410 80359 197438 123955
rect 197398 80353 197450 80359
rect 197398 80295 197450 80301
rect 197206 48459 197258 48465
rect 197206 48401 197258 48407
rect 194326 48385 194378 48391
rect 194326 48327 194378 48333
rect 200098 47281 200126 224669
rect 204502 224653 204554 224659
rect 204502 224595 204554 224601
rect 204514 224035 204542 224595
rect 204598 224579 204650 224585
rect 204598 224521 204650 224527
rect 204500 224026 204556 224035
rect 204500 223961 204556 223970
rect 204610 223443 204638 224521
rect 204694 224505 204746 224511
rect 204694 224447 204746 224453
rect 204596 223434 204652 223443
rect 204596 223369 204652 223378
rect 204706 222851 204734 224447
rect 204790 224431 204842 224437
rect 204790 224373 204842 224379
rect 204692 222842 204748 222851
rect 204692 222777 204748 222786
rect 204802 221815 204830 224373
rect 204788 221806 204844 221815
rect 204502 221767 204554 221773
rect 204788 221741 204844 221750
rect 204502 221709 204554 221715
rect 204514 221223 204542 221709
rect 204598 221693 204650 221699
rect 204598 221635 204650 221641
rect 204500 221214 204556 221223
rect 204500 221149 204556 221158
rect 204610 221075 204638 221635
rect 204694 221619 204746 221625
rect 204694 221561 204746 221567
rect 204596 221066 204652 221075
rect 204596 221001 204652 221010
rect 204706 220187 204734 221561
rect 204790 221545 204842 221551
rect 204790 221487 204842 221493
rect 204692 220178 204748 220187
rect 204692 220113 204748 220122
rect 204802 219595 204830 221487
rect 204886 221471 204938 221477
rect 204886 221413 204938 221419
rect 204788 219586 204844 219595
rect 204788 219521 204844 219530
rect 204898 219447 204926 221413
rect 204884 219438 204940 219447
rect 204884 219373 204940 219382
rect 204502 218881 204554 218887
rect 204502 218823 204554 218829
rect 204514 218559 204542 218823
rect 204598 218807 204650 218813
rect 204598 218749 204650 218755
rect 204500 218550 204556 218559
rect 204500 218485 204556 218494
rect 204610 217967 204638 218749
rect 204694 218733 204746 218739
rect 204694 218675 204746 218681
rect 204596 217958 204652 217967
rect 204596 217893 204652 217902
rect 204706 217819 204734 218675
rect 204790 218659 204842 218665
rect 204790 218601 204842 218607
rect 204692 217810 204748 217819
rect 204692 217745 204748 217754
rect 204802 216931 204830 218601
rect 204788 216922 204844 216931
rect 204788 216857 204844 216866
rect 204502 215995 204554 216001
rect 204502 215937 204554 215943
rect 204514 215895 204542 215937
rect 204598 215921 204650 215927
rect 204500 215886 204556 215895
rect 204598 215863 204650 215869
rect 204500 215821 204556 215830
rect 204610 215303 204638 215863
rect 204596 215294 204652 215303
rect 204596 215229 204652 215238
rect 203062 207411 203114 207417
rect 203062 207353 203114 207359
rect 202966 201639 203018 201645
rect 202966 201581 203018 201587
rect 200182 155611 200234 155617
rect 200182 155553 200234 155559
rect 200194 91903 200222 155553
rect 200278 123939 200330 123945
rect 200278 123881 200330 123887
rect 200182 91897 200234 91903
rect 200182 91839 200234 91845
rect 200290 80433 200318 123881
rect 201718 94931 201770 94937
rect 201718 94873 201770 94879
rect 201730 92315 201758 94873
rect 201716 92306 201772 92315
rect 201716 92241 201772 92250
rect 200278 80427 200330 80433
rect 200278 80369 200330 80375
rect 202978 48317 203006 201581
rect 203074 94493 203102 207353
rect 203158 126825 203210 126831
rect 203158 126767 203210 126773
rect 203062 94487 203114 94493
rect 203062 94429 203114 94435
rect 203170 80507 203198 126767
rect 204502 103663 204554 103669
rect 204502 103605 204554 103611
rect 204514 102083 204542 103605
rect 204598 103589 204650 103595
rect 204598 103531 204650 103537
rect 204500 102074 204556 102083
rect 204500 102009 204556 102018
rect 204610 101639 204638 103531
rect 204694 103515 204746 103521
rect 204694 103457 204746 103463
rect 204596 101630 204652 101639
rect 204596 101565 204652 101574
rect 204706 101047 204734 103457
rect 204692 101038 204748 101047
rect 204692 100973 204748 100982
rect 204886 100777 204938 100783
rect 204886 100719 204938 100725
rect 204790 100703 204842 100709
rect 204790 100645 204842 100651
rect 204598 100629 204650 100635
rect 204598 100571 204650 100577
rect 204502 100481 204554 100487
rect 204610 100455 204638 100571
rect 204694 100555 204746 100561
rect 204694 100497 204746 100503
rect 204502 100423 204554 100429
rect 204596 100446 204652 100455
rect 204514 100307 204542 100423
rect 204596 100381 204652 100390
rect 204500 100298 204556 100307
rect 204500 100233 204556 100242
rect 204706 99419 204734 100497
rect 204692 99410 204748 99419
rect 204692 99345 204748 99354
rect 204802 98827 204830 100645
rect 204788 98818 204844 98827
rect 204788 98753 204844 98762
rect 204898 98679 204926 100719
rect 204884 98670 204940 98679
rect 204884 98605 204940 98614
rect 204790 97891 204842 97897
rect 204790 97833 204842 97839
rect 204502 97817 204554 97823
rect 204500 97782 204502 97791
rect 204554 97782 204556 97791
rect 204500 97717 204556 97726
rect 204694 97743 204746 97749
rect 204694 97685 204746 97691
rect 204598 97669 204650 97675
rect 204598 97611 204650 97617
rect 204502 97595 204554 97601
rect 204502 97537 204554 97543
rect 204514 97199 204542 97537
rect 204500 97190 204556 97199
rect 204500 97125 204556 97134
rect 204610 97051 204638 97611
rect 204596 97042 204652 97051
rect 204596 96977 204652 96986
rect 204706 95571 204734 97685
rect 204802 96163 204830 97833
rect 204788 96154 204844 96163
rect 204788 96089 204844 96098
rect 204692 95562 204748 95571
rect 204692 95497 204748 95506
rect 204790 94857 204842 94863
rect 204596 94822 204652 94831
rect 204502 94783 204554 94789
rect 204790 94799 204842 94805
rect 204596 94757 204652 94766
rect 204502 94725 204554 94731
rect 204514 94535 204542 94725
rect 204610 94715 204638 94757
rect 204598 94709 204650 94715
rect 204598 94651 204650 94657
rect 204694 94635 204746 94641
rect 204694 94577 204746 94583
rect 204500 94526 204556 94535
rect 204500 94461 204556 94470
rect 204706 92907 204734 94577
rect 204802 93795 204830 94799
rect 205270 94487 205322 94493
rect 205270 94429 205322 94435
rect 205282 93943 205310 94429
rect 205268 93934 205324 93943
rect 205268 93869 205324 93878
rect 204788 93786 204844 93795
rect 204788 93721 204844 93730
rect 204692 92898 204748 92907
rect 204692 92833 204748 92842
rect 204502 92119 204554 92125
rect 204502 92061 204554 92067
rect 204514 92019 204542 92061
rect 204694 92045 204746 92051
rect 204500 92010 204556 92019
rect 204694 91987 204746 91993
rect 204500 91945 204556 91954
rect 204598 91971 204650 91977
rect 204598 91913 204650 91919
rect 204502 91823 204554 91829
rect 204502 91765 204554 91771
rect 204514 90687 204542 91765
rect 204500 90678 204556 90687
rect 204500 90613 204556 90622
rect 204610 90095 204638 91913
rect 204596 90086 204652 90095
rect 204596 90021 204652 90030
rect 204706 89651 204734 91987
rect 205366 91897 205418 91903
rect 205366 91839 205418 91845
rect 205378 91279 205406 91839
rect 205364 91270 205420 91279
rect 205364 91205 205420 91214
rect 204692 89642 204748 89651
rect 204692 89577 204748 89586
rect 204886 89233 204938 89239
rect 204886 89175 204938 89181
rect 204790 89159 204842 89165
rect 204790 89101 204842 89107
rect 204694 89085 204746 89091
rect 204500 89050 204556 89059
rect 204694 89027 204746 89033
rect 204500 88985 204556 88994
rect 204598 89011 204650 89017
rect 204514 88943 204542 88985
rect 204598 88953 204650 88959
rect 204502 88937 204554 88943
rect 204502 88879 204554 88885
rect 204610 88467 204638 88953
rect 204596 88458 204652 88467
rect 204596 88393 204652 88402
rect 204706 88023 204734 89027
rect 204692 88014 204748 88023
rect 204692 87949 204748 87958
rect 204802 87431 204830 89101
rect 204788 87422 204844 87431
rect 204788 87357 204844 87366
rect 204898 86839 204926 89175
rect 204884 86830 204940 86839
rect 204884 86765 204940 86774
rect 204886 86421 204938 86427
rect 204500 86386 204556 86395
rect 204886 86363 204938 86369
rect 204500 86321 204556 86330
rect 204790 86347 204842 86353
rect 204514 86131 204542 86321
rect 204790 86289 204842 86295
rect 204694 86273 204746 86279
rect 204694 86215 204746 86221
rect 204598 86199 204650 86205
rect 204598 86141 204650 86147
rect 204502 86125 204554 86131
rect 204502 86067 204554 86073
rect 204500 85794 204556 85803
rect 204500 85729 204556 85738
rect 204514 85021 204542 85729
rect 204610 85211 204638 86141
rect 204596 85202 204652 85211
rect 204596 85137 204652 85146
rect 204502 85015 204554 85021
rect 204502 84957 204554 84963
rect 204706 84767 204734 86215
rect 204692 84758 204748 84767
rect 204692 84693 204748 84702
rect 204802 84175 204830 86289
rect 204788 84166 204844 84175
rect 204788 84101 204844 84110
rect 204898 83583 204926 86363
rect 204884 83574 204940 83583
rect 204790 83535 204842 83541
rect 204884 83509 204940 83518
rect 204790 83477 204842 83483
rect 204694 83461 204746 83467
rect 204694 83403 204746 83409
rect 204598 83387 204650 83393
rect 204598 83329 204650 83335
rect 204502 83313 204554 83319
rect 204502 83255 204554 83261
rect 204514 83139 204542 83255
rect 204500 83130 204556 83139
rect 204500 83065 204556 83074
rect 204610 82547 204638 83329
rect 204596 82538 204652 82547
rect 204596 82473 204652 82482
rect 204502 82129 204554 82135
rect 204502 82071 204554 82077
rect 204514 81955 204542 82071
rect 204500 81946 204556 81955
rect 204500 81881 204556 81890
rect 204706 81511 204734 83403
rect 204692 81502 204748 81511
rect 204692 81437 204748 81446
rect 204802 80919 204830 83477
rect 204788 80910 204844 80919
rect 204788 80845 204844 80854
rect 204598 80649 204650 80655
rect 204598 80591 204650 80597
rect 204502 80575 204554 80581
rect 204502 80517 204554 80523
rect 203158 80501 203210 80507
rect 203158 80443 203210 80449
rect 204514 78699 204542 80517
rect 204500 78690 204556 78699
rect 204500 78625 204556 78634
rect 204610 78551 204638 80591
rect 205462 80427 205514 80433
rect 205462 80369 205514 80375
rect 204694 80353 204746 80359
rect 204694 80295 204746 80301
rect 204706 79291 204734 80295
rect 205474 80179 205502 80369
rect 205460 80170 205516 80179
rect 205460 80105 205516 80114
rect 204692 79282 204748 79291
rect 204692 79217 204748 79226
rect 204596 78542 204652 78551
rect 204596 78477 204652 78486
rect 204982 77763 205034 77769
rect 204982 77705 205034 77711
rect 204886 77689 204938 77695
rect 204596 77654 204652 77663
rect 204886 77631 204938 77637
rect 204596 77589 204652 77598
rect 204790 77615 204842 77621
rect 204502 77467 204554 77473
rect 204502 77409 204554 77415
rect 204514 77071 204542 77409
rect 204610 77399 204638 77589
rect 204790 77557 204842 77563
rect 204694 77541 204746 77547
rect 204694 77483 204746 77489
rect 204598 77393 204650 77399
rect 204598 77335 204650 77341
rect 204500 77062 204556 77071
rect 204500 76997 204556 77006
rect 204706 76923 204734 77483
rect 204692 76914 204748 76923
rect 204692 76849 204748 76858
rect 204802 76035 204830 77557
rect 204788 76026 204844 76035
rect 204788 75961 204844 75970
rect 204898 75443 204926 77631
rect 204884 75434 204940 75443
rect 204884 75369 204940 75378
rect 204994 75295 205022 77705
rect 204980 75286 205036 75295
rect 204980 75221 205036 75230
rect 204886 74877 204938 74883
rect 204886 74819 204938 74825
rect 204790 74803 204842 74809
rect 204790 74745 204842 74751
rect 204694 74729 204746 74735
rect 204694 74671 204746 74677
rect 204598 74655 204650 74661
rect 204598 74597 204650 74603
rect 204502 74581 204554 74587
rect 204502 74523 204554 74529
rect 204514 74407 204542 74523
rect 204500 74398 204556 74407
rect 204500 74333 204556 74342
rect 204610 73815 204638 74597
rect 204596 73806 204652 73815
rect 204596 73741 204652 73750
rect 204706 73667 204734 74671
rect 204692 73658 204748 73667
rect 204692 73593 204748 73602
rect 204802 72779 204830 74745
rect 204788 72770 204844 72779
rect 204788 72705 204844 72714
rect 204898 72187 204926 74819
rect 204884 72178 204940 72187
rect 204884 72113 204940 72122
rect 204790 71991 204842 71997
rect 204790 71933 204842 71939
rect 204694 71843 204746 71849
rect 204694 71785 204746 71791
rect 204598 71769 204650 71775
rect 204500 71734 204556 71743
rect 204598 71711 204650 71717
rect 204500 71669 204502 71678
rect 204554 71669 204556 71678
rect 204502 71637 204554 71643
rect 204610 71151 204638 71711
rect 204596 71142 204652 71151
rect 204596 71077 204652 71086
rect 204706 70559 204734 71785
rect 204692 70550 204748 70559
rect 204692 70485 204748 70494
rect 204802 69967 204830 71933
rect 204886 71917 204938 71923
rect 204886 71859 204938 71865
rect 204788 69958 204844 69967
rect 204788 69893 204844 69902
rect 204898 69523 204926 71859
rect 204884 69514 204940 69523
rect 204884 69449 204940 69458
rect 204886 69105 204938 69111
rect 204886 69047 204938 69053
rect 204790 69031 204842 69037
rect 204790 68973 204842 68979
rect 204694 68957 204746 68963
rect 204500 68922 204556 68931
rect 204694 68899 204746 68905
rect 204500 68857 204556 68866
rect 204598 68883 204650 68889
rect 204514 68815 204542 68857
rect 204598 68825 204650 68831
rect 204502 68809 204554 68815
rect 204502 68751 204554 68757
rect 204610 68339 204638 68825
rect 204596 68330 204652 68339
rect 204596 68265 204652 68274
rect 204706 67895 204734 68899
rect 204692 67886 204748 67895
rect 204692 67821 204748 67830
rect 204802 67303 204830 68973
rect 204788 67294 204844 67303
rect 204788 67229 204844 67238
rect 204898 66711 204926 69047
rect 204884 66702 204940 66711
rect 204884 66637 204940 66646
rect 204596 66258 204652 66267
rect 204596 66193 204652 66202
rect 204694 66219 204746 66225
rect 204502 66145 204554 66151
rect 204502 66087 204554 66093
rect 204514 65675 204542 66087
rect 204610 66077 204638 66193
rect 204694 66161 204746 66167
rect 204598 66071 204650 66077
rect 204598 66013 204650 66019
rect 204500 65666 204556 65675
rect 204500 65601 204556 65610
rect 204706 65083 204734 66161
rect 204692 65074 204748 65083
rect 204692 65009 204748 65018
rect 204502 64887 204554 64893
rect 204502 64829 204554 64835
rect 204514 64639 204542 64829
rect 204598 64813 204650 64819
rect 204598 64755 204650 64761
rect 204500 64630 204556 64639
rect 204500 64565 204556 64574
rect 204610 64047 204638 64755
rect 204596 64038 204652 64047
rect 204596 63973 204652 63982
rect 204500 63446 204556 63455
rect 204500 63381 204502 63390
rect 204554 63381 204556 63390
rect 204502 63349 204554 63355
rect 204596 63002 204652 63011
rect 204596 62937 204652 62946
rect 204610 60823 204638 62937
rect 204692 62410 204748 62419
rect 204692 62345 204748 62354
rect 204598 60817 204650 60823
rect 204500 60782 204556 60791
rect 204598 60759 204650 60765
rect 204706 60749 204734 62345
rect 204884 61818 204940 61827
rect 204884 61753 204940 61762
rect 204788 61374 204844 61383
rect 204788 61309 204844 61318
rect 204500 60717 204556 60726
rect 204694 60743 204746 60749
rect 204514 60675 204542 60717
rect 204694 60685 204746 60691
rect 204502 60669 204554 60675
rect 204502 60611 204554 60617
rect 204802 60527 204830 61309
rect 204898 60601 204926 61753
rect 204886 60595 204938 60601
rect 204886 60537 204938 60543
rect 204790 60521 204842 60527
rect 204790 60463 204842 60469
rect 204502 60447 204554 60453
rect 204502 60389 204554 60395
rect 204514 60051 204542 60389
rect 204694 60373 204746 60379
rect 204694 60315 204746 60321
rect 204596 60190 204652 60199
rect 204596 60125 204652 60134
rect 204500 60042 204556 60051
rect 204500 59977 204556 59986
rect 204610 59047 204638 60125
rect 204706 59163 204734 60315
rect 204692 59154 204748 59163
rect 204692 59089 204748 59098
rect 204598 59041 204650 59047
rect 204598 58983 204650 58989
rect 205666 53645 205694 227851
rect 205762 227291 205790 227980
rect 205748 227282 205804 227291
rect 205748 227217 205804 227226
rect 205858 226213 205886 241911
rect 205954 228327 205982 243391
rect 205940 228318 205996 228327
rect 205940 228253 205996 228262
rect 205942 228205 205994 228211
rect 205942 228147 205994 228153
rect 205846 226207 205898 226213
rect 205846 226149 205898 226155
rect 205954 226084 205982 228147
rect 206050 226139 206078 243613
rect 206134 243375 206186 243381
rect 206134 243317 206186 243323
rect 206146 229363 206174 243317
rect 206132 229354 206188 229363
rect 206132 229289 206188 229298
rect 205762 226056 205982 226084
rect 206038 226133 206090 226139
rect 206038 226075 206090 226081
rect 205762 212047 205790 226056
rect 205846 225985 205898 225991
rect 205846 225927 205898 225933
rect 205748 212038 205804 212047
rect 205748 211973 205804 211982
rect 205858 211455 205886 225927
rect 206242 214563 206270 243687
rect 206338 226287 206366 243835
rect 206422 243819 206474 243825
rect 206422 243761 206474 243767
rect 206326 226281 206378 226287
rect 206326 226223 206378 226229
rect 206326 226133 206378 226139
rect 206326 226075 206378 226081
rect 206338 214711 206366 226075
rect 206324 214702 206380 214711
rect 206324 214637 206380 214646
rect 206228 214554 206284 214563
rect 206228 214489 206284 214498
rect 206434 213675 206462 243761
rect 206420 213666 206476 213675
rect 206420 213601 206476 213610
rect 206530 212935 206558 243909
rect 206626 226435 206654 244057
rect 206818 243677 206846 244704
rect 206998 244633 207050 244639
rect 206900 244598 206956 244607
rect 206998 244575 207050 244581
rect 206900 244533 206956 244542
rect 206806 243671 206858 243677
rect 206806 243613 206858 243619
rect 206710 243597 206762 243603
rect 206710 243539 206762 243545
rect 206614 226429 206666 226435
rect 206614 226371 206666 226377
rect 206614 226281 206666 226287
rect 206614 226223 206666 226229
rect 206626 213083 206654 226223
rect 206722 216339 206750 243539
rect 206806 243523 206858 243529
rect 206806 243465 206858 243471
rect 206818 222407 206846 243465
rect 206914 243423 206942 244533
rect 206900 243414 206956 243423
rect 206900 243349 206956 243358
rect 206900 227430 206956 227439
rect 206900 227365 206956 227374
rect 206914 225071 206942 227365
rect 206900 225062 206956 225071
rect 206900 224997 206956 225006
rect 207010 224479 207038 244575
rect 207094 244559 207146 244565
rect 207094 244501 207146 244507
rect 207106 227439 207134 244501
rect 207202 243899 207230 261257
rect 207284 255402 207340 255411
rect 207284 255337 207340 255346
rect 207298 246193 207326 255337
rect 208724 247706 208780 247715
rect 208724 247641 208780 247650
rect 207286 246187 207338 246193
rect 207286 246129 207338 246135
rect 208738 245971 208766 247641
rect 210356 247114 210412 247123
rect 210356 247049 210412 247058
rect 210164 246818 210220 246827
rect 210164 246753 210220 246762
rect 210178 246119 210206 246753
rect 210260 246522 210316 246531
rect 210260 246457 210316 246466
rect 210274 246267 210302 246457
rect 210370 246383 210398 247049
rect 210356 246374 210412 246383
rect 210356 246309 210412 246318
rect 210262 246261 210314 246267
rect 210262 246203 210314 246209
rect 210166 246113 210218 246119
rect 210166 246055 210218 246061
rect 210356 246078 210412 246087
rect 210412 246036 210494 246064
rect 210356 246013 210412 246022
rect 208726 245965 208778 245971
rect 208726 245907 208778 245913
rect 210358 245817 210410 245823
rect 210356 245782 210358 245791
rect 210410 245782 210412 245791
rect 207286 245743 207338 245749
rect 210356 245717 210412 245726
rect 207286 245685 207338 245691
rect 207190 243893 207242 243899
rect 207190 243835 207242 243841
rect 207190 243671 207242 243677
rect 207190 243613 207242 243619
rect 207202 237609 207230 243613
rect 207190 237603 207242 237609
rect 207190 237545 207242 237551
rect 207298 229955 207326 245685
rect 210356 245634 210412 245643
rect 210356 245569 210412 245578
rect 210166 245373 210218 245379
rect 210166 245315 210218 245321
rect 210260 245338 210316 245347
rect 210178 245199 210206 245315
rect 210260 245273 210316 245282
rect 210164 245190 210220 245199
rect 210164 245125 210220 245134
rect 210068 245042 210124 245051
rect 210068 244977 210124 244986
rect 209972 244894 210028 244903
rect 210082 244861 210110 244977
rect 209972 244829 210028 244838
rect 210070 244855 210122 244861
rect 209986 243719 210014 244829
rect 210070 244797 210122 244803
rect 209972 243710 210028 243719
rect 209972 243645 210028 243654
rect 210274 243127 210302 245273
rect 210370 243275 210398 245569
rect 210466 243719 210494 246036
rect 210452 243710 210508 243719
rect 210452 243645 210508 243654
rect 210356 243266 210412 243275
rect 210356 243201 210412 243210
rect 210260 243118 210316 243127
rect 210260 243053 210316 243062
rect 208534 243005 208586 243011
rect 208534 242947 208586 242953
rect 208546 239131 208574 242947
rect 210658 242387 210686 264851
rect 211522 249910 211550 268213
rect 211426 249882 211550 249910
rect 210742 249221 210794 249227
rect 210742 249163 210794 249169
rect 210644 242378 210700 242387
rect 210644 242313 210700 242322
rect 208532 239122 208588 239131
rect 208532 239057 208588 239066
rect 209876 239122 209932 239131
rect 209876 239057 209932 239066
rect 209588 237642 209644 237651
rect 209588 237577 209644 237586
rect 208150 233607 208202 233613
rect 208150 233549 208202 233555
rect 208052 230982 208108 230991
rect 208052 230917 208108 230926
rect 207284 229946 207340 229955
rect 207202 229904 207284 229932
rect 207092 227430 207148 227439
rect 207092 227365 207148 227374
rect 207094 226207 207146 226213
rect 207094 226149 207146 226155
rect 206996 224470 207052 224479
rect 206996 224405 207052 224414
rect 206804 222398 206860 222407
rect 206804 222333 206860 222342
rect 206708 216330 206764 216339
rect 206708 216265 206764 216274
rect 206612 213074 206668 213083
rect 206612 213009 206668 213018
rect 206516 212926 206572 212935
rect 206516 212861 206572 212870
rect 205844 211446 205900 211455
rect 205844 211381 205900 211390
rect 207106 202723 207134 226149
rect 207092 202714 207148 202723
rect 207092 202649 207148 202658
rect 206902 80501 206954 80507
rect 206902 80443 206954 80449
rect 206914 80327 206942 80443
rect 206900 80318 206956 80327
rect 206900 80253 206956 80262
rect 207106 64912 207134 202649
rect 207010 64884 207134 64912
rect 206900 55898 206956 55907
rect 206900 55833 206956 55842
rect 205654 53639 205706 53645
rect 205654 53581 205706 53587
rect 202966 48311 203018 48317
rect 202966 48253 203018 48259
rect 200086 47275 200138 47281
rect 200086 47217 200138 47223
rect 191446 46979 191498 46985
rect 191446 46921 191498 46927
rect 149206 46757 149258 46763
rect 149206 46699 149258 46705
rect 149110 46535 149162 46541
rect 149110 46477 149162 46483
rect 148630 46461 148682 46467
rect 148630 46403 148682 46409
rect 133654 42835 133706 42841
rect 133654 42777 133706 42783
rect 136534 42835 136586 42841
rect 136534 42777 136586 42783
rect 136546 40219 136574 42777
rect 206914 42175 206942 55833
rect 207010 54089 207038 64884
rect 207202 64764 207230 229904
rect 207284 229881 207340 229890
rect 207106 64736 207230 64764
rect 206998 54083 207050 54089
rect 206998 54025 207050 54031
rect 207106 53053 207134 64736
rect 207766 60003 207818 60009
rect 207766 59945 207818 59951
rect 207284 57526 207340 57535
rect 207284 57461 207340 57470
rect 207298 53201 207326 57461
rect 207286 53195 207338 53201
rect 207286 53137 207338 53143
rect 207094 53047 207146 53053
rect 207094 52989 207146 52995
rect 207778 46615 207806 59945
rect 208066 53793 208094 230917
rect 208054 53787 208106 53793
rect 208054 53729 208106 53735
rect 208162 52979 208190 233549
rect 209204 232166 209260 232175
rect 209204 232101 209260 232110
rect 208726 138295 208778 138301
rect 208726 138237 208778 138243
rect 208630 126751 208682 126757
rect 208630 126693 208682 126699
rect 208534 106623 208586 106629
rect 208534 106565 208586 106571
rect 208438 103737 208490 103743
rect 208438 103679 208490 103685
rect 208342 97965 208394 97971
rect 208342 97907 208394 97913
rect 208246 77837 208298 77843
rect 208246 77779 208298 77785
rect 208150 52973 208202 52979
rect 208150 52915 208202 52921
rect 208054 50457 208106 50463
rect 208054 50399 208106 50405
rect 207958 50383 208010 50389
rect 207958 50325 208010 50331
rect 207862 50309 207914 50315
rect 207862 50251 207914 50257
rect 207874 49649 207902 50251
rect 207970 49797 207998 50325
rect 208066 49945 208094 50399
rect 208258 50389 208286 77779
rect 208354 53719 208382 97907
rect 208342 53713 208394 53719
rect 208342 53655 208394 53661
rect 208246 50383 208298 50389
rect 208246 50325 208298 50331
rect 208450 50315 208478 103679
rect 208438 50309 208490 50315
rect 208438 50251 208490 50257
rect 208546 50241 208574 106565
rect 208342 50235 208394 50241
rect 208342 50177 208394 50183
rect 208534 50235 208586 50241
rect 208534 50177 208586 50183
rect 208054 49939 208106 49945
rect 208054 49881 208106 49887
rect 208354 49871 208382 50177
rect 208342 49865 208394 49871
rect 208342 49807 208394 49813
rect 207958 49791 208010 49797
rect 207958 49733 208010 49739
rect 207862 49643 207914 49649
rect 207862 49585 207914 49591
rect 208642 48761 208670 126693
rect 208738 60009 208766 138237
rect 208822 135335 208874 135341
rect 208822 135277 208874 135283
rect 208726 60003 208778 60009
rect 208726 59945 208778 59951
rect 208834 59140 208862 135277
rect 208918 132597 208970 132603
rect 208918 132539 208970 132545
rect 208738 59112 208862 59140
rect 208630 48755 208682 48761
rect 208630 48697 208682 48703
rect 208534 48237 208586 48243
rect 208534 48179 208586 48185
rect 208438 46757 208490 46763
rect 208438 46699 208490 46705
rect 207766 46609 207818 46615
rect 207766 46551 207818 46557
rect 208342 46535 208394 46541
rect 208342 46477 208394 46483
rect 208354 46245 208382 46477
rect 208450 46319 208478 46699
rect 208546 46393 208574 48179
rect 208630 48163 208682 48169
rect 208630 48105 208682 48111
rect 208642 46541 208670 48105
rect 208738 46763 208766 59112
rect 208930 58992 208958 132539
rect 209014 132523 209066 132529
rect 209014 132465 209066 132471
rect 208834 58964 208958 58992
rect 208834 48169 208862 58964
rect 209026 58844 209054 132465
rect 209110 129637 209162 129643
rect 209110 129579 209162 129585
rect 208930 58816 209054 58844
rect 208930 48243 208958 58816
rect 209122 58696 209150 129579
rect 209026 58668 209150 58696
rect 209026 48835 209054 58668
rect 209218 53497 209246 232101
rect 209492 231574 209548 231583
rect 209492 231509 209548 231518
rect 209396 230538 209452 230547
rect 209396 230473 209452 230482
rect 209302 120979 209354 120985
rect 209302 120921 209354 120927
rect 209314 106333 209342 120921
rect 209302 106327 209354 106333
rect 209302 106269 209354 106275
rect 209300 56638 209356 56647
rect 209300 56573 209356 56582
rect 209314 54163 209342 56573
rect 209302 54157 209354 54163
rect 209302 54099 209354 54105
rect 209206 53491 209258 53497
rect 209206 53433 209258 53439
rect 209410 53423 209438 230473
rect 209506 54311 209534 231509
rect 209494 54305 209546 54311
rect 209494 54247 209546 54253
rect 209398 53417 209450 53423
rect 209398 53359 209450 53365
rect 209602 51647 209630 237577
rect 209780 237050 209836 237059
rect 209780 236985 209836 236994
rect 209684 236902 209740 236911
rect 209684 236837 209740 236846
rect 209698 53275 209726 236837
rect 209794 53349 209822 236985
rect 209782 53343 209834 53349
rect 209782 53285 209834 53291
rect 209686 53269 209738 53275
rect 209686 53211 209738 53217
rect 209890 51721 209918 239057
rect 210754 236203 210782 249163
rect 210934 246705 210986 246711
rect 210934 246647 210986 246653
rect 210262 236197 210314 236203
rect 210262 236139 210314 236145
rect 210742 236197 210794 236203
rect 210742 236139 210794 236145
rect 210164 234830 210220 234839
rect 210164 234765 210220 234774
rect 209974 233533 210026 233539
rect 209974 233475 210026 233481
rect 209986 54237 210014 233475
rect 210070 233459 210122 233465
rect 210070 233401 210122 233407
rect 209974 54231 210026 54237
rect 209974 54173 210026 54179
rect 209878 51715 209930 51721
rect 209878 51657 209930 51663
rect 209590 51641 209642 51647
rect 209590 51583 209642 51589
rect 210082 48983 210110 233401
rect 210178 228919 210206 234765
rect 210164 228910 210220 228919
rect 210164 228845 210220 228854
rect 210274 227841 210302 236139
rect 210946 233484 210974 246647
rect 211426 241943 211454 249882
rect 211618 249764 211646 272843
rect 212182 272013 212234 272019
rect 212182 271955 212234 271961
rect 212086 271421 212138 271427
rect 212086 271363 212138 271369
rect 211894 271347 211946 271353
rect 211894 271289 211946 271295
rect 211798 271199 211850 271205
rect 211798 271141 211850 271147
rect 211700 271090 211756 271099
rect 211700 271025 211756 271034
rect 211522 249736 211646 249764
rect 211522 242239 211550 249736
rect 211714 246859 211742 271025
rect 211702 246853 211754 246859
rect 211702 246795 211754 246801
rect 211810 246637 211838 271141
rect 211906 246785 211934 271289
rect 211988 271238 212044 271247
rect 211988 271173 212044 271182
rect 211894 246779 211946 246785
rect 211894 246721 211946 246727
rect 211798 246631 211850 246637
rect 211798 246573 211850 246579
rect 212002 246489 212030 271173
rect 212098 246711 212126 271363
rect 212086 246705 212138 246711
rect 212086 246647 212138 246653
rect 211990 246483 212042 246489
rect 211990 246425 212042 246431
rect 212194 246415 212222 271955
rect 212276 267982 212332 267991
rect 212276 267917 212332 267926
rect 212182 246409 212234 246415
rect 212182 246351 212234 246357
rect 211508 242230 211564 242239
rect 211508 242165 211564 242174
rect 211412 241934 211468 241943
rect 211412 241869 211468 241878
rect 212290 238983 212318 267917
rect 212386 265142 212414 273509
rect 212482 265729 212510 277856
rect 213238 272161 213290 272167
rect 213238 272103 213290 272109
rect 212470 265723 212522 265729
rect 212470 265665 212522 265671
rect 213250 265142 213278 272103
rect 213346 271353 213374 277870
rect 214594 274165 214622 277870
rect 215746 276755 215774 277870
rect 215734 276749 215786 276755
rect 215734 276691 215786 276697
rect 214582 274159 214634 274165
rect 214582 274101 214634 274107
rect 216118 271421 216170 271427
rect 216118 271363 216170 271369
rect 213334 271347 213386 271353
rect 213334 271289 213386 271295
rect 214966 271273 215018 271279
rect 214966 271215 215018 271221
rect 213814 270977 213866 270983
rect 213814 270919 213866 270925
rect 213826 265156 213854 270919
rect 214486 270829 214538 270835
rect 214486 270771 214538 270777
rect 213826 265128 214080 265156
rect 214498 265142 214526 270771
rect 214978 265142 215006 271215
rect 215446 271125 215498 271131
rect 215446 271067 215498 271073
rect 215458 265142 215486 271067
rect 215542 270755 215594 270761
rect 215542 270697 215594 270703
rect 215554 265156 215582 270697
rect 216130 265156 216158 271363
rect 216694 271347 216746 271353
rect 216694 271289 216746 271295
rect 215554 265128 215808 265156
rect 216130 265128 216288 265156
rect 216706 265142 216734 271289
rect 216898 265156 216926 277870
rect 217558 270755 217610 270761
rect 217558 270697 217610 270703
rect 216898 265128 217200 265156
rect 217570 265142 217598 270697
rect 218050 268393 218078 277870
rect 219312 277856 219614 277884
rect 219286 271199 219338 271205
rect 219286 271141 219338 271147
rect 218902 271125 218954 271131
rect 218902 271067 218954 271073
rect 218710 270977 218762 270983
rect 218710 270919 218762 270925
rect 218230 270829 218282 270835
rect 218230 270771 218282 270777
rect 218038 268387 218090 268393
rect 218038 268329 218090 268335
rect 218242 265156 218270 270771
rect 218722 265156 218750 270919
rect 218016 265128 218270 265156
rect 218496 265128 218750 265156
rect 218914 265142 218942 271067
rect 219298 265142 219326 271141
rect 219586 265137 219614 277856
rect 220342 271421 220394 271427
rect 220342 271363 220394 271369
rect 219766 271347 219818 271353
rect 219766 271289 219818 271295
rect 219778 265142 219806 271289
rect 220354 265156 220382 271363
rect 220450 270761 220478 277870
rect 220822 272901 220874 272907
rect 220822 272843 220874 272849
rect 220438 270755 220490 270761
rect 220438 270697 220490 270703
rect 220834 265156 220862 272843
rect 221014 272161 221066 272167
rect 221014 272103 221066 272109
rect 219574 265131 219626 265137
rect 220224 265128 220382 265156
rect 220608 265128 220862 265156
rect 221026 265142 221054 272103
rect 221494 269275 221546 269281
rect 221494 269217 221546 269223
rect 221506 265142 221534 269217
rect 221698 265285 221726 277870
rect 223030 274677 223082 274683
rect 223030 274619 223082 274625
rect 222550 268239 222602 268245
rect 222550 268181 222602 268187
rect 221974 268017 222026 268023
rect 221974 267959 222026 267965
rect 221686 265279 221738 265285
rect 221686 265221 221738 265227
rect 221986 265142 222014 267959
rect 222562 265156 222590 268181
rect 223042 265156 223070 274619
rect 223702 271495 223754 271501
rect 223702 271437 223754 271443
rect 223222 268165 223274 268171
rect 223222 268107 223274 268113
rect 222336 265128 222590 265156
rect 222816 265128 223070 265156
rect 223234 265142 223262 268107
rect 223714 265142 223742 271437
rect 224002 270835 224030 277870
rect 225250 277125 225278 277870
rect 225238 277119 225290 277125
rect 225238 277061 225290 277067
rect 226294 274307 226346 274313
rect 226294 274249 226346 274255
rect 225430 274085 225482 274091
rect 225430 274027 225482 274033
rect 225238 274011 225290 274017
rect 225238 273953 225290 273959
rect 224566 273493 224618 273499
rect 224566 273435 224618 273441
rect 224086 272013 224138 272019
rect 224086 271955 224138 271961
rect 223990 270829 224042 270835
rect 223990 270771 224042 270777
rect 224098 265142 224126 271955
rect 224578 265156 224606 273435
rect 225250 265156 225278 273953
rect 224544 265128 224606 265156
rect 225024 265128 225278 265156
rect 225442 265142 225470 274027
rect 225814 268831 225866 268837
rect 225814 268773 225866 268779
rect 225826 265142 225854 268773
rect 226306 265142 226334 274249
rect 226402 265951 226430 277870
rect 227446 275787 227498 275793
rect 227446 275729 227498 275735
rect 226966 269867 227018 269873
rect 226966 269809 227018 269815
rect 226390 265945 226442 265951
rect 226390 265887 226442 265893
rect 226978 265156 227006 269809
rect 227458 265156 227486 275729
rect 227650 270983 227678 277870
rect 228022 275195 228074 275201
rect 228022 275137 228074 275143
rect 227638 270977 227690 270983
rect 227638 270919 227690 270925
rect 227542 269497 227594 269503
rect 227542 269439 227594 269445
rect 226752 265128 227006 265156
rect 227232 265128 227486 265156
rect 227554 265142 227582 269439
rect 228034 265142 228062 275137
rect 228502 269349 228554 269355
rect 228502 269291 228554 269297
rect 228514 265142 228542 269291
rect 228802 268319 228830 277870
rect 229078 275047 229130 275053
rect 229078 274989 229130 274995
rect 228790 268313 228842 268319
rect 228790 268255 228842 268261
rect 229090 265156 229118 274989
rect 229750 273789 229802 273795
rect 229750 273731 229802 273737
rect 229558 268979 229610 268985
rect 229558 268921 229610 268927
rect 229570 265156 229598 268921
rect 228864 265128 229118 265156
rect 229344 265128 229598 265156
rect 229762 265142 229790 273731
rect 230050 266247 230078 277870
rect 230614 276453 230666 276459
rect 230614 276395 230666 276401
rect 230230 270681 230282 270687
rect 230230 270623 230282 270629
rect 230038 266241 230090 266247
rect 230038 266183 230090 266189
rect 230242 265142 230270 270623
rect 230626 265142 230654 276395
rect 231202 271131 231230 277870
rect 231958 276305 232010 276311
rect 231958 276247 232010 276253
rect 231766 273715 231818 273721
rect 231766 273657 231818 273663
rect 231190 271125 231242 271131
rect 231190 271067 231242 271073
rect 231286 270607 231338 270613
rect 231286 270549 231338 270555
rect 231298 265156 231326 270549
rect 231778 265156 231806 273657
rect 231072 265128 231326 265156
rect 231552 265128 231806 265156
rect 231970 265142 231998 276247
rect 232342 276231 232394 276237
rect 232342 276173 232394 276179
rect 232354 265142 232382 276173
rect 232450 273869 232478 277870
rect 233494 275935 233546 275941
rect 233494 275877 233546 275883
rect 232438 273863 232490 273869
rect 232438 273805 232490 273811
rect 232822 270385 232874 270391
rect 232822 270327 232874 270333
rect 232834 265142 232862 270327
rect 233506 265156 233534 275877
rect 234070 275639 234122 275645
rect 234070 275581 234122 275587
rect 233974 270237 234026 270243
rect 233974 270179 234026 270185
rect 233986 265156 234014 270179
rect 233280 265128 233534 265156
rect 233760 265128 234014 265156
rect 234082 265142 234110 275581
rect 234658 271205 234686 277870
rect 235030 275417 235082 275423
rect 235030 275359 235082 275365
rect 234646 271199 234698 271205
rect 234646 271141 234698 271147
rect 234550 270089 234602 270095
rect 234550 270031 234602 270037
rect 234562 265142 234590 270031
rect 235042 265142 235070 275359
rect 235702 269793 235754 269799
rect 235702 269735 235754 269741
rect 235714 265156 235742 269735
rect 235906 268097 235934 277870
rect 237168 277856 237470 277884
rect 235990 275343 236042 275349
rect 235990 275285 236042 275291
rect 235894 268091 235946 268097
rect 235894 268033 235946 268039
rect 236002 265156 236030 275285
rect 236758 275121 236810 275127
rect 236758 275063 236810 275069
rect 236278 269571 236330 269577
rect 236278 269513 236330 269519
rect 235488 265128 235742 265156
rect 235872 265128 236030 265156
rect 236290 265142 236318 269513
rect 236770 265142 236798 275063
rect 237142 268461 237194 268467
rect 237142 268403 237194 268409
rect 237154 265142 237182 268403
rect 237442 266543 237470 277856
rect 237814 274381 237866 274387
rect 237814 274323 237866 274329
rect 237430 266537 237482 266543
rect 237430 266479 237482 266485
rect 237826 265156 237854 274323
rect 238306 271353 238334 277870
rect 239350 274529 239402 274535
rect 239350 274471 239402 274477
rect 238486 274455 238538 274461
rect 238486 274397 238538 274403
rect 238294 271347 238346 271353
rect 238294 271289 238346 271295
rect 238294 268535 238346 268541
rect 238294 268477 238346 268483
rect 238306 265156 238334 268477
rect 237600 265128 237854 265156
rect 238080 265128 238334 265156
rect 238498 265142 238526 274397
rect 238870 268609 238922 268615
rect 238870 268551 238922 268557
rect 238882 265142 238910 268551
rect 239362 265142 239390 274471
rect 239458 273943 239486 277870
rect 241078 274751 241130 274757
rect 241078 274693 241130 274699
rect 240502 274603 240554 274609
rect 240502 274545 240554 274551
rect 239446 273937 239498 273943
rect 239446 273879 239498 273885
rect 240022 268757 240074 268763
rect 240022 268699 240074 268705
rect 240034 265156 240062 268699
rect 240514 265156 240542 274545
rect 240886 268905 240938 268911
rect 240886 268847 240938 268853
rect 240898 265156 240926 268847
rect 239808 265128 240062 265156
rect 240288 265128 240542 265156
rect 240672 265128 240926 265156
rect 241090 265142 241118 274693
rect 241858 271427 241886 277870
rect 242998 274973 243050 274979
rect 242998 274915 243050 274921
rect 242230 274825 242282 274831
rect 242230 274767 242282 274773
rect 241846 271421 241898 271427
rect 241846 271363 241898 271369
rect 241558 269053 241610 269059
rect 241558 268995 241610 269001
rect 241570 265142 241598 268995
rect 242242 265156 242270 274767
rect 242614 269127 242666 269133
rect 242614 269069 242666 269075
rect 242626 265156 242654 269069
rect 243010 265156 243038 274915
rect 243106 267949 243134 277870
rect 243766 276379 243818 276385
rect 243766 276321 243818 276327
rect 243286 269201 243338 269207
rect 243286 269143 243338 269149
rect 243094 267943 243146 267949
rect 243094 267885 243146 267891
rect 242016 265128 242270 265156
rect 242400 265128 242654 265156
rect 242880 265128 243038 265156
rect 243298 265142 243326 269143
rect 243778 265142 243806 276321
rect 244150 270459 244202 270465
rect 244150 270401 244202 270407
rect 244162 265142 244190 270401
rect 244258 266617 244286 277870
rect 244726 276157 244778 276163
rect 244726 276099 244778 276105
rect 244246 266611 244298 266617
rect 244246 266553 244298 266559
rect 244738 265156 244766 276099
rect 245398 276083 245450 276089
rect 245398 276025 245450 276031
rect 245302 270311 245354 270317
rect 245302 270253 245354 270259
rect 245314 265156 245342 270253
rect 244608 265128 244766 265156
rect 245088 265128 245342 265156
rect 245410 265142 245438 276025
rect 245506 272907 245534 277870
rect 246358 276009 246410 276015
rect 246358 275951 246410 275957
rect 245494 272901 245546 272907
rect 245494 272843 245546 272849
rect 245878 270163 245930 270169
rect 245878 270105 245930 270111
rect 245890 265142 245918 270105
rect 246370 265142 246398 275951
rect 246658 271427 246686 277870
rect 247906 277421 247934 277870
rect 247894 277415 247946 277421
rect 247894 277357 247946 277363
rect 247414 275861 247466 275867
rect 247414 275803 247466 275809
rect 246646 271421 246698 271427
rect 246646 271363 246698 271369
rect 247030 269941 247082 269947
rect 247030 269883 247082 269889
rect 247042 265156 247070 269883
rect 247426 265156 247454 275803
rect 248086 275713 248138 275719
rect 248086 275655 248138 275661
rect 247606 269719 247658 269725
rect 247606 269661 247658 269667
rect 246816 265128 247070 265156
rect 247200 265128 247454 265156
rect 247618 265142 247646 269661
rect 248098 265142 248126 275655
rect 249058 272167 249086 277870
rect 249142 275565 249194 275571
rect 249142 275507 249194 275513
rect 249046 272161 249098 272167
rect 249046 272103 249098 272109
rect 248566 269645 248618 269651
rect 248566 269587 248618 269593
rect 248578 265142 248606 269587
rect 249154 265156 249182 275507
rect 249812 274050 249868 274059
rect 249812 273985 249868 273994
rect 249622 269423 249674 269429
rect 249622 269365 249674 269371
rect 249634 265156 249662 269365
rect 248928 265128 249182 265156
rect 249408 265128 249662 265156
rect 249826 265142 249854 273985
rect 250210 270761 250238 277870
rect 251170 277856 251376 277884
rect 251554 277856 252528 277884
rect 250676 274198 250732 274207
rect 250676 274133 250732 274142
rect 250198 270755 250250 270761
rect 250198 270697 250250 270703
rect 250292 268130 250348 268139
rect 250292 268065 250348 268074
rect 250306 265142 250334 268065
rect 250690 265142 250718 274133
rect 251170 266913 251198 277856
rect 251554 272001 251582 277856
rect 252404 274494 252460 274503
rect 252404 274429 252460 274438
rect 251828 274346 251884 274355
rect 251828 274281 251884 274290
rect 251266 271973 251582 272001
rect 251266 269281 251294 271973
rect 251254 269275 251306 269281
rect 251254 269217 251306 269223
rect 251350 269275 251402 269281
rect 251350 269217 251402 269223
rect 251158 266907 251210 266913
rect 251158 266849 251210 266855
rect 251362 265156 251390 269217
rect 251842 265156 251870 274281
rect 252020 268426 252076 268435
rect 252020 268361 252076 268370
rect 251136 265128 251390 265156
rect 251616 265128 251870 265156
rect 252034 265142 252062 268361
rect 252418 265142 252446 274429
rect 253762 271427 253790 277870
rect 254132 274790 254188 274799
rect 254132 274725 254188 274734
rect 253940 274642 253996 274651
rect 253940 274577 253996 274586
rect 253750 271421 253802 271427
rect 253750 271363 253802 271369
rect 253364 269166 253420 269175
rect 253364 269101 253420 269110
rect 252884 268722 252940 268731
rect 252884 268657 252940 268666
rect 252898 265142 252926 268657
rect 253378 265156 253406 269101
rect 253954 265156 253982 274577
rect 253344 265128 253406 265156
rect 253728 265128 253982 265156
rect 254146 265142 254174 274725
rect 255860 268574 255916 268583
rect 255860 268509 255916 268518
rect 254612 268278 254668 268287
rect 254612 268213 254668 268222
rect 254626 265142 254654 268213
rect 255092 267834 255148 267843
rect 255092 267769 255148 267778
rect 255106 265142 255134 267769
rect 255670 265205 255722 265211
rect 255456 265153 255670 265156
rect 255456 265147 255722 265153
rect 255456 265128 255710 265147
rect 219574 265073 219626 265079
rect 255874 265008 255902 268509
rect 256162 268023 256190 277870
rect 256820 273754 256876 273763
rect 256820 273689 256876 273698
rect 256150 268017 256202 268023
rect 256150 267959 256202 267965
rect 256628 267834 256684 267843
rect 256628 267769 256684 267778
rect 256642 265156 256670 267769
rect 256368 265128 256670 265156
rect 256834 265142 256862 273689
rect 257314 270983 257342 277870
rect 257302 270977 257354 270983
rect 257302 270919 257354 270925
rect 257506 265156 257534 278448
rect 267778 278457 267902 278476
rect 268162 278457 268190 278541
rect 287254 278525 287306 278531
rect 293986 278499 294014 278596
rect 299542 278599 299594 278605
rect 299542 278541 299594 278547
rect 330166 278599 330218 278605
rect 330166 278541 330218 278547
rect 332758 278599 332810 278605
rect 332758 278541 332810 278547
rect 348790 278599 348842 278605
rect 348790 278541 348842 278547
rect 350326 278599 350378 278605
rect 383828 278638 383884 278647
rect 368564 278573 368620 278582
rect 380662 278599 380714 278605
rect 350326 278541 350378 278547
rect 299554 278499 299582 278541
rect 287254 278467 287306 278473
rect 293972 278490 294028 278499
rect 257588 278425 257644 278434
rect 267766 278451 267914 278457
rect 267818 278448 267862 278451
rect 267766 278393 267818 278399
rect 267862 278393 267914 278399
rect 268150 278451 268202 278457
rect 268150 278393 268202 278399
rect 266038 278081 266090 278087
rect 265776 278029 266038 278032
rect 265776 278023 266090 278029
rect 265776 278004 266078 278023
rect 258562 274905 258590 277870
rect 258550 274899 258602 274905
rect 258550 274841 258602 274847
rect 257878 273567 257930 273573
rect 257878 273509 257930 273515
rect 257890 265156 257918 273509
rect 259412 273310 259468 273319
rect 259412 273245 259468 273254
rect 258358 272161 258410 272167
rect 258358 272103 258410 272109
rect 258370 265156 258398 272103
rect 258932 270498 258988 270507
rect 258932 270433 258988 270442
rect 258550 267869 258602 267875
rect 258550 267811 258602 267817
rect 257232 265128 257534 265156
rect 257664 265128 257918 265156
rect 258144 265128 258398 265156
rect 258562 265142 258590 267811
rect 258946 265142 258974 270433
rect 259426 265142 259454 273245
rect 259714 268245 259742 277870
rect 260962 270835 260990 277870
rect 262128 277856 262430 277884
rect 261620 274938 261676 274947
rect 261620 274873 261676 274882
rect 260950 270829 261002 270835
rect 260660 270794 260716 270803
rect 260950 270771 261002 270777
rect 260660 270729 260716 270738
rect 260564 269018 260620 269027
rect 260564 268953 260620 268962
rect 259702 268239 259754 268245
rect 259702 268181 259754 268187
rect 260086 268239 260138 268245
rect 260086 268181 260138 268187
rect 260098 265156 260126 268181
rect 260578 265156 260606 268953
rect 259872 265128 260126 265156
rect 260352 265128 260606 265156
rect 260674 265142 260702 270729
rect 261140 269758 261196 269767
rect 261140 269693 261196 269702
rect 261154 265142 261182 269693
rect 261634 265142 261662 274873
rect 262004 269906 262060 269915
rect 262004 269841 262060 269850
rect 262018 265156 262046 269841
rect 262402 267135 262430 277856
rect 262868 276418 262924 276427
rect 262868 276353 262924 276362
rect 262678 273641 262730 273647
rect 262678 273583 262730 273589
rect 262390 267129 262442 267135
rect 262390 267071 262442 267077
rect 262690 265156 262718 273583
rect 261984 265128 262046 265156
rect 262464 265128 262718 265156
rect 262882 265142 262910 276353
rect 263362 274683 263390 277870
rect 264404 275530 264460 275539
rect 264404 275465 264460 275474
rect 263350 274677 263402 274683
rect 263350 274619 263402 274625
rect 263348 273902 263404 273911
rect 263348 273837 263404 273846
rect 263362 265142 263390 273837
rect 263732 267982 263788 267991
rect 263732 267917 263788 267926
rect 263746 265142 263774 267917
rect 264418 265156 264446 275465
rect 264514 271353 264542 277870
rect 265940 275382 265996 275391
rect 265940 275317 265996 275326
rect 264502 271347 264554 271353
rect 264502 271289 264554 271295
rect 265460 271090 265516 271099
rect 265460 271025 265516 271034
rect 264884 269610 264940 269619
rect 264884 269545 264940 269554
rect 264898 265156 264926 269545
rect 265076 268278 265132 268287
rect 265076 268213 265132 268222
rect 264192 265128 264446 265156
rect 264672 265128 264926 265156
rect 265090 265142 265118 268213
rect 265474 265142 265502 271025
rect 265954 265142 265982 275317
rect 266612 269462 266668 269471
rect 266612 269397 266668 269406
rect 266626 265156 266654 269397
rect 266818 268171 266846 277870
rect 267092 275234 267148 275243
rect 267092 275169 267148 275178
rect 266806 268165 266858 268171
rect 266806 268107 266858 268113
rect 267106 265156 267134 275169
rect 267188 275086 267244 275095
rect 267188 275021 267244 275030
rect 266400 265128 266654 265156
rect 266880 265128 267134 265156
rect 267202 265142 267230 275021
rect 267862 272901 267914 272907
rect 267862 272843 267914 272849
rect 267874 271501 267902 272843
rect 268066 272019 268094 277870
rect 269218 274683 269246 277870
rect 269396 276122 269452 276131
rect 269396 276057 269452 276066
rect 269206 274677 269258 274683
rect 269206 274619 269258 274625
rect 267958 272013 268010 272019
rect 267958 271955 268010 271961
rect 268054 272013 268106 272019
rect 268054 271955 268106 271961
rect 267970 271501 267998 271955
rect 267862 271495 267914 271501
rect 267862 271437 267914 271443
rect 267958 271495 268010 271501
rect 267958 271437 268010 271443
rect 268726 271125 268778 271131
rect 268726 271067 268778 271073
rect 268148 270054 268204 270063
rect 268148 269989 268204 269998
rect 267668 269314 267724 269323
rect 267668 269249 267724 269258
rect 267682 265142 267710 269249
rect 267764 267834 267820 267843
rect 267764 267769 267820 267778
rect 255874 264980 255936 265008
rect 267778 264989 267806 267769
rect 267862 265205 267914 265211
rect 267862 265147 267914 265153
rect 267766 264983 267818 264989
rect 267766 264925 267818 264931
rect 212470 264909 212522 264915
rect 267874 264883 267902 265147
rect 268162 265142 268190 269989
rect 268738 265156 268766 271067
rect 269204 267982 269260 267991
rect 269204 267917 269260 267926
rect 269218 265156 269246 267917
rect 268512 265128 268766 265156
rect 268992 265128 269246 265156
rect 269410 265142 269438 276057
rect 270262 275491 270314 275497
rect 270262 275433 270314 275439
rect 269878 271051 269930 271057
rect 269878 270993 269930 270999
rect 269890 265142 269918 270993
rect 270274 265142 270302 275433
rect 270370 272907 270398 277870
rect 270838 275269 270890 275275
rect 270838 275211 270890 275217
rect 270358 272901 270410 272907
rect 270358 272843 270410 272849
rect 270454 272901 270506 272907
rect 270454 272843 270506 272849
rect 270466 271131 270494 272843
rect 270454 271125 270506 271131
rect 270454 271067 270506 271073
rect 270850 265156 270878 275211
rect 271318 274233 271370 274239
rect 271318 274175 271370 274181
rect 271414 274233 271466 274239
rect 271414 274175 271466 274181
rect 270934 270533 270986 270539
rect 270934 270475 270986 270481
rect 270720 265128 270878 265156
rect 270946 265156 270974 270475
rect 271330 265156 271358 274175
rect 271426 272907 271454 274175
rect 271618 273499 271646 277870
rect 272470 274159 272522 274165
rect 272470 274101 272522 274107
rect 271510 273493 271562 273499
rect 271510 273435 271562 273441
rect 271606 273493 271658 273499
rect 271606 273435 271658 273441
rect 271522 272907 271550 273435
rect 271414 272901 271466 272907
rect 271414 272843 271466 272849
rect 271510 272901 271562 272907
rect 271510 272843 271562 272849
rect 271990 268683 272042 268689
rect 271990 268625 272042 268631
rect 270946 265128 271200 265156
rect 271330 265128 271632 265156
rect 272002 265142 272030 268625
rect 272482 265142 272510 274101
rect 272770 268689 272798 277870
rect 273622 277119 273674 277125
rect 273622 277061 273674 277067
rect 272758 268683 272810 268689
rect 272758 268625 272810 268631
rect 272662 268387 272714 268393
rect 272662 268329 272714 268335
rect 272674 265156 272702 268329
rect 273142 265279 273194 265285
rect 273142 265221 273194 265227
rect 273154 265156 273182 265221
rect 273634 265156 273662 277061
rect 274018 271501 274046 277870
rect 274678 273863 274730 273869
rect 274678 273805 274730 273811
rect 274006 271495 274058 271501
rect 274006 271437 274058 271443
rect 274198 268313 274250 268319
rect 274198 268255 274250 268261
rect 272674 265128 272928 265156
rect 273154 265128 273408 265156
rect 273634 265128 273792 265156
rect 274210 265142 274238 268255
rect 274690 265142 274718 273805
rect 275170 271501 275198 277870
rect 276418 274239 276446 277870
rect 276406 274233 276458 274239
rect 276406 274175 276458 274181
rect 275254 273937 275306 273943
rect 275254 273879 275306 273885
rect 275158 271495 275210 271501
rect 275158 271437 275210 271443
rect 274870 268091 274922 268097
rect 274870 268033 274922 268039
rect 274882 265156 274910 268033
rect 275266 265156 275294 273879
rect 277570 272907 277598 277870
rect 278818 272907 278846 277870
rect 279478 273493 279530 273499
rect 279478 273435 279530 273441
rect 277558 272901 277610 272907
rect 277558 272843 277610 272849
rect 278806 272901 278858 272907
rect 278806 272843 278858 272849
rect 278998 272013 279050 272019
rect 278998 271955 279050 271961
rect 277270 271421 277322 271427
rect 277270 271363 277322 271369
rect 276406 271199 276458 271205
rect 276406 271141 276458 271147
rect 275734 267943 275786 267949
rect 275734 267885 275786 267891
rect 275746 265156 275774 267885
rect 276212 267834 276268 267843
rect 276212 267769 276268 267778
rect 276226 267727 276254 267769
rect 276214 267721 276266 267727
rect 276214 267663 276266 267669
rect 274882 265128 275136 265156
rect 275266 265128 275520 265156
rect 275746 265128 276000 265156
rect 276418 265142 276446 271141
rect 276790 270755 276842 270761
rect 276790 270697 276842 270703
rect 276502 265205 276554 265211
rect 276502 265147 276554 265153
rect 276514 264883 276542 265147
rect 276802 265142 276830 270697
rect 277282 265142 277310 271363
rect 278518 271347 278570 271353
rect 278518 271289 278570 271295
rect 277462 270977 277514 270983
rect 277462 270919 277514 270925
rect 277474 265156 277502 270919
rect 277942 270829 277994 270835
rect 277942 270771 277994 270777
rect 277954 265156 277982 270771
rect 277474 265128 277728 265156
rect 277954 265128 278208 265156
rect 278530 265142 278558 271289
rect 279010 265142 279038 271955
rect 279490 265142 279518 273435
rect 279670 271495 279722 271501
rect 279670 271437 279722 271443
rect 279682 265156 279710 271437
rect 279970 267579 279998 277870
rect 281122 274017 281150 277870
rect 281110 274011 281162 274017
rect 281110 273953 281162 273959
rect 281206 273493 281258 273499
rect 281206 273435 281258 273441
rect 280054 272901 280106 272907
rect 280054 272843 280106 272849
rect 280726 272901 280778 272907
rect 280726 272843 280778 272849
rect 279958 267573 280010 267579
rect 279958 267515 280010 267521
rect 280066 265156 280094 272843
rect 279682 265128 279936 265156
rect 280066 265128 280320 265156
rect 280738 265142 280766 272843
rect 281218 265142 281246 273435
rect 282370 272907 282398 277870
rect 282454 273567 282506 273573
rect 282454 273509 282506 273515
rect 282466 272907 282494 273509
rect 282358 272901 282410 272907
rect 282358 272843 282410 272849
rect 282454 272901 282506 272907
rect 282454 272843 282506 272849
rect 282742 271421 282794 271427
rect 282742 271363 282794 271369
rect 282166 271051 282218 271057
rect 282166 270993 282218 270999
rect 281686 270977 281738 270983
rect 281686 270919 281738 270925
rect 281698 265142 281726 270919
rect 282178 265156 282206 270993
rect 282754 265156 282782 271363
rect 282934 271347 282986 271353
rect 282934 271289 282986 271295
rect 282048 265128 282206 265156
rect 282528 265128 282782 265156
rect 282946 265142 282974 271289
rect 283414 271273 283466 271279
rect 283414 271215 283466 271221
rect 283426 265142 283454 271215
rect 283522 268393 283550 277870
rect 284674 274091 284702 277870
rect 284950 275269 285002 275275
rect 284950 275211 285002 275217
rect 284662 274085 284714 274091
rect 284662 274027 284714 274033
rect 283798 271495 283850 271501
rect 283798 271437 283850 271443
rect 283510 268387 283562 268393
rect 283510 268329 283562 268335
rect 283810 265142 283838 271437
rect 284470 271199 284522 271205
rect 284470 271141 284522 271147
rect 284482 265156 284510 271141
rect 284962 265156 284990 275211
rect 285826 273499 285854 277870
rect 287074 274165 287102 277870
rect 287062 274159 287114 274165
rect 287062 274101 287114 274107
rect 286678 274085 286730 274091
rect 286678 274027 286730 274033
rect 285814 273493 285866 273499
rect 285814 273435 285866 273441
rect 285910 273493 285962 273499
rect 285910 273435 285962 273441
rect 285526 272013 285578 272019
rect 285526 271955 285578 271961
rect 285046 267943 285098 267949
rect 285046 267885 285098 267891
rect 284256 265128 284510 265156
rect 284736 265128 284990 265156
rect 285058 265142 285086 267885
rect 285538 265142 285566 271955
rect 285922 271205 285950 273435
rect 285910 271199 285962 271205
rect 285910 271141 285962 271147
rect 286006 268017 286058 268023
rect 286006 267959 286058 267965
rect 286018 265142 286046 267959
rect 286690 265156 286718 274027
rect 287062 268165 287114 268171
rect 287062 268107 287114 268113
rect 287074 265156 287102 268107
rect 286464 265128 286718 265156
rect 286848 265128 287102 265156
rect 287266 265142 287294 278467
rect 293782 278451 293834 278457
rect 293972 278425 294028 278434
rect 299540 278490 299596 278499
rect 299540 278425 299596 278434
rect 299732 278490 299788 278499
rect 299732 278425 299734 278434
rect 293782 278393 293834 278399
rect 299786 278425 299788 278434
rect 300404 278490 300460 278499
rect 300404 278425 300406 278434
rect 299734 278393 299786 278399
rect 300458 278425 300460 278434
rect 315284 278490 315340 278499
rect 315284 278425 315340 278434
rect 300406 278393 300458 278399
rect 293206 278377 293258 278383
rect 293206 278319 293258 278325
rect 290806 278303 290858 278309
rect 290806 278245 290858 278251
rect 288226 268837 288254 277870
rect 288406 277859 288458 277865
rect 288406 277801 288458 277807
rect 288214 268831 288266 268837
rect 288214 268773 288266 268779
rect 287734 267647 287786 267653
rect 287734 267589 287786 267595
rect 287746 265142 287774 267589
rect 288418 265156 288446 277801
rect 289270 276897 289322 276903
rect 289270 276839 289322 276845
rect 288790 267425 288842 267431
rect 288790 267367 288842 267373
rect 288802 265156 288830 267367
rect 289282 265156 289310 276839
rect 289474 270983 289502 277870
rect 289942 277785 289994 277791
rect 289942 277727 289994 277733
rect 289462 270977 289514 270983
rect 289462 270919 289514 270925
rect 289462 267277 289514 267283
rect 289462 267219 289514 267225
rect 288240 265128 288446 265156
rect 288576 265128 288830 265156
rect 289056 265128 289310 265156
rect 289474 265142 289502 267219
rect 289954 265142 289982 277727
rect 290626 268319 290654 277870
rect 290614 268313 290666 268319
rect 290614 268255 290666 268261
rect 290326 267499 290378 267505
rect 290326 267441 290378 267447
rect 290338 265142 290366 267441
rect 290818 265156 290846 278245
rect 291478 277933 291530 277939
rect 291478 277875 291530 277881
rect 291490 265156 291518 277875
rect 291874 274313 291902 277870
rect 292054 277489 292106 277495
rect 292054 277431 292106 277437
rect 291862 274307 291914 274313
rect 291862 274249 291914 274255
rect 291670 267351 291722 267357
rect 291670 267293 291722 267299
rect 290784 265128 290846 265156
rect 291264 265128 291518 265156
rect 291682 265142 291710 267293
rect 292066 265142 292094 277431
rect 292534 271125 292586 271131
rect 292534 271067 292586 271073
rect 292546 265142 292574 271067
rect 293026 271057 293054 277870
rect 293014 271051 293066 271057
rect 293014 270993 293066 270999
rect 293218 265156 293246 278319
rect 293590 267203 293642 267209
rect 293590 267145 293642 267151
rect 293602 265156 293630 267145
rect 292992 265128 293246 265156
rect 293376 265128 293630 265156
rect 293794 265142 293822 278393
rect 299542 278377 299594 278383
rect 299540 278342 299542 278351
rect 300310 278377 300362 278383
rect 299594 278342 299596 278351
rect 299540 278277 299596 278286
rect 300308 278342 300310 278351
rect 300362 278342 300364 278351
rect 300308 278277 300364 278286
rect 303380 278342 303436 278351
rect 303380 278277 303436 278286
rect 294742 278229 294794 278235
rect 294742 278171 294794 278177
rect 299542 278229 299594 278235
rect 299830 278229 299882 278235
rect 299594 278177 299830 278180
rect 299542 278171 299882 278177
rect 294288 277856 294590 277884
rect 294262 270977 294314 270983
rect 294262 270919 294314 270925
rect 294274 265142 294302 270919
rect 294562 268097 294590 277856
rect 294550 268091 294602 268097
rect 294550 268033 294602 268039
rect 294754 265142 294782 278171
rect 299554 278152 299870 278171
rect 299926 278155 299978 278161
rect 299926 278097 299978 278103
rect 299830 278081 299882 278087
rect 299938 278032 299966 278097
rect 299882 278029 299966 278032
rect 299830 278023 299966 278029
rect 300406 278081 300458 278087
rect 300406 278023 300458 278029
rect 299494 278007 299546 278013
rect 299494 277949 299546 277955
rect 299638 278007 299690 278013
rect 299842 278004 299966 278023
rect 300310 278007 300362 278013
rect 299638 277949 299690 277955
rect 300310 277949 300362 277955
rect 299506 277884 299534 277949
rect 299650 277907 299678 277949
rect 299636 277898 299692 277907
rect 295426 269873 295454 277870
rect 295798 277711 295850 277717
rect 295798 277653 295850 277659
rect 295414 269867 295466 269873
rect 295414 269809 295466 269815
rect 295318 267055 295370 267061
rect 295318 266997 295370 267003
rect 295330 265156 295358 266997
rect 295810 265156 295838 277653
rect 296470 277637 296522 277643
rect 296470 277579 296522 277585
rect 295990 266981 296042 266987
rect 295990 266923 296042 266929
rect 295104 265128 295358 265156
rect 295584 265128 295838 265156
rect 296002 265142 296030 266923
rect 296482 265142 296510 277579
rect 296674 271427 296702 277870
rect 297526 277563 297578 277569
rect 297526 277505 297578 277511
rect 296662 271421 296714 271427
rect 296662 271363 296714 271369
rect 296854 266833 296906 266839
rect 296854 266775 296906 266781
rect 296866 265142 296894 266775
rect 297538 265156 297566 277505
rect 297826 274313 297854 277870
rect 298198 277341 298250 277347
rect 298198 277283 298250 277289
rect 297814 274307 297866 274313
rect 297814 274249 297866 274255
rect 298004 268574 298060 268583
rect 298004 268509 298060 268518
rect 298018 267991 298046 268509
rect 298210 268079 298238 277283
rect 298978 275793 299006 277870
rect 299506 277856 299582 277884
rect 299554 277759 299582 277856
rect 299636 277833 299692 277842
rect 299540 277750 299596 277759
rect 299540 277685 299596 277694
rect 299062 277267 299114 277273
rect 299062 277209 299114 277215
rect 298966 275787 299018 275793
rect 298966 275729 299018 275735
rect 298210 268051 298334 268079
rect 298004 267982 298060 267991
rect 298196 267982 298252 267991
rect 298004 267917 298060 267926
rect 298114 267940 298196 267968
rect 297812 267834 297868 267843
rect 297812 267769 297868 267778
rect 297826 267653 297854 267769
rect 298006 267721 298058 267727
rect 298114 267709 298142 267940
rect 298196 267917 298252 267926
rect 298058 267681 298142 267709
rect 298006 267663 298058 267669
rect 297814 267647 297866 267653
rect 297814 267589 297866 267595
rect 298006 266759 298058 266765
rect 298006 266701 298058 266707
rect 298018 265156 298046 266701
rect 298306 265156 298334 268051
rect 298388 267834 298444 267843
rect 298388 267769 298444 267778
rect 298402 267653 298430 267769
rect 298390 267647 298442 267653
rect 298390 267589 298442 267595
rect 298582 266685 298634 266691
rect 298582 266627 298634 266633
rect 297312 265128 297566 265156
rect 297792 265128 298046 265156
rect 298224 265128 298334 265156
rect 298594 265142 298622 266627
rect 299074 265142 299102 277209
rect 300130 271353 300158 277870
rect 300322 277759 300350 277949
rect 300418 277907 300446 278023
rect 300404 277898 300460 277907
rect 300404 277833 300460 277842
rect 300308 277750 300364 277759
rect 300308 277685 300364 277694
rect 300214 277119 300266 277125
rect 300214 277061 300266 277067
rect 300118 271347 300170 271353
rect 300118 271289 300170 271295
rect 299734 266463 299786 266469
rect 299734 266405 299786 266411
rect 299746 265156 299774 266405
rect 300226 265156 300254 277061
rect 301282 277051 301310 277870
rect 302544 277856 302654 277884
rect 301270 277045 301322 277051
rect 301270 276987 301322 276993
rect 300790 276971 300842 276977
rect 300790 276913 300842 276919
rect 300310 266389 300362 266395
rect 300310 266331 300362 266337
rect 299520 265128 299774 265156
rect 300000 265128 300254 265156
rect 300322 265142 300350 266331
rect 300802 265142 300830 276913
rect 301846 276823 301898 276829
rect 301846 276765 301898 276771
rect 301270 266315 301322 266321
rect 301270 266257 301322 266263
rect 301282 265142 301310 266257
rect 301858 265156 301886 276765
rect 302518 271051 302570 271057
rect 302518 270993 302570 270999
rect 302326 266167 302378 266173
rect 302326 266109 302378 266115
rect 302338 265156 302366 266109
rect 301632 265128 301886 265156
rect 302112 265128 302366 265156
rect 302530 265142 302558 270993
rect 302626 269503 302654 277856
rect 302614 269497 302666 269503
rect 302614 269439 302666 269445
rect 302998 266093 303050 266099
rect 302998 266035 303050 266041
rect 303010 265142 303038 266035
rect 303394 265142 303422 278277
rect 304532 278194 304588 278203
rect 304532 278129 304588 278138
rect 303682 271279 303710 277870
rect 303670 271273 303722 271279
rect 303670 271215 303722 271221
rect 304054 266019 304106 266025
rect 304054 265961 304106 265967
rect 304066 265156 304094 265961
rect 304546 265156 304574 278129
rect 305204 278046 305260 278055
rect 305204 277981 305260 277990
rect 304930 274017 304958 277870
rect 304918 274011 304970 274017
rect 304918 273953 304970 273959
rect 304726 265871 304778 265877
rect 304726 265813 304778 265819
rect 303840 265128 304094 265156
rect 304320 265128 304574 265156
rect 304738 265142 304766 265813
rect 305218 265156 305246 277981
rect 306356 277898 306412 277907
rect 306082 275201 306110 277870
rect 306356 277833 306412 277842
rect 306070 275195 306122 275201
rect 306070 275137 306122 275143
rect 305590 265797 305642 265803
rect 305590 265739 305642 265745
rect 305136 265128 305246 265156
rect 305602 265142 305630 265739
rect 306370 265156 306398 277833
rect 307124 277750 307180 277759
rect 307124 277685 307180 277694
rect 306742 265649 306794 265655
rect 306742 265591 306794 265597
rect 306754 265156 306782 265591
rect 307138 265156 307166 277685
rect 307330 271501 307358 277870
rect 308372 277602 308428 277611
rect 308372 277537 308428 277546
rect 307318 271495 307370 271501
rect 307318 271437 307370 271443
rect 308182 271347 308234 271353
rect 308182 271289 308234 271295
rect 308194 270983 308222 271289
rect 308182 270977 308234 270983
rect 308182 270919 308234 270925
rect 307798 270533 307850 270539
rect 307798 270475 307850 270481
rect 307318 265575 307370 265581
rect 307318 265517 307370 265523
rect 306048 265128 306398 265156
rect 306528 265128 306782 265156
rect 306912 265128 307166 265156
rect 307330 265142 307358 265517
rect 307810 265142 307838 270475
rect 308086 265205 308138 265211
rect 308386 265156 308414 277537
rect 308482 271279 308510 277870
rect 309524 277454 309580 277463
rect 309524 277389 309580 277398
rect 308854 273863 308906 273869
rect 308854 273805 308906 273811
rect 308470 271273 308522 271279
rect 308470 271215 308522 271221
rect 308866 265156 308894 273805
rect 309334 265501 309386 265507
rect 309334 265443 309386 265449
rect 309346 265156 309374 265443
rect 308086 265147 308138 265153
rect 308098 264883 308126 265147
rect 308256 265128 308414 265156
rect 308640 265128 308894 265156
rect 309120 265128 309374 265156
rect 309538 265142 309566 277389
rect 309730 269355 309758 277870
rect 310882 273499 310910 277870
rect 310964 277306 311020 277315
rect 310964 277241 311020 277250
rect 310870 273493 310922 273499
rect 310870 273435 310922 273441
rect 310294 270681 310346 270687
rect 310294 270623 310346 270629
rect 310390 270681 310442 270687
rect 310390 270623 310442 270629
rect 310306 269873 310334 270623
rect 310294 269867 310346 269873
rect 310294 269809 310346 269815
rect 309718 269349 309770 269355
rect 309718 269291 309770 269297
rect 309910 265427 309962 265433
rect 309910 265369 309962 265375
rect 309922 265142 309950 265369
rect 310402 265142 310430 270623
rect 310978 265156 311006 277241
rect 311542 275787 311594 275793
rect 311542 275729 311594 275735
rect 311554 265156 311582 275729
rect 312130 271427 312158 277870
rect 312308 277158 312364 277167
rect 312308 277093 312364 277102
rect 312118 271421 312170 271427
rect 312118 271363 312170 271369
rect 311926 267573 311978 267579
rect 311926 267515 311978 267521
rect 311638 265353 311690 265359
rect 311638 265295 311690 265301
rect 310848 265128 311006 265156
rect 311328 265128 311582 265156
rect 311650 265142 311678 265295
rect 311938 265063 311966 267515
rect 312322 265156 312350 277093
rect 313282 275053 313310 277870
rect 314434 275275 314462 277870
rect 314710 277193 314762 277199
rect 314710 277135 314762 277141
rect 314722 276755 314750 277135
rect 314710 276749 314762 276755
rect 314710 276691 314762 276697
rect 314422 275269 314474 275275
rect 314422 275211 314474 275217
rect 313270 275047 313322 275053
rect 313270 274989 313322 274995
rect 314518 273493 314570 273499
rect 314518 273435 314570 273441
rect 313654 271495 313706 271501
rect 313654 271437 313706 271443
rect 312598 269497 312650 269503
rect 312598 269439 312650 269445
rect 312144 265128 312350 265156
rect 312610 265142 312638 269439
rect 312694 267795 312746 267801
rect 312694 267737 312746 267743
rect 311926 265057 311978 265063
rect 311926 264999 311978 265005
rect 312706 264989 312734 267737
rect 313270 265279 313322 265285
rect 313270 265221 313322 265227
rect 313282 265156 313310 265221
rect 313666 265156 313694 271437
rect 314420 270054 314476 270063
rect 314038 270015 314090 270021
rect 314420 269989 314422 269998
rect 314038 269957 314090 269963
rect 314474 269989 314476 269998
rect 314422 269957 314474 269963
rect 313846 269349 313898 269355
rect 313846 269291 313898 269297
rect 313056 265128 313310 265156
rect 313440 265128 313694 265156
rect 313858 265142 313886 269291
rect 314050 268985 314078 269957
rect 313942 268979 313994 268985
rect 313942 268921 313994 268927
rect 314038 268979 314090 268985
rect 314038 268921 314090 268927
rect 313954 268837 313982 268921
rect 313942 268831 313994 268837
rect 313942 268773 313994 268779
rect 314530 265156 314558 273435
rect 315298 270951 315326 278425
rect 329110 278007 329162 278013
rect 329110 277949 329162 277955
rect 315696 277856 315998 277884
rect 315382 273567 315434 273573
rect 315382 273509 315434 273515
rect 315284 270942 315340 270951
rect 315284 270877 315340 270886
rect 314806 270829 314858 270835
rect 314806 270771 314858 270777
rect 314352 265128 314558 265156
rect 314818 265142 314846 270771
rect 315394 265156 315422 273509
rect 315970 271131 315998 277856
rect 316450 277856 316752 277884
rect 317794 277856 318000 277884
rect 315958 271125 316010 271131
rect 315958 271067 316010 271073
rect 316450 268837 316478 277856
rect 316630 275269 316682 275275
rect 316630 275211 316682 275217
rect 316438 268831 316490 268837
rect 316438 268773 316490 268779
rect 315970 268236 316574 268264
rect 315970 268097 315998 268236
rect 316546 268171 316574 268236
rect 316534 268165 316586 268171
rect 316162 268097 316478 268116
rect 316534 268107 316586 268113
rect 315958 268091 316010 268097
rect 315958 268033 316010 268039
rect 316162 268091 316490 268097
rect 316162 268088 316438 268091
rect 316162 268023 316190 268088
rect 316438 268033 316490 268039
rect 316150 268017 316202 268023
rect 315860 267982 315916 267991
rect 316150 267959 316202 267965
rect 315860 267917 315916 267926
rect 315874 265156 315902 267917
rect 316642 265304 316670 275211
rect 316918 275195 316970 275201
rect 316918 275137 316970 275143
rect 316724 268870 316780 268879
rect 316724 268805 316780 268814
rect 316354 265276 316670 265304
rect 316354 265156 316382 265276
rect 316738 265156 316766 268805
rect 315168 265128 315422 265156
rect 315648 265128 315902 265156
rect 316080 265128 316382 265156
rect 316464 265128 316766 265156
rect 316930 265142 316958 275137
rect 317494 270755 317546 270761
rect 317494 270697 317546 270703
rect 317506 270655 317534 270697
rect 317492 270646 317548 270655
rect 317684 270646 317740 270655
rect 317492 270581 317548 270590
rect 317602 270604 317684 270632
rect 317602 265156 317630 270604
rect 317684 270581 317740 270590
rect 317686 268831 317738 268837
rect 317686 268773 317738 268779
rect 317698 268583 317726 268773
rect 317684 268574 317740 268583
rect 317684 268509 317740 268518
rect 317794 267949 317822 277856
rect 318644 276270 318700 276279
rect 318644 276205 318700 276214
rect 317974 275047 318026 275053
rect 317974 274989 318026 274995
rect 317876 268574 317932 268583
rect 317876 268509 317932 268518
rect 317890 267991 317918 268509
rect 317876 267982 317932 267991
rect 317782 267943 317834 267949
rect 317876 267917 317932 267926
rect 317782 267885 317834 267891
rect 317986 265156 318014 274989
rect 318164 270350 318220 270359
rect 318164 270285 318220 270294
rect 318068 269906 318124 269915
rect 318068 269841 318124 269850
rect 318082 267991 318110 269841
rect 318068 267982 318124 267991
rect 318068 267917 318124 267926
rect 317376 265128 317630 265156
rect 317856 265128 318014 265156
rect 318178 265142 318206 270285
rect 318658 265142 318686 276205
rect 319138 271205 319166 277870
rect 320098 277856 320400 277884
rect 319796 275974 319852 275983
rect 319796 275909 319852 275918
rect 319414 271347 319466 271353
rect 319414 271289 319466 271295
rect 319126 271199 319178 271205
rect 319126 271141 319178 271147
rect 318932 270202 318988 270211
rect 318932 270137 318988 270146
rect 318946 265156 318974 270137
rect 319426 267801 319454 271289
rect 319702 270829 319754 270835
rect 319702 270771 319754 270777
rect 319714 269915 319742 270771
rect 319700 269906 319756 269915
rect 319700 269841 319756 269850
rect 319414 267795 319466 267801
rect 319414 267737 319466 267743
rect 319318 265279 319370 265285
rect 319370 265239 319454 265267
rect 319318 265221 319370 265227
rect 318946 265128 319152 265156
rect 319426 265137 319454 265239
rect 319414 265131 319466 265137
rect 319414 265073 319466 265079
rect 319810 265008 319838 275909
rect 320098 273795 320126 277856
rect 320852 275826 320908 275835
rect 320852 275761 320908 275770
rect 320086 273789 320138 273795
rect 320086 273731 320138 273737
rect 320374 271347 320426 271353
rect 320374 271289 320426 271295
rect 320278 271051 320330 271057
rect 320278 270993 320330 270999
rect 320180 270054 320236 270063
rect 320180 269989 320236 269998
rect 320194 265156 320222 269989
rect 320290 265211 320318 270993
rect 319968 265128 320222 265156
rect 320278 265205 320330 265211
rect 320278 265147 320330 265153
rect 320386 265142 320414 271289
rect 320566 267573 320618 267579
rect 320566 267515 320618 267521
rect 320578 265063 320606 267515
rect 320866 265142 320894 275761
rect 321538 272019 321566 277870
rect 321908 276862 321964 276871
rect 321908 276797 321964 276806
rect 321526 272013 321578 272019
rect 321526 271955 321578 271961
rect 321622 272013 321674 272019
rect 321622 271955 321674 271961
rect 321634 271501 321662 271955
rect 321622 271495 321674 271501
rect 321622 271437 321674 271443
rect 321526 267573 321578 267579
rect 321526 267515 321578 267521
rect 321538 265156 321566 267515
rect 321922 265156 321950 276797
rect 322102 276527 322154 276533
rect 322102 276469 322154 276475
rect 322006 271125 322058 271131
rect 322006 271067 322058 271073
rect 322018 270835 322046 271067
rect 322114 271057 322142 276469
rect 322582 275491 322634 275497
rect 322582 275433 322634 275439
rect 322594 273573 322622 275433
rect 322582 273567 322634 273573
rect 322582 273509 322634 273515
rect 322678 273567 322730 273573
rect 322678 273509 322730 273515
rect 322102 271051 322154 271057
rect 322102 270993 322154 270999
rect 322690 270983 322718 273509
rect 322786 271131 322814 277870
rect 323362 277856 323952 277884
rect 324898 277856 325200 277884
rect 322868 275678 322924 275687
rect 322868 275613 322924 275622
rect 322774 271125 322826 271131
rect 322774 271067 322826 271073
rect 322678 270977 322730 270983
rect 322678 270919 322730 270925
rect 322006 270829 322058 270835
rect 322006 270771 322058 270777
rect 322390 267943 322442 267949
rect 322390 267885 322442 267891
rect 322402 267801 322430 267885
rect 322390 267795 322442 267801
rect 322390 267737 322442 267743
rect 322486 267795 322538 267801
rect 322486 267737 322538 267743
rect 322498 265156 322526 267737
rect 322882 265156 322910 275613
rect 322966 270977 323018 270983
rect 322966 270919 323018 270925
rect 322978 268097 323006 270919
rect 323362 269873 323390 277856
rect 324692 276566 324748 276575
rect 324692 276501 324748 276510
rect 324118 271421 324170 271427
rect 324118 271363 324170 271369
rect 323350 269867 323402 269873
rect 323350 269809 323402 269815
rect 323446 269867 323498 269873
rect 323446 269809 323498 269815
rect 322966 268091 323018 268097
rect 322966 268033 323018 268039
rect 323062 268091 323114 268097
rect 323062 268033 323114 268039
rect 321360 265128 321566 265156
rect 321696 265128 321950 265156
rect 322176 265128 322526 265156
rect 322608 265128 322910 265156
rect 323074 265142 323102 268033
rect 323458 265142 323486 269809
rect 324130 265156 324158 271363
rect 324500 271238 324556 271247
rect 324500 271173 324556 271182
rect 324514 268023 324542 271173
rect 324502 268017 324554 268023
rect 324502 267959 324554 267965
rect 324598 268017 324650 268023
rect 324598 267959 324650 267965
rect 324610 265156 324638 267959
rect 323904 265128 324158 265156
rect 324384 265128 324638 265156
rect 324706 265142 324734 276501
rect 324898 270983 324926 277856
rect 325282 276820 325982 276848
rect 324982 276675 325034 276681
rect 324982 276617 325034 276623
rect 324886 270977 324938 270983
rect 324886 270919 324938 270925
rect 324994 265452 325022 276617
rect 325282 273573 325310 276820
rect 325556 276714 325612 276723
rect 325556 276649 325612 276658
rect 325462 276453 325514 276459
rect 325462 276395 325514 276401
rect 325474 276131 325502 276395
rect 325460 276122 325516 276131
rect 325460 276057 325516 276066
rect 325462 273715 325514 273721
rect 325462 273657 325514 273663
rect 325474 273573 325502 273657
rect 325270 273567 325322 273573
rect 325270 273509 325322 273515
rect 325462 273567 325514 273573
rect 325462 273509 325514 273515
rect 325570 271427 325598 276649
rect 325954 276607 325982 276820
rect 325846 276601 325898 276607
rect 325846 276543 325898 276549
rect 325942 276601 325994 276607
rect 325942 276543 325994 276549
rect 325652 276122 325708 276131
rect 325652 276057 325708 276066
rect 325558 271421 325610 271427
rect 325558 271363 325610 271369
rect 325666 271353 325694 276057
rect 325654 271347 325706 271353
rect 325654 271289 325706 271295
rect 325268 270942 325324 270951
rect 325268 270877 325324 270886
rect 325282 270655 325310 270877
rect 325858 270780 325886 276543
rect 326338 270983 326366 277870
rect 327202 277856 327504 277884
rect 327202 276533 327230 277856
rect 328054 277193 328106 277199
rect 328054 277135 328106 277141
rect 328150 277193 328202 277199
rect 328150 277135 328202 277141
rect 327382 276749 327434 276755
rect 327382 276691 327434 276697
rect 327190 276527 327242 276533
rect 327190 276469 327242 276475
rect 326326 270977 326378 270983
rect 326326 270919 326378 270925
rect 325858 270752 326174 270780
rect 325654 270681 325706 270687
rect 325268 270646 325324 270655
rect 325268 270581 325324 270590
rect 325460 270646 325516 270655
rect 325654 270623 325706 270629
rect 325460 270581 325516 270590
rect 325474 270021 325502 270581
rect 325462 270015 325514 270021
rect 325462 269957 325514 269963
rect 325558 270015 325610 270021
rect 325558 269957 325610 269963
rect 325570 269873 325598 269957
rect 325666 269873 325694 270623
rect 325558 269867 325610 269873
rect 325558 269809 325610 269815
rect 325654 269867 325706 269873
rect 325654 269809 325706 269815
rect 324898 265424 325022 265452
rect 325090 269124 325310 269152
rect 312694 264983 312746 264989
rect 319584 264980 319838 265008
rect 320566 265057 320618 265063
rect 320566 264999 320618 265005
rect 312694 264925 312746 264931
rect 267860 264874 267916 264883
rect 212522 264857 212784 264860
rect 212470 264851 212784 264857
rect 212482 264832 212784 264851
rect 267860 264809 267916 264818
rect 276500 264874 276556 264883
rect 276500 264809 276556 264818
rect 308084 264874 308140 264883
rect 324898 264860 324926 265424
rect 325090 264989 325118 269124
rect 325282 268985 325310 269124
rect 325174 268979 325226 268985
rect 325174 268921 325226 268927
rect 325270 268979 325322 268985
rect 325270 268921 325322 268927
rect 325186 268560 325214 268921
rect 325186 268532 325310 268560
rect 325282 265156 325310 268532
rect 325748 267982 325804 267991
rect 325748 267917 325804 267926
rect 325282 265128 325680 265156
rect 325762 264989 325790 267917
rect 326146 265008 326174 270752
rect 327188 269906 327244 269915
rect 327188 269841 327244 269850
rect 327202 268985 327230 269841
rect 327094 268979 327146 268985
rect 327094 268921 327146 268927
rect 327190 268979 327242 268985
rect 327190 268921 327242 268927
rect 326722 268125 327038 268153
rect 326722 267727 326750 268125
rect 327010 268097 327038 268125
rect 326902 268091 326954 268097
rect 326902 268033 326954 268039
rect 326998 268091 327050 268097
rect 326998 268033 327050 268039
rect 326914 267949 326942 268033
rect 327106 267991 327134 268921
rect 327092 267982 327148 267991
rect 326806 267943 326858 267949
rect 326806 267885 326858 267891
rect 326902 267943 326954 267949
rect 327092 267917 327148 267926
rect 326902 267885 326954 267891
rect 326818 267727 326846 267885
rect 326710 267721 326762 267727
rect 326710 267663 326762 267669
rect 326806 267721 326858 267727
rect 326806 267663 326858 267669
rect 327286 265205 327338 265211
rect 327286 265147 327338 265153
rect 325078 264983 325130 264989
rect 325078 264925 325130 264931
rect 325750 264983 325802 264989
rect 326112 264980 326174 265008
rect 326230 265057 326282 265063
rect 326282 265005 326496 265008
rect 326230 264999 326496 265005
rect 326242 264980 326496 264999
rect 326722 264989 326928 265008
rect 327298 264989 327326 265147
rect 327394 265142 327422 276691
rect 327958 267647 328010 267653
rect 327958 267589 328010 267595
rect 327970 265729 327998 267589
rect 327862 265723 327914 265729
rect 327862 265665 327914 265671
rect 327958 265723 328010 265729
rect 327958 265665 328010 265671
rect 327874 265142 327902 265665
rect 328066 265156 328094 277135
rect 328162 276607 328190 277135
rect 328150 276601 328202 276607
rect 328150 276543 328202 276549
rect 328738 274091 328766 277870
rect 328726 274085 328778 274091
rect 328726 274027 328778 274033
rect 328628 271238 328684 271247
rect 328628 271173 328684 271182
rect 328436 270942 328492 270951
rect 328436 270877 328492 270886
rect 328342 270681 328394 270687
rect 328342 270623 328394 270629
rect 328354 270391 328382 270623
rect 328342 270385 328394 270391
rect 328342 270327 328394 270333
rect 328450 269915 328478 270877
rect 328642 270613 328670 271173
rect 329012 270942 329068 270951
rect 329012 270877 329068 270886
rect 328534 270607 328586 270613
rect 328534 270549 328586 270555
rect 328630 270607 328682 270613
rect 328630 270549 328682 270555
rect 328546 270391 328574 270549
rect 328534 270385 328586 270391
rect 328534 270327 328586 270333
rect 328436 269906 328492 269915
rect 328436 269841 328492 269850
rect 329026 268097 329054 270877
rect 329014 268091 329066 268097
rect 329014 268033 329066 268039
rect 328630 268017 328682 268023
rect 328630 267959 328682 267965
rect 328642 267579 328670 267959
rect 328630 267573 328682 267579
rect 328630 267515 328682 267521
rect 328066 265128 328224 265156
rect 328450 265137 328704 265156
rect 329122 265142 329150 277949
rect 329782 272013 329834 272019
rect 329782 271955 329834 271961
rect 329494 271125 329546 271131
rect 329494 271067 329546 271073
rect 329686 271125 329738 271131
rect 329686 271067 329738 271073
rect 329398 265205 329450 265211
rect 329398 265147 329450 265153
rect 328438 265131 328704 265137
rect 328490 265128 328704 265131
rect 328438 265073 328490 265079
rect 329410 264989 329438 265147
rect 329506 264989 329534 271067
rect 329698 270687 329726 271067
rect 329794 270687 329822 271955
rect 329986 271427 330014 277870
rect 329974 271421 330026 271427
rect 329974 271363 330026 271369
rect 329686 270681 329738 270687
rect 329686 270623 329738 270629
rect 329782 270681 329834 270687
rect 329782 270623 329834 270629
rect 329974 266241 330026 266247
rect 329974 266183 330026 266189
rect 329590 265945 329642 265951
rect 329590 265887 329642 265893
rect 329602 265142 329630 265887
rect 329986 265142 330014 266183
rect 330178 265156 330206 278541
rect 331318 278155 331370 278161
rect 331318 278097 331370 278103
rect 331138 270391 331166 277870
rect 331126 270385 331178 270391
rect 331126 270327 331178 270333
rect 330646 266537 330698 266543
rect 330646 266479 330698 266485
rect 330658 265156 330686 266479
rect 330178 265128 330432 265156
rect 330658 265128 330912 265156
rect 331330 265142 331358 278097
rect 332182 277415 332234 277421
rect 332182 277357 332234 277363
rect 331702 266611 331754 266617
rect 331702 266553 331754 266559
rect 331714 265142 331742 266553
rect 332194 265142 332222 277357
rect 332290 270613 332318 277870
rect 332564 270942 332620 270951
rect 332564 270877 332620 270886
rect 332278 270607 332330 270613
rect 332278 270549 332330 270555
rect 332578 270317 332606 270877
rect 332566 270311 332618 270317
rect 332566 270253 332618 270259
rect 332374 266907 332426 266913
rect 332374 266849 332426 266855
rect 332386 265156 332414 266849
rect 332770 265156 332798 278541
rect 335542 278525 335594 278531
rect 335594 278473 335856 278476
rect 335542 278467 335856 278473
rect 335554 278448 335856 278467
rect 334390 278081 334442 278087
rect 334390 278023 334442 278029
rect 333142 274899 333194 274905
rect 333142 274841 333194 274847
rect 333154 265156 333182 274841
rect 333442 271501 333470 277870
rect 333334 271495 333386 271501
rect 333334 271437 333386 271443
rect 333430 271495 333482 271501
rect 333430 271437 333482 271443
rect 333346 271131 333374 271437
rect 333334 271125 333386 271131
rect 333334 271067 333386 271073
rect 333910 267129 333962 267135
rect 333910 267071 333962 267077
rect 332386 265128 332640 265156
rect 332770 265128 333024 265156
rect 333154 265128 333456 265156
rect 333922 265142 333950 267071
rect 334402 265142 334430 278023
rect 334486 274677 334538 274683
rect 334486 274619 334538 274625
rect 334498 265156 334526 274619
rect 334594 273573 334622 277870
rect 335638 274233 335690 274239
rect 335638 274175 335690 274181
rect 334582 273567 334634 273573
rect 334582 273509 334634 273515
rect 334966 268683 335018 268689
rect 334966 268625 335018 268631
rect 334978 265156 335006 268625
rect 334498 265128 334752 265156
rect 334978 265128 335232 265156
rect 335650 265142 335678 274175
rect 336994 272019 337022 277870
rect 338242 276311 338270 277870
rect 339106 277856 339408 277884
rect 338806 277045 338858 277051
rect 338806 276987 338858 276993
rect 338230 276305 338282 276311
rect 338230 276247 338282 276253
rect 337942 274307 337994 274313
rect 337942 274249 337994 274255
rect 337078 274159 337130 274165
rect 337078 274101 337130 274107
rect 336982 272013 337034 272019
rect 336982 271955 337034 271961
rect 336694 271125 336746 271131
rect 336694 271067 336746 271073
rect 336884 271090 336940 271099
rect 336706 270613 336734 271067
rect 336884 271025 336886 271034
rect 336938 271025 336940 271034
rect 336886 270993 336938 270999
rect 336694 270607 336746 270613
rect 336694 270549 336746 270555
rect 336406 268979 336458 268985
rect 336406 268921 336458 268927
rect 336118 268017 336170 268023
rect 336214 268017 336266 268023
rect 336118 267959 336170 267965
rect 336212 267982 336214 267991
rect 336418 267991 336446 268921
rect 336502 268387 336554 268393
rect 336502 268329 336554 268335
rect 336266 267982 336268 267991
rect 336130 265142 336158 267959
rect 336212 267917 336268 267926
rect 336404 267982 336460 267991
rect 336404 267917 336460 267926
rect 336514 265142 336542 268329
rect 337090 265156 337118 274101
rect 337954 269744 337982 274249
rect 338708 270350 338764 270359
rect 338050 270308 338708 270336
rect 338050 269915 338078 270308
rect 338708 270285 338764 270294
rect 338036 269906 338092 269915
rect 338036 269841 338092 269850
rect 337954 269716 338078 269744
rect 337462 268313 337514 268319
rect 337462 268255 337514 268261
rect 337474 265452 337502 268255
rect 337846 268165 337898 268171
rect 337846 268107 337898 268113
rect 336960 265128 337118 265156
rect 337426 265424 337502 265452
rect 337426 265142 337454 265424
rect 337858 265142 337886 268107
rect 338050 265156 338078 269716
rect 338326 267499 338378 267505
rect 338326 267441 338378 267447
rect 338338 266617 338366 267441
rect 338326 266611 338378 266617
rect 338326 266553 338378 266559
rect 338818 265156 338846 276987
rect 338902 274011 338954 274017
rect 338902 273953 338954 273959
rect 338050 265128 338256 265156
rect 338736 265128 338846 265156
rect 338914 265156 338942 273953
rect 338998 270385 339050 270391
rect 338998 270327 339050 270333
rect 339010 270243 339038 270327
rect 338998 270237 339050 270243
rect 338998 270179 339050 270185
rect 339106 265729 339134 277856
rect 340642 273573 340670 277870
rect 341794 276237 341822 277870
rect 342754 277865 342960 277884
rect 342742 277859 342960 277865
rect 342794 277856 342960 277859
rect 342742 277801 342794 277807
rect 341782 276231 341834 276237
rect 341782 276173 341834 276179
rect 340630 273567 340682 273573
rect 340630 273509 340682 273515
rect 343510 273567 343562 273573
rect 343510 273509 343562 273515
rect 343030 272013 343082 272019
rect 343030 271955 343082 271961
rect 342646 271495 342698 271501
rect 342646 271437 342698 271443
rect 341974 271421 342026 271427
rect 341974 271363 342026 271369
rect 339382 271347 339434 271353
rect 339382 271289 339434 271295
rect 339188 270942 339244 270951
rect 339188 270877 339244 270886
rect 339202 270317 339230 270877
rect 339190 270311 339242 270317
rect 339190 270253 339242 270259
rect 339094 265723 339146 265729
rect 339094 265665 339146 265671
rect 339394 265156 339422 271289
rect 340918 271273 340970 271279
rect 340918 271215 340970 271221
rect 340438 270829 340490 270835
rect 340438 270771 340490 270777
rect 339862 270607 339914 270613
rect 339862 270549 339914 270555
rect 339874 265156 339902 270549
rect 338914 265128 339168 265156
rect 339394 265128 339648 265156
rect 339874 265128 340032 265156
rect 340450 265142 340478 270771
rect 340930 265142 340958 271215
rect 341494 270977 341546 270983
rect 341494 270919 341546 270925
rect 341506 265156 341534 270919
rect 341986 265156 342014 271363
rect 341506 265128 341760 265156
rect 341986 265128 342240 265156
rect 342658 265142 342686 271437
rect 342742 270829 342794 270835
rect 342742 270771 342794 270777
rect 342754 270095 342782 270771
rect 342742 270089 342794 270095
rect 342742 270031 342794 270037
rect 343042 265142 343070 271955
rect 343522 265142 343550 273509
rect 344194 265156 344222 277870
rect 344662 273567 344714 273573
rect 344662 273509 344714 273515
rect 344674 265156 344702 273509
rect 345346 271353 345374 277870
rect 346486 276305 346538 276311
rect 346486 276247 346538 276253
rect 345718 271495 345770 271501
rect 345718 271437 345770 271443
rect 345334 271347 345386 271353
rect 345334 271289 345386 271295
rect 345238 271199 345290 271205
rect 345238 271141 345290 271147
rect 344758 270977 344810 270983
rect 344758 270919 344810 270925
rect 343968 265128 344222 265156
rect 344448 265128 344702 265156
rect 344770 265142 344798 270919
rect 345250 265142 345278 271141
rect 345730 265142 345758 271437
rect 346390 271273 346442 271279
rect 346390 271215 346442 271221
rect 346402 265156 346430 271215
rect 346176 265128 346430 265156
rect 346498 265156 346526 276247
rect 346594 267431 346622 277870
rect 347746 273573 347774 277870
rect 348406 276231 348458 276237
rect 348406 276173 348458 276179
rect 347734 273567 347786 273573
rect 347734 273509 347786 273515
rect 347926 272013 347978 272019
rect 347926 271955 347978 271961
rect 347446 271421 347498 271427
rect 347446 271363 347498 271369
rect 347254 271347 347306 271353
rect 347254 271289 347306 271295
rect 346582 267425 346634 267431
rect 346582 267367 346634 267373
rect 347266 265156 347294 271289
rect 346498 265128 346560 265156
rect 346992 265128 347294 265156
rect 347458 265142 347486 271363
rect 347938 265142 347966 271955
rect 348310 270607 348362 270613
rect 348310 270549 348362 270555
rect 348322 270169 348350 270549
rect 348310 270163 348362 270169
rect 348310 270105 348362 270111
rect 348418 265156 348446 276173
rect 348692 272570 348748 272579
rect 348692 272505 348748 272514
rect 348706 271247 348734 272505
rect 348692 271238 348748 271247
rect 348692 271173 348748 271182
rect 348598 268683 348650 268689
rect 348598 268625 348650 268631
rect 348610 268097 348638 268625
rect 348598 268091 348650 268097
rect 348598 268033 348650 268039
rect 348802 265452 348830 278541
rect 348994 275941 349022 277870
rect 350050 276903 350078 277870
rect 350038 276897 350090 276903
rect 350038 276839 350090 276845
rect 349174 276749 349226 276755
rect 349174 276691 349226 276697
rect 348982 275935 349034 275941
rect 348982 275877 349034 275883
rect 348288 265128 348446 265156
rect 348754 265424 348830 265452
rect 348754 265142 348782 265424
rect 349186 265142 349214 276691
rect 350338 265156 350366 278541
rect 364162 278309 364464 278328
rect 364150 278303 364464 278309
rect 364202 278300 364464 278303
rect 365782 278303 365834 278309
rect 364150 278245 364202 278251
rect 365782 278245 365834 278251
rect 352918 278155 352970 278161
rect 352918 278097 352970 278103
rect 351094 276527 351146 276533
rect 351094 276469 351146 276475
rect 350710 265723 350762 265729
rect 350710 265665 350762 265671
rect 350722 265156 350750 265665
rect 351106 265156 351134 276469
rect 351298 270983 351326 277870
rect 352246 273937 352298 273943
rect 352246 273879 352298 273885
rect 351286 270977 351338 270983
rect 351286 270919 351338 270925
rect 351766 268979 351818 268985
rect 351766 268921 351818 268927
rect 351286 267129 351338 267135
rect 351286 267071 351338 267077
rect 350064 265128 350366 265156
rect 350496 265128 350750 265156
rect 350976 265128 351134 265156
rect 351298 265142 351326 267071
rect 351778 265142 351806 268921
rect 352258 265142 352286 273879
rect 352450 270391 352478 277870
rect 352726 270607 352778 270613
rect 352726 270549 352778 270555
rect 352438 270385 352490 270391
rect 352438 270327 352490 270333
rect 352738 270169 352766 270549
rect 352726 270163 352778 270169
rect 352726 270105 352778 270111
rect 352930 265156 352958 278097
rect 353494 278081 353546 278087
rect 353494 278023 353546 278029
rect 353302 267573 353354 267579
rect 353302 267515 353354 267521
rect 353314 265156 353342 267515
rect 352704 265128 352958 265156
rect 353088 265128 353342 265156
rect 353506 265142 353534 278023
rect 355510 278007 355562 278013
rect 355510 277949 355562 277955
rect 353698 267283 353726 277870
rect 354454 273715 354506 273721
rect 354454 273657 354506 273663
rect 353974 268313 354026 268319
rect 353974 268255 354026 268261
rect 353686 267277 353738 267283
rect 353686 267219 353738 267225
rect 353986 265142 354014 268255
rect 354466 265142 354494 273657
rect 354850 271205 354878 277870
rect 354838 271199 354890 271205
rect 354838 271141 354890 271147
rect 355030 267425 355082 267431
rect 355030 267367 355082 267373
rect 355042 265156 355070 267367
rect 355522 265156 355550 277949
rect 356950 277933 357002 277939
rect 356950 277875 357002 277881
rect 356098 275645 356126 277870
rect 356854 277859 356906 277865
rect 356854 277801 356906 277807
rect 356086 275639 356138 275645
rect 356086 275581 356138 275587
rect 356182 273863 356234 273869
rect 356182 273805 356234 273811
rect 355606 270385 355658 270391
rect 355606 270327 355658 270333
rect 355618 268245 355646 270327
rect 355606 268239 355658 268245
rect 355606 268181 355658 268187
rect 355702 268017 355754 268023
rect 355702 267959 355754 267965
rect 354816 265128 355070 265156
rect 355296 265128 355550 265156
rect 355714 265142 355742 267959
rect 356194 265142 356222 273805
rect 356866 272852 356894 277801
rect 356962 273573 356990 277875
rect 357058 277856 357264 277884
rect 357058 277791 357086 277856
rect 357046 277785 357098 277791
rect 357046 277727 357098 277733
rect 358294 274307 358346 274313
rect 358294 274249 358346 274255
rect 356950 273567 357002 273573
rect 356950 273509 357002 273515
rect 356866 272824 356990 272852
rect 356566 267277 356618 267283
rect 356566 267219 356618 267225
rect 356578 265142 356606 267219
rect 356962 265452 356990 272824
rect 357622 270237 357674 270243
rect 357622 270179 357674 270185
rect 357634 268467 357662 270179
rect 357622 268461 357674 268467
rect 357622 268403 357674 268409
rect 357718 268461 357770 268467
rect 357718 268403 357770 268409
rect 357238 268387 357290 268393
rect 357238 268329 357290 268335
rect 357250 267505 357278 268329
rect 357238 267499 357290 267505
rect 357238 267441 357290 267447
rect 357334 267499 357386 267505
rect 357334 267441 357386 267447
rect 357346 267135 357374 267441
rect 357334 267129 357386 267135
rect 357334 267071 357386 267077
rect 356962 265424 357038 265452
rect 357010 265142 357038 265424
rect 357730 265156 357758 268403
rect 357814 267129 357866 267135
rect 357814 267071 357866 267077
rect 357504 265128 357758 265156
rect 357826 265142 357854 267071
rect 358306 265142 358334 274249
rect 358402 271501 358430 277870
rect 358774 277785 358826 277791
rect 358774 277727 358826 277733
rect 358676 272422 358732 272431
rect 358676 272357 358732 272366
rect 358690 272135 358718 272357
rect 358676 272126 358732 272135
rect 358676 272061 358732 272070
rect 358486 272013 358538 272019
rect 358486 271955 358538 271961
rect 358498 271501 358526 271955
rect 358390 271495 358442 271501
rect 358390 271437 358442 271443
rect 358486 271495 358538 271501
rect 358486 271437 358538 271443
rect 358486 270607 358538 270613
rect 358486 270549 358538 270555
rect 358498 269577 358526 270549
rect 358486 269571 358538 269577
rect 358486 269513 358538 269519
rect 358582 269571 358634 269577
rect 358582 269513 358634 269519
rect 358594 268467 358622 269513
rect 358582 268461 358634 268467
rect 358582 268403 358634 268409
rect 358390 268239 358442 268245
rect 358390 268181 358442 268187
rect 358402 267875 358430 268181
rect 358390 267869 358442 267875
rect 358390 267811 358442 267817
rect 358786 265142 358814 277727
rect 359650 270835 359678 277870
rect 360502 274159 360554 274165
rect 360502 274101 360554 274107
rect 360022 274085 360074 274091
rect 360022 274027 360074 274033
rect 359638 270829 359690 270835
rect 359638 270771 359690 270777
rect 358870 268387 358922 268393
rect 358870 268329 358922 268335
rect 359446 268387 359498 268393
rect 359446 268329 359498 268335
rect 358882 267875 358910 268329
rect 358870 267869 358922 267875
rect 358870 267811 358922 267817
rect 359458 265156 359486 268329
rect 359830 266907 359882 266913
rect 359830 266849 359882 266855
rect 359842 265156 359870 266849
rect 359232 265128 359486 265156
rect 359616 265128 359870 265156
rect 360034 265142 360062 274027
rect 360514 265142 360542 274101
rect 360802 266617 360830 277870
rect 361558 276601 361610 276607
rect 361558 276543 361610 276549
rect 360982 268313 361034 268319
rect 360982 268255 361034 268261
rect 360790 266611 360842 266617
rect 360790 266553 360842 266559
rect 360994 265142 361022 268255
rect 361570 265156 361598 276543
rect 362050 271279 362078 277870
rect 363202 275423 363230 277870
rect 363766 277415 363818 277421
rect 363766 277357 363818 277363
rect 363190 275417 363242 275423
rect 363190 275359 363242 275365
rect 362038 271273 362090 271279
rect 362038 271215 362090 271221
rect 362038 270829 362090 270835
rect 362038 270771 362090 270777
rect 362050 265156 362078 270771
rect 363094 270089 363146 270095
rect 363094 270031 363146 270037
rect 362230 266611 362282 266617
rect 362230 266553 362282 266559
rect 361344 265128 361598 265156
rect 361824 265128 362078 265156
rect 362242 265142 362270 266553
rect 362710 266537 362762 266543
rect 362710 266479 362762 266485
rect 362722 265142 362750 266479
rect 363106 265142 363134 270031
rect 363778 265156 363806 277357
rect 364822 277045 364874 277051
rect 364822 276987 364874 276993
rect 364246 275639 364298 275645
rect 364246 275581 364298 275587
rect 363862 270977 363914 270983
rect 363862 270919 363914 270925
rect 363874 267357 363902 270919
rect 363862 267351 363914 267357
rect 363862 267293 363914 267299
rect 364258 265156 364286 275581
rect 364342 274233 364394 274239
rect 364342 274175 364394 274181
rect 363552 265128 363806 265156
rect 364032 265128 364286 265156
rect 364354 265142 364382 274175
rect 364834 265142 364862 276987
rect 365602 276311 365630 277870
rect 365794 276681 365822 278245
rect 366466 277856 366768 277884
rect 365782 276675 365834 276681
rect 365782 276617 365834 276623
rect 365590 276305 365642 276311
rect 365590 276247 365642 276253
rect 365878 273937 365930 273943
rect 365878 273879 365930 273885
rect 365110 273789 365162 273795
rect 365110 273731 365162 273737
rect 365206 273789 365258 273795
rect 365206 273731 365258 273737
rect 365122 271279 365150 273731
rect 365110 271273 365162 271279
rect 365110 271215 365162 271221
rect 365218 270835 365246 273731
rect 365890 273647 365918 273879
rect 365782 273641 365834 273647
rect 365782 273583 365834 273589
rect 365878 273641 365930 273647
rect 365878 273583 365930 273589
rect 365794 272019 365822 273583
rect 365782 272013 365834 272019
rect 365782 271955 365834 271961
rect 366166 271347 366218 271353
rect 366166 271289 366218 271295
rect 365206 270829 365258 270835
rect 365206 270771 365258 270777
rect 365302 270829 365354 270835
rect 365302 270771 365354 270777
rect 365314 265142 365342 270771
rect 366178 270243 366206 271289
rect 366166 270237 366218 270243
rect 366166 270179 366218 270185
rect 366466 269799 366494 277856
rect 366934 276749 366986 276755
rect 366934 276691 366986 276697
rect 367030 276749 367082 276755
rect 367030 276691 367082 276697
rect 366946 276533 366974 276691
rect 366934 276527 366986 276533
rect 366934 276469 366986 276475
rect 367042 270835 367070 276691
rect 367906 273573 367934 277870
rect 368578 275423 368606 278573
rect 380854 278599 380906 278605
rect 380714 278559 380854 278587
rect 380662 278541 380714 278547
rect 380854 278541 380906 278547
rect 381238 278599 381290 278605
rect 393826 278605 394128 278624
rect 383828 278573 383884 278582
rect 390262 278599 390314 278605
rect 381238 278541 381290 278547
rect 368852 278490 368908 278499
rect 368852 278425 368908 278434
rect 368866 278309 368894 278425
rect 380278 278377 380330 278383
rect 380662 278377 380714 278383
rect 380330 278337 380662 278365
rect 380278 278319 380330 278325
rect 380662 278319 380714 278325
rect 368854 278303 368906 278309
rect 368854 278245 368906 278251
rect 378262 278303 378314 278309
rect 378262 278245 378314 278251
rect 369622 278155 369674 278161
rect 369622 278097 369674 278103
rect 368566 275417 368618 275423
rect 368566 275359 368618 275365
rect 368086 274899 368138 274905
rect 368086 274841 368138 274847
rect 367894 273567 367946 273573
rect 367894 273509 367946 273515
rect 367030 270829 367082 270835
rect 367030 270771 367082 270777
rect 367126 270829 367178 270835
rect 367126 270771 367178 270777
rect 366454 269793 366506 269799
rect 366454 269735 366506 269741
rect 366550 269793 366602 269799
rect 366550 269735 366602 269741
rect 366358 268461 366410 268467
rect 366358 268403 366410 268409
rect 365974 266241 366026 266247
rect 365974 266183 366026 266189
rect 365986 265156 366014 266183
rect 366370 265156 366398 268403
rect 365760 265128 366014 265156
rect 366144 265128 366398 265156
rect 366562 265142 366590 269735
rect 367030 265945 367082 265951
rect 367030 265887 367082 265893
rect 367042 265142 367070 265887
rect 367138 265137 367166 270771
rect 367510 270237 367562 270243
rect 367510 270179 367562 270185
rect 367522 265142 367550 270179
rect 368098 265156 368126 274841
rect 369044 271978 369100 271987
rect 369044 271913 369100 271922
rect 369058 271099 369086 271913
rect 369154 271205 369182 277870
rect 369526 275935 369578 275941
rect 369526 275877 369578 275883
rect 369142 271199 369194 271205
rect 369142 271141 369194 271147
rect 369238 271199 369290 271205
rect 369238 271141 369290 271147
rect 369044 271090 369100 271099
rect 369044 271025 369100 271034
rect 369250 270835 369278 271141
rect 369238 270829 369290 270835
rect 369238 270771 369290 270777
rect 368278 267499 368330 267505
rect 368278 267441 368330 267447
rect 368374 267499 368426 267505
rect 368374 267441 368426 267447
rect 368290 267357 368318 267441
rect 368278 267351 368330 267357
rect 368278 267293 368330 267299
rect 368386 265729 368414 267441
rect 368374 265723 368426 265729
rect 368374 265665 368426 265671
rect 368566 265723 368618 265729
rect 368566 265665 368618 265671
rect 368578 265156 368606 265665
rect 369334 265279 369386 265285
rect 369334 265221 369386 265227
rect 367126 265131 367178 265137
rect 367872 265128 368126 265156
rect 368352 265128 368606 265156
rect 369346 265137 369374 265221
rect 369334 265131 369386 265137
rect 367126 265073 367178 265079
rect 369334 265073 369386 265079
rect 369538 265008 369566 275877
rect 369634 265142 369662 278097
rect 370306 275349 370334 277870
rect 370294 275343 370346 275349
rect 370294 275285 370346 275291
rect 370966 274677 371018 274683
rect 370966 274619 371018 274625
rect 370294 273937 370346 273943
rect 370294 273879 370346 273885
rect 369718 265353 369770 265359
rect 369718 265295 369770 265301
rect 341026 264989 341328 265008
rect 326710 264983 326928 264989
rect 325750 264925 325802 264931
rect 326762 264980 326928 264983
rect 327286 264983 327338 264989
rect 326710 264925 326762 264931
rect 327286 264925 327338 264931
rect 329398 264983 329450 264989
rect 329398 264925 329450 264931
rect 329494 264983 329546 264989
rect 329494 264925 329546 264931
rect 341014 264983 341328 264989
rect 341066 264980 341328 264983
rect 369264 264980 369566 265008
rect 341014 264925 341066 264931
rect 369730 264915 369758 265295
rect 370306 265156 370334 273879
rect 370388 271682 370444 271691
rect 370388 271617 370444 271626
rect 370402 271353 370430 271617
rect 370390 271347 370442 271353
rect 370390 271289 370442 271295
rect 370486 271347 370538 271353
rect 370486 271289 370538 271295
rect 370498 270507 370526 271289
rect 370678 270829 370730 270835
rect 370678 270771 370730 270777
rect 370690 270613 370718 270771
rect 370678 270607 370730 270613
rect 370678 270549 370730 270555
rect 370774 270607 370826 270613
rect 370774 270549 370826 270555
rect 370484 270498 370540 270507
rect 370484 270433 370540 270442
rect 370676 270498 370732 270507
rect 370676 270433 370732 270442
rect 370690 265729 370718 270433
rect 370678 265723 370730 265729
rect 370678 265665 370730 265671
rect 370786 265156 370814 270549
rect 370868 270498 370924 270507
rect 370868 270433 370924 270442
rect 370882 268171 370910 270433
rect 370870 268165 370922 268171
rect 370870 268107 370922 268113
rect 370080 265128 370334 265156
rect 370560 265128 370814 265156
rect 370978 265142 371006 274619
rect 371554 270983 371582 277870
rect 372034 276487 372254 276515
rect 372034 276459 372062 276487
rect 372022 276453 372074 276459
rect 372022 276395 372074 276401
rect 372118 276453 372170 276459
rect 372118 276395 372170 276401
rect 371542 270977 371594 270983
rect 371542 270919 371594 270925
rect 371444 270498 371500 270507
rect 371732 270498 371788 270507
rect 371444 270433 371500 270442
rect 371554 270456 371732 270484
rect 371458 270021 371486 270433
rect 371446 270015 371498 270021
rect 371446 269957 371498 269963
rect 371554 269892 371582 270456
rect 371732 270433 371788 270442
rect 371266 269864 371582 269892
rect 371266 269027 371294 269864
rect 371252 269018 371308 269027
rect 371252 268953 371308 268962
rect 371444 269018 371500 269027
rect 371444 268953 371500 268962
rect 371458 268837 371486 268953
rect 371446 268831 371498 268837
rect 371446 268773 371498 268779
rect 371542 268831 371594 268837
rect 371542 268773 371594 268779
rect 371554 268708 371582 268773
rect 371074 268680 371582 268708
rect 371074 268541 371102 268680
rect 371062 268535 371114 268541
rect 371062 268477 371114 268483
rect 371350 268535 371402 268541
rect 371350 268477 371402 268483
rect 371362 265142 371390 268477
rect 371542 268091 371594 268097
rect 371542 268033 371594 268039
rect 371638 268091 371690 268097
rect 371638 268033 371690 268039
rect 371554 264915 371582 268033
rect 371650 267875 371678 268033
rect 371638 267869 371690 267875
rect 371638 267811 371690 267817
rect 372130 265156 372158 276395
rect 372226 276311 372254 276487
rect 372214 276305 372266 276311
rect 372214 276247 372266 276253
rect 372598 275343 372650 275349
rect 372598 275285 372650 275291
rect 372610 274387 372638 275285
rect 372598 274381 372650 274387
rect 372598 274323 372650 274329
rect 372706 271427 372734 277870
rect 373570 277856 373872 277884
rect 372982 275417 373034 275423
rect 372982 275359 373034 275365
rect 372790 274455 372842 274461
rect 372790 274397 372842 274403
rect 372886 274455 372938 274461
rect 372886 274397 372938 274403
rect 372802 272135 372830 274397
rect 372788 272126 372844 272135
rect 372788 272061 372844 272070
rect 372694 271421 372746 271427
rect 372694 271363 372746 271369
rect 372502 268165 372554 268171
rect 372502 268107 372554 268113
rect 372514 265156 372542 268107
rect 372898 265156 372926 274397
rect 372994 274387 373022 275359
rect 373364 274938 373420 274947
rect 373364 274873 373420 274882
rect 372982 274381 373034 274387
rect 372982 274323 373034 274329
rect 372980 273606 373036 273615
rect 372980 273541 373036 273550
rect 373172 273606 373228 273615
rect 373172 273541 373228 273550
rect 372994 270951 373022 273541
rect 373186 273023 373214 273541
rect 373378 273023 373406 274873
rect 373172 273014 373228 273023
rect 373172 272949 373228 272958
rect 373364 273014 373420 273023
rect 373364 272949 373420 272958
rect 373462 270977 373514 270983
rect 372980 270942 373036 270951
rect 373462 270919 373514 270925
rect 372980 270877 373036 270886
rect 373474 270613 373502 270919
rect 373570 270835 373598 277856
rect 375106 277495 375134 277870
rect 375094 277489 375146 277495
rect 375094 277431 375146 277437
rect 375190 277489 375242 277495
rect 375190 277431 375242 277437
rect 374132 276418 374188 276427
rect 374132 276353 374188 276362
rect 374324 276418 374380 276427
rect 374324 276353 374380 276362
rect 374146 273573 374174 276353
rect 374338 274017 374366 276353
rect 375202 274683 375230 277431
rect 375574 275417 375626 275423
rect 375574 275359 375626 275365
rect 375190 274677 375242 274683
rect 375190 274619 375242 274625
rect 374326 274011 374378 274017
rect 374326 273953 374378 273959
rect 374134 273567 374186 273573
rect 374134 273509 374186 273515
rect 374422 271495 374474 271501
rect 374422 271437 374474 271443
rect 374710 271495 374762 271501
rect 374710 271437 374762 271443
rect 374038 271421 374090 271427
rect 373844 271386 373900 271395
rect 374038 271363 374090 271369
rect 373844 271321 373900 271330
rect 373654 271199 373706 271205
rect 373654 271141 373706 271147
rect 373666 270835 373694 271141
rect 373558 270829 373610 270835
rect 373558 270771 373610 270777
rect 373654 270829 373706 270835
rect 373654 270771 373706 270777
rect 373462 270607 373514 270613
rect 373462 270549 373514 270555
rect 373558 270607 373610 270613
rect 373558 270549 373610 270555
rect 372994 268837 373214 268856
rect 372982 268831 373214 268837
rect 373034 268828 373214 268831
rect 372982 268773 373034 268779
rect 373186 268689 373214 268828
rect 373366 268831 373418 268837
rect 373366 268773 373418 268779
rect 373078 268683 373130 268689
rect 373078 268625 373130 268631
rect 373174 268683 373226 268689
rect 373174 268625 373226 268631
rect 372982 268609 373034 268615
rect 372982 268551 373034 268557
rect 373090 268560 373118 268625
rect 372994 267875 373022 268551
rect 373090 268541 373214 268560
rect 373090 268535 373226 268541
rect 373090 268532 373174 268535
rect 373174 268477 373226 268483
rect 372982 267869 373034 267875
rect 372982 267811 373034 267817
rect 373378 265156 373406 268773
rect 371856 265128 372158 265156
rect 372288 265128 372542 265156
rect 372672 265128 372926 265156
rect 373152 265128 373406 265156
rect 373570 265142 373598 270549
rect 373858 270391 373886 271321
rect 373846 270385 373898 270391
rect 373846 270327 373898 270333
rect 374050 265142 374078 271363
rect 374434 271205 374462 271437
rect 374422 271199 374474 271205
rect 374422 271141 374474 271147
rect 374722 265156 374750 271437
rect 375094 270385 375146 270391
rect 375094 270327 375146 270333
rect 375106 265156 375134 270327
rect 375586 265156 375614 275359
rect 375958 274677 376010 274683
rect 375958 274619 376010 274625
rect 375670 273937 375722 273943
rect 375670 273879 375722 273885
rect 375682 273467 375710 273879
rect 375668 273458 375724 273467
rect 375668 273393 375724 273402
rect 375860 273458 375916 273467
rect 375860 273393 375916 273402
rect 375874 272875 375902 273393
rect 375860 272866 375916 272875
rect 375860 272801 375916 272810
rect 375766 270015 375818 270021
rect 375766 269957 375818 269963
rect 374448 265128 374750 265156
rect 374880 265128 375134 265156
rect 375360 265128 375614 265156
rect 375778 265142 375806 269957
rect 375970 265211 375998 274619
rect 376148 272718 376204 272727
rect 376148 272653 376204 272662
rect 376162 270835 376190 272653
rect 376258 271205 376286 277870
rect 376630 276897 376682 276903
rect 376630 276839 376682 276845
rect 376340 272126 376396 272135
rect 376340 272061 376396 272070
rect 376354 271205 376382 272061
rect 376246 271199 376298 271205
rect 376246 271141 376298 271147
rect 376342 271199 376394 271205
rect 376342 271141 376394 271147
rect 376150 270829 376202 270835
rect 376150 270771 376202 270777
rect 376054 267721 376106 267727
rect 376054 267663 376106 267669
rect 376066 265211 376094 267663
rect 375958 265205 376010 265211
rect 375958 265147 376010 265153
rect 376054 265205 376106 265211
rect 376054 265147 376106 265153
rect 376642 265142 376670 276839
rect 377506 275127 377534 277870
rect 378274 277019 378302 278245
rect 380194 278161 380702 278180
rect 380182 278155 380714 278161
rect 380234 278152 380662 278155
rect 380182 278097 380234 278103
rect 380662 278097 380714 278103
rect 378370 277856 378672 277884
rect 378260 277010 378316 277019
rect 378260 276945 378316 276954
rect 377494 275121 377546 275127
rect 377494 275063 377546 275069
rect 377686 275121 377738 275127
rect 377686 275063 377738 275069
rect 377300 273162 377356 273171
rect 377300 273097 377356 273106
rect 377314 272135 377342 273097
rect 377300 272126 377356 272135
rect 377300 272061 377356 272070
rect 377590 270829 377642 270835
rect 377590 270771 377642 270777
rect 377014 268683 377066 268689
rect 377014 268625 377066 268631
rect 377110 268683 377162 268689
rect 377110 268625 377162 268631
rect 377026 268116 377054 268625
rect 377122 268467 377150 268625
rect 377110 268461 377162 268467
rect 377110 268403 377162 268409
rect 377206 268461 377258 268467
rect 377206 268403 377258 268409
rect 377108 268278 377164 268287
rect 377218 268264 377246 268403
rect 377164 268236 377246 268264
rect 377108 268213 377164 268222
rect 377026 268088 377534 268116
rect 377218 267903 377438 267931
rect 377218 267653 377246 267903
rect 377302 267869 377354 267875
rect 377410 267843 377438 267903
rect 377506 267875 377534 268088
rect 377494 267869 377546 267875
rect 377302 267811 377354 267817
rect 377396 267834 377452 267843
rect 377314 267653 377342 267811
rect 377494 267811 377546 267817
rect 377396 267769 377452 267778
rect 377206 267647 377258 267653
rect 377206 267589 377258 267595
rect 377302 267647 377354 267653
rect 377302 267589 377354 267595
rect 377206 265649 377258 265655
rect 377206 265591 377258 265597
rect 377218 265156 377246 265591
rect 377602 265304 377630 270771
rect 377698 267505 377726 275063
rect 378068 274938 378124 274947
rect 378068 274873 378124 274882
rect 378082 273763 378110 274873
rect 378370 274683 378398 277856
rect 378742 277415 378794 277421
rect 378742 277357 378794 277363
rect 378838 277415 378890 277421
rect 379906 277403 379934 277870
rect 380578 277856 381072 277884
rect 379906 277375 380030 277403
rect 378838 277357 378890 277363
rect 378754 277051 378782 277357
rect 378646 277045 378698 277051
rect 378452 277010 378508 277019
rect 378646 276987 378698 276993
rect 378742 277045 378794 277051
rect 378742 276987 378794 276993
rect 378452 276945 378508 276954
rect 378466 276459 378494 276945
rect 378658 276903 378686 276987
rect 378550 276897 378602 276903
rect 378550 276839 378602 276845
rect 378646 276897 378698 276903
rect 378646 276839 378698 276845
rect 378562 276552 378590 276839
rect 378850 276681 378878 277357
rect 378838 276675 378890 276681
rect 378838 276617 378890 276623
rect 378934 276675 378986 276681
rect 378934 276617 378986 276623
rect 378946 276552 378974 276617
rect 378562 276524 378974 276552
rect 379030 276601 379082 276607
rect 380002 276552 380030 277375
rect 379030 276543 379082 276549
rect 379042 276459 379070 276543
rect 379906 276524 380030 276552
rect 378454 276453 378506 276459
rect 378454 276395 378506 276401
rect 379030 276453 379082 276459
rect 379030 276395 379082 276401
rect 379606 276453 379658 276459
rect 379606 276395 379658 276401
rect 378754 275784 379070 275812
rect 378754 275645 378782 275784
rect 378742 275639 378794 275645
rect 378742 275581 378794 275587
rect 378838 275639 378890 275645
rect 378838 275581 378890 275587
rect 378850 275423 378878 275581
rect 378838 275417 378890 275423
rect 378838 275359 378890 275365
rect 378934 275417 378986 275423
rect 378934 275359 378986 275365
rect 378946 275072 378974 275359
rect 378466 275044 378782 275072
rect 378358 274677 378410 274683
rect 378358 274619 378410 274625
rect 378466 273888 378494 275044
rect 378754 274905 378782 275044
rect 378850 275044 378974 275072
rect 378646 274899 378698 274905
rect 378646 274841 378698 274847
rect 378742 274899 378794 274905
rect 378742 274841 378794 274847
rect 378658 274683 378686 274841
rect 378646 274677 378698 274683
rect 378646 274619 378698 274625
rect 378850 274480 378878 275044
rect 378658 274461 378878 274480
rect 379042 274461 379070 275784
rect 378646 274455 378878 274461
rect 378698 274452 378878 274455
rect 379030 274455 379082 274461
rect 378646 274397 378698 274403
rect 379030 274397 379082 274403
rect 378646 274307 378698 274313
rect 378646 274249 378698 274255
rect 378742 274307 378794 274313
rect 378742 274249 378794 274255
rect 378658 274017 378686 274249
rect 378550 274011 378602 274017
rect 378550 273953 378602 273959
rect 378646 274011 378698 274017
rect 378646 273953 378698 273959
rect 378178 273860 378494 273888
rect 378562 273888 378590 273953
rect 378754 273888 378782 274249
rect 378562 273860 378782 273888
rect 378068 273754 378124 273763
rect 378068 273689 378124 273698
rect 378178 273629 378206 273860
rect 378260 273754 378316 273763
rect 378260 273689 378316 273698
rect 377890 273601 378206 273629
rect 377782 267943 377834 267949
rect 377782 267885 377834 267891
rect 377794 267505 377822 267885
rect 377686 267499 377738 267505
rect 377686 267441 377738 267447
rect 377782 267499 377834 267505
rect 377782 267441 377834 267447
rect 377088 265128 377246 265156
rect 377506 265276 377630 265304
rect 376438 265057 376490 265063
rect 376176 265005 376438 265008
rect 376176 264999 376490 265005
rect 377506 265008 377534 265276
rect 377890 265142 377918 273601
rect 378070 273567 378122 273573
rect 378070 273509 378122 273515
rect 378082 273171 378110 273509
rect 378068 273162 378124 273171
rect 377974 273123 378026 273129
rect 378068 273097 378124 273106
rect 377974 273065 378026 273071
rect 377986 271076 378014 273065
rect 378274 272907 378302 273689
rect 378358 273567 378410 273573
rect 378358 273509 378410 273515
rect 378262 272901 378314 272907
rect 378262 272843 378314 272849
rect 378370 272611 378398 273509
rect 378454 273197 378506 273203
rect 378454 273139 378506 273145
rect 378466 272704 378494 273139
rect 378742 273049 378794 273055
rect 378658 272997 378742 273000
rect 378658 272991 378794 272997
rect 378658 272972 378782 272991
rect 378658 272907 378686 272972
rect 378646 272901 378698 272907
rect 378646 272843 378698 272849
rect 378934 272901 378986 272907
rect 378934 272843 378986 272849
rect 378838 272827 378890 272833
rect 378838 272769 378890 272775
rect 378466 272685 378782 272704
rect 378466 272679 378794 272685
rect 378466 272676 378742 272679
rect 378742 272621 378794 272627
rect 378358 272605 378410 272611
rect 378358 272547 378410 272553
rect 378550 272605 378602 272611
rect 378550 272547 378602 272553
rect 378562 272315 378590 272547
rect 378550 272309 378602 272315
rect 378550 272251 378602 272257
rect 378742 272235 378794 272241
rect 378082 272195 378742 272223
rect 378082 271205 378110 272195
rect 378742 272177 378794 272183
rect 378070 271199 378122 271205
rect 378070 271141 378122 271147
rect 378166 271199 378218 271205
rect 378166 271141 378218 271147
rect 378178 271076 378206 271141
rect 377986 271048 378206 271076
rect 378370 271048 378686 271076
rect 378370 270951 378398 271048
rect 378356 270942 378412 270951
rect 378356 270877 378412 270886
rect 378548 270942 378604 270951
rect 378548 270877 378604 270886
rect 378562 270507 378590 270877
rect 378658 270632 378686 271048
rect 378850 270835 378878 272769
rect 378946 272241 378974 272843
rect 378934 272235 378986 272241
rect 378934 272177 378986 272183
rect 378838 270829 378890 270835
rect 378838 270771 378890 270777
rect 378934 270829 378986 270835
rect 378934 270771 378986 270777
rect 378946 270632 378974 270771
rect 378658 270604 378974 270632
rect 379126 270607 379178 270613
rect 379126 270549 379178 270555
rect 378548 270498 378604 270507
rect 378548 270433 378604 270442
rect 378836 270498 378892 270507
rect 378836 270433 378892 270442
rect 378850 270336 378878 270433
rect 378562 270308 378878 270336
rect 379030 270385 379082 270391
rect 379030 270327 379082 270333
rect 378358 268979 378410 268985
rect 378358 268921 378410 268927
rect 378370 267949 378398 268921
rect 378562 268615 378590 270308
rect 378838 270237 378890 270243
rect 378838 270179 378890 270185
rect 378742 268979 378794 268985
rect 378742 268921 378794 268927
rect 378754 268837 378782 268921
rect 378742 268831 378794 268837
rect 378742 268773 378794 268779
rect 378850 268763 378878 270179
rect 378934 270089 378986 270095
rect 378934 270031 378986 270037
rect 378646 268757 378698 268763
rect 378646 268699 378698 268705
rect 378838 268757 378890 268763
rect 378838 268699 378890 268705
rect 378658 268615 378686 268699
rect 378550 268609 378602 268615
rect 378550 268551 378602 268557
rect 378646 268609 378698 268615
rect 378646 268551 378698 268557
rect 378562 268421 378878 268449
rect 378562 268171 378590 268421
rect 378646 268387 378698 268393
rect 378646 268329 378698 268335
rect 378658 268171 378686 268329
rect 378850 268264 378878 268421
rect 378946 268393 378974 270031
rect 379042 269892 379070 270327
rect 379138 270095 379166 270549
rect 379220 270498 379276 270507
rect 379220 270433 379276 270442
rect 379412 270498 379468 270507
rect 379412 270433 379468 270442
rect 379234 270391 379262 270433
rect 379222 270385 379274 270391
rect 379222 270327 379274 270333
rect 379318 270237 379370 270243
rect 379234 270197 379318 270225
rect 379126 270089 379178 270095
rect 379126 270031 379178 270037
rect 379042 269864 379166 269892
rect 379138 269799 379166 269864
rect 379030 269793 379082 269799
rect 379030 269735 379082 269741
rect 379126 269793 379178 269799
rect 379126 269735 379178 269741
rect 379042 268837 379070 269735
rect 379030 268831 379082 268837
rect 379030 268773 379082 268779
rect 378934 268387 378986 268393
rect 378934 268329 378986 268335
rect 379234 268264 379262 270197
rect 379318 270179 379370 270185
rect 378850 268236 379262 268264
rect 378550 268165 378602 268171
rect 378550 268107 378602 268113
rect 378646 268165 378698 268171
rect 378646 268107 378698 268113
rect 379426 268079 379454 270433
rect 378754 268051 379454 268079
rect 378358 267943 378410 267949
rect 378358 267885 378410 267891
rect 378454 267869 378506 267875
rect 378754 267820 378782 268051
rect 379318 267943 379370 267949
rect 379318 267885 379370 267891
rect 378454 267811 378506 267817
rect 378466 267727 378494 267811
rect 378562 267792 378782 267820
rect 378454 267721 378506 267727
rect 378454 267663 378506 267669
rect 378358 265427 378410 265433
rect 378178 265387 378358 265415
rect 378178 265359 378206 265387
rect 378358 265369 378410 265375
rect 378166 265353 378218 265359
rect 378166 265295 378218 265301
rect 378562 265156 378590 267792
rect 379330 267727 379358 267885
rect 379318 267721 379370 267727
rect 378658 267681 379262 267709
rect 378658 267357 378686 267681
rect 379234 267635 379262 267681
rect 379318 267663 379370 267669
rect 379414 267721 379466 267727
rect 379414 267663 379466 267669
rect 379426 267635 379454 267663
rect 378754 267607 379070 267635
rect 379234 267607 379454 267635
rect 378646 267351 378698 267357
rect 378646 267293 378698 267299
rect 378754 267061 378782 267607
rect 379042 267505 379070 267607
rect 378934 267499 378986 267505
rect 378934 267441 378986 267447
rect 379030 267499 379082 267505
rect 379030 267441 379082 267447
rect 378946 267080 378974 267441
rect 379510 267351 379562 267357
rect 379042 267311 379510 267339
rect 379042 267209 379070 267311
rect 379510 267293 379562 267299
rect 379618 267228 379646 276395
rect 379906 276237 379934 276524
rect 379894 276231 379946 276237
rect 379894 276173 379946 276179
rect 379990 276231 380042 276237
rect 379990 276173 380042 276179
rect 380002 275423 380030 276173
rect 379990 275417 380042 275423
rect 379990 275359 380042 275365
rect 380374 272679 380426 272685
rect 380374 272621 380426 272627
rect 380386 272537 380414 272621
rect 380278 272531 380330 272537
rect 380278 272473 380330 272479
rect 380374 272531 380426 272537
rect 380374 272473 380426 272479
rect 379990 272235 380042 272241
rect 379990 272177 380042 272183
rect 380002 272135 380030 272177
rect 379988 272126 380044 272135
rect 379988 272061 380044 272070
rect 380180 272126 380236 272135
rect 380180 272061 380236 272070
rect 380194 272019 380222 272061
rect 380290 272019 380318 272473
rect 380182 272013 380234 272019
rect 380182 271955 380234 271961
rect 380278 272013 380330 272019
rect 380278 271955 380330 271961
rect 380578 271691 380606 277856
rect 380950 275417 381002 275423
rect 380950 275359 381002 275365
rect 380758 272901 380810 272907
rect 380758 272843 380810 272849
rect 380854 272901 380906 272907
rect 380854 272843 380906 272849
rect 380770 272685 380798 272843
rect 380758 272679 380810 272685
rect 380758 272621 380810 272627
rect 380564 271682 380620 271691
rect 380564 271617 380620 271626
rect 379798 270607 379850 270613
rect 379798 270549 379850 270555
rect 379810 269027 379838 270549
rect 379796 269018 379852 269027
rect 379796 268953 379852 268962
rect 379988 269018 380044 269027
rect 379988 268953 380044 268962
rect 380276 269018 380332 269027
rect 380276 268953 380332 268962
rect 379030 267203 379082 267209
rect 379030 267145 379082 267151
rect 379126 267203 379178 267209
rect 379126 267145 379178 267151
rect 379330 267200 379646 267228
rect 378742 267055 378794 267061
rect 378742 266997 378794 267003
rect 378838 267055 378890 267061
rect 378946 267052 379070 267080
rect 378838 266997 378890 267003
rect 378850 265951 378878 266997
rect 378838 265945 378890 265951
rect 378838 265887 378890 265893
rect 378934 265945 378986 265951
rect 378934 265887 378986 265893
rect 378946 265655 378974 265887
rect 379042 265655 379070 267052
rect 378934 265649 378986 265655
rect 378934 265591 378986 265597
rect 379030 265649 379082 265655
rect 379030 265591 379082 265597
rect 378934 265501 378986 265507
rect 378754 265461 378934 265489
rect 378754 265433 378782 265461
rect 378934 265443 378986 265449
rect 378742 265427 378794 265433
rect 378742 265369 378794 265375
rect 379138 265156 379166 267145
rect 379330 265452 379358 267200
rect 380002 265711 380030 268953
rect 378384 265128 378590 265156
rect 378864 265128 379166 265156
rect 379282 265424 379358 265452
rect 379426 265683 380030 265711
rect 379282 265142 379310 265424
rect 379426 265285 379454 265683
rect 379894 265501 379946 265507
rect 379522 265461 379894 265489
rect 379414 265279 379466 265285
rect 379414 265221 379466 265227
rect 379522 265211 379550 265461
rect 379894 265443 379946 265449
rect 379702 265427 379754 265433
rect 379990 265427 380042 265433
rect 379754 265387 379990 265415
rect 379702 265369 379754 265375
rect 379990 265369 380042 265375
rect 379606 265353 379658 265359
rect 380182 265353 380234 265359
rect 379658 265313 380182 265341
rect 379606 265295 379658 265301
rect 380182 265295 380234 265301
rect 379990 265279 380042 265285
rect 379810 265239 379990 265267
rect 379510 265205 379562 265211
rect 379810 265156 379838 265239
rect 379990 265221 380042 265227
rect 380290 265156 380318 268953
rect 380866 265156 380894 272843
rect 379510 265147 379562 265153
rect 379680 265128 379838 265156
rect 380112 265128 380318 265156
rect 380592 265128 380894 265156
rect 380962 265142 380990 275359
rect 381250 272519 381278 278541
rect 383062 278525 383114 278531
rect 383114 278473 383376 278476
rect 383062 278467 383376 278473
rect 383074 278448 383376 278467
rect 381910 278377 381962 278383
rect 381962 278325 382320 278328
rect 381910 278319 382320 278325
rect 381922 278300 382320 278319
rect 382402 277116 383198 277144
rect 381622 274381 381674 274387
rect 381622 274323 381674 274329
rect 381634 272685 381662 274323
rect 382402 273795 382430 277116
rect 383060 277010 383116 277019
rect 383170 276996 383198 277116
rect 383252 277010 383308 277019
rect 383170 276968 383252 276996
rect 383060 276945 383116 276954
rect 383252 276945 383308 276954
rect 383074 276311 383102 276945
rect 382966 276305 383018 276311
rect 382966 276247 383018 276253
rect 383062 276305 383114 276311
rect 383062 276247 383114 276253
rect 382978 275072 383006 276247
rect 382978 275044 383294 275072
rect 383266 274947 383294 275044
rect 382676 274938 382732 274947
rect 382676 274873 382732 274882
rect 383252 274938 383308 274947
rect 383252 274873 383308 274882
rect 382390 273789 382442 273795
rect 382390 273731 382442 273737
rect 382486 273789 382538 273795
rect 382486 273731 382538 273737
rect 382196 273606 382252 273615
rect 382196 273541 382252 273550
rect 381334 272679 381386 272685
rect 381334 272621 381386 272627
rect 381622 272679 381674 272685
rect 381622 272621 381674 272627
rect 381154 272491 381278 272519
rect 381154 265211 381182 272491
rect 381236 272422 381292 272431
rect 381236 272357 381292 272366
rect 381142 265205 381194 265211
rect 381142 265147 381194 265153
rect 381250 265156 381278 272357
rect 381346 271691 381374 272621
rect 382210 272579 382238 273541
rect 382004 272570 382060 272579
rect 382004 272505 382060 272514
rect 382196 272570 382252 272579
rect 382196 272505 382252 272514
rect 381428 272422 381484 272431
rect 381428 272357 381484 272366
rect 381442 272241 381470 272357
rect 381430 272235 381482 272241
rect 381430 272177 381482 272183
rect 381526 272235 381578 272241
rect 381526 272177 381578 272183
rect 381332 271682 381388 271691
rect 381332 271617 381388 271626
rect 381538 271279 381566 272177
rect 381526 271273 381578 271279
rect 381910 271273 381962 271279
rect 381526 271215 381578 271221
rect 381620 271238 381676 271247
rect 381620 271173 381676 271182
rect 381908 271238 381910 271247
rect 381962 271238 381964 271247
rect 381908 271173 381964 271182
rect 381634 265156 381662 271173
rect 382018 265156 382046 272505
rect 382498 272241 382526 273731
rect 382690 272241 382718 274873
rect 382774 274381 382826 274387
rect 382774 274323 382826 274329
rect 382486 272235 382538 272241
rect 382486 272177 382538 272183
rect 382678 272235 382730 272241
rect 382678 272177 382730 272183
rect 382390 268535 382442 268541
rect 382390 268477 382442 268483
rect 382486 268535 382538 268541
rect 382486 268477 382538 268483
rect 382402 265156 382430 268477
rect 382498 267653 382526 268477
rect 382486 267647 382538 267653
rect 382486 267589 382538 267595
rect 382786 267505 382814 274323
rect 383542 274307 383594 274313
rect 383542 274249 383594 274255
rect 382882 274008 383294 274036
rect 382882 271691 382910 274008
rect 382964 273902 383020 273911
rect 382964 273837 383020 273846
rect 382978 273615 383006 273837
rect 383266 273795 383294 274008
rect 383554 273943 383582 274249
rect 383446 273937 383498 273943
rect 383446 273879 383498 273885
rect 383542 273937 383594 273943
rect 383542 273879 383594 273885
rect 383158 273789 383210 273795
rect 383158 273731 383210 273737
rect 383254 273789 383306 273795
rect 383254 273731 383306 273737
rect 382964 273606 383020 273615
rect 382964 273541 383020 273550
rect 382868 271682 382924 271691
rect 382868 271617 382924 271626
rect 383060 271682 383116 271691
rect 383060 271617 383116 271626
rect 383074 271057 383102 271617
rect 383170 271057 383198 273731
rect 383348 272866 383404 272875
rect 383348 272801 383404 272810
rect 383252 272274 383308 272283
rect 383252 272209 383308 272218
rect 383062 271051 383114 271057
rect 383062 270993 383114 270999
rect 383158 271051 383210 271057
rect 383158 270993 383210 270999
rect 383062 267647 383114 267653
rect 383062 267589 383114 267595
rect 382774 267499 382826 267505
rect 382774 267441 382826 267447
rect 383074 267357 383102 267589
rect 383062 267351 383114 267357
rect 383062 267293 383114 267299
rect 383266 265156 383294 272209
rect 381250 265128 381408 265156
rect 381634 265128 381888 265156
rect 382018 265128 382320 265156
rect 382402 265128 382704 265156
rect 383184 265128 383294 265156
rect 383362 265156 383390 272801
rect 383458 271247 383486 273879
rect 383444 271238 383500 271247
rect 383444 271173 383500 271182
rect 383842 265156 383870 278573
rect 390262 278541 390314 278547
rect 393814 278599 394128 278605
rect 393866 278596 394128 278599
rect 393814 278541 393866 278547
rect 389014 278377 389066 278383
rect 389066 278325 389328 278328
rect 389014 278319 389328 278325
rect 387766 278303 387818 278309
rect 389026 278300 389328 278319
rect 387766 278245 387818 278251
rect 384610 275349 384638 277870
rect 385474 277856 385776 277884
rect 385174 277489 385226 277495
rect 385174 277431 385226 277437
rect 385186 276311 385214 277431
rect 385174 276305 385226 276311
rect 385174 276247 385226 276253
rect 384982 276231 385034 276237
rect 384982 276173 385034 276179
rect 384994 275941 385022 276173
rect 384886 275935 384938 275941
rect 384886 275877 384938 275883
rect 384982 275935 385034 275941
rect 384982 275877 385034 275883
rect 384790 275417 384842 275423
rect 384790 275359 384842 275365
rect 384598 275343 384650 275349
rect 384598 275285 384650 275291
rect 384802 274905 384830 275359
rect 384898 274905 384926 275877
rect 384790 274899 384842 274905
rect 384790 274841 384842 274847
rect 384886 274899 384938 274905
rect 384886 274841 384938 274847
rect 385078 274307 385130 274313
rect 385078 274249 385130 274255
rect 384404 273458 384460 273467
rect 384404 273393 384460 273402
rect 383362 265128 383616 265156
rect 383842 265128 384096 265156
rect 384418 265142 384446 273393
rect 384884 272570 384940 272579
rect 384884 272505 384940 272514
rect 384898 265142 384926 272505
rect 378946 265017 379166 265045
rect 376176 264980 376478 264999
rect 377506 264980 377568 265008
rect 378946 264920 378974 265017
rect 379138 264989 379166 265017
rect 379030 264983 379082 264989
rect 379030 264925 379082 264931
rect 379126 264983 379178 264989
rect 379126 264925 379178 264931
rect 349846 264909 349898 264915
rect 324898 264832 325200 264860
rect 349584 264857 349846 264860
rect 369046 264909 369098 264915
rect 349584 264851 349898 264857
rect 368784 264857 369046 264860
rect 368784 264851 369098 264857
rect 369718 264909 369770 264915
rect 369718 264851 369770 264857
rect 371542 264909 371594 264915
rect 371542 264851 371594 264857
rect 378932 264911 378988 264920
rect 349584 264832 349886 264851
rect 368784 264832 369086 264851
rect 378932 264846 378988 264855
rect 379042 264860 379070 264925
rect 385090 264920 385118 274249
rect 385364 273458 385420 273467
rect 385364 273393 385420 273402
rect 385378 265142 385406 273393
rect 385474 267653 385502 277856
rect 387010 276607 387038 277870
rect 386998 276601 387050 276607
rect 386998 276543 387050 276549
rect 387668 273014 387724 273023
rect 387668 272949 387724 272958
rect 387572 272866 387628 272875
rect 387572 272801 387628 272810
rect 387586 272759 387614 272801
rect 387574 272753 387626 272759
rect 387574 272695 387626 272701
rect 386422 272679 386474 272685
rect 386422 272621 386474 272627
rect 386518 272679 386570 272685
rect 386518 272621 386570 272627
rect 385940 272422 385996 272431
rect 385940 272357 385996 272366
rect 385556 271238 385612 271247
rect 385556 271173 385612 271182
rect 385462 267647 385514 267653
rect 385462 267589 385514 267595
rect 385570 265156 385598 271173
rect 385954 265156 385982 272357
rect 386434 271247 386462 272621
rect 386420 271238 386476 271247
rect 386420 271173 386476 271182
rect 386530 267949 386558 272621
rect 386612 272274 386668 272283
rect 386612 272209 386668 272218
rect 386518 267943 386570 267949
rect 386518 267885 386570 267891
rect 385570 265128 385824 265156
rect 385954 265128 386208 265156
rect 386626 265142 386654 272209
rect 387682 271099 387710 272949
rect 387476 271090 387532 271099
rect 387476 271025 387532 271034
rect 387668 271090 387724 271099
rect 387668 271025 387724 271034
rect 386902 270829 386954 270835
rect 386902 270771 386954 270777
rect 386914 265156 386942 270771
rect 387382 270015 387434 270021
rect 387382 269957 387434 269963
rect 387394 269577 387422 269957
rect 387286 269571 387338 269577
rect 387286 269513 387338 269519
rect 387382 269571 387434 269577
rect 387382 269513 387434 269519
rect 387298 268097 387326 269513
rect 387190 268091 387242 268097
rect 387190 268033 387242 268039
rect 387286 268091 387338 268097
rect 387286 268033 387338 268039
rect 387202 267653 387230 268033
rect 387190 267647 387242 267653
rect 387190 267589 387242 267595
rect 387490 265156 387518 271025
rect 387574 270089 387626 270095
rect 387574 270031 387626 270037
rect 387586 268985 387614 270031
rect 387574 268979 387626 268985
rect 387574 268921 387626 268927
rect 387778 265156 387806 278245
rect 390274 278161 390302 278541
rect 440662 278525 440714 278531
rect 397460 278490 397516 278499
rect 397460 278425 397462 278434
rect 397514 278425 397516 278434
rect 417428 278490 417484 278499
rect 417428 278425 417430 278434
rect 397462 278393 397514 278399
rect 417482 278425 417484 278434
rect 428852 278490 428908 278499
rect 429044 278490 429100 278499
rect 428908 278448 429044 278476
rect 428852 278425 428908 278434
rect 429044 278425 429100 278434
rect 440660 278490 440662 278499
rect 489622 278525 489674 278531
rect 440714 278490 440716 278499
rect 440660 278425 440716 278434
rect 489620 278490 489622 278499
rect 495382 278525 495434 278531
rect 489674 278490 489676 278499
rect 489620 278425 489676 278434
rect 495380 278490 495382 278499
rect 501334 278525 501386 278531
rect 495434 278490 495436 278499
rect 495380 278425 495436 278434
rect 501332 278490 501334 278499
rect 625078 278525 625130 278531
rect 501386 278490 501388 278499
rect 501332 278425 501388 278434
rect 525524 278490 525580 278499
rect 525524 278425 525526 278434
rect 417430 278393 417482 278399
rect 525578 278425 525580 278434
rect 551252 278490 551308 278499
rect 551252 278425 551254 278434
rect 525526 278393 525578 278399
rect 551306 278425 551308 278434
rect 610484 278490 610540 278499
rect 610484 278425 610486 278434
rect 551254 278393 551306 278399
rect 610538 278425 610540 278434
rect 610772 278490 610828 278499
rect 610772 278425 610774 278434
rect 610486 278393 610538 278399
rect 610826 278425 610828 278434
rect 625076 278490 625078 278499
rect 631030 278525 631082 278531
rect 625130 278490 625132 278499
rect 625076 278425 625132 278434
rect 631028 278490 631030 278499
rect 631082 278490 631084 278499
rect 631028 278425 631084 278434
rect 610774 278393 610826 278399
rect 467540 278342 467596 278351
rect 440674 278309 440798 278328
rect 396694 278303 396746 278309
rect 396694 278245 396746 278251
rect 440662 278303 440810 278309
rect 440714 278300 440758 278303
rect 440662 278245 440714 278251
rect 467596 278300 467856 278328
rect 490210 278309 490512 278328
rect 490198 278303 490512 278309
rect 467540 278277 467596 278286
rect 440758 278245 440810 278251
rect 490250 278300 490512 278303
rect 490198 278245 490250 278251
rect 396214 278229 396266 278235
rect 396266 278177 396528 278180
rect 396214 278171 396528 278177
rect 390166 278155 390218 278161
rect 390166 278097 390218 278103
rect 390262 278155 390314 278161
rect 396226 278152 396528 278171
rect 390262 278097 390314 278103
rect 387874 277856 388176 277884
rect 387874 272685 387902 277856
rect 390178 276681 390206 278097
rect 390166 276675 390218 276681
rect 390166 276617 390218 276623
rect 390562 274313 390590 277870
rect 390550 274307 390602 274313
rect 390550 274249 390602 274255
rect 391714 273795 391742 277870
rect 391702 273789 391754 273795
rect 391702 273731 391754 273737
rect 391414 272827 391466 272833
rect 391414 272769 391466 272775
rect 387862 272679 387914 272685
rect 387862 272621 387914 272627
rect 389684 272422 389740 272431
rect 389684 272357 389740 272366
rect 388148 271978 388204 271987
rect 388148 271913 388204 271922
rect 389588 271978 389644 271987
rect 389588 271913 389644 271922
rect 388054 270829 388106 270835
rect 388054 270771 388106 270777
rect 387862 267351 387914 267357
rect 387862 267293 387914 267299
rect 387874 267209 387902 267293
rect 387862 267203 387914 267209
rect 387862 267145 387914 267151
rect 386914 265128 387120 265156
rect 387490 265128 387600 265156
rect 387778 265128 387936 265156
rect 385076 264911 385132 264920
rect 388066 264915 388094 270771
rect 388162 265156 388190 271913
rect 389396 271830 389452 271839
rect 389396 271765 389452 271774
rect 388724 271238 388780 271247
rect 388724 271173 388780 271182
rect 388738 270983 388766 271173
rect 388630 270977 388682 270983
rect 388630 270919 388682 270925
rect 388726 270977 388778 270983
rect 388726 270919 388778 270925
rect 388642 270891 388670 270919
rect 388642 270863 388862 270891
rect 388834 270613 388862 270863
rect 388726 270607 388778 270613
rect 388726 270549 388778 270555
rect 388822 270607 388874 270613
rect 388822 270549 388874 270555
rect 388628 270498 388684 270507
rect 388738 270484 388766 270549
rect 388820 270498 388876 270507
rect 388738 270456 388820 270484
rect 388628 270433 388684 270442
rect 388820 270433 388876 270442
rect 388642 268985 388670 270433
rect 388630 268979 388682 268985
rect 388630 268921 388682 268927
rect 388918 268979 388970 268985
rect 388918 268921 388970 268927
rect 388930 268287 388958 268921
rect 388724 268278 388780 268287
rect 388724 268213 388780 268222
rect 388916 268278 388972 268287
rect 388916 268213 388972 268222
rect 388738 267949 388766 268213
rect 388726 267943 388778 267949
rect 388726 267885 388778 267891
rect 388820 267834 388876 267843
rect 388820 267769 388876 267778
rect 389012 267834 389068 267843
rect 389012 267769 389068 267778
rect 389300 267834 389356 267843
rect 389300 267769 389356 267778
rect 388834 267487 388862 267769
rect 389026 267653 389054 267769
rect 389110 267721 389162 267727
rect 389110 267663 389162 267669
rect 389206 267721 389258 267727
rect 389206 267663 389258 267669
rect 389014 267647 389066 267653
rect 389014 267589 389066 267595
rect 389014 267499 389066 267505
rect 388834 267459 389014 267487
rect 389014 267441 389066 267447
rect 388534 267203 388586 267209
rect 388534 267145 388586 267151
rect 388546 265211 388574 267145
rect 389122 266987 389150 267663
rect 389014 266981 389066 266987
rect 389014 266923 389066 266929
rect 389110 266981 389162 266987
rect 389110 266923 389162 266929
rect 388822 265353 388874 265359
rect 388822 265295 388874 265301
rect 388534 265205 388586 265211
rect 388162 265128 388416 265156
rect 388534 265147 388586 265153
rect 388834 265142 388862 265295
rect 389026 265211 389054 266923
rect 389218 266839 389246 267663
rect 389314 266839 389342 267769
rect 389206 266833 389258 266839
rect 389206 266775 389258 266781
rect 389302 266833 389354 266839
rect 389302 266775 389354 266781
rect 389014 265205 389066 265211
rect 389410 265156 389438 271765
rect 389602 265359 389630 271913
rect 389590 265353 389642 265359
rect 389590 265295 389642 265301
rect 389014 265147 389066 265153
rect 389232 265128 389438 265156
rect 389698 265142 389726 272357
rect 390934 272309 390986 272315
rect 390934 272251 390986 272257
rect 390836 271830 390892 271839
rect 390836 271765 390892 271774
rect 389876 271534 389932 271543
rect 389876 271469 389932 271478
rect 389782 265353 389834 265359
rect 389782 265295 389834 265301
rect 389794 264989 389822 265295
rect 389890 265156 389918 271469
rect 390166 268979 390218 268985
rect 390166 268921 390218 268927
rect 390178 267875 390206 268921
rect 390454 268461 390506 268467
rect 390454 268403 390506 268409
rect 390466 267949 390494 268403
rect 390358 267943 390410 267949
rect 390358 267885 390410 267891
rect 390454 267943 390506 267949
rect 390454 267885 390506 267891
rect 390166 267869 390218 267875
rect 390166 267811 390218 267817
rect 390262 267869 390314 267875
rect 390262 267811 390314 267817
rect 390274 267505 390302 267811
rect 390370 267653 390398 267885
rect 390358 267647 390410 267653
rect 390358 267589 390410 267595
rect 390262 267499 390314 267505
rect 390262 267441 390314 267447
rect 390454 265205 390506 265211
rect 389890 265128 390144 265156
rect 390850 265156 390878 271765
rect 390454 265147 390506 265153
rect 390262 265131 390314 265137
rect 390262 265073 390314 265079
rect 390274 264989 390302 265073
rect 390466 265063 390494 265147
rect 390624 265128 390878 265156
rect 390946 265142 390974 272251
rect 391426 265142 391454 272769
rect 391894 272605 391946 272611
rect 391894 272547 391946 272553
rect 391906 265142 391934 272547
rect 392470 272383 392522 272389
rect 392470 272325 392522 272331
rect 392482 272135 392510 272325
rect 392566 272309 392618 272315
rect 392566 272251 392618 272257
rect 392468 272126 392524 272135
rect 392468 272061 392524 272070
rect 392086 270755 392138 270761
rect 392086 270697 392138 270703
rect 392098 265156 392126 270697
rect 392578 265156 392606 272251
rect 392962 265507 392990 277870
rect 394582 273419 394634 273425
rect 394582 273361 394634 273367
rect 394100 273014 394156 273023
rect 394100 272949 394156 272958
rect 393140 272866 393196 272875
rect 393140 272801 393196 272810
rect 392950 265501 393002 265507
rect 392950 265443 393002 265449
rect 392098 265128 392352 265156
rect 392578 265128 392736 265156
rect 393154 265142 393182 272801
rect 393814 272309 393866 272315
rect 393814 272251 393866 272257
rect 393622 271125 393674 271131
rect 393622 271067 393674 271073
rect 393634 265142 393662 271067
rect 393826 270803 393854 272251
rect 393812 270794 393868 270803
rect 393812 270729 393868 270738
rect 394114 265142 394142 272949
rect 394594 272611 394622 273361
rect 394870 273271 394922 273277
rect 394870 273213 394922 273219
rect 394582 272605 394634 272611
rect 394292 272570 394348 272579
rect 394582 272547 394634 272553
rect 394292 272505 394348 272514
rect 394306 272463 394334 272505
rect 394198 272457 394250 272463
rect 394198 272399 394250 272405
rect 394294 272457 394346 272463
rect 394294 272399 394346 272405
rect 394210 265156 394238 272399
rect 394882 271871 394910 273213
rect 395254 272013 395306 272019
rect 395254 271955 395306 271961
rect 394870 271865 394922 271871
rect 394870 271807 394922 271813
rect 394966 271865 395018 271871
rect 394966 271807 395018 271813
rect 394486 271125 394538 271131
rect 394484 271090 394486 271099
rect 394538 271090 394540 271099
rect 394484 271025 394540 271034
rect 394484 270942 394540 270951
rect 394978 270909 395006 271807
rect 395156 271534 395212 271543
rect 395156 271469 395212 271478
rect 395062 271199 395114 271205
rect 395062 271141 395114 271147
rect 395074 270909 395102 271141
rect 394484 270877 394540 270886
rect 394966 270903 395018 270909
rect 394498 270761 394526 270877
rect 394966 270845 395018 270851
rect 395062 270903 395114 270909
rect 395062 270845 395114 270851
rect 394486 270755 394538 270761
rect 394486 270697 394538 270703
rect 395170 265156 395198 271469
rect 394210 265128 394464 265156
rect 394944 265128 395198 265156
rect 395266 265156 395294 271955
rect 395362 268541 395390 277870
rect 396706 277019 396734 278245
rect 474740 278194 474796 278203
rect 474796 278152 475056 278180
rect 636514 278161 636720 278180
rect 636502 278155 636720 278161
rect 474740 278129 474796 278138
rect 636554 278152 636720 278155
rect 636502 278097 636554 278103
rect 415318 278081 415370 278087
rect 481844 278046 481900 278055
rect 415370 278029 415632 278032
rect 415318 278023 415632 278029
rect 415330 278004 415632 278023
rect 422338 278013 422640 278032
rect 422326 278007 422640 278013
rect 422378 278004 422640 278007
rect 646004 278046 646060 278055
rect 481900 278004 482160 278032
rect 481844 277981 481900 277990
rect 646060 278004 646320 278032
rect 646004 277981 646060 277990
rect 422326 277949 422378 277955
rect 436630 277933 436682 277939
rect 397474 277856 397776 277884
rect 398626 277856 398928 277884
rect 396692 277010 396748 277019
rect 396692 276945 396748 276954
rect 397474 275127 397502 277856
rect 397462 275121 397514 275127
rect 397462 275063 397514 275069
rect 398626 274535 398654 277856
rect 398902 276453 398954 276459
rect 398902 276395 398954 276401
rect 398914 275349 398942 276395
rect 398806 275343 398858 275349
rect 398806 275285 398858 275291
rect 398902 275343 398954 275349
rect 398902 275285 398954 275291
rect 398818 275127 398846 275285
rect 398806 275121 398858 275127
rect 398806 275063 398858 275069
rect 398614 274529 398666 274535
rect 398614 274471 398666 274477
rect 398902 274455 398954 274461
rect 398902 274397 398954 274403
rect 398914 274239 398942 274397
rect 400066 274387 400094 277870
rect 401218 276533 401246 277870
rect 401206 276527 401258 276533
rect 401206 276469 401258 276475
rect 400054 274381 400106 274387
rect 400054 274323 400106 274329
rect 398902 274233 398954 274239
rect 398902 274175 398954 274181
rect 397364 273606 397420 273615
rect 396214 273567 396266 273573
rect 397364 273541 397366 273550
rect 396214 273509 396266 273515
rect 397418 273541 397420 273550
rect 397366 273509 397418 273515
rect 395828 272718 395884 272727
rect 395828 272653 395884 272662
rect 395446 271199 395498 271205
rect 395446 271141 395498 271147
rect 395458 270835 395486 271141
rect 395446 270829 395498 270835
rect 395446 270771 395498 270777
rect 395636 270794 395692 270803
rect 395636 270729 395692 270738
rect 395446 268979 395498 268985
rect 395446 268921 395498 268927
rect 395458 268541 395486 268921
rect 395350 268535 395402 268541
rect 395350 268477 395402 268483
rect 395446 268535 395498 268541
rect 395446 268477 395498 268483
rect 395650 267505 395678 270729
rect 395638 267499 395690 267505
rect 395638 267441 395690 267447
rect 395734 265501 395786 265507
rect 395734 265443 395786 265449
rect 395746 265359 395774 265443
rect 395734 265353 395786 265359
rect 395734 265295 395786 265301
rect 395266 265128 395376 265156
rect 395842 265142 395870 272653
rect 395924 270794 395980 270803
rect 395924 270729 395980 270738
rect 395938 265359 395966 270729
rect 395926 265353 395978 265359
rect 395926 265295 395978 265301
rect 396226 265142 396254 273509
rect 400630 273197 400682 273203
rect 397364 273162 397420 273171
rect 397364 273097 397420 273106
rect 397556 273162 397612 273171
rect 400630 273139 400682 273145
rect 397556 273097 397612 273106
rect 399670 273123 399722 273129
rect 397270 272753 397322 272759
rect 397270 272695 397322 272701
rect 396886 272605 396938 272611
rect 396886 272547 396938 272553
rect 396980 272570 397036 272579
rect 396898 272019 396926 272547
rect 396980 272505 397036 272514
rect 396886 272013 396938 272019
rect 396886 271955 396938 271961
rect 396884 271238 396940 271247
rect 396884 271173 396940 271182
rect 396898 265156 396926 271173
rect 396672 265128 396926 265156
rect 396994 265156 397022 272505
rect 397282 271691 397310 272695
rect 397378 272611 397406 273097
rect 397366 272605 397418 272611
rect 397366 272547 397418 272553
rect 397570 272431 397598 273097
rect 399670 273065 399722 273071
rect 398614 273049 398666 273055
rect 398614 272991 398666 272997
rect 398038 272975 398090 272981
rect 398038 272917 398090 272923
rect 397556 272422 397612 272431
rect 397556 272357 397612 272366
rect 397268 271682 397324 271691
rect 397268 271617 397324 271626
rect 397844 270942 397900 270951
rect 397844 270877 397900 270886
rect 397556 267834 397612 267843
rect 397556 267769 397612 267778
rect 397570 265655 397598 267769
rect 397558 265649 397610 265655
rect 397558 265591 397610 265597
rect 397858 265156 397886 270877
rect 398050 265156 398078 272917
rect 398420 272570 398476 272579
rect 398420 272505 398476 272514
rect 396994 265128 397152 265156
rect 397488 265128 397886 265156
rect 397968 265128 398078 265156
rect 398434 265142 398462 272505
rect 398626 265156 398654 272991
rect 398806 272679 398858 272685
rect 398806 272621 398858 272627
rect 398818 272019 398846 272621
rect 398710 272013 398762 272019
rect 398710 271955 398762 271961
rect 398806 272013 398858 272019
rect 398806 271955 398858 271961
rect 398722 271779 398750 271955
rect 398722 271751 398942 271779
rect 398914 270835 398942 271751
rect 399476 271090 399532 271099
rect 399476 271025 399532 271034
rect 398902 270829 398954 270835
rect 398902 270771 398954 270777
rect 398806 268979 398858 268985
rect 398806 268921 398858 268927
rect 398818 268763 398846 268921
rect 398806 268757 398858 268763
rect 398806 268699 398858 268705
rect 398722 267607 399038 267635
rect 398722 267505 398750 267607
rect 398710 267499 398762 267505
rect 398710 267441 398762 267447
rect 398806 267499 398858 267505
rect 398806 267441 398858 267447
rect 398818 266765 398846 267441
rect 398902 267055 398954 267061
rect 398902 266997 398954 267003
rect 398806 266759 398858 266765
rect 398806 266701 398858 266707
rect 398914 265951 398942 266997
rect 399010 266765 399038 267607
rect 398998 266759 399050 266765
rect 398998 266701 399050 266707
rect 398806 265945 398858 265951
rect 398806 265887 398858 265893
rect 398902 265945 398954 265951
rect 398902 265887 398954 265893
rect 398818 265729 398846 265887
rect 398806 265723 398858 265729
rect 398806 265665 398858 265671
rect 398626 265128 398880 265156
rect 399382 265131 399434 265137
rect 399382 265073 399434 265079
rect 390454 265057 390506 265063
rect 390454 264999 390506 265005
rect 399394 264989 399422 265073
rect 389782 264983 389834 264989
rect 389782 264925 389834 264931
rect 390262 264983 390314 264989
rect 390262 264925 390314 264931
rect 399382 264983 399434 264989
rect 399382 264925 399434 264931
rect 379124 264874 379180 264883
rect 379042 264832 379124 264860
rect 308084 264809 308140 264818
rect 385076 264846 385132 264855
rect 388054 264909 388106 264915
rect 399490 264860 399518 271025
rect 399682 265142 399710 273065
rect 400148 272422 400204 272431
rect 400148 272357 400204 272366
rect 399862 267647 399914 267653
rect 399862 267589 399914 267595
rect 399874 264989 399902 267589
rect 400162 265142 400190 272357
rect 400642 265142 400670 273139
rect 402358 272531 402410 272537
rect 402358 272473 402410 272479
rect 401876 271682 401932 271691
rect 401876 271617 401932 271626
rect 401302 270903 401354 270909
rect 401302 270845 401354 270851
rect 401204 270794 401260 270803
rect 401204 270729 401260 270738
rect 401218 265156 401246 270729
rect 400992 265128 401246 265156
rect 401314 265156 401342 270845
rect 401314 265128 401472 265156
rect 401890 265142 401918 271617
rect 402370 265142 402398 272473
rect 402466 268615 402494 277870
rect 403618 277717 403646 277870
rect 403606 277711 403658 277717
rect 403606 277653 403658 277659
rect 403124 273902 403180 273911
rect 403124 273837 403180 273846
rect 403138 273795 403166 273837
rect 403126 273789 403178 273795
rect 403126 273731 403178 273737
rect 404086 273419 404138 273425
rect 404086 273361 404138 273367
rect 403990 273345 404042 273351
rect 403990 273287 404042 273293
rect 402740 272126 402796 272135
rect 402740 272061 402796 272070
rect 402454 268609 402506 268615
rect 402454 268551 402506 268557
rect 402754 265142 402782 272061
rect 403186 271751 403742 271779
rect 403186 271723 403214 271751
rect 403174 271717 403226 271723
rect 403174 271659 403226 271665
rect 403030 271643 403082 271649
rect 403030 271585 403082 271591
rect 403042 267653 403070 271585
rect 403126 271569 403178 271575
rect 403318 271569 403370 271575
rect 403126 271511 403178 271517
rect 403234 271517 403318 271520
rect 403234 271511 403370 271517
rect 403030 267647 403082 267653
rect 403030 267589 403082 267595
rect 403138 267061 403166 271511
rect 403234 271501 403358 271511
rect 403222 271495 403358 271501
rect 403274 271492 403358 271495
rect 403222 271437 403274 271443
rect 403414 271347 403466 271353
rect 403414 271289 403466 271295
rect 403426 270909 403454 271289
rect 403414 270903 403466 270909
rect 403414 270845 403466 270851
rect 403222 268757 403274 268763
rect 403222 268699 403274 268705
rect 403126 267055 403178 267061
rect 403126 266997 403178 267003
rect 403234 265156 403262 268699
rect 403714 268615 403742 271751
rect 404002 268763 404030 273287
rect 403990 268757 404042 268763
rect 403990 268699 404042 268705
rect 403702 268609 403754 268615
rect 403702 268551 403754 268557
rect 403702 268461 403754 268467
rect 403702 268403 403754 268409
rect 403714 268287 403742 268403
rect 403700 268278 403756 268287
rect 403700 268213 403756 268222
rect 403892 268278 403948 268287
rect 403892 268213 403948 268222
rect 403906 265156 403934 268213
rect 403200 265128 403262 265156
rect 403680 265128 403934 265156
rect 404098 265142 404126 273361
rect 404770 266987 404798 277870
rect 406018 274609 406046 277870
rect 406978 277856 407184 277884
rect 408130 277856 408432 277884
rect 488948 277898 489004 277907
rect 436682 277881 436944 277884
rect 436630 277875 436944 277881
rect 406006 274603 406058 274609
rect 406006 274545 406058 274551
rect 405910 272087 405962 272093
rect 405910 272029 405962 272035
rect 404950 270829 405002 270835
rect 404950 270771 405002 270777
rect 404852 268278 404908 268287
rect 404852 268213 404908 268222
rect 404758 266981 404810 266987
rect 404758 266923 404810 266929
rect 404866 265156 404894 268213
rect 404496 265128 404894 265156
rect 404962 265142 404990 270771
rect 405716 268278 405772 268287
rect 405538 268236 405716 268264
rect 405538 265156 405566 268236
rect 405716 268213 405772 268222
rect 405922 265156 405950 272029
rect 406678 271865 406730 271871
rect 406678 271807 406730 271813
rect 406102 268461 406154 268467
rect 406102 268403 406154 268409
rect 406114 268287 406142 268403
rect 406100 268278 406156 268287
rect 406100 268213 406156 268222
rect 405408 265128 405566 265156
rect 405792 265128 405950 265156
rect 406690 265142 406718 271807
rect 406978 265063 407006 277856
rect 407542 271939 407594 271945
rect 407542 271881 407594 271887
rect 407060 271682 407116 271691
rect 407060 271617 407116 271626
rect 407074 271247 407102 271617
rect 407060 271238 407116 271247
rect 407060 271173 407116 271182
rect 407062 265501 407114 265507
rect 407062 265443 407114 265449
rect 407074 265063 407102 265443
rect 407554 265142 407582 271881
rect 408130 268541 408158 277856
rect 408982 274381 409034 274387
rect 408982 274323 409034 274329
rect 408994 274239 409022 274323
rect 408982 274233 409034 274239
rect 408982 274175 409034 274181
rect 408214 273271 408266 273277
rect 408214 273213 408266 273219
rect 408118 268535 408170 268541
rect 408118 268477 408170 268483
rect 408226 266987 408254 273213
rect 408596 272718 408652 272727
rect 408596 272653 408652 272662
rect 408500 272570 408556 272579
rect 408500 272505 408556 272514
rect 408404 272422 408460 272431
rect 408404 272357 408460 272366
rect 408418 271691 408446 272357
rect 408514 271839 408542 272505
rect 408610 272135 408638 272653
rect 408596 272126 408652 272135
rect 408596 272061 408652 272070
rect 408500 271830 408556 271839
rect 408500 271765 408556 271774
rect 409270 271791 409322 271797
rect 409270 271733 409322 271739
rect 408404 271682 408460 271691
rect 408404 271617 408460 271626
rect 408214 266981 408266 266987
rect 408214 266923 408266 266929
rect 408694 266981 408746 266987
rect 408694 266923 408746 266929
rect 408214 266759 408266 266765
rect 408214 266701 408266 266707
rect 408406 266759 408458 266765
rect 408406 266701 408458 266707
rect 408226 265507 408254 266701
rect 408214 265501 408266 265507
rect 408214 265443 408266 265449
rect 408418 265341 408446 266701
rect 408322 265313 408446 265341
rect 408322 265119 408350 265313
rect 408226 265091 408350 265119
rect 406966 265057 407018 265063
rect 406966 264999 407018 265005
rect 407062 265057 407114 265063
rect 407062 264999 407114 265005
rect 399862 264983 399914 264989
rect 399862 264925 399914 264931
rect 406484 264911 406540 264920
rect 388054 264851 388106 264857
rect 399264 264832 399518 264860
rect 406272 264855 406484 264860
rect 407252 264911 407308 264920
rect 406272 264846 406540 264855
rect 407184 264855 407252 264860
rect 407184 264846 407308 264855
rect 407732 264911 407788 264920
rect 408116 264911 408172 264920
rect 407788 264855 408000 264860
rect 407732 264846 408000 264855
rect 408226 264897 408254 265091
rect 408706 264897 408734 266923
rect 409282 265142 409310 271733
rect 409570 268911 409598 277870
rect 410818 277643 410846 277870
rect 410806 277637 410858 277643
rect 410806 277579 410858 277585
rect 411970 273647 411998 277870
rect 413218 274757 413246 277870
rect 413206 274751 413258 274757
rect 413206 274693 413258 274699
rect 411958 273641 412010 273647
rect 411958 273583 412010 273589
rect 412246 272827 412298 272833
rect 412246 272769 412298 272775
rect 409654 271939 409706 271945
rect 409654 271881 409706 271887
rect 409666 271279 409694 271881
rect 409654 271273 409706 271279
rect 409654 271215 409706 271221
rect 409558 268905 409610 268911
rect 409558 268847 409610 268853
rect 409942 268609 409994 268615
rect 409942 268551 409994 268557
rect 409954 265156 409982 268551
rect 410998 267647 411050 267653
rect 410998 267589 411050 267595
rect 409954 265128 410208 265156
rect 411010 265142 411038 267589
rect 411958 267055 412010 267061
rect 411958 266997 412010 267003
rect 411970 265142 411998 266997
rect 409570 264980 409776 265008
rect 411202 264980 411504 265008
rect 409570 264920 409598 264980
rect 411202 264920 411230 264980
rect 408172 264869 408254 264897
rect 408610 264869 408734 264897
rect 408788 264911 408844 264920
rect 408610 264860 408638 264869
rect 408116 264846 408172 264855
rect 406272 264832 406526 264846
rect 407184 264832 407294 264846
rect 407746 264832 408000 264846
rect 408480 264832 408638 264860
rect 409556 264911 409612 264920
rect 408844 264855 408912 264860
rect 408788 264846 408912 264855
rect 410804 264911 410860 264920
rect 409556 264846 409612 264855
rect 410688 264855 410804 264860
rect 410688 264846 410860 264855
rect 411188 264911 411244 264920
rect 411188 264846 411244 264855
rect 408802 264832 408912 264846
rect 410688 264832 410846 264846
rect 379124 264809 379180 264818
rect 412148 247262 412204 247271
rect 412148 247197 412204 247206
rect 223124 246818 223180 246827
rect 223124 246753 223180 246762
rect 224852 246818 224908 246827
rect 224852 246753 224908 246762
rect 225332 246818 225388 246827
rect 228116 246818 228172 246827
rect 225332 246753 225388 246762
rect 227446 246779 227498 246785
rect 212276 238974 212332 238983
rect 212276 238909 212332 238918
rect 211892 236606 211948 236615
rect 211892 236541 211948 236550
rect 211316 236458 211372 236467
rect 211316 236393 211372 236402
rect 211330 233484 211358 236393
rect 211796 233498 211852 233507
rect 210370 233456 211200 233484
rect 211330 233456 211796 233484
rect 210262 227835 210314 227841
rect 210262 227777 210314 227783
rect 210262 227613 210314 227619
rect 210262 227555 210314 227561
rect 210274 187437 210302 227555
rect 210262 187431 210314 187437
rect 210262 187373 210314 187379
rect 210262 187135 210314 187141
rect 210262 187077 210314 187083
rect 210164 161570 210220 161579
rect 210164 161505 210220 161514
rect 210178 158471 210206 161505
rect 210164 158462 210220 158471
rect 210164 158397 210220 158406
rect 210274 147033 210302 187077
rect 210262 147027 210314 147033
rect 210262 146969 210314 146975
rect 210262 146583 210314 146589
rect 210262 146525 210314 146531
rect 210164 141590 210220 141599
rect 210164 141525 210220 141534
rect 210178 138491 210206 141525
rect 210164 138482 210220 138491
rect 210164 138417 210220 138426
rect 210164 129158 210220 129167
rect 210164 129093 210220 129102
rect 210178 126207 210206 129093
rect 210164 126198 210220 126207
rect 210164 126133 210220 126142
rect 210164 121166 210220 121175
rect 210164 121101 210220 121110
rect 210178 113775 210206 121101
rect 210274 120985 210302 146525
rect 210262 120979 210314 120985
rect 210262 120921 210314 120927
rect 210164 113766 210220 113775
rect 210164 113701 210220 113710
rect 210166 106327 210218 106333
rect 210166 106269 210218 106275
rect 210178 86797 210206 106269
rect 210370 106204 210398 233456
rect 211906 233484 211934 236541
rect 212276 236310 212332 236319
rect 212276 236245 212332 236254
rect 212180 233646 212236 233655
rect 212180 233581 212236 233590
rect 212194 233484 212222 233581
rect 211906 233456 212222 233484
rect 212290 233484 212318 236245
rect 212386 235135 212414 246494
rect 212770 240865 212798 246494
rect 213142 245447 213194 245453
rect 213142 245389 213194 245395
rect 212758 240859 212810 240865
rect 212758 240801 212810 240807
rect 212660 236754 212716 236763
rect 212660 236689 212716 236698
rect 212372 235126 212428 235135
rect 212372 235061 212428 235070
rect 212564 233498 212620 233507
rect 212290 233470 212564 233484
rect 212304 233456 212564 233470
rect 211796 233433 211852 233442
rect 212674 233484 212702 236689
rect 213046 236197 213098 236203
rect 213046 236139 213098 236145
rect 212852 233498 212908 233507
rect 212674 233470 212852 233484
rect 212688 233456 212852 233470
rect 212564 233433 212620 233442
rect 213058 233470 213086 236139
rect 213154 233539 213182 245389
rect 213250 243719 213278 246494
rect 213696 246480 213950 246508
rect 213236 243710 213292 243719
rect 213236 243645 213292 243654
rect 213526 243301 213578 243307
rect 213526 243243 213578 243249
rect 213538 233613 213566 243243
rect 213922 241605 213950 246480
rect 214066 246212 214094 246494
rect 214198 246335 214250 246341
rect 214198 246277 214250 246283
rect 214066 246184 214142 246212
rect 213910 241599 213962 241605
rect 213910 241541 213962 241547
rect 214114 234987 214142 246184
rect 214100 234978 214156 234987
rect 214100 234913 214156 234922
rect 214210 233928 214238 246277
rect 214294 244929 214346 244935
rect 214294 244871 214346 244877
rect 214114 233900 214238 233928
rect 213526 233607 213578 233613
rect 213526 233549 213578 233555
rect 213142 233533 213194 233539
rect 213538 233484 213566 233549
rect 213910 233533 213962 233539
rect 213194 233481 213408 233484
rect 213142 233475 213408 233481
rect 213154 233456 213408 233475
rect 213538 233456 213792 233484
rect 214114 233484 214142 233900
rect 214306 233507 214334 244871
rect 214498 239755 214526 246494
rect 214978 243275 215006 246494
rect 214964 243266 215020 243275
rect 214964 243201 215020 243210
rect 215458 241827 215486 246494
rect 215808 246480 215966 246508
rect 216288 246480 216542 246508
rect 215446 241821 215498 241827
rect 215446 241763 215498 241769
rect 214486 239749 214538 239755
rect 214486 239691 214538 239697
rect 215938 239237 215966 246480
rect 216514 244935 216542 246480
rect 216598 245225 216650 245231
rect 216598 245167 216650 245173
rect 216502 244929 216554 244935
rect 216502 244871 216554 244877
rect 215926 239231 215978 239237
rect 215926 239173 215978 239179
rect 215828 238234 215884 238243
rect 215828 238169 215884 238178
rect 215252 238086 215308 238095
rect 215252 238021 215308 238030
rect 214868 237938 214924 237947
rect 214868 237873 214924 237882
rect 214772 237642 214828 237651
rect 214772 237577 214828 237586
rect 214786 236615 214814 237577
rect 214772 236606 214828 236615
rect 214772 236541 214828 236550
rect 213962 233481 214142 233484
rect 213910 233475 214142 233481
rect 213922 233456 214142 233475
rect 212852 233433 212908 233442
rect 214114 233336 214142 233456
rect 214292 233498 214348 233507
rect 214348 233456 214512 233484
rect 214882 233470 214910 237873
rect 215266 233470 215294 238021
rect 215842 233484 215870 238169
rect 216212 237642 216268 237651
rect 216212 237577 216268 237586
rect 216226 233484 216254 237577
rect 216610 233484 216638 245167
rect 216706 241161 216734 246494
rect 217186 243127 217214 246494
rect 217172 243118 217228 243127
rect 217172 243053 217228 243062
rect 217570 241901 217598 246494
rect 218016 246480 218270 246508
rect 218496 246480 218750 246508
rect 217558 241895 217610 241901
rect 217558 241837 217610 241843
rect 216694 241155 216746 241161
rect 216694 241097 216746 241103
rect 217078 238565 217130 238571
rect 217078 238507 217130 238513
rect 216692 237790 216748 237799
rect 216692 237725 216748 237734
rect 215616 233456 215870 233484
rect 216000 233456 216254 233484
rect 216384 233456 216638 233484
rect 216706 233470 216734 237725
rect 217090 233470 217118 238507
rect 218038 238343 218090 238349
rect 218038 238285 218090 238291
rect 217462 236419 217514 236425
rect 217462 236361 217514 236367
rect 217474 233470 217502 236361
rect 218050 233484 218078 238285
rect 218242 235283 218270 246480
rect 218722 241753 218750 246480
rect 218914 242979 218942 246494
rect 218900 242970 218956 242979
rect 218900 242905 218956 242914
rect 218710 241747 218762 241753
rect 218710 241689 218762 241695
rect 219298 241679 219326 246494
rect 219286 241673 219338 241679
rect 219286 241615 219338 241621
rect 219286 240711 219338 240717
rect 219286 240653 219338 240659
rect 218806 240341 218858 240347
rect 218806 240283 218858 240289
rect 218422 240193 218474 240199
rect 218422 240135 218474 240141
rect 218228 235274 218284 235283
rect 218228 235209 218284 235218
rect 218434 233484 218462 240135
rect 218818 233484 218846 240283
rect 218902 239231 218954 239237
rect 218902 239173 218954 239179
rect 217824 233456 218078 233484
rect 218208 233456 218462 233484
rect 218592 233456 218846 233484
rect 218914 233470 218942 239173
rect 219298 233470 219326 240653
rect 219670 240563 219722 240569
rect 219670 240505 219722 240511
rect 219682 233470 219710 240505
rect 219778 235727 219806 246494
rect 220224 246480 220478 246508
rect 220608 246480 220862 246508
rect 221040 246480 221342 246508
rect 220246 240637 220298 240643
rect 220246 240579 220298 240585
rect 219764 235718 219820 235727
rect 219764 235653 219820 235662
rect 220258 233484 220286 240579
rect 220450 240495 220478 246480
rect 220834 242831 220862 246480
rect 220820 242822 220876 242831
rect 220820 242757 220876 242766
rect 220438 240489 220490 240495
rect 220438 240431 220490 240437
rect 220630 240415 220682 240421
rect 220630 240357 220682 240363
rect 220642 233484 220670 240357
rect 221014 237381 221066 237387
rect 221014 237323 221066 237329
rect 221026 233484 221054 237323
rect 221110 237307 221162 237313
rect 221110 237249 221162 237255
rect 220032 233456 220286 233484
rect 220416 233456 220670 233484
rect 220800 233456 221054 233484
rect 221122 233470 221150 237249
rect 221314 235579 221342 246480
rect 221396 242082 221452 242091
rect 221396 242017 221452 242026
rect 221410 241827 221438 242017
rect 221398 241821 221450 241827
rect 221398 241763 221450 241769
rect 221506 241087 221534 246494
rect 221986 242683 222014 246494
rect 222336 246480 222590 246508
rect 222816 246480 223070 246508
rect 221972 242674 222028 242683
rect 221972 242609 222028 242618
rect 222562 241531 222590 246480
rect 222550 241525 222602 241531
rect 222550 241467 222602 241473
rect 221494 241081 221546 241087
rect 221494 241023 221546 241029
rect 221782 240119 221834 240125
rect 221782 240061 221834 240067
rect 221494 237677 221546 237683
rect 221494 237619 221546 237625
rect 221300 235570 221356 235579
rect 221300 235505 221356 235514
rect 221506 233470 221534 237619
rect 221794 236425 221822 240061
rect 221878 238047 221930 238053
rect 221878 237989 221930 237995
rect 221782 236419 221834 236425
rect 221782 236361 221834 236367
rect 221890 233470 221918 237989
rect 222838 237899 222890 237905
rect 222838 237841 222890 237847
rect 221974 237603 222026 237609
rect 221974 237545 222026 237551
rect 221986 233484 222014 237545
rect 222850 233484 222878 237841
rect 223042 235431 223070 246480
rect 223138 245527 223166 246753
rect 223126 245521 223178 245527
rect 223126 245463 223178 245469
rect 223234 239977 223262 246494
rect 223510 243079 223562 243085
rect 223510 243021 223562 243027
rect 223522 242239 223550 243021
rect 223714 242239 223742 246494
rect 223990 242561 224042 242567
rect 223988 242526 223990 242535
rect 224042 242526 224044 242535
rect 223988 242461 224044 242470
rect 223508 242230 223564 242239
rect 223508 242165 223564 242174
rect 223700 242230 223756 242239
rect 223700 242165 223756 242174
rect 224098 240791 224126 246494
rect 224530 246212 224558 246494
rect 224482 246184 224558 246212
rect 224086 240785 224138 240791
rect 224086 240727 224138 240733
rect 223222 239971 223274 239977
rect 223222 239913 223274 239919
rect 223222 238121 223274 238127
rect 223222 238063 223274 238069
rect 223028 235422 223084 235431
rect 223028 235357 223084 235366
rect 223234 233484 223262 238063
rect 223318 237973 223370 237979
rect 223318 237915 223370 237921
rect 221986 233456 222240 233484
rect 222624 233456 222878 233484
rect 223008 233456 223262 233484
rect 223330 233470 223358 237915
rect 223702 237825 223754 237831
rect 223702 237767 223754 237773
rect 223714 233470 223742 237767
rect 224086 237011 224138 237017
rect 224086 236953 224138 236959
rect 224098 233470 224126 236953
rect 224482 235875 224510 246184
rect 224866 245749 224894 246753
rect 225346 246563 225374 246753
rect 227446 246721 227498 246727
rect 227926 246779 227978 246785
rect 228116 246753 228172 246762
rect 228308 246818 228364 246827
rect 228308 246753 228364 246762
rect 228596 246818 228652 246827
rect 246164 246818 246220 246827
rect 228596 246753 228652 246762
rect 231862 246779 231914 246785
rect 227926 246721 227978 246727
rect 227062 246705 227114 246711
rect 227062 246647 227114 246653
rect 226486 246631 226538 246637
rect 226486 246573 226538 246579
rect 226966 246631 227018 246637
rect 226966 246573 227018 246579
rect 225334 246557 225386 246563
rect 225024 246480 225278 246508
rect 225334 246499 225386 246505
rect 224854 245743 224906 245749
rect 224854 245685 224906 245691
rect 225250 241013 225278 246480
rect 225238 241007 225290 241013
rect 225238 240949 225290 240955
rect 225442 240939 225470 246494
rect 225430 240933 225482 240939
rect 225430 240875 225482 240881
rect 225142 239749 225194 239755
rect 225142 239691 225194 239697
rect 224566 238787 224618 238793
rect 224566 238729 224618 238735
rect 224468 235866 224524 235875
rect 224468 235801 224524 235810
rect 224578 233484 224606 238729
rect 225046 236863 225098 236869
rect 225046 236805 225098 236811
rect 225058 233484 225086 236805
rect 224448 233456 224606 233484
rect 224832 233456 225086 233484
rect 225154 233484 225182 239691
rect 225526 237159 225578 237165
rect 225526 237101 225578 237107
rect 225154 233456 225216 233484
rect 225538 233470 225566 237101
rect 225826 236171 225854 246494
rect 226306 241235 226334 246494
rect 226498 245601 226526 246573
rect 226752 246480 226814 246508
rect 226486 245595 226538 245601
rect 226486 245537 226538 245543
rect 226786 243455 226814 246480
rect 226978 245823 227006 246573
rect 226966 245817 227018 245823
rect 226966 245759 227018 245765
rect 227074 245675 227102 246647
rect 227170 246480 227232 246508
rect 227062 245669 227114 245675
rect 227062 245611 227114 245617
rect 227060 243710 227116 243719
rect 227060 243645 227062 243654
rect 227114 243645 227116 243654
rect 227062 243613 227114 243619
rect 226774 243449 226826 243455
rect 226774 243391 226826 243397
rect 227060 243118 227116 243127
rect 227060 243053 227116 243062
rect 227074 242789 227102 243053
rect 227062 242783 227114 242789
rect 227062 242725 227114 242731
rect 226294 241229 226346 241235
rect 226294 241171 226346 241177
rect 227170 239903 227198 246480
rect 227458 245823 227486 246721
rect 227830 246705 227882 246711
rect 227830 246647 227882 246653
rect 227842 246563 227870 246647
rect 227830 246557 227882 246563
rect 227830 246499 227882 246505
rect 227446 245817 227498 245823
rect 227446 245759 227498 245765
rect 227348 243710 227404 243719
rect 227266 243668 227348 243696
rect 227266 242387 227294 243668
rect 227348 243645 227404 243654
rect 227348 243266 227404 243275
rect 227348 243201 227404 243210
rect 227362 243085 227390 243201
rect 227350 243079 227402 243085
rect 227350 243021 227402 243027
rect 227348 242970 227404 242979
rect 227554 242956 227582 246494
rect 227938 246341 227966 246721
rect 227926 246335 227978 246341
rect 227926 246277 227978 246283
rect 227554 242928 227966 242956
rect 227348 242905 227404 242914
rect 227362 242715 227390 242905
rect 227830 242857 227882 242863
rect 227636 242822 227692 242831
rect 227830 242799 227882 242805
rect 227636 242757 227638 242766
rect 227690 242757 227692 242766
rect 227638 242725 227690 242731
rect 227350 242709 227402 242715
rect 227734 242709 227786 242715
rect 227350 242651 227402 242657
rect 227540 242674 227596 242683
rect 227540 242609 227596 242618
rect 227732 242674 227734 242683
rect 227786 242674 227788 242683
rect 227732 242609 227788 242618
rect 227554 242387 227582 242609
rect 227842 242512 227870 242799
rect 227650 242484 227870 242512
rect 227252 242378 227308 242387
rect 227252 242313 227308 242322
rect 227540 242378 227596 242387
rect 227540 242313 227596 242322
rect 227650 242239 227678 242484
rect 227636 242230 227692 242239
rect 227636 242165 227692 242174
rect 227158 239897 227210 239903
rect 227158 239839 227210 239845
rect 227734 238935 227786 238941
rect 227734 238877 227786 238883
rect 226294 238713 226346 238719
rect 226294 238655 226346 238661
rect 225910 236271 225962 236277
rect 225910 236213 225962 236219
rect 225812 236162 225868 236171
rect 225812 236097 225868 236106
rect 225922 233470 225950 236213
rect 226306 233470 226334 238655
rect 227254 238639 227306 238645
rect 227254 238581 227306 238587
rect 226870 238491 226922 238497
rect 226870 238433 226922 238439
rect 226882 233484 226910 238433
rect 227266 233484 227294 238581
rect 227444 238234 227500 238243
rect 227500 238192 227678 238220
rect 227444 238169 227500 238178
rect 227650 238095 227678 238192
rect 227636 238086 227692 238095
rect 227636 238021 227692 238030
rect 227350 237455 227402 237461
rect 227350 237397 227402 237403
rect 226656 233456 226910 233484
rect 227040 233456 227294 233484
rect 214292 233433 214348 233442
rect 227362 233336 227390 237397
rect 227444 237050 227500 237059
rect 227500 237008 227678 237036
rect 227444 236985 227500 236994
rect 227650 236763 227678 237008
rect 227636 236754 227692 236763
rect 227636 236689 227692 236698
rect 227746 233470 227774 238877
rect 227938 234723 227966 242928
rect 228034 239755 228062 246494
rect 228130 245749 228158 246753
rect 228322 246119 228350 246753
rect 228310 246113 228362 246119
rect 228310 246055 228362 246061
rect 228118 245743 228170 245749
rect 228118 245685 228170 245691
rect 228514 243529 228542 246494
rect 228610 244861 228638 246753
rect 246164 246753 246220 246762
rect 246452 246818 246508 246827
rect 246452 246753 246508 246762
rect 247316 246818 247372 246827
rect 247316 246753 247372 246762
rect 247796 246818 247852 246827
rect 248180 246818 248236 246827
rect 247796 246753 247852 246762
rect 247894 246779 247946 246785
rect 231862 246721 231914 246727
rect 231382 246631 231434 246637
rect 231382 246573 231434 246579
rect 228864 246480 229214 246508
rect 229344 246480 229598 246508
rect 228598 244855 228650 244861
rect 228598 244797 228650 244803
rect 228502 243523 228554 243529
rect 228502 243465 228554 243471
rect 229186 241772 229214 246480
rect 229270 246261 229322 246267
rect 229270 246203 229322 246209
rect 229282 245897 229310 246203
rect 229270 245891 229322 245897
rect 229270 245833 229322 245839
rect 229186 241744 229406 241772
rect 229174 241599 229226 241605
rect 229174 241541 229226 241547
rect 228022 239749 228074 239755
rect 228022 239691 228074 239697
rect 229078 239675 229130 239681
rect 229078 239617 229130 239623
rect 228118 239009 228170 239015
rect 228118 238951 228170 238957
rect 227926 234717 227978 234723
rect 227926 234659 227978 234665
rect 228130 233470 228158 238951
rect 228502 237751 228554 237757
rect 228502 237693 228554 237699
rect 228514 233470 228542 237693
rect 229090 233484 229118 239617
rect 229186 233780 229214 241541
rect 229186 233752 229262 233780
rect 228864 233456 229118 233484
rect 229234 233470 229262 233752
rect 229378 233484 229406 241744
rect 229570 236023 229598 246480
rect 229762 243381 229790 246494
rect 229750 243375 229802 243381
rect 229750 243317 229802 243323
rect 229942 239749 229994 239755
rect 229942 239691 229994 239697
rect 229556 236014 229612 236023
rect 229556 235949 229612 235958
rect 229378 233456 229632 233484
rect 229954 233470 229982 239691
rect 230242 239681 230270 246494
rect 230326 239897 230378 239903
rect 230326 239839 230378 239845
rect 230230 239675 230282 239681
rect 230230 239617 230282 239623
rect 230338 233470 230366 239839
rect 230626 234797 230654 246494
rect 230818 246480 231072 246508
rect 230710 241229 230762 241235
rect 230710 241171 230762 241177
rect 230614 234791 230666 234797
rect 230614 234733 230666 234739
rect 230722 233470 230750 241171
rect 230818 237757 230846 246480
rect 230902 246409 230954 246415
rect 230902 246351 230954 246357
rect 230914 246267 230942 246351
rect 230902 246261 230954 246267
rect 230902 246203 230954 246209
rect 231394 245601 231422 246573
rect 231552 246480 231806 246508
rect 231382 245595 231434 245601
rect 231382 245537 231434 245543
rect 231778 243677 231806 246480
rect 231874 245823 231902 246721
rect 232150 246705 232202 246711
rect 232150 246647 232202 246653
rect 231862 245817 231914 245823
rect 231862 245759 231914 245765
rect 231862 245373 231914 245379
rect 231862 245315 231914 245321
rect 231874 245157 231902 245315
rect 231862 245151 231914 245157
rect 231862 245093 231914 245099
rect 231670 243671 231722 243677
rect 231670 243613 231722 243619
rect 231766 243671 231818 243677
rect 231766 243613 231818 243619
rect 231682 242979 231710 243613
rect 231668 242970 231724 242979
rect 231668 242905 231724 242914
rect 231190 241007 231242 241013
rect 231190 240949 231242 240955
rect 230902 240933 230954 240939
rect 230902 240875 230954 240881
rect 230806 237751 230858 237757
rect 230806 237693 230858 237699
rect 230914 233484 230942 240875
rect 231202 233484 231230 240949
rect 231574 240785 231626 240791
rect 231574 240727 231626 240733
rect 231586 233484 231614 240727
rect 231970 239015 231998 246494
rect 232162 245675 232190 246647
rect 232150 245669 232202 245675
rect 232150 245611 232202 245617
rect 232354 240051 232382 246494
rect 232534 241525 232586 241531
rect 232534 241467 232586 241473
rect 232342 240045 232394 240051
rect 232342 239987 232394 239993
rect 232150 239971 232202 239977
rect 232150 239913 232202 239919
rect 231958 239009 232010 239015
rect 231958 238951 232010 238957
rect 230914 233456 231072 233484
rect 231202 233456 231456 233484
rect 231586 233456 231840 233484
rect 232162 233470 232190 239913
rect 232546 233470 232574 241467
rect 232834 238941 232862 246494
rect 233280 246480 233534 246508
rect 233506 241827 233534 246480
rect 233602 246480 233760 246508
rect 233494 241821 233546 241827
rect 233494 241763 233546 241769
rect 232918 241081 232970 241087
rect 232918 241023 232970 241029
rect 232822 238935 232874 238941
rect 232822 238877 232874 238883
rect 232930 233470 232958 241023
rect 233302 240859 233354 240865
rect 233302 240801 233354 240807
rect 233314 233484 233342 240801
rect 233398 240489 233450 240495
rect 233398 240431 233450 240437
rect 233280 233456 233342 233484
rect 233410 233484 233438 240431
rect 233602 237461 233630 246480
rect 233782 241673 233834 241679
rect 233782 241615 233834 241621
rect 233590 237455 233642 237461
rect 233590 237397 233642 237403
rect 233794 233484 233822 241615
rect 234082 238645 234110 246494
rect 234562 241901 234590 246494
rect 234454 241895 234506 241901
rect 234454 241837 234506 241843
rect 234550 241895 234602 241901
rect 234550 241837 234602 241843
rect 234358 241747 234410 241753
rect 234358 241689 234410 241695
rect 234070 238639 234122 238645
rect 234070 238581 234122 238587
rect 233410 233456 233664 233484
rect 233794 233456 234048 233484
rect 234370 233470 234398 241689
rect 234466 233484 234494 241837
rect 235042 238497 235070 246494
rect 235488 246480 235550 246508
rect 235126 244337 235178 244343
rect 235126 244279 235178 244285
rect 235030 238491 235082 238497
rect 235030 238433 235082 238439
rect 234466 233456 234768 233484
rect 235138 233470 235166 244279
rect 235522 239385 235550 246480
rect 235618 246480 235872 246508
rect 235510 239379 235562 239385
rect 235510 239321 235562 239327
rect 235618 238719 235646 246480
rect 236182 246039 236234 246045
rect 236182 245981 236234 245987
rect 236194 245601 236222 245981
rect 236182 245595 236234 245601
rect 236182 245537 236234 245543
rect 236290 243603 236318 246494
rect 236278 243597 236330 243603
rect 236278 243539 236330 243545
rect 236566 240267 236618 240273
rect 236566 240209 236618 240215
rect 235606 238713 235658 238719
rect 235606 238655 235658 238661
rect 236470 236641 236522 236647
rect 236470 236583 236522 236589
rect 235702 235901 235754 235907
rect 235702 235843 235754 235849
rect 235714 233484 235742 235843
rect 236086 235457 236138 235463
rect 236086 235399 236138 235405
rect 236098 233484 236126 235399
rect 236482 233484 236510 236583
rect 235488 233456 235742 233484
rect 235872 233456 236126 233484
rect 236256 233456 236510 233484
rect 236578 233470 236606 240209
rect 236770 236277 236798 246494
rect 237154 239459 237182 246494
rect 237346 246480 237600 246508
rect 238080 246480 238334 246508
rect 237142 239453 237194 239459
rect 237142 239395 237194 239401
rect 237346 237165 237374 246480
rect 238306 242197 238334 246480
rect 238294 242191 238346 242197
rect 238294 242133 238346 242139
rect 237430 241747 237482 241753
rect 237430 241689 237482 241695
rect 237334 237159 237386 237165
rect 237334 237101 237386 237107
rect 236758 236271 236810 236277
rect 236758 236213 236810 236219
rect 236950 236271 237002 236277
rect 236950 236213 237002 236219
rect 236962 233470 236990 236213
rect 237442 233484 237470 241689
rect 238390 241155 238442 241161
rect 238390 241097 238442 241103
rect 237526 241081 237578 241087
rect 237526 241023 237578 241029
rect 237538 240125 237566 241023
rect 237814 240859 237866 240865
rect 237814 240801 237866 240807
rect 237718 240785 237770 240791
rect 237718 240727 237770 240733
rect 237730 240347 237758 240727
rect 237718 240341 237770 240347
rect 237718 240283 237770 240289
rect 237826 240199 237854 240801
rect 237814 240193 237866 240199
rect 237814 240135 237866 240141
rect 237526 240119 237578 240125
rect 237526 240061 237578 240067
rect 237910 240119 237962 240125
rect 237910 240061 237962 240067
rect 237922 233484 237950 240061
rect 238198 240045 238250 240051
rect 238198 239987 238250 239993
rect 238294 240045 238346 240051
rect 238294 239987 238346 239993
rect 238210 234395 238238 239987
rect 238196 234386 238252 234395
rect 238196 234321 238252 234330
rect 238306 233484 238334 239987
rect 237360 233456 237470 233484
rect 237696 233456 237950 233484
rect 238080 233456 238334 233484
rect 238402 233484 238430 241097
rect 238498 239163 238526 246494
rect 238594 246480 238896 246508
rect 238486 239157 238538 239163
rect 238486 239099 238538 239105
rect 238594 236869 238622 246480
rect 239362 243751 239390 246494
rect 239458 246480 239808 246508
rect 239350 243745 239402 243751
rect 239350 243687 239402 243693
rect 238966 242117 239018 242123
rect 238966 242059 239018 242065
rect 238978 241827 239006 242059
rect 238966 241821 239018 241827
rect 238966 241763 239018 241769
rect 239158 241451 239210 241457
rect 239158 241393 239210 241399
rect 238966 240341 239018 240347
rect 238966 240283 239018 240289
rect 238870 240267 238922 240273
rect 238870 240209 238922 240215
rect 238678 239379 238730 239385
rect 238678 239321 238730 239327
rect 238582 236863 238634 236869
rect 238582 236805 238634 236811
rect 238690 234543 238718 239321
rect 238774 237455 238826 237461
rect 238774 237397 238826 237403
rect 238676 234534 238732 234543
rect 238676 234469 238732 234478
rect 238402 233456 238464 233484
rect 238786 233470 238814 237397
rect 238882 236647 238910 240209
rect 238870 236641 238922 236647
rect 238870 236583 238922 236589
rect 238978 236277 239006 240283
rect 239060 238086 239116 238095
rect 239060 238021 239116 238030
rect 239074 237535 239102 238021
rect 239062 237529 239114 237535
rect 239062 237471 239114 237477
rect 239062 236789 239114 236795
rect 239060 236754 239062 236763
rect 239114 236754 239116 236763
rect 239060 236689 239116 236698
rect 238966 236271 239018 236277
rect 238966 236213 239018 236219
rect 239170 233470 239198 241393
rect 239458 238793 239486 246480
rect 240274 246212 240302 246494
rect 240418 246480 240672 246508
rect 240274 246184 240350 246212
rect 240322 240717 240350 246184
rect 240310 240711 240362 240717
rect 240310 240653 240362 240659
rect 240118 239009 240170 239015
rect 240118 238951 240170 238957
rect 239446 238787 239498 238793
rect 239446 238729 239498 238735
rect 239542 238787 239594 238793
rect 239542 238729 239594 238735
rect 239554 233470 239582 238729
rect 240130 233484 240158 238951
rect 240418 237017 240446 246480
rect 241090 241901 241118 246494
rect 241078 241895 241130 241901
rect 241078 241837 241130 241843
rect 240980 240454 241036 240463
rect 240886 240415 240938 240421
rect 240980 240389 241036 240398
rect 240886 240357 240938 240363
rect 240502 238935 240554 238941
rect 240502 238877 240554 238883
rect 240406 237011 240458 237017
rect 240406 236953 240458 236959
rect 240514 233484 240542 238877
rect 240898 233484 240926 240357
rect 239904 233456 240158 233484
rect 240288 233456 240542 233484
rect 240672 233456 240926 233484
rect 240994 233470 241022 240389
rect 241364 238234 241420 238243
rect 241364 238169 241420 238178
rect 241378 233470 241406 238169
rect 241570 237831 241598 246494
rect 242016 246480 242078 246508
rect 241940 242378 241996 242387
rect 241940 242313 241942 242322
rect 241994 242313 241996 242322
rect 241942 242281 241994 242287
rect 241748 240602 241804 240611
rect 241748 240537 241804 240546
rect 241654 239157 241706 239163
rect 241654 239099 241706 239105
rect 241558 237825 241610 237831
rect 241558 237767 241610 237773
rect 241666 234871 241694 239099
rect 241654 234865 241706 234871
rect 241654 234807 241706 234813
rect 241762 233470 241790 240537
rect 241846 239453 241898 239459
rect 241846 239395 241898 239401
rect 241858 235093 241886 239395
rect 242050 235167 242078 246480
rect 242146 246480 242400 246508
rect 242626 246480 242880 246508
rect 242146 237979 242174 246480
rect 242324 242378 242380 242387
rect 242324 242313 242326 242322
rect 242378 242313 242380 242322
rect 242326 242281 242378 242287
rect 242324 238530 242380 238539
rect 242324 238465 242380 238474
rect 242134 237973 242186 237979
rect 242134 237915 242186 237921
rect 242038 235161 242090 235167
rect 242038 235103 242090 235109
rect 241846 235087 241898 235093
rect 241846 235029 241898 235035
rect 242338 233484 242366 238465
rect 242626 238127 242654 246480
rect 243188 241046 243244 241055
rect 243188 240981 243244 240990
rect 242708 240750 242764 240759
rect 242708 240685 242764 240694
rect 242614 238121 242666 238127
rect 242614 238063 242666 238069
rect 242722 233484 242750 240685
rect 243092 237346 243148 237355
rect 243092 237281 243148 237290
rect 243106 233484 243134 237281
rect 242112 233456 242366 233484
rect 242496 233456 242750 233484
rect 242880 233456 243134 233484
rect 243202 233470 243230 240981
rect 243298 235019 243326 246494
rect 243572 238678 243628 238687
rect 243572 238613 243628 238622
rect 243286 235013 243338 235019
rect 243286 234955 243338 234961
rect 243586 233470 243614 238613
rect 243778 237905 243806 246494
rect 244176 246480 244478 246508
rect 244450 242271 244478 246480
rect 244594 246212 244622 246494
rect 244834 246480 245088 246508
rect 244594 246184 244670 246212
rect 244438 242265 244490 242271
rect 244438 242207 244490 242213
rect 244532 241194 244588 241203
rect 244532 241129 244588 241138
rect 244150 240711 244202 240717
rect 244150 240653 244202 240659
rect 243766 237899 243818 237905
rect 243766 237841 243818 237847
rect 243956 237494 244012 237503
rect 243956 237429 244012 237438
rect 243970 233470 243998 237429
rect 244162 234945 244190 240653
rect 244150 234939 244202 234945
rect 244150 234881 244202 234887
rect 244546 233484 244574 241129
rect 244642 239977 244670 246184
rect 244726 241303 244778 241309
rect 244726 241245 244778 241251
rect 244630 239971 244682 239977
rect 244630 239913 244682 239919
rect 244738 233780 244766 241245
rect 244834 238053 244862 246480
rect 245410 243825 245438 246494
rect 245398 243819 245450 243825
rect 245398 243761 245450 243767
rect 245396 241786 245452 241795
rect 245396 241721 245452 241730
rect 244822 238047 244874 238053
rect 244822 237989 244874 237995
rect 245300 237198 245356 237207
rect 245300 237133 245356 237142
rect 244320 233456 244574 233484
rect 244690 233752 244766 233780
rect 244690 233470 244718 233752
rect 245314 233484 245342 237133
rect 245088 233456 245342 233484
rect 245410 233470 245438 241721
rect 245890 237683 245918 246494
rect 246178 245453 246206 246753
rect 246262 245891 246314 245897
rect 246262 245833 246314 245839
rect 246166 245447 246218 245453
rect 246166 245389 246218 245395
rect 246274 245379 246302 245833
rect 246262 245373 246314 245379
rect 246262 245315 246314 245321
rect 246070 239971 246122 239977
rect 246070 239913 246122 239919
rect 245878 237677 245930 237683
rect 245878 237619 245930 237625
rect 245782 237603 245834 237609
rect 245782 237545 245834 237551
rect 245794 233470 245822 237545
rect 246082 235389 246110 239913
rect 246166 237677 246218 237683
rect 246166 237619 246218 237625
rect 246070 235383 246122 235389
rect 246070 235325 246122 235331
rect 246178 233470 246206 237619
rect 246370 235241 246398 246494
rect 246466 245675 246494 246753
rect 247330 246563 247358 246753
rect 247318 246557 247370 246563
rect 246562 246480 246816 246508
rect 247318 246499 247370 246505
rect 246454 245669 246506 245675
rect 246454 245611 246506 245617
rect 246562 237313 246590 246480
rect 247186 246212 247214 246494
rect 247186 246184 247262 246212
rect 246740 241638 246796 241647
rect 246740 241573 246796 241582
rect 246550 237307 246602 237313
rect 246550 237249 246602 237255
rect 246358 235235 246410 235241
rect 246358 235177 246410 235183
rect 246754 233484 246782 241573
rect 247126 237825 247178 237831
rect 247126 237767 247178 237773
rect 247138 233484 247166 237767
rect 247234 237387 247262 246184
rect 247318 242561 247370 242567
rect 247316 242526 247318 242535
rect 247370 242526 247372 242535
rect 247316 242461 247372 242470
rect 247618 241328 247646 246494
rect 247810 246415 247838 246753
rect 248372 246818 248428 246827
rect 248180 246753 248182 246762
rect 247894 246721 247946 246727
rect 248234 246753 248236 246762
rect 248278 246779 248330 246785
rect 248182 246721 248234 246727
rect 260948 246818 261004 246827
rect 248372 246753 248428 246762
rect 251926 246779 251978 246785
rect 248278 246721 248330 246727
rect 247798 246409 247850 246415
rect 247798 246351 247850 246357
rect 247906 245897 247934 246721
rect 248182 246631 248234 246637
rect 248182 246573 248234 246579
rect 247894 245891 247946 245897
rect 247894 245833 247946 245839
rect 247798 242857 247850 242863
rect 247798 242799 247850 242805
rect 247810 242535 247838 242799
rect 247796 242526 247852 242535
rect 247796 242461 247852 242470
rect 247618 241300 247838 241328
rect 247700 240158 247756 240167
rect 247700 240093 247756 240102
rect 247714 238220 247742 240093
rect 247522 238192 247742 238220
rect 247222 237381 247274 237387
rect 247222 237323 247274 237329
rect 247522 233484 247550 238192
rect 247606 237751 247658 237757
rect 247606 237693 247658 237699
rect 246528 233456 246782 233484
rect 246912 233456 247166 233484
rect 247296 233456 247550 233484
rect 247618 233470 247646 237693
rect 247810 235315 247838 241300
rect 248098 240495 248126 246494
rect 248194 245823 248222 246573
rect 248290 246045 248318 246721
rect 248278 246039 248330 246045
rect 248278 245981 248330 245987
rect 248182 245817 248234 245823
rect 248182 245759 248234 245765
rect 248386 245453 248414 246753
rect 260948 246753 261004 246762
rect 269204 246818 269260 246827
rect 281300 246818 281356 246827
rect 269204 246753 269260 246762
rect 276886 246779 276938 246785
rect 251926 246721 251978 246727
rect 248374 245447 248426 245453
rect 248374 245389 248426 245395
rect 248086 240489 248138 240495
rect 248086 240431 248138 240437
rect 248374 240489 248426 240495
rect 248374 240431 248426 240437
rect 247988 240010 248044 240019
rect 247988 239945 248044 239954
rect 247798 235309 247850 235315
rect 247798 235251 247850 235257
rect 248002 233470 248030 239945
rect 248386 233470 248414 240431
rect 248578 239755 248606 246494
rect 248674 246480 248928 246508
rect 249046 246483 249098 246489
rect 248674 240643 248702 246480
rect 249408 246480 249662 246508
rect 249046 246425 249098 246431
rect 249058 245601 249086 246425
rect 249142 246113 249194 246119
rect 249142 246055 249194 246061
rect 249046 245595 249098 245601
rect 249046 245537 249098 245543
rect 249154 245379 249182 246055
rect 249634 245379 249662 246480
rect 249142 245373 249194 245379
rect 249142 245315 249194 245321
rect 249622 245373 249674 245379
rect 249622 245315 249674 245321
rect 248662 240637 248714 240643
rect 248662 240579 248714 240585
rect 249826 240569 249854 246494
rect 250306 245305 250334 246494
rect 250294 245299 250346 245305
rect 250294 245241 250346 245247
rect 250690 240939 250718 246494
rect 251136 246480 251390 246508
rect 251616 246480 251870 246508
rect 251362 245749 251390 246480
rect 251734 245965 251786 245971
rect 251734 245907 251786 245913
rect 251350 245743 251402 245749
rect 251350 245685 251402 245691
rect 251746 245527 251774 245907
rect 251734 245521 251786 245527
rect 251734 245463 251786 245469
rect 251842 241901 251870 246480
rect 251938 245897 251966 246721
rect 252118 246631 252170 246637
rect 252118 246573 252170 246579
rect 258658 246628 258960 246656
rect 251926 245891 251978 245897
rect 251926 245833 251978 245839
rect 251830 241895 251882 241901
rect 251830 241837 251882 241843
rect 250678 240933 250730 240939
rect 250678 240875 250730 240881
rect 252034 240791 252062 246494
rect 252130 245823 252158 246573
rect 252118 245817 252170 245823
rect 252118 245759 252170 245765
rect 252418 245527 252446 246494
rect 252406 245521 252458 245527
rect 252406 245463 252458 245469
rect 252790 241673 252842 241679
rect 252790 241615 252842 241621
rect 252310 240933 252362 240939
rect 252310 240875 252362 240881
rect 252022 240785 252074 240791
rect 252022 240727 252074 240733
rect 251542 240711 251594 240717
rect 251542 240653 251594 240659
rect 250582 240637 250634 240643
rect 250582 240579 250634 240585
rect 249814 240563 249866 240569
rect 249814 240505 249866 240511
rect 250198 240563 250250 240569
rect 250198 240505 250250 240511
rect 249718 239971 249770 239977
rect 249718 239913 249770 239919
rect 248566 239749 248618 239755
rect 248566 239691 248618 239697
rect 248950 238639 249002 238645
rect 248950 238581 249002 238587
rect 248962 233484 248990 238581
rect 249334 237899 249386 237905
rect 249334 237841 249386 237847
rect 249346 233484 249374 237841
rect 249730 233484 249758 239913
rect 249814 237973 249866 237979
rect 249814 237915 249866 237921
rect 248736 233456 248990 233484
rect 249120 233456 249374 233484
rect 249504 233456 249758 233484
rect 249826 233470 249854 237915
rect 250210 233470 250238 240505
rect 250594 233470 250622 240579
rect 251158 238047 251210 238053
rect 251158 237989 251210 237995
rect 251170 233484 251198 237989
rect 251554 233484 251582 240653
rect 251926 238121 251978 238127
rect 251926 238063 251978 238069
rect 251938 233484 251966 238063
rect 252322 233484 252350 240875
rect 252406 238195 252458 238201
rect 252406 238137 252458 238143
rect 250944 233456 251198 233484
rect 251328 233456 251582 233484
rect 251712 233456 251966 233484
rect 252048 233456 252350 233484
rect 252418 233470 252446 238137
rect 252802 233470 252830 241615
rect 252898 240865 252926 246494
rect 253344 246480 253406 246508
rect 253378 245453 253406 246480
rect 253474 246480 253728 246508
rect 253366 245447 253418 245453
rect 253366 245389 253418 245395
rect 252886 240859 252938 240865
rect 252886 240801 252938 240807
rect 253474 238349 253502 246480
rect 254146 245749 254174 246494
rect 254134 245743 254186 245749
rect 254134 245685 254186 245691
rect 253750 241229 253802 241235
rect 253750 241171 253802 241177
rect 253462 238343 253514 238349
rect 253462 238285 253514 238291
rect 253366 238269 253418 238275
rect 253366 238211 253418 238217
rect 253378 233484 253406 238211
rect 253762 233484 253790 241171
rect 254230 241155 254282 241161
rect 254230 241097 254282 241103
rect 254134 238491 254186 238497
rect 254134 238433 254186 238439
rect 254146 233484 254174 238433
rect 253152 233456 253406 233484
rect 253536 233456 253790 233484
rect 253920 233456 254174 233484
rect 254242 233470 254270 241097
rect 254626 241087 254654 246494
rect 255106 245823 255134 246494
rect 255202 246480 255456 246508
rect 255682 246480 255936 246508
rect 255094 245817 255146 245823
rect 255094 245759 255146 245765
rect 254998 241525 255050 241531
rect 254998 241467 255050 241473
rect 254614 241081 254666 241087
rect 254614 241023 254666 241029
rect 254614 238417 254666 238423
rect 254614 238359 254666 238365
rect 254626 233470 254654 238359
rect 255010 233470 255038 241467
rect 255202 238571 255230 246480
rect 255478 240785 255530 240791
rect 255478 240727 255530 240733
rect 255490 240347 255518 240727
rect 255478 240341 255530 240347
rect 255478 240283 255530 240289
rect 255682 238941 255710 246480
rect 256354 244047 256382 246494
rect 256342 244041 256394 244047
rect 256342 243983 256394 243989
rect 255958 241377 256010 241383
rect 255958 241319 256010 241325
rect 255670 238935 255722 238941
rect 255670 238877 255722 238883
rect 255190 238565 255242 238571
rect 255190 238507 255242 238513
rect 255574 238565 255626 238571
rect 255574 238507 255626 238513
rect 255586 233484 255614 238507
rect 255970 233484 255998 241319
rect 256438 239897 256490 239903
rect 256438 239839 256490 239845
rect 256246 238713 256298 238719
rect 256246 238655 256298 238661
rect 256258 233484 256286 238655
rect 255360 233456 255614 233484
rect 255744 233456 255998 233484
rect 256128 233456 256286 233484
rect 256450 233470 256478 239839
rect 256834 239015 256862 246494
rect 257232 246480 257342 246508
rect 257206 239823 257258 239829
rect 257206 239765 257258 239771
rect 256822 239009 256874 239015
rect 256822 238951 256874 238957
rect 256822 238861 256874 238867
rect 256822 238803 256874 238809
rect 256834 233470 256862 238803
rect 257218 233470 257246 239765
rect 257314 235537 257342 246480
rect 257410 246480 257664 246508
rect 258144 246480 258398 246508
rect 257410 238793 257438 246480
rect 258370 244195 258398 246480
rect 258358 244189 258410 244195
rect 258358 244131 258410 244137
rect 258562 241457 258590 246494
rect 258550 241451 258602 241457
rect 258550 241393 258602 241399
rect 257686 241007 257738 241013
rect 257686 240949 257738 240955
rect 257698 240421 257726 240949
rect 257878 240637 257930 240643
rect 257878 240579 257930 240585
rect 257686 240415 257738 240421
rect 257686 240357 257738 240363
rect 257890 239977 257918 240579
rect 257878 239971 257930 239977
rect 257878 239913 257930 239919
rect 258658 239089 258686 246628
rect 259126 246483 259178 246489
rect 259126 246425 259178 246431
rect 259138 246045 259166 246425
rect 259126 246039 259178 246045
rect 259126 245981 259178 245987
rect 259028 240898 259084 240907
rect 259028 240833 259084 240842
rect 258646 239083 258698 239089
rect 258646 239025 258698 239031
rect 258934 239083 258986 239089
rect 258934 239025 258986 239031
rect 257398 238787 257450 238793
rect 257398 238729 257450 238735
rect 257782 238787 257834 238793
rect 257782 238729 257834 238735
rect 257302 235531 257354 235537
rect 257302 235473 257354 235479
rect 257794 233484 257822 238729
rect 258644 238382 258700 238391
rect 258550 238343 258602 238349
rect 258644 238317 258700 238326
rect 258550 238285 258602 238291
rect 258166 236567 258218 236573
rect 258166 236509 258218 236515
rect 258178 233484 258206 236509
rect 258562 233484 258590 238285
rect 257568 233456 257822 233484
rect 257952 233456 258206 233484
rect 258336 233456 258590 233484
rect 258658 233470 258686 238317
rect 258946 235685 258974 239025
rect 258934 235679 258986 235685
rect 258934 235621 258986 235627
rect 259042 233470 259070 240833
rect 259124 238086 259180 238095
rect 259124 238021 259180 238030
rect 259138 237535 259166 238021
rect 259126 237529 259178 237535
rect 259126 237471 259178 237477
rect 259426 237461 259454 246494
rect 259872 246480 260126 246508
rect 260352 246480 260606 246508
rect 260098 243973 260126 246480
rect 260374 246113 260426 246119
rect 260374 246055 260426 246061
rect 260278 245151 260330 245157
rect 260278 245093 260330 245099
rect 260290 244861 260318 245093
rect 260278 244855 260330 244861
rect 260278 244797 260330 244803
rect 260086 243967 260138 243973
rect 260086 243909 260138 243915
rect 260386 243159 260414 246055
rect 260374 243153 260426 243159
rect 260374 243095 260426 243101
rect 259604 239862 259660 239871
rect 259604 239797 259660 239806
rect 259414 237455 259466 237461
rect 259414 237397 259466 237403
rect 259126 236789 259178 236795
rect 259124 236754 259126 236763
rect 259178 236754 259180 236763
rect 259124 236689 259180 236698
rect 259618 233484 259646 239797
rect 260374 239009 260426 239015
rect 260374 238951 260426 238957
rect 259990 238935 260042 238941
rect 259990 238877 260042 238883
rect 260002 233484 260030 238877
rect 260386 233484 260414 238951
rect 260578 235611 260606 246480
rect 260674 240051 260702 246494
rect 260758 246409 260810 246415
rect 260758 246351 260810 246357
rect 260770 244269 260798 246351
rect 260854 246261 260906 246267
rect 260854 246203 260906 246209
rect 260758 244263 260810 244269
rect 260758 244205 260810 244211
rect 260866 243011 260894 246203
rect 260962 244787 260990 246753
rect 260950 244781 261002 244787
rect 260950 244723 261002 244729
rect 261154 244121 261182 246494
rect 261142 244115 261194 244121
rect 261142 244057 261194 244063
rect 260854 243005 260906 243011
rect 260854 242947 260906 242953
rect 261236 241342 261292 241351
rect 261236 241277 261292 241286
rect 260662 240045 260714 240051
rect 260662 239987 260714 239993
rect 260758 240045 260810 240051
rect 260758 239987 260810 239993
rect 260770 239755 260798 239987
rect 260758 239749 260810 239755
rect 260758 239691 260810 239697
rect 260758 236715 260810 236721
rect 260758 236657 260810 236663
rect 260566 235605 260618 235611
rect 260566 235547 260618 235553
rect 260770 233484 260798 236657
rect 260854 234643 260906 234649
rect 260854 234585 260906 234591
rect 259440 233456 259646 233484
rect 259776 233456 260030 233484
rect 260160 233456 260414 233484
rect 260544 233456 260798 233484
rect 260866 233470 260894 234585
rect 261250 233470 261278 241277
rect 261634 240125 261662 246494
rect 261970 246212 261998 246494
rect 261922 246184 261998 246212
rect 262210 246480 262464 246508
rect 261814 245151 261866 245157
rect 261814 245093 261866 245099
rect 261622 240119 261674 240125
rect 261622 240061 261674 240067
rect 261826 233484 261854 245093
rect 261922 235759 261950 246184
rect 262210 241753 262238 246480
rect 262882 244713 262910 246494
rect 262870 244707 262922 244713
rect 262870 244649 262922 244655
rect 262198 241747 262250 241753
rect 262198 241689 262250 241695
rect 263362 240791 263390 246494
rect 263446 245077 263498 245083
rect 263446 245019 263498 245025
rect 263350 240785 263402 240791
rect 263350 240727 263402 240733
rect 262964 240306 263020 240315
rect 262006 240267 262058 240273
rect 262964 240241 263020 240250
rect 262006 240209 262058 240215
rect 261910 235753 261962 235759
rect 261910 235695 261962 235701
rect 262018 233484 262046 240209
rect 262342 233755 262394 233761
rect 262342 233697 262394 233703
rect 261648 233456 261854 233484
rect 261984 233456 262046 233484
rect 262354 233470 262382 233697
rect 262978 233484 263006 240241
rect 263062 236419 263114 236425
rect 263062 236361 263114 236367
rect 262752 233456 263006 233484
rect 263074 233470 263102 236361
rect 263458 233470 263486 245019
rect 263746 235833 263774 246494
rect 263938 246480 264192 246508
rect 264418 246480 264672 246508
rect 263830 245003 263882 245009
rect 263830 244945 263882 244951
rect 263734 235827 263786 235833
rect 263734 235769 263786 235775
rect 263842 233470 263870 244945
rect 263938 240199 263966 246480
rect 264310 241821 264362 241827
rect 264310 241763 264362 241769
rect 263926 240193 263978 240199
rect 263926 240135 263978 240141
rect 264022 240193 264074 240199
rect 264022 240135 264074 240141
rect 264034 236573 264062 240135
rect 264022 236567 264074 236573
rect 264022 236509 264074 236515
rect 264322 233484 264350 241763
rect 264418 240347 264446 246480
rect 264790 243301 264842 243307
rect 264790 243243 264842 243249
rect 264406 240341 264458 240347
rect 264406 240283 264458 240289
rect 264802 233484 264830 243243
rect 264886 236049 264938 236055
rect 264886 235991 264938 235997
rect 264192 233456 264350 233484
rect 264576 233456 264830 233484
rect 264898 233484 264926 235991
rect 265090 235981 265118 246494
rect 265270 243079 265322 243085
rect 265270 243021 265322 243027
rect 265078 235975 265130 235981
rect 265078 235917 265130 235923
rect 264898 233456 264960 233484
rect 265282 233470 265310 243021
rect 265474 235463 265502 246494
rect 265954 244639 265982 246494
rect 266146 246480 266400 246508
rect 266818 246480 266880 246508
rect 265942 244633 265994 244639
rect 265942 244575 265994 244581
rect 266038 242931 266090 242937
rect 266038 242873 266090 242879
rect 265654 236123 265706 236129
rect 265654 236065 265706 236071
rect 265462 235457 265514 235463
rect 265462 235399 265514 235405
rect 265666 233470 265694 236065
rect 266050 233470 266078 242873
rect 266146 235907 266174 246480
rect 266614 242857 266666 242863
rect 266614 242799 266666 242805
rect 266134 235901 266186 235907
rect 266134 235843 266186 235849
rect 266626 233484 266654 242799
rect 266818 235907 266846 246480
rect 267202 244343 267230 246494
rect 267696 246480 267998 246508
rect 268176 246480 268382 246508
rect 268512 246480 268766 246508
rect 267970 246249 267998 246480
rect 268054 246409 268106 246415
rect 268106 246357 268286 246360
rect 268054 246351 268286 246357
rect 268066 246341 268286 246351
rect 268066 246335 268298 246341
rect 268066 246332 268246 246335
rect 268246 246277 268298 246283
rect 267970 246221 268286 246249
rect 268150 246187 268202 246193
rect 268150 246129 268202 246135
rect 267490 245703 267902 245731
rect 267490 245675 267518 245703
rect 267478 245669 267530 245675
rect 267478 245611 267530 245617
rect 267478 245003 267530 245009
rect 267478 244945 267530 244951
rect 267490 244565 267518 244945
rect 267478 244559 267530 244565
rect 267478 244501 267530 244507
rect 267190 244337 267242 244343
rect 267190 244279 267242 244285
rect 267874 244177 267902 245703
rect 267958 244855 268010 244861
rect 267958 244797 268010 244803
rect 268054 244855 268106 244861
rect 268054 244797 268106 244803
rect 267970 244491 267998 244797
rect 268066 244565 268094 244797
rect 268054 244559 268106 244565
rect 268054 244501 268106 244507
rect 267958 244485 268010 244491
rect 267958 244427 268010 244433
rect 268162 244269 268190 246129
rect 268258 244269 268286 246221
rect 268150 244263 268202 244269
rect 268150 244205 268202 244211
rect 268246 244263 268298 244269
rect 268246 244205 268298 244211
rect 267874 244149 268190 244177
rect 268162 243899 268190 244149
rect 268054 243893 268106 243899
rect 268054 243835 268106 243841
rect 268150 243893 268202 243899
rect 268150 243835 268202 243841
rect 267956 243710 268012 243719
rect 267956 243645 268012 243654
rect 267382 243227 267434 243233
rect 267382 243169 267434 243175
rect 266806 235901 266858 235907
rect 266806 235843 266858 235849
rect 266998 234569 267050 234575
rect 266998 234511 267050 234517
rect 267010 233484 267038 234511
rect 267394 233484 267422 243169
rect 267766 242709 267818 242715
rect 267766 242651 267818 242657
rect 267778 242535 267806 242651
rect 267970 242535 267998 243645
rect 268066 242789 268094 243835
rect 268244 242970 268300 242979
rect 268244 242905 268300 242914
rect 268054 242783 268106 242789
rect 268054 242725 268106 242731
rect 268258 242715 268286 242905
rect 268246 242709 268298 242715
rect 268246 242651 268298 242657
rect 268150 242561 268202 242567
rect 267764 242526 267820 242535
rect 267764 242461 267820 242470
rect 267956 242526 268012 242535
rect 268150 242503 268202 242509
rect 267956 242461 268012 242470
rect 267956 241786 268012 241795
rect 267956 241721 268012 241730
rect 267668 241490 267724 241499
rect 267586 241448 267668 241476
rect 267586 241351 267614 241448
rect 267668 241425 267724 241434
rect 267572 241342 267628 241351
rect 267572 241277 267628 241286
rect 267764 241342 267820 241351
rect 267764 241277 267820 241286
rect 267778 239871 267806 241277
rect 267764 239862 267820 239871
rect 267764 239797 267820 239806
rect 267970 239723 267998 241721
rect 267956 239714 268012 239723
rect 267956 239649 268012 239658
rect 267478 234421 267530 234427
rect 267478 234363 267530 234369
rect 266400 233456 266654 233484
rect 266784 233456 267038 233484
rect 267168 233456 267422 233484
rect 267490 233470 267518 234363
rect 268162 233484 268190 242503
rect 268246 239749 268298 239755
rect 268246 239691 268298 239697
rect 267888 233456 268190 233484
rect 268258 233470 268286 239691
rect 268354 236499 268382 246480
rect 268630 246409 268682 246415
rect 268630 246351 268682 246357
rect 268534 246261 268586 246267
rect 268534 246203 268586 246209
rect 268438 245595 268490 245601
rect 268438 245537 268490 245543
rect 268342 236493 268394 236499
rect 268342 236435 268394 236441
rect 268450 234649 268478 245537
rect 268546 243011 268574 246203
rect 268642 243159 268670 246351
rect 268630 243153 268682 243159
rect 268630 243095 268682 243101
rect 268534 243005 268586 243011
rect 268534 242947 268586 242953
rect 268738 239977 268766 246480
rect 268822 246483 268874 246489
rect 268992 246480 269150 246508
rect 268822 246425 268874 246431
rect 268834 246119 268862 246425
rect 268822 246113 268874 246119
rect 268822 246055 268874 246061
rect 268918 246113 268970 246119
rect 268918 246055 268970 246061
rect 268726 239971 268778 239977
rect 268726 239913 268778 239919
rect 268438 234643 268490 234649
rect 268438 234585 268490 234591
rect 268822 234125 268874 234131
rect 268822 234067 268874 234073
rect 268834 233484 268862 234067
rect 268930 233761 268958 246055
rect 269014 245669 269066 245675
rect 269014 245611 269066 245617
rect 269026 236425 269054 245611
rect 269014 236419 269066 236425
rect 269014 236361 269066 236367
rect 268918 233755 268970 233761
rect 268918 233697 268970 233703
rect 269122 233613 269150 246480
rect 269218 244491 269246 246753
rect 276886 246721 276938 246727
rect 280822 246779 280874 246785
rect 280822 246721 280874 246727
rect 280918 246779 280970 246785
rect 281300 246753 281356 246762
rect 284948 246818 285004 246827
rect 284948 246753 284950 246762
rect 280918 246721 280970 246727
rect 269206 244485 269258 244491
rect 269206 244427 269258 244433
rect 269206 242635 269258 242641
rect 269206 242577 269258 242583
rect 269110 233607 269162 233613
rect 269110 233549 269162 233555
rect 269218 233484 269246 242577
rect 269302 241599 269354 241605
rect 269302 241541 269354 241547
rect 269314 239829 269342 241541
rect 269410 239829 269438 246494
rect 269494 245077 269546 245083
rect 269494 245019 269546 245025
rect 269302 239823 269354 239829
rect 269302 239765 269354 239771
rect 269398 239823 269450 239829
rect 269398 239765 269450 239771
rect 269506 236721 269534 245019
rect 269890 243011 269918 246494
rect 269878 243005 269930 243011
rect 269878 242947 269930 242953
rect 269686 242709 269738 242715
rect 269686 242651 269738 242657
rect 269494 236715 269546 236721
rect 269494 236657 269546 236663
rect 269590 234051 269642 234057
rect 269590 233993 269642 233999
rect 269602 233484 269630 233993
rect 268608 233456 268862 233484
rect 268992 233456 269246 233484
rect 269376 233456 269630 233484
rect 269698 233470 269726 242651
rect 270274 239681 270302 246494
rect 270720 246480 270878 246508
rect 270850 243159 270878 246480
rect 270946 246480 271200 246508
rect 270838 243153 270890 243159
rect 270838 243095 270890 243101
rect 270946 239755 270974 246480
rect 271030 240785 271082 240791
rect 271030 240727 271082 240733
rect 270934 239749 270986 239755
rect 270934 239691 270986 239697
rect 270262 239675 270314 239681
rect 270262 239617 270314 239623
rect 270070 233755 270122 233761
rect 270070 233697 270122 233703
rect 270082 233470 270110 233697
rect 270646 233681 270698 233687
rect 270646 233623 270698 233629
rect 270658 233484 270686 233623
rect 271042 233484 271070 240727
rect 271414 236271 271466 236277
rect 271414 236213 271466 236219
rect 271426 233484 271454 236213
rect 271618 234353 271646 246494
rect 271894 242339 271946 242345
rect 271894 242281 271946 242287
rect 271906 240051 271934 242281
rect 272002 241827 272030 246494
rect 271990 241821 272042 241827
rect 271990 241763 272042 241769
rect 271894 240045 271946 240051
rect 271894 239987 271946 239993
rect 272278 239675 272330 239681
rect 272278 239617 272330 239623
rect 271798 239601 271850 239607
rect 271798 239543 271850 239549
rect 271606 234347 271658 234353
rect 271606 234289 271658 234295
rect 271810 233484 271838 239543
rect 271894 237011 271946 237017
rect 271894 236953 271946 236959
rect 270480 233456 270686 233484
rect 270816 233456 271070 233484
rect 271200 233456 271454 233484
rect 271584 233456 271838 233484
rect 271906 233470 271934 236953
rect 272290 233470 272318 239617
rect 272482 239385 272510 246494
rect 272928 246480 273182 246508
rect 273408 246480 273566 246508
rect 273792 246480 274046 246508
rect 273046 244707 273098 244713
rect 273046 244649 273098 244655
rect 273058 244343 273086 244649
rect 273046 244337 273098 244343
rect 273046 244279 273098 244285
rect 273154 241901 273182 246480
rect 273142 241895 273194 241901
rect 273142 241837 273194 241843
rect 272470 239379 272522 239385
rect 272470 239321 272522 239327
rect 273430 239231 273482 239237
rect 273430 239173 273482 239179
rect 272662 239157 272714 239163
rect 272662 239099 272714 239105
rect 272674 233470 272702 239099
rect 273238 237381 273290 237387
rect 273238 237323 273290 237329
rect 273250 233484 273278 237323
rect 273442 233780 273470 239173
rect 273538 236351 273566 246480
rect 273622 241821 273674 241827
rect 273622 241763 273674 241769
rect 273526 236345 273578 236351
rect 273526 236287 273578 236293
rect 273634 235463 273662 241763
rect 274018 240347 274046 246480
rect 274102 246483 274154 246489
rect 274102 246425 274154 246431
rect 274114 244639 274142 246425
rect 274102 244633 274154 244639
rect 274102 244575 274154 244581
rect 274102 241451 274154 241457
rect 274102 241393 274154 241399
rect 274006 240341 274058 240347
rect 274006 240283 274058 240289
rect 274114 239903 274142 241393
rect 274210 239903 274238 246494
rect 274486 241081 274538 241087
rect 274486 241023 274538 241029
rect 274102 239897 274154 239903
rect 274102 239839 274154 239845
rect 274198 239897 274250 239903
rect 274198 239839 274250 239845
rect 274006 237233 274058 237239
rect 274006 237175 274058 237181
rect 273622 235457 273674 235463
rect 273622 235399 273674 235405
rect 273024 233456 273278 233484
rect 273394 233752 273470 233780
rect 273394 233470 273422 233752
rect 274018 233484 274046 237175
rect 274102 236715 274154 236721
rect 274102 236657 274154 236663
rect 273792 233456 274046 233484
rect 274114 233470 274142 236657
rect 274498 233470 274526 241023
rect 274690 240051 274718 246494
rect 275136 246480 275390 246508
rect 275520 246480 275774 246508
rect 276000 246480 276254 246508
rect 275362 240421 275390 246480
rect 275350 240415 275402 240421
rect 275350 240357 275402 240363
rect 274678 240045 274730 240051
rect 274678 239987 274730 239993
rect 275746 239311 275774 246480
rect 276022 244707 276074 244713
rect 276022 244649 276074 244655
rect 276034 242937 276062 244649
rect 276022 242931 276074 242937
rect 276022 242873 276074 242879
rect 276226 239755 276254 246480
rect 276310 239823 276362 239829
rect 276310 239765 276362 239771
rect 276214 239749 276266 239755
rect 276214 239691 276266 239697
rect 276214 239453 276266 239459
rect 276214 239395 276266 239401
rect 275734 239305 275786 239311
rect 275734 239247 275786 239253
rect 275254 238935 275306 238941
rect 275254 238877 275306 238883
rect 275266 237535 275294 238877
rect 275254 237529 275306 237535
rect 275254 237471 275306 237477
rect 275446 237455 275498 237461
rect 275446 237397 275498 237403
rect 274870 236789 274922 236795
rect 274870 236731 274922 236737
rect 274882 233470 274910 236731
rect 275458 233484 275486 237397
rect 275830 237307 275882 237313
rect 275830 237249 275882 237255
rect 275842 233484 275870 237249
rect 276226 233484 276254 239395
rect 275232 233456 275486 233484
rect 275616 233456 275870 233484
rect 276000 233456 276254 233484
rect 276322 233470 276350 239765
rect 276418 236647 276446 246494
rect 276694 239823 276746 239829
rect 276694 239765 276746 239771
rect 276406 236641 276458 236647
rect 276406 236583 276458 236589
rect 276706 233470 276734 239765
rect 276802 236943 276830 246494
rect 276898 244565 276926 246721
rect 276982 246557 277034 246563
rect 276982 246499 277034 246505
rect 276886 244559 276938 244565
rect 276886 244501 276938 244507
rect 276994 242493 277022 246499
rect 276982 242487 277034 242493
rect 276982 242429 277034 242435
rect 277078 239527 277130 239533
rect 277078 239469 277130 239475
rect 276790 236937 276842 236943
rect 276790 236879 276842 236885
rect 277090 233470 277118 239469
rect 277282 234205 277310 246494
rect 277474 246480 277728 246508
rect 278208 246480 278462 246508
rect 278544 246480 278750 246508
rect 277366 246409 277418 246415
rect 277366 246351 277418 246357
rect 277378 245971 277406 246351
rect 277366 245965 277418 245971
rect 277366 245907 277418 245913
rect 277474 240125 277502 246480
rect 277750 246113 277802 246119
rect 277750 246055 277802 246061
rect 277558 245965 277610 245971
rect 277558 245907 277610 245913
rect 277570 245009 277598 245907
rect 277762 245601 277790 246055
rect 278038 245965 278090 245971
rect 278038 245907 278090 245913
rect 277654 245595 277706 245601
rect 277654 245537 277706 245543
rect 277750 245595 277802 245601
rect 277750 245537 277802 245543
rect 277666 245472 277694 245537
rect 277666 245444 277982 245472
rect 277954 245083 277982 245444
rect 277942 245077 277994 245083
rect 277942 245019 277994 245025
rect 277558 245003 277610 245009
rect 277558 244945 277610 244951
rect 278050 244861 278078 245907
rect 278038 244855 278090 244861
rect 278038 244797 278090 244803
rect 278134 244855 278186 244861
rect 278134 244797 278186 244803
rect 278146 244732 278174 244797
rect 278050 244704 278174 244732
rect 278050 244639 278078 244704
rect 278038 244633 278090 244639
rect 278038 244575 278090 244581
rect 278134 244633 278186 244639
rect 278134 244575 278186 244581
rect 277750 244559 277802 244565
rect 277750 244501 277802 244507
rect 277762 242845 277790 244501
rect 277846 244485 277898 244491
rect 277846 244427 277898 244433
rect 277858 243307 277886 244427
rect 277846 243301 277898 243307
rect 277846 243243 277898 243249
rect 278146 243085 278174 244575
rect 278134 243079 278186 243085
rect 278134 243021 278186 243027
rect 278038 242931 278090 242937
rect 278038 242873 278090 242879
rect 278050 242845 278078 242873
rect 277762 242817 278078 242845
rect 278326 242783 278378 242789
rect 278146 242743 278326 242771
rect 278146 242715 278174 242743
rect 278326 242725 278378 242731
rect 278134 242709 278186 242715
rect 278134 242651 278186 242657
rect 278230 241821 278282 241827
rect 278230 241763 278282 241769
rect 277654 241747 277706 241753
rect 277654 241689 277706 241695
rect 277556 240454 277612 240463
rect 277556 240389 277612 240398
rect 277462 240119 277514 240125
rect 277462 240061 277514 240067
rect 277570 239871 277598 240389
rect 277666 240199 277694 241689
rect 278132 241194 278188 241203
rect 278132 241129 278188 241138
rect 277748 241046 277804 241055
rect 277748 240981 277804 240990
rect 277762 240736 277790 240981
rect 278036 240750 278092 240759
rect 277762 240708 278036 240736
rect 278036 240685 278092 240694
rect 277654 240193 277706 240199
rect 277654 240135 277706 240141
rect 277750 240193 277802 240199
rect 277750 240135 277802 240141
rect 277556 239862 277612 239871
rect 277556 239797 277612 239806
rect 277762 239681 277790 240135
rect 278146 239723 278174 241129
rect 278242 240273 278270 241763
rect 278230 240267 278282 240273
rect 278230 240209 278282 240215
rect 278132 239714 278188 239723
rect 277750 239675 277802 239681
rect 277750 239617 277802 239623
rect 278038 239675 278090 239681
rect 278132 239649 278188 239658
rect 278038 239617 278090 239623
rect 277654 239601 277706 239607
rect 277654 239543 277706 239549
rect 277270 234199 277322 234205
rect 277270 234141 277322 234147
rect 277666 233484 277694 239543
rect 278050 233484 278078 239617
rect 278434 239015 278462 246480
rect 278422 239009 278474 239015
rect 278422 238951 278474 238957
rect 278518 237159 278570 237165
rect 278518 237101 278570 237107
rect 278422 236419 278474 236425
rect 278422 236361 278474 236367
rect 278434 233484 278462 236361
rect 277440 233456 277694 233484
rect 277824 233456 278078 233484
rect 278208 233456 278462 233484
rect 278530 233470 278558 237101
rect 278722 236573 278750 246480
rect 278804 239566 278860 239575
rect 278804 239501 278860 239510
rect 278818 239237 278846 239501
rect 278806 239231 278858 239237
rect 278806 239173 278858 239179
rect 278902 239231 278954 239237
rect 278902 239173 278954 239179
rect 278710 236567 278762 236573
rect 278710 236509 278762 236515
rect 278914 233470 278942 239173
rect 279010 233484 279038 246494
rect 279094 243005 279146 243011
rect 279094 242947 279146 242953
rect 279106 242863 279134 242947
rect 279094 242857 279146 242863
rect 279094 242799 279146 242805
rect 279490 240199 279518 246494
rect 279682 246480 279936 246508
rect 280320 246480 280478 246508
rect 279478 240193 279530 240199
rect 279478 240135 279530 240141
rect 279682 239237 279710 246480
rect 280150 239971 280202 239977
rect 280150 239913 280202 239919
rect 280246 239971 280298 239977
rect 280246 239913 280298 239919
rect 279670 239231 279722 239237
rect 279670 239173 279722 239179
rect 279382 239009 279434 239015
rect 279382 238951 279434 238957
rect 279478 239009 279530 239015
rect 279478 238951 279530 238957
rect 279394 236740 279422 238951
rect 279490 238349 279518 238951
rect 279478 238343 279530 238349
rect 279478 238285 279530 238291
rect 279394 236712 279518 236740
rect 279490 233484 279518 236712
rect 279766 234199 279818 234205
rect 279766 234141 279818 234147
rect 279778 233484 279806 234141
rect 280162 233484 280190 239913
rect 280258 239575 280286 239913
rect 280244 239566 280300 239575
rect 280244 239501 280300 239510
rect 280450 239237 280478 246480
rect 280534 239749 280586 239755
rect 280534 239691 280586 239697
rect 280438 239231 280490 239237
rect 280438 239173 280490 239179
rect 280546 233484 280574 239691
rect 280738 237165 280766 246494
rect 280834 246489 280862 246721
rect 280930 246563 280958 246721
rect 281314 246711 281342 246753
rect 285002 246753 285004 246762
rect 285236 246818 285292 246827
rect 285236 246753 285292 246762
rect 287540 246818 287596 246827
rect 307412 246818 307468 246827
rect 287540 246753 287596 246762
rect 288310 246779 288362 246785
rect 284950 246721 285002 246727
rect 281302 246705 281354 246711
rect 281302 246647 281354 246653
rect 280918 246557 280970 246563
rect 280918 246499 280970 246505
rect 280822 246483 280874 246489
rect 280822 246425 280874 246431
rect 280822 246335 280874 246341
rect 280822 246277 280874 246283
rect 280834 242863 280862 246277
rect 280822 242857 280874 242863
rect 280822 242799 280874 242805
rect 281110 240415 281162 240421
rect 281110 240357 281162 240363
rect 280726 237159 280778 237165
rect 280726 237101 280778 237107
rect 279010 233456 279312 233484
rect 279490 233456 279648 233484
rect 279778 233456 280032 233484
rect 280162 233456 280416 233484
rect 280546 233456 280752 233484
rect 281122 233470 281150 240357
rect 281218 236425 281246 246494
rect 281398 240785 281450 240791
rect 281398 240727 281450 240733
rect 281410 240421 281438 240727
rect 281398 240415 281450 240421
rect 281398 240357 281450 240363
rect 281494 239897 281546 239903
rect 281494 239839 281546 239845
rect 281206 236419 281258 236425
rect 281206 236361 281258 236367
rect 281506 233470 281534 239839
rect 281698 238941 281726 246494
rect 281794 246480 282048 246508
rect 282528 246480 282782 246508
rect 281794 239681 281822 246480
rect 282262 240785 282314 240791
rect 282262 240727 282314 240733
rect 282166 240193 282218 240199
rect 282166 240135 282218 240141
rect 282178 239681 282206 240135
rect 281782 239675 281834 239681
rect 281782 239617 281834 239623
rect 282166 239675 282218 239681
rect 282166 239617 282218 239623
rect 282274 239089 282302 240727
rect 282262 239083 282314 239089
rect 282262 239025 282314 239031
rect 281686 238935 281738 238941
rect 281686 238877 281738 238883
rect 282754 236869 282782 246480
rect 282946 239607 282974 246494
rect 283222 243301 283274 243307
rect 283222 243243 283274 243249
rect 282934 239601 282986 239607
rect 282934 239543 282986 239549
rect 283030 239601 283082 239607
rect 283030 239543 283082 239549
rect 283042 239311 283070 239543
rect 283030 239305 283082 239311
rect 283030 239247 283082 239253
rect 282742 236863 282794 236869
rect 282742 236805 282794 236811
rect 281590 236345 281642 236351
rect 281590 236287 281642 236293
rect 281602 233484 281630 236287
rect 282454 234643 282506 234649
rect 282454 234585 282506 234591
rect 282466 233484 282494 234585
rect 282838 234495 282890 234501
rect 282838 234437 282890 234443
rect 282850 233484 282878 234437
rect 283234 233484 283262 243243
rect 283318 236345 283370 236351
rect 283318 236287 283370 236293
rect 281602 233456 281856 233484
rect 282240 233456 282494 233484
rect 282624 233456 282878 233484
rect 282960 233456 283262 233484
rect 283330 233470 283358 236287
rect 283426 234247 283454 246494
rect 283702 242413 283754 242419
rect 283702 242355 283754 242361
rect 283412 234238 283468 234247
rect 283412 234173 283468 234182
rect 283714 233470 283742 242355
rect 283810 239533 283838 246494
rect 284256 246480 284414 246508
rect 283990 242487 284042 242493
rect 283990 242429 284042 242435
rect 284002 241901 284030 242429
rect 283894 241895 283946 241901
rect 283894 241837 283946 241843
rect 283990 241895 284042 241901
rect 283990 241837 284042 241843
rect 283906 239533 283934 241837
rect 283798 239527 283850 239533
rect 283798 239469 283850 239475
rect 283894 239527 283946 239533
rect 283894 239469 283946 239475
rect 284086 239305 284138 239311
rect 284086 239247 284138 239253
rect 284098 239089 284126 239247
rect 284086 239083 284138 239089
rect 284086 239025 284138 239031
rect 284386 236203 284414 246480
rect 284482 246480 284736 246508
rect 284962 246480 285072 246508
rect 284482 239829 284510 246480
rect 284470 239823 284522 239829
rect 284470 239765 284522 239771
rect 284374 236197 284426 236203
rect 284374 236139 284426 236145
rect 284662 234273 284714 234279
rect 284662 234215 284714 234221
rect 284278 234199 284330 234205
rect 284278 234141 284330 234147
rect 284290 233484 284318 234141
rect 284674 233484 284702 234215
rect 284962 234099 284990 246480
rect 285250 243899 285278 246753
rect 287554 246711 287582 246753
rect 288694 246779 288746 246785
rect 288362 246739 288446 246767
rect 288310 246721 288362 246727
rect 287542 246705 287594 246711
rect 287074 246628 287280 246656
rect 287542 246647 287594 246653
rect 288418 246637 288446 246739
rect 288694 246721 288746 246727
rect 292246 246779 292298 246785
rect 292246 246721 292298 246727
rect 295702 246779 295754 246785
rect 307412 246753 307468 246762
rect 307892 246818 307948 246827
rect 308084 246818 308140 246827
rect 307892 246753 307948 246762
rect 308002 246776 308084 246804
rect 295702 246721 295754 246727
rect 288406 246631 288458 246637
rect 285552 246480 285854 246508
rect 285238 243893 285290 243899
rect 285238 243835 285290 243841
rect 285622 240267 285674 240273
rect 285622 240209 285674 240215
rect 285044 239714 285100 239723
rect 285044 239649 285100 239658
rect 285058 236351 285086 239649
rect 285634 239385 285662 240209
rect 285526 239379 285578 239385
rect 285526 239321 285578 239327
rect 285622 239379 285674 239385
rect 285622 239321 285674 239327
rect 285238 236863 285290 236869
rect 285238 236805 285290 236811
rect 285250 236425 285278 236805
rect 285238 236419 285290 236425
rect 285238 236361 285290 236367
rect 285046 236345 285098 236351
rect 285046 236287 285098 236293
rect 284948 234090 285004 234099
rect 284948 234025 285004 234034
rect 285142 233977 285194 233983
rect 285142 233919 285194 233925
rect 285046 233829 285098 233835
rect 285046 233771 285098 233777
rect 285058 233484 285086 233771
rect 284064 233456 284318 233484
rect 284448 233456 284702 233484
rect 284832 233456 285086 233484
rect 285154 233470 285182 233919
rect 285538 233470 285566 239321
rect 285826 237165 285854 246480
rect 286018 239459 286046 246494
rect 286450 246212 286478 246494
rect 286402 246184 286478 246212
rect 286594 246480 286848 246508
rect 286006 239453 286058 239459
rect 286006 239395 286058 239401
rect 285814 237159 285866 237165
rect 285814 237101 285866 237107
rect 286402 237091 286430 246184
rect 286486 242487 286538 242493
rect 286486 242429 286538 242435
rect 286390 237085 286442 237091
rect 286390 237027 286442 237033
rect 285910 236863 285962 236869
rect 285910 236805 285962 236811
rect 285922 233470 285950 236805
rect 286498 233484 286526 242429
rect 286594 237313 286622 246480
rect 286870 240415 286922 240421
rect 286870 240357 286922 240363
rect 286582 237307 286634 237313
rect 286582 237249 286634 237255
rect 286882 233484 286910 240357
rect 287074 239163 287102 246628
rect 288406 246573 288458 246579
rect 287362 246480 287760 246508
rect 288240 246480 288446 246508
rect 287362 246249 287390 246480
rect 287170 246221 287390 246249
rect 287842 246295 288062 246323
rect 287062 239157 287114 239163
rect 287062 239099 287114 239105
rect 287170 237461 287198 246221
rect 287842 246193 287870 246295
rect 288034 246267 288062 246295
rect 287926 246261 287978 246267
rect 287926 246203 287978 246209
rect 288022 246261 288074 246267
rect 288022 246203 288074 246209
rect 287350 246187 287402 246193
rect 287350 246129 287402 246135
rect 287830 246187 287882 246193
rect 287938 246175 287966 246203
rect 288118 246187 288170 246193
rect 287938 246147 288118 246175
rect 287830 246129 287882 246135
rect 288118 246129 288170 246135
rect 287362 244861 287390 246129
rect 287254 244855 287306 244861
rect 287254 244797 287306 244803
rect 287350 244855 287402 244861
rect 287350 244797 287402 244803
rect 287266 239575 287294 244797
rect 287458 244713 287966 244732
rect 287446 244707 287978 244713
rect 287498 244704 287926 244707
rect 287446 244649 287498 244655
rect 287926 244649 287978 244655
rect 287830 244559 287882 244565
rect 287554 244519 287830 244547
rect 287446 244263 287498 244269
rect 287446 244205 287498 244211
rect 287458 240273 287486 244205
rect 287554 243011 287582 244519
rect 287830 244501 287882 244507
rect 287746 244445 287966 244473
rect 287746 244343 287774 244445
rect 287734 244337 287786 244343
rect 287734 244279 287786 244285
rect 287938 244269 287966 244445
rect 287926 244263 287978 244269
rect 287926 244205 287978 244211
rect 288118 243893 288170 243899
rect 288118 243835 288170 243841
rect 288130 243719 288158 243835
rect 288116 243710 288172 243719
rect 287938 243668 288062 243696
rect 287542 243005 287594 243011
rect 287734 243005 287786 243011
rect 287542 242947 287594 242953
rect 287636 242970 287692 242979
rect 287734 242947 287786 242953
rect 287636 242905 287692 242914
rect 287650 242715 287678 242905
rect 287542 242709 287594 242715
rect 287542 242651 287594 242657
rect 287638 242709 287690 242715
rect 287638 242651 287690 242657
rect 287446 240267 287498 240273
rect 287446 240209 287498 240215
rect 287350 240045 287402 240051
rect 287350 239987 287402 239993
rect 287252 239566 287308 239575
rect 287252 239501 287308 239510
rect 287362 239311 287390 239987
rect 287350 239305 287402 239311
rect 287350 239247 287402 239253
rect 287158 237455 287210 237461
rect 287158 237397 287210 237403
rect 287254 237455 287306 237461
rect 287254 237397 287306 237403
rect 287266 233484 287294 237397
rect 287350 233903 287402 233909
rect 287350 233845 287402 233851
rect 286272 233456 286526 233484
rect 286656 233456 286910 233484
rect 287040 233456 287294 233484
rect 287362 233470 287390 233845
rect 287554 233484 287582 242651
rect 287746 242567 287774 242947
rect 287734 242561 287786 242567
rect 287734 242503 287786 242509
rect 287828 242526 287884 242535
rect 287938 242512 287966 243668
rect 288034 243548 288062 243668
rect 288116 243645 288172 243654
rect 288308 243710 288364 243719
rect 288308 243645 288364 243654
rect 288322 243548 288350 243645
rect 288034 243520 288350 243548
rect 288310 242931 288362 242937
rect 288310 242873 288362 242879
rect 288214 242783 288266 242789
rect 288214 242725 288266 242731
rect 288022 242709 288074 242715
rect 288022 242651 288074 242657
rect 288034 242535 288062 242651
rect 288118 242561 288170 242567
rect 287884 242484 287966 242512
rect 288020 242526 288076 242535
rect 287828 242461 287884 242470
rect 288118 242503 288170 242509
rect 288020 242461 288076 242470
rect 287638 241081 287690 241087
rect 287638 241023 287690 241029
rect 287650 240051 287678 241023
rect 287830 240267 287882 240273
rect 287830 240209 287882 240215
rect 287926 240267 287978 240273
rect 287926 240209 287978 240215
rect 287842 240125 287870 240209
rect 287830 240119 287882 240125
rect 287830 240061 287882 240067
rect 287638 240045 287690 240051
rect 287638 239987 287690 239993
rect 287938 237461 287966 240209
rect 288130 239723 288158 242503
rect 288116 239714 288172 239723
rect 288116 239649 288172 239658
rect 288118 238343 288170 238349
rect 288118 238285 288170 238291
rect 287926 237455 287978 237461
rect 287926 237397 287978 237403
rect 288130 237017 288158 238285
rect 288118 237011 288170 237017
rect 288118 236953 288170 236959
rect 288118 236345 288170 236351
rect 288118 236287 288170 236293
rect 287554 233456 287760 233484
rect 288130 233470 288158 236287
rect 288226 233835 288254 242725
rect 288322 241087 288350 242873
rect 288310 241081 288362 241087
rect 288310 241023 288362 241029
rect 288418 237165 288446 246480
rect 288562 246212 288590 246494
rect 288706 246415 288734 246721
rect 289056 246628 289310 246656
rect 292258 246637 292286 246721
rect 289174 246483 289226 246489
rect 289174 246425 289226 246431
rect 288694 246409 288746 246415
rect 288694 246351 288746 246357
rect 288514 246184 288590 246212
rect 288406 237159 288458 237165
rect 288406 237101 288458 237107
rect 288514 236795 288542 246184
rect 289186 244991 289214 246425
rect 288802 244963 289214 244991
rect 288802 244861 288830 244963
rect 288790 244855 288842 244861
rect 288790 244797 288842 244803
rect 288886 244855 288938 244861
rect 288886 244797 288938 244803
rect 288598 242931 288650 242937
rect 288598 242873 288650 242879
rect 288610 241901 288638 242873
rect 288898 242863 288926 244797
rect 288886 242857 288938 242863
rect 288886 242799 288938 242805
rect 288982 242857 289034 242863
rect 288982 242799 289034 242805
rect 288598 241895 288650 241901
rect 288598 241837 288650 241843
rect 288694 241895 288746 241901
rect 288694 241837 288746 241843
rect 288502 236789 288554 236795
rect 288502 236731 288554 236737
rect 288214 233829 288266 233835
rect 288214 233771 288266 233777
rect 288706 233484 288734 241837
rect 288994 236869 289022 242799
rect 289282 237239 289310 246628
rect 292246 246631 292298 246637
rect 292246 246573 292298 246579
rect 294838 246557 294890 246563
rect 289474 240051 289502 246494
rect 289762 246480 289968 246508
rect 289652 241786 289708 241795
rect 289652 241721 289708 241730
rect 289666 241203 289694 241721
rect 289652 241194 289708 241203
rect 289652 241129 289708 241138
rect 289462 240045 289514 240051
rect 289462 239987 289514 239993
rect 289462 239897 289514 239903
rect 289462 239839 289514 239845
rect 289270 237233 289322 237239
rect 289270 237175 289322 237181
rect 289076 237050 289132 237059
rect 289076 236985 289132 236994
rect 288982 236863 289034 236869
rect 288982 236805 289034 236811
rect 289090 233484 289118 236985
rect 289270 236567 289322 236573
rect 289270 236509 289322 236515
rect 289282 233909 289310 236509
rect 289270 233903 289322 233909
rect 289270 233845 289322 233851
rect 289474 233484 289502 239839
rect 289762 236721 289790 246480
rect 290038 244337 290090 244343
rect 290038 244279 290090 244285
rect 289844 241194 289900 241203
rect 289844 241129 289900 241138
rect 289858 240759 289886 241129
rect 290050 241087 290078 244279
rect 290038 241081 290090 241087
rect 290038 241023 290090 241029
rect 289844 240750 289900 240759
rect 289844 240685 289900 240694
rect 290338 237387 290366 246494
rect 290626 246480 290784 246508
rect 291264 246480 291518 246508
rect 290518 240045 290570 240051
rect 290518 239987 290570 239993
rect 290326 237381 290378 237387
rect 290326 237323 290378 237329
rect 289750 236715 289802 236721
rect 289750 236657 289802 236663
rect 289940 233942 289996 233951
rect 289940 233877 289996 233886
rect 289844 233498 289900 233507
rect 288480 233456 288734 233484
rect 288864 233456 289118 233484
rect 289248 233456 289502 233484
rect 289584 233456 289844 233484
rect 289954 233470 289982 233877
rect 290530 233484 290558 239987
rect 290626 237313 290654 246480
rect 290710 240193 290762 240199
rect 290710 240135 290762 240141
rect 290806 240193 290858 240199
rect 290806 240135 290858 240141
rect 290722 237313 290750 240135
rect 290818 239459 290846 240135
rect 291382 239749 291434 239755
rect 291382 239691 291434 239697
rect 291190 239675 291242 239681
rect 291190 239617 291242 239623
rect 290806 239453 290858 239459
rect 290806 239395 290858 239401
rect 290902 239453 290954 239459
rect 290902 239395 290954 239401
rect 290914 239237 290942 239395
rect 291202 239256 291230 239617
rect 291394 239607 291422 239691
rect 291490 239681 291518 246480
rect 291682 239829 291710 246494
rect 291958 241081 292010 241087
rect 291958 241023 292010 241029
rect 291670 239823 291722 239829
rect 291670 239765 291722 239771
rect 291478 239675 291530 239681
rect 291478 239617 291530 239623
rect 291382 239601 291434 239607
rect 291382 239543 291434 239549
rect 291202 239237 291326 239256
rect 290902 239231 290954 239237
rect 291202 239231 291338 239237
rect 291202 239228 291286 239231
rect 290902 239173 290954 239179
rect 291286 239173 291338 239179
rect 290806 239083 290858 239089
rect 290806 239025 290858 239031
rect 290614 237307 290666 237313
rect 290614 237249 290666 237255
rect 290710 237307 290762 237313
rect 290710 237249 290762 237255
rect 290708 236310 290764 236319
rect 290818 236277 290846 239025
rect 291970 237535 291998 241023
rect 292066 237535 292094 246494
rect 292150 239527 292202 239533
rect 292150 239469 292202 239475
rect 291958 237529 292010 237535
rect 291958 237471 292010 237477
rect 292054 237529 292106 237535
rect 292054 237471 292106 237477
rect 291766 236863 291818 236869
rect 291766 236805 291818 236811
rect 291670 236789 291722 236795
rect 291670 236731 291722 236737
rect 291286 236493 291338 236499
rect 291286 236435 291338 236441
rect 290708 236245 290710 236254
rect 290762 236245 290764 236254
rect 290806 236271 290858 236277
rect 290710 236213 290762 236219
rect 290806 236213 290858 236219
rect 290902 233533 290954 233539
rect 290352 233456 290558 233484
rect 290688 233481 290902 233484
rect 291298 233484 291326 236435
rect 291682 233484 291710 236731
rect 290688 233475 290954 233481
rect 290688 233456 290942 233475
rect 291072 233456 291326 233484
rect 291456 233456 291710 233484
rect 291778 233470 291806 236805
rect 292162 233470 292190 239469
rect 292244 239270 292300 239279
rect 292244 239205 292300 239214
rect 292258 239015 292286 239205
rect 292246 239009 292298 239015
rect 292246 238951 292298 238957
rect 292546 237461 292574 246494
rect 292992 246480 293246 246508
rect 293110 243153 293162 243159
rect 293110 243095 293162 243101
rect 293122 239427 293150 243095
rect 293218 239681 293246 246480
rect 293314 246480 293376 246508
rect 293808 246480 294014 246508
rect 293206 239675 293258 239681
rect 293206 239617 293258 239623
rect 293314 239459 293342 246480
rect 293398 243153 293450 243159
rect 293398 243095 293450 243101
rect 293410 242937 293438 243095
rect 293782 243079 293834 243085
rect 293782 243021 293834 243027
rect 293878 243079 293930 243085
rect 293878 243021 293930 243027
rect 293398 242931 293450 242937
rect 293398 242873 293450 242879
rect 293590 242931 293642 242937
rect 293590 242873 293642 242879
rect 293398 240045 293450 240051
rect 293398 239987 293450 239993
rect 293410 239459 293438 239987
rect 293302 239453 293354 239459
rect 293108 239418 293164 239427
rect 293302 239395 293354 239401
rect 293398 239453 293450 239459
rect 293398 239395 293450 239401
rect 293108 239353 293164 239362
rect 292534 237455 292586 237461
rect 292534 237397 292586 237403
rect 293494 236715 293546 236721
rect 293494 236657 293546 236663
rect 292534 233903 292586 233909
rect 292534 233845 292586 233851
rect 292546 233470 292574 233845
rect 293110 233829 293162 233835
rect 293110 233771 293162 233777
rect 293122 233484 293150 233771
rect 293506 233484 293534 236657
rect 292896 233456 293150 233484
rect 293280 233456 293534 233484
rect 293602 233484 293630 242873
rect 293794 239723 293822 243021
rect 293780 239714 293836 239723
rect 293780 239649 293836 239658
rect 293780 239566 293836 239575
rect 293780 239501 293836 239510
rect 293794 238349 293822 239501
rect 293686 238343 293738 238349
rect 293686 238285 293738 238291
rect 293782 238343 293834 238349
rect 293782 238285 293834 238291
rect 293698 238220 293726 238285
rect 293890 238220 293918 243021
rect 293986 239015 294014 246480
rect 294178 246480 294288 246508
rect 294466 246480 294768 246508
rect 294838 246499 294890 246505
rect 294178 239404 294206 246480
rect 294358 243153 294410 243159
rect 294358 243095 294410 243101
rect 294370 242993 294398 243095
rect 294466 243085 294494 246480
rect 294850 244288 294878 246499
rect 295104 246480 295358 246508
rect 294562 244260 294878 244288
rect 294454 243079 294506 243085
rect 294454 243021 294506 243027
rect 294562 242993 294590 244260
rect 294370 242965 294590 242993
rect 294454 239823 294506 239829
rect 294454 239765 294506 239771
rect 294466 239459 294494 239765
rect 294742 239749 294794 239755
rect 294742 239691 294794 239697
rect 294454 239453 294506 239459
rect 294178 239385 294302 239404
rect 294454 239395 294506 239401
rect 294178 239379 294314 239385
rect 294178 239376 294262 239379
rect 294262 239321 294314 239327
rect 294358 239305 294410 239311
rect 294358 239247 294410 239253
rect 293974 239009 294026 239015
rect 293974 238951 294026 238957
rect 293698 238192 293918 238220
rect 293974 237307 294026 237313
rect 293974 237249 294026 237255
rect 294070 237307 294122 237313
rect 294070 237249 294122 237255
rect 293602 233456 293664 233484
rect 293986 233470 294014 237249
rect 294082 236319 294110 237249
rect 294068 236310 294124 236319
rect 294068 236245 294124 236254
rect 294370 233470 294398 239247
rect 294754 233470 294782 239691
rect 295330 237461 295358 246480
rect 295426 246480 295584 246508
rect 295426 240199 295454 246480
rect 295714 244343 295742 246721
rect 295702 244337 295754 244343
rect 295702 244279 295754 244285
rect 295604 241194 295660 241203
rect 295604 241129 295660 241138
rect 295618 241032 295646 241129
rect 295892 241046 295948 241055
rect 295618 241004 295892 241032
rect 295892 240981 295948 240990
rect 295414 240193 295466 240199
rect 295414 240135 295466 240141
rect 295702 240045 295754 240051
rect 295702 239987 295754 239993
rect 295606 239971 295658 239977
rect 295606 239913 295658 239919
rect 295318 237455 295370 237461
rect 295318 237397 295370 237403
rect 295222 236937 295274 236943
rect 295222 236879 295274 236885
rect 294838 236641 294890 236647
rect 294838 236583 294890 236589
rect 294850 233484 294878 236583
rect 295234 233484 295262 236879
rect 295618 233484 295646 239913
rect 295714 239279 295742 239987
rect 296002 239459 296030 246494
rect 296086 239971 296138 239977
rect 296086 239913 296138 239919
rect 295990 239453 296042 239459
rect 295990 239395 296042 239401
rect 295700 239270 295756 239279
rect 295700 239205 295756 239214
rect 295798 236641 295850 236647
rect 295798 236583 295850 236589
rect 295810 233951 295838 236583
rect 295796 233942 295852 233951
rect 295796 233877 295852 233886
rect 296098 233507 296126 239913
rect 296482 237313 296510 246494
rect 296662 239897 296714 239903
rect 296662 239839 296714 239845
rect 296674 239237 296702 239839
rect 296566 239231 296618 239237
rect 296566 239173 296618 239179
rect 296662 239231 296714 239237
rect 296662 239173 296714 239179
rect 296470 237307 296522 237313
rect 296470 237249 296522 237255
rect 296182 236419 296234 236425
rect 296182 236361 296234 236367
rect 296084 233498 296140 233507
rect 294850 233456 295104 233484
rect 295234 233456 295488 233484
rect 295618 233456 295872 233484
rect 289844 233433 289900 233442
rect 296194 233470 296222 236361
rect 296578 233470 296606 239173
rect 296866 237017 296894 246494
rect 297058 246480 297312 246508
rect 297634 246480 297792 246508
rect 298224 246480 298430 246508
rect 298608 246480 299006 246508
rect 297058 240347 297086 246480
rect 297430 244337 297482 244343
rect 297430 244279 297482 244285
rect 297442 242863 297470 244279
rect 297430 242857 297482 242863
rect 297430 242799 297482 242805
rect 297634 240440 297662 246480
rect 298210 243381 298334 243400
rect 297814 243375 297866 243381
rect 297814 243317 297866 243323
rect 298198 243375 298334 243381
rect 298250 243372 298334 243375
rect 298198 243317 298250 243323
rect 297826 242863 297854 243317
rect 298306 243307 298334 243372
rect 298294 243301 298346 243307
rect 298196 243266 298252 243275
rect 297922 243224 298196 243252
rect 297922 243127 297950 243224
rect 298294 243243 298346 243249
rect 298196 243201 298252 243210
rect 298402 243141 298430 246480
rect 298498 243381 298910 243400
rect 298486 243375 298910 243381
rect 298538 243372 298910 243375
rect 298486 243317 298538 243323
rect 298582 243227 298634 243233
rect 298678 243227 298730 243233
rect 298634 243187 298678 243215
rect 298582 243169 298634 243175
rect 298678 243169 298730 243175
rect 298882 243159 298910 243372
rect 298870 243153 298922 243159
rect 297908 243118 297964 243127
rect 298402 243113 298718 243141
rect 297908 243053 297964 243062
rect 298018 243039 298622 243067
rect 297910 242931 297962 242937
rect 297910 242873 297962 242879
rect 297814 242857 297866 242863
rect 297814 242799 297866 242805
rect 297922 242364 297950 242873
rect 298018 242493 298046 243039
rect 298594 243011 298622 243039
rect 298582 243005 298634 243011
rect 298582 242947 298634 242953
rect 298006 242487 298058 242493
rect 298006 242429 298058 242435
rect 298102 242487 298154 242493
rect 298102 242429 298154 242435
rect 298114 242364 298142 242429
rect 297922 242336 298142 242364
rect 298690 241476 298718 243113
rect 298870 243095 298922 243101
rect 298498 241448 298718 241476
rect 298004 240454 298060 240463
rect 297634 240412 297854 240440
rect 297046 240341 297098 240347
rect 297046 240283 297098 240289
rect 297826 239533 297854 240412
rect 298004 240389 298060 240398
rect 298018 239871 298046 240389
rect 298198 240193 298250 240199
rect 298198 240135 298250 240141
rect 298004 239862 298060 239871
rect 298210 239829 298238 240135
rect 298004 239797 298060 239806
rect 298198 239823 298250 239829
rect 298198 239765 298250 239771
rect 297814 239527 297866 239533
rect 297814 239469 297866 239475
rect 297430 238935 297482 238941
rect 297430 238877 297482 238883
rect 296854 237011 296906 237017
rect 296854 236953 296906 236959
rect 296950 236271 297002 236277
rect 296950 236213 297002 236219
rect 296962 233470 296990 236213
rect 297046 233607 297098 233613
rect 297046 233549 297098 233555
rect 297058 233484 297086 233549
rect 297442 233484 297470 238877
rect 297814 236345 297866 236351
rect 297814 236287 297866 236293
rect 297826 233484 297854 236287
rect 298388 234238 298444 234247
rect 298388 234173 298444 234182
rect 297058 233456 297312 233484
rect 297442 233456 297696 233484
rect 297826 233456 298080 233484
rect 298402 233470 298430 234173
rect 298498 233687 298526 241448
rect 298978 241328 299006 246480
rect 298594 241300 299006 241328
rect 298594 233761 298622 241300
rect 299074 238941 299102 246494
rect 299520 246480 299582 246508
rect 300000 246480 300254 246508
rect 299446 243375 299498 243381
rect 299446 243317 299498 243323
rect 299458 242937 299486 243317
rect 299446 242931 299498 242937
rect 299446 242873 299498 242879
rect 299554 242715 299582 246480
rect 299638 242931 299690 242937
rect 299638 242873 299690 242879
rect 299650 242789 299678 242873
rect 299638 242783 299690 242789
rect 299638 242725 299690 242731
rect 299542 242709 299594 242715
rect 299542 242651 299594 242657
rect 299734 242709 299786 242715
rect 299734 242651 299786 242657
rect 299062 238935 299114 238941
rect 299062 238877 299114 238883
rect 299542 237085 299594 237091
rect 299542 237027 299594 237033
rect 298774 236197 298826 236203
rect 298774 236139 298826 236145
rect 298582 233755 298634 233761
rect 298582 233697 298634 233703
rect 298486 233681 298538 233687
rect 298486 233623 298538 233629
rect 298786 233470 298814 236139
rect 299156 234090 299212 234099
rect 299156 234025 299212 234034
rect 299170 233470 299198 234025
rect 299554 233484 299582 237027
rect 299638 236937 299690 236943
rect 299638 236879 299690 236885
rect 299520 233456 299582 233484
rect 299650 233484 299678 236879
rect 299746 236721 299774 242651
rect 300022 239083 300074 239089
rect 300022 239025 300074 239031
rect 299734 236715 299786 236721
rect 299734 236657 299786 236663
rect 300034 233484 300062 239025
rect 300226 237313 300254 246480
rect 300214 237307 300266 237313
rect 300214 237249 300266 237255
rect 300322 234057 300350 246494
rect 300598 237159 300650 237165
rect 300598 237101 300650 237107
rect 300310 234051 300362 234057
rect 300310 233993 300362 233999
rect 299650 233456 299904 233484
rect 300034 233456 300288 233484
rect 300610 233470 300638 237101
rect 300802 236425 300830 246494
rect 301282 242641 301310 246494
rect 301632 246480 301886 246508
rect 301270 242635 301322 242641
rect 301270 242577 301322 242583
rect 301858 239829 301886 246480
rect 301954 246480 302112 246508
rect 301846 239823 301898 239829
rect 301846 239765 301898 239771
rect 301076 239714 301132 239723
rect 301076 239649 301132 239658
rect 300982 237233 301034 237239
rect 300982 237175 301034 237181
rect 300790 236419 300842 236425
rect 300790 236361 300842 236367
rect 300994 233470 301022 237175
rect 301090 233484 301118 239649
rect 301846 239601 301898 239607
rect 301846 239543 301898 239549
rect 301462 237381 301514 237387
rect 301462 237323 301514 237329
rect 301474 233484 301502 237323
rect 301858 233484 301886 239543
rect 301954 234131 301982 246480
rect 302530 239607 302558 246494
rect 303010 239681 303038 246494
rect 303394 243085 303422 246494
rect 303840 246480 304094 246508
rect 303382 243079 303434 243085
rect 303382 243021 303434 243027
rect 303670 239971 303722 239977
rect 303670 239913 303722 239919
rect 302806 239675 302858 239681
rect 302806 239617 302858 239623
rect 302998 239675 303050 239681
rect 302998 239617 303050 239623
rect 302518 239601 302570 239607
rect 302518 239543 302570 239549
rect 302422 237529 302474 237535
rect 302422 237471 302474 237477
rect 301942 234125 301994 234131
rect 301942 234067 301994 234073
rect 302434 233484 302462 237471
rect 301090 233456 301392 233484
rect 301474 233456 301728 233484
rect 301858 233456 302112 233484
rect 302434 233456 302496 233484
rect 302818 233470 302846 239617
rect 303682 239385 303710 239913
rect 303574 239379 303626 239385
rect 303574 239321 303626 239327
rect 303670 239379 303722 239385
rect 303670 239321 303722 239327
rect 303190 239009 303242 239015
rect 303190 238951 303242 238957
rect 303202 233470 303230 238951
rect 303586 233470 303614 239321
rect 304066 237535 304094 246480
rect 304306 246212 304334 246494
rect 304258 246184 304334 246212
rect 304150 239453 304202 239459
rect 304150 239395 304202 239401
rect 304054 237529 304106 237535
rect 304054 237471 304106 237477
rect 303670 237455 303722 237461
rect 303670 237397 303722 237403
rect 303682 233484 303710 237397
rect 304162 233484 304190 239395
rect 304258 234427 304286 246184
rect 304738 239015 304766 246494
rect 305122 243233 305150 246494
rect 305110 243227 305162 243233
rect 305110 243169 305162 243175
rect 305014 239527 305066 239533
rect 305014 239469 305066 239475
rect 304726 239009 304778 239015
rect 304726 238951 304778 238957
rect 304438 237011 304490 237017
rect 304438 236953 304490 236959
rect 304246 234421 304298 234427
rect 304246 234363 304298 234369
rect 304450 233484 304478 236953
rect 303682 233456 303936 233484
rect 304162 233456 304320 233484
rect 304450 233456 304704 233484
rect 305026 233470 305054 239469
rect 305300 239418 305356 239427
rect 305300 239353 305356 239362
rect 305314 233484 305342 239353
rect 305602 233761 305630 246494
rect 305698 246480 306048 246508
rect 305698 234575 305726 246480
rect 306514 246212 306542 246494
rect 306466 246184 306542 246212
rect 306658 246480 306912 246508
rect 305782 242783 305834 242789
rect 305782 242725 305834 242731
rect 305794 242641 305822 242725
rect 305782 242635 305834 242641
rect 305782 242577 305834 242583
rect 305782 238935 305834 238941
rect 305782 238877 305834 238883
rect 305686 234569 305738 234575
rect 305686 234511 305738 234517
rect 305590 233755 305642 233761
rect 305590 233697 305642 233703
rect 305314 233456 305424 233484
rect 305794 233470 305822 238877
rect 305878 237307 305930 237313
rect 305878 237249 305930 237255
rect 305974 237307 306026 237313
rect 305974 237249 306026 237255
rect 305890 233484 305918 237249
rect 305986 236795 306014 237249
rect 306466 236795 306494 246184
rect 306658 244565 306686 246480
rect 307330 244713 307358 246494
rect 307426 244713 307454 246753
rect 307510 246409 307562 246415
rect 307510 246351 307562 246357
rect 307702 246409 307754 246415
rect 307702 246351 307754 246357
rect 307318 244707 307370 244713
rect 307318 244649 307370 244655
rect 307414 244707 307466 244713
rect 307414 244649 307466 244655
rect 307522 244565 307550 246351
rect 307714 246193 307742 246351
rect 307702 246187 307754 246193
rect 307702 246129 307754 246135
rect 306646 244559 306698 244565
rect 306646 244501 306698 244507
rect 307510 244559 307562 244565
rect 307510 244501 307562 244507
rect 307702 242857 307754 242863
rect 307702 242799 307754 242805
rect 307714 242535 307742 242799
rect 307700 242526 307756 242535
rect 306646 242487 306698 242493
rect 307700 242461 307756 242470
rect 306646 242429 306698 242435
rect 306658 240125 306686 242429
rect 306646 240119 306698 240125
rect 306646 240061 306698 240067
rect 307810 239977 307838 246494
rect 307906 246193 307934 246753
rect 308002 246415 308030 246776
rect 311156 246818 311212 246827
rect 308084 246753 308140 246762
rect 309238 246779 309290 246785
rect 309238 246721 309290 246727
rect 309334 246779 309386 246785
rect 309334 246721 309386 246727
rect 309430 246779 309482 246785
rect 328340 246818 328396 246827
rect 311156 246753 311212 246762
rect 313750 246779 313802 246785
rect 309430 246721 309482 246727
rect 308256 246480 308414 246508
rect 308640 246480 308894 246508
rect 307990 246409 308042 246415
rect 307990 246351 308042 246357
rect 307894 246187 307946 246193
rect 307894 246129 307946 246135
rect 308086 243893 308138 243899
rect 308086 243835 308138 243841
rect 308098 243275 308126 243835
rect 307892 243266 307948 243275
rect 307892 243201 307948 243210
rect 308084 243266 308140 243275
rect 308084 243201 308140 243210
rect 307906 242535 307934 243201
rect 308278 242857 308330 242863
rect 308084 242822 308140 242831
rect 308084 242757 308140 242766
rect 308276 242822 308278 242831
rect 308330 242822 308332 242831
rect 308276 242757 308332 242766
rect 308098 242715 308126 242757
rect 308086 242709 308138 242715
rect 308086 242651 308138 242657
rect 307892 242526 307948 242535
rect 307892 242461 307948 242470
rect 307894 241895 307946 241901
rect 307894 241837 307946 241843
rect 307798 239971 307850 239977
rect 307798 239913 307850 239919
rect 307906 239829 307934 241837
rect 306646 239823 306698 239829
rect 306646 239765 306698 239771
rect 307894 239823 307946 239829
rect 307894 239765 307946 239771
rect 305974 236789 306026 236795
rect 305974 236731 306026 236737
rect 306454 236789 306506 236795
rect 306454 236731 306506 236737
rect 306262 236419 306314 236425
rect 306262 236361 306314 236367
rect 306274 233484 306302 236361
rect 306658 233484 306686 239765
rect 307606 239675 307658 239681
rect 307606 239617 307658 239623
rect 307222 239601 307274 239607
rect 307222 239543 307274 239549
rect 305890 233456 306144 233484
rect 306274 233456 306528 233484
rect 306658 233456 306912 233484
rect 307234 233470 307262 239543
rect 307618 233470 307646 239617
rect 308182 239009 308234 239015
rect 308182 238951 308234 238957
rect 307990 237529 308042 237535
rect 307990 237471 308042 237477
rect 308002 233470 308030 237471
rect 308194 233484 308222 238951
rect 308386 236129 308414 246480
rect 308866 239607 308894 246480
rect 308962 246480 309120 246508
rect 308962 244639 308990 246480
rect 309250 244639 309278 246721
rect 309346 246341 309374 246721
rect 309334 246335 309386 246341
rect 309334 246277 309386 246283
rect 309442 244861 309470 246721
rect 309430 244855 309482 244861
rect 309430 244797 309482 244803
rect 308950 244633 309002 244639
rect 308950 244575 309002 244581
rect 309238 244633 309290 244639
rect 309238 244575 309290 244581
rect 309538 239681 309566 246494
rect 309814 239971 309866 239977
rect 309814 239913 309866 239919
rect 309526 239675 309578 239681
rect 309526 239617 309578 239623
rect 308854 239601 308906 239607
rect 308854 239543 308906 239549
rect 308950 236789 309002 236795
rect 308950 236731 309002 236737
rect 308374 236123 308426 236129
rect 308374 236065 308426 236071
rect 308710 233755 308762 233761
rect 308710 233697 308762 233703
rect 308194 233456 308352 233484
rect 308722 233470 308750 233697
rect 308962 233484 308990 236731
rect 309430 234347 309482 234353
rect 309430 234289 309482 234295
rect 308962 233456 309120 233484
rect 309442 233470 309470 234289
rect 309826 233470 309854 239913
rect 309922 236055 309950 246494
rect 310416 246480 310718 246508
rect 310294 239675 310346 239681
rect 310294 239617 310346 239623
rect 310198 239601 310250 239607
rect 310198 239543 310250 239549
rect 309910 236049 309962 236055
rect 309910 235991 309962 235997
rect 310210 233470 310238 239543
rect 310306 233484 310334 239617
rect 310690 233484 310718 246480
rect 310834 246212 310862 246494
rect 311170 246489 311198 246753
rect 313750 246721 313802 246727
rect 314038 246779 314090 246785
rect 328532 246818 328588 246827
rect 328396 246776 328478 246804
rect 328340 246753 328396 246762
rect 314038 246721 314090 246727
rect 311734 246705 311786 246711
rect 311734 246647 311786 246653
rect 311746 246563 311774 246647
rect 313762 246637 313790 246721
rect 313942 246705 313994 246711
rect 313942 246647 313994 246653
rect 312310 246631 312362 246637
rect 312310 246573 312362 246579
rect 313750 246631 313802 246637
rect 313750 246573 313802 246579
rect 311734 246557 311786 246563
rect 311158 246483 311210 246489
rect 311158 246425 311210 246431
rect 311266 246480 311328 246508
rect 311458 246480 311664 246508
rect 311734 246499 311786 246505
rect 310786 246184 310862 246212
rect 310786 244491 310814 246184
rect 310774 244485 310826 244491
rect 310774 244427 310826 244433
rect 311266 233484 311294 246480
rect 311458 236573 311486 246480
rect 311830 244855 311882 244861
rect 311830 244797 311882 244803
rect 311842 244713 311870 244797
rect 311830 244707 311882 244713
rect 311830 244649 311882 244655
rect 311926 244707 311978 244713
rect 311926 244649 311978 244655
rect 311938 244417 311966 244649
rect 312022 244559 312074 244565
rect 312022 244501 312074 244507
rect 311926 244411 311978 244417
rect 311926 244353 311978 244359
rect 311734 241895 311786 241901
rect 311734 241837 311786 241843
rect 311746 241679 311774 241837
rect 311734 241673 311786 241679
rect 311734 241615 311786 241621
rect 311638 241599 311690 241605
rect 311638 241541 311690 241547
rect 311650 239903 311678 241541
rect 311638 239897 311690 239903
rect 311638 239839 311690 239845
rect 311638 239009 311690 239015
rect 311638 238951 311690 238957
rect 311446 236567 311498 236573
rect 311446 236509 311498 236515
rect 310306 233456 310560 233484
rect 310690 233456 310944 233484
rect 311266 233456 311328 233484
rect 311650 233470 311678 238951
rect 312034 233470 312062 244501
rect 312130 239829 312158 246494
rect 312322 246415 312350 246573
rect 312310 246409 312362 246415
rect 312310 246351 312362 246357
rect 312406 244485 312458 244491
rect 312406 244427 312458 244433
rect 312118 239823 312170 239829
rect 312118 239765 312170 239771
rect 312418 233470 312446 244427
rect 312610 240273 312638 246494
rect 312802 246480 313056 246508
rect 313186 246480 313440 246508
rect 313654 246483 313706 246489
rect 312598 240267 312650 240273
rect 312598 240209 312650 240215
rect 312802 237059 312830 246480
rect 313186 240347 313214 246480
rect 313654 246425 313706 246431
rect 313270 246409 313322 246415
rect 313666 246397 313694 246425
rect 313322 246369 313694 246397
rect 313270 246351 313322 246357
rect 313366 243893 313418 243899
rect 313366 243835 313418 243841
rect 313174 240341 313226 240347
rect 313174 240283 313226 240289
rect 312788 237050 312844 237059
rect 312788 236985 312844 236994
rect 312982 236049 313034 236055
rect 312982 235991 313034 235997
rect 312994 233484 313022 235991
rect 313378 233484 313406 243835
rect 313654 240341 313706 240347
rect 313654 240283 313706 240289
rect 313666 236647 313694 240283
rect 313750 239971 313802 239977
rect 313750 239913 313802 239919
rect 313654 236641 313706 236647
rect 313654 236583 313706 236589
rect 313762 233484 313790 239913
rect 313858 239237 313886 246494
rect 313954 246415 313982 246647
rect 313942 246409 313994 246415
rect 313942 246351 313994 246357
rect 314050 244639 314078 246721
rect 314038 244633 314090 244639
rect 314038 244575 314090 244581
rect 314338 243011 314366 246494
rect 314326 243005 314378 243011
rect 314326 242947 314378 242953
rect 314614 240267 314666 240273
rect 314614 240209 314666 240215
rect 314230 240119 314282 240125
rect 314230 240061 314282 240067
rect 313846 239231 313898 239237
rect 313846 239173 313898 239179
rect 313846 236641 313898 236647
rect 313846 236583 313898 236589
rect 312768 233456 313022 233484
rect 313152 233456 313406 233484
rect 313536 233456 313790 233484
rect 313858 233470 313886 236583
rect 314242 233470 314270 240061
rect 314626 233470 314654 240209
rect 314818 239385 314846 246494
rect 314914 246480 315168 246508
rect 315394 246480 315648 246508
rect 314914 244343 314942 246480
rect 314902 244337 314954 244343
rect 314902 244279 314954 244285
rect 315190 239823 315242 239829
rect 315190 239765 315242 239771
rect 314806 239379 314858 239385
rect 314806 239321 314858 239327
rect 315202 233484 315230 239765
rect 315394 236721 315422 246480
rect 315574 240415 315626 240421
rect 315574 240357 315626 240363
rect 315382 236715 315434 236721
rect 315382 236657 315434 236663
rect 315586 233484 315614 240357
rect 316066 240199 316094 246494
rect 316464 246480 316574 246508
rect 316944 246480 317246 246508
rect 317376 246480 317438 246508
rect 316054 240193 316106 240199
rect 316054 240135 316106 240141
rect 316150 240193 316202 240199
rect 316150 240135 316202 240141
rect 316162 239977 316190 240135
rect 316150 239971 316202 239977
rect 316150 239913 316202 239919
rect 316246 238861 316298 238867
rect 316246 238803 316298 238809
rect 316054 237455 316106 237461
rect 316054 237397 316106 237403
rect 315958 236197 316010 236203
rect 315958 236139 316010 236145
rect 315970 233484 315998 236139
rect 314976 233456 315230 233484
rect 315360 233456 315614 233484
rect 315744 233456 315998 233484
rect 316066 233470 316094 237397
rect 316258 237165 316286 238803
rect 316342 238639 316394 238645
rect 316342 238581 316394 238587
rect 316438 238639 316490 238645
rect 316438 238581 316490 238587
rect 316246 237159 316298 237165
rect 316246 237101 316298 237107
rect 316354 237017 316382 238581
rect 316342 237011 316394 237017
rect 316342 236953 316394 236959
rect 316450 233470 316478 238581
rect 316546 233983 316574 246480
rect 317218 246415 317246 246480
rect 317206 246409 317258 246415
rect 317206 246351 317258 246357
rect 316822 244781 316874 244787
rect 316918 244781 316970 244787
rect 316874 244741 316918 244769
rect 316822 244723 316874 244729
rect 316918 244723 316970 244729
rect 317026 244713 317150 244732
rect 317014 244707 317162 244713
rect 317066 244704 317110 244707
rect 317014 244649 317066 244655
rect 317110 244649 317162 244655
rect 317206 244189 317258 244195
rect 317206 244131 317258 244137
rect 316822 243967 316874 243973
rect 316822 243909 316874 243915
rect 316834 243085 316862 243909
rect 316918 243301 316970 243307
rect 316918 243243 316970 243249
rect 316822 243079 316874 243085
rect 316822 243021 316874 243027
rect 316930 242493 316958 243243
rect 317218 243233 317246 244131
rect 317206 243227 317258 243233
rect 317206 243169 317258 243175
rect 317410 242937 317438 246480
rect 317602 246480 317856 246508
rect 317986 246480 318192 246508
rect 318466 246480 318672 246508
rect 317494 246409 317546 246415
rect 317494 246351 317546 246357
rect 317398 242931 317450 242937
rect 317398 242873 317450 242879
rect 317506 242493 317534 246351
rect 316918 242487 316970 242493
rect 316918 242429 316970 242435
rect 317014 242487 317066 242493
rect 317014 242429 317066 242435
rect 317494 242487 317546 242493
rect 317494 242429 317546 242435
rect 316822 237381 316874 237387
rect 316822 237323 316874 237329
rect 316534 233977 316586 233983
rect 316534 233919 316586 233925
rect 316834 233470 316862 237323
rect 317026 233687 317054 242429
rect 317494 241525 317546 241531
rect 317494 241467 317546 241473
rect 317506 241309 317534 241467
rect 317494 241303 317546 241309
rect 317494 241245 317546 241251
rect 317398 238861 317450 238867
rect 317398 238803 317450 238809
rect 317014 233681 317066 233687
rect 317014 233623 317066 233629
rect 317410 233484 317438 238803
rect 317602 236499 317630 246480
rect 317878 241599 317930 241605
rect 317878 241541 317930 241547
rect 317782 239897 317834 239903
rect 317782 239839 317834 239845
rect 317590 236493 317642 236499
rect 317590 236435 317642 236441
rect 317794 233484 317822 239839
rect 317184 233456 317438 233484
rect 317568 233456 317822 233484
rect 317890 233484 317918 241541
rect 317986 234279 318014 246480
rect 318262 241451 318314 241457
rect 318262 241393 318314 241399
rect 318274 239163 318302 241393
rect 318262 239157 318314 239163
rect 318262 239099 318314 239105
rect 318166 238787 318218 238793
rect 318166 238729 318218 238735
rect 318070 238565 318122 238571
rect 318070 238507 318122 238513
rect 318082 236573 318110 238507
rect 318178 237239 318206 238729
rect 318262 238713 318314 238719
rect 318262 238655 318314 238661
rect 318166 237233 318218 237239
rect 318166 237175 318218 237181
rect 318274 237091 318302 238655
rect 318466 237313 318494 246480
rect 318550 238935 318602 238941
rect 318550 238877 318602 238883
rect 318454 237307 318506 237313
rect 318454 237249 318506 237255
rect 318262 237085 318314 237091
rect 318262 237027 318314 237033
rect 318070 236567 318122 236573
rect 318070 236509 318122 236515
rect 317974 234273 318026 234279
rect 317974 234215 318026 234221
rect 318562 233484 318590 238877
rect 318646 238713 318698 238719
rect 318646 238655 318698 238661
rect 317890 233456 317952 233484
rect 318288 233456 318590 233484
rect 318658 233470 318686 238655
rect 319030 238639 319082 238645
rect 319030 238581 319082 238587
rect 319042 233470 319070 238581
rect 319138 234205 319166 246494
rect 319330 246480 319584 246508
rect 319968 246480 320222 246508
rect 319330 236943 319358 246480
rect 319714 245009 319838 245028
rect 319702 245003 319838 245009
rect 319754 245000 319838 245003
rect 319702 244945 319754 244951
rect 319606 244633 319658 244639
rect 319606 244575 319658 244581
rect 319618 244343 319646 244575
rect 319810 244343 319838 245000
rect 319606 244337 319658 244343
rect 319606 244279 319658 244285
rect 319798 244337 319850 244343
rect 319798 244279 319850 244285
rect 320194 242419 320222 246480
rect 320386 242789 320414 246494
rect 320578 246480 320880 246508
rect 320374 242783 320426 242789
rect 320374 242725 320426 242731
rect 320182 242413 320234 242419
rect 320182 242355 320234 242361
rect 320470 241451 320522 241457
rect 320470 241393 320522 241399
rect 319606 238565 319658 238571
rect 319606 238507 319658 238513
rect 319318 236937 319370 236943
rect 319318 236879 319370 236885
rect 319126 234199 319178 234205
rect 319126 234141 319178 234147
rect 319618 233484 319646 238507
rect 319700 238086 319756 238095
rect 319700 238021 319756 238030
rect 319714 237059 319742 238021
rect 319990 237529 320042 237535
rect 319990 237471 320042 237477
rect 319700 237050 319756 237059
rect 319700 236985 319756 236994
rect 319700 236754 319756 236763
rect 319700 236689 319756 236698
rect 319714 236129 319742 236689
rect 319702 236123 319754 236129
rect 319702 236065 319754 236071
rect 320002 233484 320030 237471
rect 320374 236493 320426 236499
rect 320374 236435 320426 236441
rect 320386 233484 320414 236435
rect 319392 233456 319646 233484
rect 319776 233456 320030 233484
rect 320160 233456 320414 233484
rect 320482 233470 320510 241393
rect 320578 233909 320606 246480
rect 321238 244781 321290 244787
rect 321238 244723 321290 244729
rect 321250 244195 321278 244723
rect 321238 244189 321290 244195
rect 321238 244131 321290 244137
rect 321346 243159 321374 246494
rect 321442 246480 321696 246508
rect 321922 246480 322176 246508
rect 321334 243153 321386 243159
rect 321334 243095 321386 243101
rect 320854 239675 320906 239681
rect 320854 239617 320906 239623
rect 320566 233903 320618 233909
rect 320566 233845 320618 233851
rect 320866 233470 320894 239617
rect 321238 239231 321290 239237
rect 321238 239173 321290 239179
rect 321250 233470 321278 239173
rect 321442 233835 321470 246480
rect 321814 237307 321866 237313
rect 321814 237249 321866 237255
rect 321430 233829 321482 233835
rect 321430 233771 321482 233777
rect 321826 233484 321854 237249
rect 321922 234501 321950 246480
rect 322594 242641 322622 246494
rect 322786 246480 323088 246508
rect 322582 242635 322634 242641
rect 322582 242577 322634 242583
rect 322678 239749 322730 239755
rect 322678 239691 322730 239697
rect 322198 239379 322250 239385
rect 322198 239321 322250 239327
rect 321910 234495 321962 234501
rect 321910 234437 321962 234443
rect 322210 233484 322238 239321
rect 322486 236419 322538 236425
rect 322486 236361 322538 236367
rect 322498 233484 322526 236361
rect 321600 233456 321854 233484
rect 321984 233456 322238 233484
rect 322368 233456 322526 233484
rect 322690 233470 322718 239691
rect 322786 234649 322814 246480
rect 323458 242567 323486 246494
rect 323650 246480 323904 246508
rect 324130 246480 324384 246508
rect 323446 242561 323498 242567
rect 323446 242503 323498 242509
rect 323062 239601 323114 239607
rect 323062 239543 323114 239549
rect 322774 234643 322826 234649
rect 322774 234585 322826 234591
rect 323074 233470 323102 239543
rect 323446 239453 323498 239459
rect 323446 239395 323498 239401
rect 323458 233470 323486 239395
rect 323650 239015 323678 246480
rect 323638 239009 323690 239015
rect 323638 238951 323690 238957
rect 323734 238861 323786 238867
rect 323926 238861 323978 238867
rect 323786 238809 323926 238812
rect 323734 238803 323978 238809
rect 323746 238784 323966 238803
rect 324130 237165 324158 246480
rect 324706 239681 324734 246494
rect 325186 241901 325214 246494
rect 325474 246480 325680 246508
rect 325858 246480 326112 246508
rect 326496 246480 326750 246508
rect 325174 241895 325226 241901
rect 325174 241837 325226 241843
rect 325270 241895 325322 241901
rect 325270 241837 325322 241843
rect 325282 239829 325310 241837
rect 325270 239823 325322 239829
rect 325270 239765 325322 239771
rect 324694 239675 324746 239681
rect 324694 239617 324746 239623
rect 325474 239108 325502 246480
rect 324406 239083 324458 239089
rect 324406 239025 324458 239031
rect 325186 239080 325502 239108
rect 324214 238787 324266 238793
rect 324214 238729 324266 238735
rect 324118 237159 324170 237165
rect 324118 237101 324170 237107
rect 324022 236715 324074 236721
rect 324022 236657 324074 236663
rect 324034 233484 324062 236657
rect 324226 236203 324254 238729
rect 324214 236197 324266 236203
rect 324214 236139 324266 236145
rect 324418 233484 324446 239025
rect 324790 236863 324842 236869
rect 324790 236805 324842 236811
rect 324802 233484 324830 236805
rect 325186 233484 325214 239080
rect 325858 237017 325886 246480
rect 326722 241383 326750 246480
rect 326914 241531 326942 246494
rect 326902 241525 326954 241531
rect 327190 241525 327242 241531
rect 326902 241467 326954 241473
rect 327010 241473 327190 241476
rect 327010 241467 327242 241473
rect 327010 241457 327230 241467
rect 326998 241451 327230 241457
rect 327050 241448 327230 241451
rect 326998 241393 327050 241399
rect 326710 241377 326762 241383
rect 326710 241319 326762 241325
rect 326230 239823 326282 239829
rect 326230 239765 326282 239771
rect 325846 237011 325898 237017
rect 325846 236953 325898 236959
rect 325654 236789 325706 236795
rect 325654 236731 325706 236737
rect 325270 236641 325322 236647
rect 325270 236583 325322 236589
rect 323808 233456 324062 233484
rect 324192 233456 324446 233484
rect 324576 233456 324830 233484
rect 324912 233456 325214 233484
rect 325282 233470 325310 236583
rect 325666 233470 325694 236731
rect 326242 233484 326270 239765
rect 326998 239749 327050 239755
rect 326998 239691 327050 239697
rect 326614 239305 326666 239311
rect 326614 239247 326666 239253
rect 326626 233484 326654 239247
rect 327010 233484 327038 239691
rect 327394 239533 327422 246494
rect 327874 241013 327902 246494
rect 327970 246480 328224 246508
rect 327970 241827 327998 246480
rect 328450 246415 328478 246776
rect 328532 246753 328588 246762
rect 328916 246818 328972 246827
rect 328916 246753 328972 246762
rect 329300 246818 329356 246827
rect 329300 246753 329356 246762
rect 342548 246818 342604 246827
rect 342548 246753 342604 246762
rect 348596 246818 348652 246827
rect 348596 246753 348652 246762
rect 349076 246818 349132 246827
rect 349076 246753 349132 246762
rect 349652 246818 349708 246827
rect 349652 246753 349708 246762
rect 366452 246818 366508 246827
rect 366452 246753 366508 246762
rect 366836 246818 366892 246827
rect 366836 246753 366892 246762
rect 367316 246818 367372 246827
rect 367316 246753 367372 246762
rect 369524 246818 369580 246827
rect 370292 246818 370348 246827
rect 369524 246753 369580 246762
rect 370210 246776 370292 246804
rect 328546 246545 328574 246753
rect 328930 246563 328958 246753
rect 328918 246557 328970 246563
rect 328546 246517 328622 246545
rect 328438 246409 328490 246415
rect 328162 246332 328382 246360
rect 328594 246397 328622 246517
rect 328704 246480 328862 246508
rect 328918 246499 328970 246505
rect 328594 246369 328670 246397
rect 328438 246351 328490 246357
rect 328162 246193 328190 246332
rect 328354 246267 328382 246332
rect 328246 246261 328298 246267
rect 328246 246203 328298 246209
rect 328342 246261 328394 246267
rect 328342 246203 328394 246209
rect 328150 246187 328202 246193
rect 328150 246129 328202 246135
rect 328258 243973 328286 246203
rect 328642 244861 328670 246369
rect 328630 244855 328682 244861
rect 328630 244797 328682 244803
rect 328246 243967 328298 243973
rect 328246 243909 328298 243915
rect 328340 242970 328396 242979
rect 328340 242905 328396 242914
rect 328532 242970 328588 242979
rect 328532 242905 328588 242914
rect 328354 242641 328382 242905
rect 328436 242822 328492 242831
rect 328546 242808 328574 242905
rect 328492 242780 328574 242808
rect 328436 242757 328492 242766
rect 328726 242709 328778 242715
rect 328724 242674 328726 242683
rect 328778 242674 328780 242683
rect 328342 242635 328394 242641
rect 328724 242609 328780 242618
rect 328342 242577 328394 242583
rect 327958 241821 328010 241827
rect 327958 241763 328010 241769
rect 327862 241007 327914 241013
rect 327862 240949 327914 240955
rect 327958 241007 328010 241013
rect 327958 240949 328010 240955
rect 327970 239903 327998 240949
rect 327958 239897 328010 239903
rect 327958 239839 328010 239845
rect 328246 239897 328298 239903
rect 328246 239839 328298 239845
rect 327382 239527 327434 239533
rect 327382 239469 327434 239475
rect 327862 237159 327914 237165
rect 327862 237101 327914 237107
rect 327478 237011 327530 237017
rect 327478 236953 327530 236959
rect 327094 236937 327146 236943
rect 327094 236879 327146 236885
rect 326016 233456 326270 233484
rect 326400 233456 326654 233484
rect 326784 233456 327038 233484
rect 327106 233470 327134 236879
rect 327490 233470 327518 236953
rect 327874 233470 327902 237101
rect 328258 233484 328286 239839
rect 328834 238793 328862 246480
rect 328918 241377 328970 241383
rect 328918 241319 328970 241325
rect 328822 238787 328874 238793
rect 328822 238729 328874 238735
rect 328438 237973 328490 237979
rect 328438 237915 328490 237921
rect 328534 237973 328586 237979
rect 328534 237915 328586 237921
rect 328450 237184 328478 237915
rect 328546 237313 328574 237915
rect 328534 237307 328586 237313
rect 328534 237249 328586 237255
rect 328726 237307 328778 237313
rect 328726 237249 328778 237255
rect 328450 237156 328574 237184
rect 328546 236721 328574 237156
rect 328738 237091 328766 237249
rect 328726 237085 328778 237091
rect 328726 237027 328778 237033
rect 328822 237085 328874 237091
rect 328822 237027 328874 237033
rect 328534 236715 328586 236721
rect 328534 236657 328586 236663
rect 328342 236641 328394 236647
rect 328342 236583 328394 236589
rect 328354 236277 328382 236583
rect 328342 236271 328394 236277
rect 328342 236213 328394 236219
rect 328834 233484 328862 237027
rect 328224 233456 328286 233484
rect 328608 233456 328862 233484
rect 328930 233484 328958 241319
rect 329122 240051 329150 246494
rect 329314 244195 329342 246753
rect 330646 246557 330698 246563
rect 329302 244189 329354 244195
rect 329302 244131 329354 244137
rect 329302 241821 329354 241827
rect 329302 241763 329354 241769
rect 329110 240045 329162 240051
rect 329110 239987 329162 239993
rect 328930 233456 328992 233484
rect 329314 233470 329342 241763
rect 329602 241013 329630 246494
rect 329686 246187 329738 246193
rect 329686 246129 329738 246135
rect 329698 244787 329726 246129
rect 329686 244781 329738 244787
rect 329686 244723 329738 244729
rect 329986 241753 330014 246494
rect 330178 246480 330432 246508
rect 330646 246499 330698 246505
rect 329974 241747 330026 241753
rect 329974 241689 330026 241695
rect 330178 241605 330206 246480
rect 330658 245823 330686 246499
rect 330850 246480 330912 246508
rect 330646 245817 330698 245823
rect 330646 245759 330698 245765
rect 330742 245817 330794 245823
rect 330742 245759 330794 245765
rect 330754 245527 330782 245759
rect 330742 245521 330794 245527
rect 330742 245463 330794 245469
rect 330166 241599 330218 241605
rect 330166 241541 330218 241547
rect 330262 241599 330314 241605
rect 330262 241541 330314 241547
rect 329590 241007 329642 241013
rect 329590 240949 329642 240955
rect 330274 240144 330302 241541
rect 330742 241007 330794 241013
rect 330742 240949 330794 240955
rect 329986 240116 330302 240144
rect 329986 233484 330014 240116
rect 330070 240045 330122 240051
rect 330070 239987 330122 239993
rect 329712 233456 330014 233484
rect 330082 233470 330110 239987
rect 330646 238787 330698 238793
rect 330646 238729 330698 238735
rect 330550 238047 330602 238053
rect 330550 237989 330602 237995
rect 330562 236795 330590 237989
rect 330454 236789 330506 236795
rect 330454 236731 330506 236737
rect 330550 236789 330602 236795
rect 330550 236731 330602 236737
rect 330466 236351 330494 236731
rect 330454 236345 330506 236351
rect 330454 236287 330506 236293
rect 330658 233484 330686 238729
rect 330754 237313 330782 240949
rect 330742 237307 330794 237313
rect 330742 237249 330794 237255
rect 330850 237239 330878 246480
rect 331030 245373 331082 245379
rect 331030 245315 331082 245321
rect 331042 245231 331070 245315
rect 331030 245225 331082 245231
rect 331030 245167 331082 245173
rect 331030 241747 331082 241753
rect 331030 241689 331082 241695
rect 330934 238491 330986 238497
rect 330934 238433 330986 238439
rect 330946 238275 330974 238433
rect 330934 238269 330986 238275
rect 330934 238211 330986 238217
rect 330838 237233 330890 237239
rect 330838 237175 330890 237181
rect 331042 233484 331070 241689
rect 331330 239015 331358 246494
rect 331510 241451 331562 241457
rect 331510 241393 331562 241399
rect 331318 239009 331370 239015
rect 331318 238951 331370 238957
rect 331126 238491 331178 238497
rect 331126 238433 331178 238439
rect 330432 233456 330686 233484
rect 330816 233456 331070 233484
rect 331138 233484 331166 238433
rect 331138 233456 331200 233484
rect 331522 233470 331550 241393
rect 331714 239977 331742 246494
rect 331702 239971 331754 239977
rect 331702 239913 331754 239919
rect 332194 238719 332222 246494
rect 332386 246480 332640 246508
rect 332770 246480 333024 246508
rect 332278 241377 332330 241383
rect 332278 241319 332330 241325
rect 332182 238713 332234 238719
rect 332182 238655 332234 238661
rect 331798 237307 331850 237313
rect 331798 237249 331850 237255
rect 331810 236869 331838 237249
rect 331798 236863 331850 236869
rect 331798 236805 331850 236811
rect 331894 236863 331946 236869
rect 331894 236805 331946 236811
rect 331906 233470 331934 236805
rect 332290 233470 332318 241319
rect 332386 238645 332414 246480
rect 332770 239163 332798 246480
rect 332950 239527 333002 239533
rect 332950 239469 333002 239475
rect 332758 239157 332810 239163
rect 332758 239099 332810 239105
rect 332374 238639 332426 238645
rect 332374 238581 332426 238587
rect 332854 237233 332906 237239
rect 332854 237175 332906 237181
rect 332866 233484 332894 237175
rect 332962 233780 332990 239469
rect 333442 238571 333470 246494
rect 333634 246480 333936 246508
rect 333634 241013 333662 246480
rect 333622 241007 333674 241013
rect 333622 240949 333674 240955
rect 333718 241007 333770 241013
rect 333718 240949 333770 240955
rect 333622 238639 333674 238645
rect 333622 238581 333674 238587
rect 333430 238565 333482 238571
rect 333430 238507 333482 238513
rect 332962 233752 333038 233780
rect 332640 233456 332894 233484
rect 333010 233470 333038 233752
rect 333634 233484 333662 238581
rect 333408 233456 333662 233484
rect 333730 233470 333758 240949
rect 334102 238713 334154 238719
rect 334102 238655 334154 238661
rect 334114 233470 334142 238655
rect 334402 237535 334430 246494
rect 334498 246480 334752 246508
rect 334978 246480 335232 246508
rect 334498 241309 334526 246480
rect 334486 241303 334538 241309
rect 334486 241245 334538 241251
rect 334486 239971 334538 239977
rect 334486 239913 334538 239919
rect 334390 237529 334442 237535
rect 334390 237471 334442 237477
rect 334498 233470 334526 239913
rect 334870 238565 334922 238571
rect 334870 238507 334922 238513
rect 334882 233484 334910 238507
rect 334978 236499 335006 246480
rect 335350 244041 335402 244047
rect 335350 243983 335402 243989
rect 334966 236493 335018 236499
rect 334966 236435 335018 236441
rect 334964 235126 335020 235135
rect 334964 235061 335020 235070
rect 334848 233456 334910 233484
rect 334978 233484 335006 235061
rect 335362 233484 335390 243983
rect 335650 236573 335678 246494
rect 336130 241531 336158 246494
rect 336310 243227 336362 243233
rect 336310 243169 336362 243175
rect 336118 241525 336170 241531
rect 336118 241467 336170 241473
rect 335638 236567 335690 236573
rect 335638 236509 335690 236515
rect 335926 235531 335978 235537
rect 335926 235473 335978 235479
rect 334978 233456 335232 233484
rect 335362 233456 335616 233484
rect 335938 233470 335966 235473
rect 336322 233470 336350 243169
rect 336514 241679 336542 246494
rect 336960 246480 337022 246508
rect 336502 241673 336554 241679
rect 336502 241615 336554 241621
rect 336994 238423 337022 246480
rect 337186 246480 337440 246508
rect 337078 243079 337130 243085
rect 337078 243021 337130 243027
rect 336982 238417 337034 238423
rect 336982 238359 337034 238365
rect 336694 235679 336746 235685
rect 336694 235621 336746 235627
rect 336706 233470 336734 235621
rect 337090 233484 337118 243021
rect 337186 239237 337214 246480
rect 337558 244115 337610 244121
rect 337558 244057 337610 244063
rect 337174 239231 337226 239237
rect 337174 239173 337226 239179
rect 337174 235605 337226 235611
rect 337174 235547 337226 235553
rect 337056 233456 337118 233484
rect 337186 233484 337214 235547
rect 337570 233484 337598 244057
rect 337858 241161 337886 246494
rect 338134 244929 338186 244935
rect 338134 244871 338186 244877
rect 338146 244195 338174 244871
rect 338134 244189 338186 244195
rect 338134 244131 338186 244137
rect 338132 242970 338188 242979
rect 338132 242905 338188 242914
rect 338146 242863 338174 242905
rect 338134 242857 338186 242863
rect 338134 242799 338186 242805
rect 337846 241155 337898 241161
rect 337846 241097 337898 241103
rect 338242 237979 338270 246494
rect 338422 245151 338474 245157
rect 338422 245093 338474 245099
rect 338434 244935 338462 245093
rect 338422 244929 338474 244935
rect 338422 244871 338474 244877
rect 338326 244633 338378 244639
rect 338326 244575 338378 244581
rect 338230 237973 338282 237979
rect 338230 237915 338282 237921
rect 338134 235753 338186 235759
rect 338134 235695 338186 235701
rect 337186 233456 337440 233484
rect 337570 233456 337824 233484
rect 338146 233470 338174 235695
rect 338338 233484 338366 244575
rect 338516 243118 338572 243127
rect 338516 243053 338572 243062
rect 338530 242091 338558 243053
rect 338516 242082 338572 242091
rect 338516 242017 338572 242026
rect 338722 238275 338750 246494
rect 338914 246480 339168 246508
rect 339394 246480 339648 246508
rect 339862 246483 339914 246489
rect 338806 242635 338858 242641
rect 338806 242577 338858 242583
rect 338818 242091 338846 242577
rect 338804 242082 338860 242091
rect 338804 242017 338860 242026
rect 338914 239385 338942 246480
rect 339190 242857 339242 242863
rect 339190 242799 339242 242805
rect 339202 242683 339230 242799
rect 338996 242674 339052 242683
rect 338996 242609 339052 242618
rect 339188 242674 339244 242683
rect 339188 242609 339244 242618
rect 338902 239379 338954 239385
rect 338902 239321 338954 239327
rect 338710 238269 338762 238275
rect 338710 238211 338762 238217
rect 338518 237529 338570 237535
rect 338518 237471 338570 237477
rect 338530 237387 338558 237471
rect 338518 237381 338570 237387
rect 338518 237323 338570 237329
rect 338902 235827 338954 235833
rect 338902 235769 338954 235775
rect 338338 233456 338544 233484
rect 338914 233470 338942 235769
rect 339010 233484 339038 242609
rect 339394 241235 339422 246480
rect 340032 246480 340286 246508
rect 339862 246425 339914 246431
rect 339670 246187 339722 246193
rect 339670 246129 339722 246135
rect 339766 246187 339818 246193
rect 339766 246129 339818 246135
rect 339682 245305 339710 246129
rect 339670 245299 339722 245305
rect 339670 245241 339722 245247
rect 339478 245151 339530 245157
rect 339478 245093 339530 245099
rect 339490 244935 339518 245093
rect 339478 244929 339530 244935
rect 339478 244871 339530 244877
rect 339574 244855 339626 244861
rect 339574 244797 339626 244803
rect 339586 244639 339614 244797
rect 339574 244633 339626 244639
rect 339574 244575 339626 244581
rect 339778 243973 339806 246129
rect 339874 246064 339902 246425
rect 339958 246261 340010 246267
rect 340150 246261 340202 246267
rect 340010 246209 340150 246212
rect 339958 246203 340202 246209
rect 339970 246184 340190 246203
rect 339874 246036 340190 246064
rect 339958 245003 340010 245009
rect 339874 244963 339958 244991
rect 339874 244417 339902 244963
rect 339958 244945 340010 244951
rect 339958 244707 340010 244713
rect 339958 244649 340010 244655
rect 339862 244411 339914 244417
rect 339862 244353 339914 244359
rect 339766 243967 339818 243973
rect 339766 243909 339818 243915
rect 339862 242783 339914 242789
rect 339862 242725 339914 242731
rect 339382 241229 339434 241235
rect 339382 241171 339434 241177
rect 339670 241155 339722 241161
rect 339670 241097 339722 241103
rect 339682 236869 339710 241097
rect 339764 238086 339820 238095
rect 339764 238021 339820 238030
rect 339778 237059 339806 238021
rect 339764 237050 339820 237059
rect 339764 236985 339820 236994
rect 339670 236863 339722 236869
rect 339670 236805 339722 236811
rect 339764 236754 339820 236763
rect 339764 236689 339820 236698
rect 339778 236129 339806 236689
rect 339874 236425 339902 242725
rect 339862 236419 339914 236425
rect 339862 236361 339914 236367
rect 339766 236123 339818 236129
rect 339766 236065 339818 236071
rect 339382 235975 339434 235981
rect 339382 235917 339434 235923
rect 339394 233484 339422 235917
rect 339970 233484 339998 244649
rect 340162 244639 340190 246036
rect 340150 244633 340202 244639
rect 340150 244575 340202 244581
rect 340258 242789 340286 246480
rect 340246 242783 340298 242789
rect 340246 242725 340298 242731
rect 340450 238201 340478 246494
rect 340726 243301 340778 243307
rect 340726 243243 340778 243249
rect 340438 238195 340490 238201
rect 340438 238137 340490 238143
rect 340342 235901 340394 235907
rect 340342 235843 340394 235849
rect 339010 233456 339264 233484
rect 339394 233456 339648 233484
rect 339970 233456 340032 233484
rect 340354 233470 340382 235843
rect 340738 233470 340766 243243
rect 340930 239681 340958 246494
rect 341204 242822 341260 242831
rect 341204 242757 341260 242766
rect 340918 239675 340970 239681
rect 340918 239617 340970 239623
rect 341108 235274 341164 235283
rect 341108 235209 341164 235218
rect 341122 233470 341150 235209
rect 341218 233484 341246 242757
rect 341314 239607 341342 246494
rect 341506 246480 341760 246508
rect 341986 246480 342240 246508
rect 341302 239601 341354 239607
rect 341302 239543 341354 239549
rect 341506 238127 341534 246480
rect 341986 239459 342014 246480
rect 342562 244713 342590 246753
rect 342742 246557 342794 246563
rect 347254 246557 347306 246563
rect 342742 246499 342794 246505
rect 342550 244707 342602 244713
rect 342550 244649 342602 244655
rect 342068 242378 342124 242387
rect 342068 242313 342124 242322
rect 341974 239453 342026 239459
rect 341974 239395 342026 239401
rect 341494 238121 341546 238127
rect 341494 238063 341546 238069
rect 341588 235718 341644 235727
rect 341588 235653 341644 235662
rect 341602 233484 341630 235653
rect 342082 233484 342110 242313
rect 342658 240939 342686 246494
rect 342754 243307 342782 246499
rect 342742 243301 342794 243307
rect 342742 243243 342794 243249
rect 342932 242230 342988 242239
rect 342932 242165 342988 242174
rect 342646 240933 342698 240939
rect 342646 240875 342698 240881
rect 342742 238121 342794 238127
rect 342740 238086 342742 238095
rect 342794 238086 342796 238095
rect 342740 238021 342796 238030
rect 342754 237563 342878 237591
rect 342754 237535 342782 237563
rect 342742 237529 342794 237535
rect 342742 237471 342794 237477
rect 342850 237387 342878 237563
rect 342838 237381 342890 237387
rect 342838 237323 342890 237329
rect 342548 235570 342604 235579
rect 342548 235505 342604 235514
rect 341218 233456 341472 233484
rect 341602 233456 341856 233484
rect 342082 233456 342240 233484
rect 342562 233470 342590 235505
rect 342946 233470 342974 242165
rect 343042 236647 343070 246494
rect 343412 242674 343468 242683
rect 343412 242609 343468 242618
rect 343030 236641 343082 236647
rect 343030 236583 343082 236589
rect 343316 235422 343372 235431
rect 343316 235357 343372 235366
rect 343330 233470 343358 235357
rect 343426 233484 343454 242609
rect 343522 238053 343550 246494
rect 343714 246480 343968 246508
rect 344194 246480 344448 246508
rect 343714 239089 343742 246480
rect 344194 240865 344222 246480
rect 344276 242082 344332 242091
rect 344276 242017 344332 242026
rect 344182 240859 344234 240865
rect 344182 240801 344234 240807
rect 343702 239083 343754 239089
rect 343702 239025 343754 239031
rect 343510 238047 343562 238053
rect 343510 237989 343562 237995
rect 343796 235866 343852 235875
rect 343796 235801 343852 235810
rect 343810 233484 343838 235801
rect 344290 233484 344318 242017
rect 344770 237313 344798 246494
rect 345142 243449 345194 243455
rect 345142 243391 345194 243397
rect 344758 237307 344810 237313
rect 344758 237249 344810 237255
rect 344756 236162 344812 236171
rect 344756 236097 344812 236106
rect 343426 233456 343680 233484
rect 343810 233456 344064 233484
rect 344290 233456 344448 233484
rect 344770 233470 344798 236097
rect 345154 233470 345182 243391
rect 345250 236795 345278 246494
rect 345622 243523 345674 243529
rect 345622 243465 345674 243471
rect 345238 236789 345290 236795
rect 345238 236731 345290 236737
rect 345526 234717 345578 234723
rect 345526 234659 345578 234665
rect 345538 233470 345566 234659
rect 345634 233484 345662 243465
rect 345730 240717 345758 246494
rect 345922 246480 346176 246508
rect 346306 246480 346560 246508
rect 347254 246499 347306 246505
rect 345718 240711 345770 240717
rect 345718 240653 345770 240659
rect 345922 236277 345950 246480
rect 346306 240569 346334 246480
rect 346390 243375 346442 243381
rect 346390 243317 346442 243323
rect 346294 240563 346346 240569
rect 346294 240505 346346 240511
rect 345910 236271 345962 236277
rect 345910 236213 345962 236219
rect 346004 236014 346060 236023
rect 346004 235949 346060 235958
rect 346018 233484 346046 235949
rect 346402 233484 346430 243317
rect 346978 236351 347006 246494
rect 347266 246415 347294 246499
rect 347254 246409 347306 246415
rect 347254 246351 347306 246357
rect 347350 243671 347402 243677
rect 347350 243613 347402 243619
rect 346966 236345 347018 236351
rect 346966 236287 347018 236293
rect 346966 234791 347018 234797
rect 346966 234733 347018 234739
rect 345634 233456 345888 233484
rect 346018 233456 346272 233484
rect 346402 233456 346656 233484
rect 346978 233470 347006 234733
rect 347362 233470 347390 243613
rect 347458 236721 347486 246494
rect 347830 242117 347882 242123
rect 347830 242059 347882 242065
rect 347446 236715 347498 236721
rect 347446 236657 347498 236663
rect 347732 234386 347788 234395
rect 347732 234321 347788 234330
rect 347746 233470 347774 234321
rect 347842 233484 347870 242059
rect 347938 239829 347966 246494
rect 348288 246480 348350 246508
rect 348214 246335 348266 246341
rect 348214 246277 348266 246283
rect 348226 246193 348254 246277
rect 348214 246187 348266 246193
rect 348214 246129 348266 246135
rect 348322 240643 348350 246480
rect 348610 246415 348638 246753
rect 348768 246480 349022 246508
rect 349090 246489 349118 246753
rect 349666 246563 349694 246753
rect 366466 246563 366494 246753
rect 349654 246557 349706 246563
rect 366454 246557 366506 246563
rect 349654 246499 349706 246505
rect 348598 246409 348650 246415
rect 348598 246351 348650 246357
rect 348406 246187 348458 246193
rect 348502 246187 348554 246193
rect 348458 246147 348502 246175
rect 348406 246129 348458 246135
rect 348502 246129 348554 246135
rect 348514 245888 348926 245916
rect 348514 245749 348542 245888
rect 348502 245743 348554 245749
rect 348502 245685 348554 245691
rect 348598 245743 348650 245749
rect 348598 245685 348650 245691
rect 348610 245620 348638 245685
rect 348514 245592 348638 245620
rect 348514 245527 348542 245592
rect 348502 245521 348554 245527
rect 348502 245463 348554 245469
rect 348694 245447 348746 245453
rect 348694 245389 348746 245395
rect 348706 244861 348734 245389
rect 348898 244935 348926 245888
rect 348886 244929 348938 244935
rect 348886 244871 348938 244877
rect 348694 244855 348746 244861
rect 348694 244797 348746 244803
rect 348598 242043 348650 242049
rect 348598 241985 348650 241991
rect 348310 240637 348362 240643
rect 348310 240579 348362 240585
rect 347926 239823 347978 239829
rect 347926 239765 347978 239771
rect 348418 238941 348542 238960
rect 348406 238935 348554 238941
rect 348458 238932 348502 238935
rect 348406 238877 348458 238883
rect 348502 238877 348554 238883
rect 348212 234978 348268 234987
rect 348212 234913 348268 234922
rect 348226 233484 348254 234913
rect 348610 233484 348638 241985
rect 348994 239311 349022 246480
rect 349078 246483 349130 246489
rect 349078 246425 349130 246431
rect 348982 239305 349034 239311
rect 348982 239247 349034 239253
rect 349186 237905 349214 246494
rect 349366 246187 349418 246193
rect 349366 246129 349418 246135
rect 349378 244269 349406 246129
rect 349366 244263 349418 244269
rect 349366 244205 349418 244211
rect 349270 243597 349322 243603
rect 349270 243539 349322 243545
rect 349174 237899 349226 237905
rect 349174 237841 349226 237847
rect 349172 234534 349228 234543
rect 349172 234469 349228 234478
rect 347842 233456 348096 233484
rect 348226 233456 348480 233484
rect 348610 233456 348864 233484
rect 349186 233470 349214 234469
rect 349282 233484 349310 243539
rect 349570 239755 349598 246494
rect 349762 246480 350064 246508
rect 350242 246480 350496 246508
rect 350722 246480 350976 246508
rect 349558 239749 349610 239755
rect 349558 239691 349610 239697
rect 349762 236943 349790 246480
rect 349942 246409 349994 246415
rect 349942 246351 349994 246357
rect 349954 244639 349982 246351
rect 349942 244633 349994 244639
rect 349942 244575 349994 244581
rect 350038 242191 350090 242197
rect 350038 242133 350090 242139
rect 349750 236937 349802 236943
rect 349750 236879 349802 236885
rect 349942 235087 349994 235093
rect 349942 235029 349994 235035
rect 349282 233456 349584 233484
rect 349954 233470 349982 235029
rect 350050 233484 350078 242133
rect 350242 240495 350270 246480
rect 350230 240489 350282 240495
rect 350230 240431 350282 240437
rect 350722 237017 350750 246480
rect 350806 243745 350858 243751
rect 350806 243687 350858 243693
rect 350710 237011 350762 237017
rect 350710 236953 350762 236959
rect 350422 234865 350474 234871
rect 350422 234807 350474 234813
rect 350434 233484 350462 234807
rect 350818 233484 350846 243687
rect 351298 240019 351326 246494
rect 351490 246480 351792 246508
rect 351970 246480 352272 246508
rect 352450 246480 352704 246508
rect 352834 246480 353088 246508
rect 351284 240010 351340 240019
rect 351284 239945 351340 239954
rect 351380 239122 351436 239131
rect 351380 239057 351436 239066
rect 351094 239009 351146 239015
rect 351094 238951 351146 238957
rect 351106 238867 351134 238951
rect 351094 238861 351146 238867
rect 351094 238803 351146 238809
rect 351190 238861 351242 238867
rect 351190 238803 351242 238809
rect 351202 238497 351230 238803
rect 351190 238491 351242 238497
rect 351190 238433 351242 238439
rect 351394 238423 351422 239057
rect 351382 238417 351434 238423
rect 351382 238359 351434 238365
rect 351490 237165 351518 246480
rect 351574 244189 351626 244195
rect 351574 244131 351626 244137
rect 351586 237165 351614 244131
rect 351766 241969 351818 241975
rect 351766 241911 351818 241917
rect 351478 237159 351530 237165
rect 351478 237101 351530 237107
rect 351574 237159 351626 237165
rect 351574 237101 351626 237107
rect 351382 234939 351434 234945
rect 351382 234881 351434 234887
rect 350050 233456 350304 233484
rect 350434 233456 350688 233484
rect 350818 233456 351072 233484
rect 351394 233470 351422 234881
rect 351778 233470 351806 241911
rect 351970 237757 351998 246480
rect 352244 242822 352300 242831
rect 352244 242757 352300 242766
rect 351958 237751 352010 237757
rect 351958 237693 352010 237699
rect 352150 235161 352202 235167
rect 352150 235103 352202 235109
rect 352162 233470 352190 235103
rect 352258 233484 352286 242757
rect 352450 239903 352478 246480
rect 352834 240167 352862 246480
rect 353014 242265 353066 242271
rect 353014 242207 353066 242213
rect 352820 240158 352876 240167
rect 352820 240093 352876 240102
rect 352438 239897 352490 239903
rect 352438 239839 352490 239845
rect 352630 235013 352682 235019
rect 352630 234955 352682 234961
rect 352642 233484 352670 234955
rect 353026 233484 353054 242207
rect 353506 237091 353534 246494
rect 353686 243819 353738 243825
rect 353686 243761 353738 243767
rect 353494 237085 353546 237091
rect 353494 237027 353546 237033
rect 353590 235383 353642 235389
rect 353590 235325 353642 235331
rect 352258 233456 352512 233484
rect 352642 233456 352896 233484
rect 353026 233456 353280 233484
rect 353602 233470 353630 235325
rect 353698 233484 353726 243761
rect 353986 237831 354014 246494
rect 354466 241647 354494 246494
rect 354562 246480 354816 246508
rect 355042 246480 355296 246508
rect 354562 241827 354590 246480
rect 354644 243118 354700 243127
rect 354644 243053 354700 243062
rect 354550 241821 354602 241827
rect 354550 241763 354602 241769
rect 354452 241638 354508 241647
rect 354452 241573 354508 241582
rect 353974 237825 354026 237831
rect 353974 237767 354026 237773
rect 354358 235235 354410 235241
rect 354358 235177 354410 235183
rect 353698 233456 354000 233484
rect 354370 233470 354398 235177
rect 354658 233780 354686 243053
rect 355042 237683 355070 246480
rect 355222 242339 355274 242345
rect 355222 242281 355274 242287
rect 355030 237677 355082 237683
rect 355030 237619 355082 237625
rect 354838 235309 354890 235315
rect 354838 235251 354890 235257
rect 354658 233752 354734 233780
rect 354706 233470 354734 233752
rect 354850 233484 354878 235251
rect 355234 233484 355262 242281
rect 355714 241605 355742 246494
rect 355798 245521 355850 245527
rect 355798 245463 355850 245469
rect 355702 241599 355754 241605
rect 355702 241541 355754 241547
rect 354850 233456 355104 233484
rect 355234 233456 355488 233484
rect 355810 233470 355838 245463
rect 355894 245225 355946 245231
rect 355894 245167 355946 245173
rect 355906 233484 355934 245167
rect 356194 237609 356222 246494
rect 356278 245891 356330 245897
rect 356278 245833 356330 245839
rect 356182 237603 356234 237609
rect 356182 237545 356234 237551
rect 356290 233484 356318 245833
rect 356578 240051 356606 246494
rect 356770 246480 357024 246508
rect 357250 246480 357504 246508
rect 356770 241795 356798 246480
rect 357142 245817 357194 245823
rect 357142 245759 357194 245765
rect 356756 241786 356812 241795
rect 356756 241721 356812 241730
rect 356566 240045 356618 240051
rect 356566 239987 356618 239993
rect 356662 235457 356714 235463
rect 356662 235399 356714 235405
rect 356674 233484 356702 235399
rect 357154 233484 357182 245759
rect 357250 238793 357278 246480
rect 357430 245743 357482 245749
rect 357430 245685 357482 245691
rect 357238 238787 357290 238793
rect 357238 238729 357290 238735
rect 357442 233484 357470 245685
rect 357826 237207 357854 246494
rect 358006 244929 358058 244935
rect 358006 244871 358058 244877
rect 357812 237198 357868 237207
rect 357812 237133 357868 237142
rect 355906 233456 356208 233484
rect 356290 233456 356592 233484
rect 356674 233456 356928 233484
rect 357154 233456 357312 233484
rect 357442 233456 357696 233484
rect 358018 233470 358046 244871
rect 358306 241753 358334 246494
rect 358390 243301 358442 243307
rect 358390 243243 358442 243249
rect 358294 241747 358346 241753
rect 358294 241689 358346 241695
rect 358402 233470 358430 243243
rect 358786 238867 358814 246494
rect 358978 246480 359232 246508
rect 359362 246480 359616 246508
rect 358978 241203 359006 246480
rect 359362 241457 359390 246480
rect 359350 241451 359402 241457
rect 359350 241393 359402 241399
rect 358964 241194 359020 241203
rect 358964 241129 359020 241138
rect 358774 238861 358826 238867
rect 358774 238803 358826 238809
rect 358870 238417 358922 238423
rect 358870 238359 358922 238365
rect 358774 237159 358826 237165
rect 358774 237101 358826 237107
rect 358786 233470 358814 237101
rect 358882 233484 358910 238359
rect 359830 237899 359882 237905
rect 359830 237841 359882 237847
rect 359252 236606 359308 236615
rect 359252 236541 359308 236550
rect 359266 233484 359294 236541
rect 358882 233456 359136 233484
rect 359266 233456 359520 233484
rect 296084 233433 296140 233442
rect 359842 233336 359870 237841
rect 360034 237503 360062 246494
rect 360514 241161 360542 246494
rect 360706 246480 361008 246508
rect 361090 246480 361344 246508
rect 361666 246480 361824 246508
rect 360598 241821 360650 241827
rect 360598 241763 360650 241769
rect 360502 241155 360554 241161
rect 360502 241097 360554 241103
rect 360214 239157 360266 239163
rect 360214 239099 360266 239105
rect 360020 237494 360076 237503
rect 360020 237429 360076 237438
rect 360226 233470 360254 239099
rect 360610 233470 360638 241763
rect 360706 238687 360734 246480
rect 361090 241383 361118 246480
rect 361558 241673 361610 241679
rect 361558 241615 361610 241621
rect 361078 241377 361130 241383
rect 361078 241319 361130 241325
rect 360982 239231 361034 239237
rect 360982 239173 361034 239179
rect 360692 238678 360748 238687
rect 360692 238613 360748 238622
rect 360886 238565 360938 238571
rect 360886 238507 360938 238513
rect 360898 237387 360926 238507
rect 360886 237381 360938 237387
rect 360886 237323 360938 237329
rect 360994 233470 361022 239173
rect 361570 233484 361598 241615
rect 361666 241055 361694 246480
rect 361942 241303 361994 241309
rect 361942 241245 361994 241251
rect 361652 241046 361708 241055
rect 361652 240981 361708 240990
rect 361954 233484 361982 241245
rect 362242 237239 362270 246494
rect 362326 241451 362378 241457
rect 362326 241393 362378 241399
rect 362230 237233 362282 237239
rect 362230 237175 362282 237181
rect 362338 233484 362366 241393
rect 362422 241229 362474 241235
rect 362422 241171 362474 241177
rect 361344 233456 361598 233484
rect 361728 233456 361982 233484
rect 362112 233456 362366 233484
rect 362434 233470 362462 241171
rect 362722 237355 362750 246494
rect 363106 240759 363134 246494
rect 363298 246480 363552 246508
rect 363874 246480 364032 246508
rect 363190 241747 363242 241753
rect 363190 241689 363242 241695
rect 363092 240750 363148 240759
rect 363092 240685 363148 240694
rect 362708 237346 362764 237355
rect 362708 237281 362764 237290
rect 362806 237233 362858 237239
rect 362806 237175 362858 237181
rect 362818 233470 362846 237175
rect 363202 233470 363230 241689
rect 363298 238645 363326 246480
rect 363766 241525 363818 241531
rect 363766 241467 363818 241473
rect 363286 238639 363338 238645
rect 363286 238581 363338 238587
rect 363778 233484 363806 241467
rect 363874 238539 363902 246480
rect 364150 241377 364202 241383
rect 364150 241319 364202 241325
rect 363860 238530 363916 238539
rect 363860 238465 363916 238474
rect 364162 233484 364190 241319
rect 364354 241013 364382 246494
rect 364534 241155 364586 241161
rect 364534 241097 364586 241103
rect 364342 241007 364394 241013
rect 364342 240949 364394 240955
rect 364546 233484 364574 241097
rect 364630 240711 364682 240717
rect 364630 240653 364682 240659
rect 363552 233456 363806 233484
rect 363936 233456 364190 233484
rect 364320 233456 364574 233484
rect 364642 233470 364670 240653
rect 364834 240611 364862 246494
rect 365014 240933 365066 240939
rect 365014 240875 365066 240881
rect 364820 240602 364876 240611
rect 364820 240537 364876 240546
rect 365026 233470 365054 240875
rect 365314 238719 365342 246494
rect 365760 246480 365822 246508
rect 365398 240637 365450 240643
rect 365398 240579 365450 240585
rect 365302 238713 365354 238719
rect 365302 238655 365354 238661
rect 365410 233470 365438 240579
rect 365794 238243 365822 246480
rect 365890 246480 366144 246508
rect 366454 246499 366506 246505
rect 365890 239977 365918 246480
rect 366358 241007 366410 241013
rect 366358 240949 366410 240955
rect 365974 240563 366026 240569
rect 365974 240505 366026 240511
rect 365878 239971 365930 239977
rect 365878 239913 365930 239919
rect 365780 238234 365836 238243
rect 365780 238169 365836 238178
rect 365986 233484 366014 240505
rect 366370 233484 366398 240949
rect 366562 240463 366590 246494
rect 366850 245897 366878 246753
rect 367330 246545 367358 246753
rect 367414 246557 367466 246563
rect 367330 246517 367414 246545
rect 367990 246557 368042 246563
rect 367414 246499 367466 246505
rect 366838 245891 366890 245897
rect 366838 245833 366890 245839
rect 366742 240489 366794 240495
rect 366548 240454 366604 240463
rect 366742 240431 366794 240437
rect 366548 240389 366604 240398
rect 366754 233484 366782 240431
rect 366838 238861 366890 238867
rect 366838 238803 366890 238809
rect 365760 233456 366014 233484
rect 366144 233456 366398 233484
rect 366528 233456 366782 233484
rect 366850 233470 366878 238803
rect 367042 238497 367070 246494
rect 367222 246483 367274 246489
rect 367222 246425 367274 246431
rect 367234 245749 367262 246425
rect 367522 245971 367550 246494
rect 367872 246480 367934 246508
rect 368470 246557 368522 246563
rect 367990 246499 368042 246505
rect 367510 245965 367562 245971
rect 367510 245907 367562 245913
rect 367222 245743 367274 245749
rect 367222 245685 367274 245691
rect 367906 244565 367934 246480
rect 368002 245823 368030 246499
rect 368098 246480 368352 246508
rect 368470 246499 368522 246505
rect 368098 246045 368126 246480
rect 368482 246415 368510 246499
rect 368470 246409 368522 246415
rect 368470 246351 368522 246357
rect 368086 246039 368138 246045
rect 368086 245981 368138 245987
rect 367990 245817 368042 245823
rect 367990 245759 368042 245765
rect 367894 244559 367946 244565
rect 367894 244501 367946 244507
rect 368770 244491 368798 246494
rect 369250 245675 369278 246494
rect 369538 246415 369566 246753
rect 369526 246409 369578 246415
rect 369526 246351 369578 246357
rect 369238 245669 369290 245675
rect 369238 245611 369290 245617
rect 368758 244485 368810 244491
rect 368758 244427 368810 244433
rect 367222 240859 367274 240865
rect 367222 240801 367274 240807
rect 367030 238491 367082 238497
rect 367030 238433 367082 238439
rect 367234 233470 367262 240801
rect 367604 240454 367660 240463
rect 367604 240389 367660 240398
rect 367618 233470 367646 240389
rect 368470 238491 368522 238497
rect 368470 238433 368522 238439
rect 367942 233755 367994 233761
rect 367942 233697 367994 233703
rect 367954 233470 367982 233697
rect 368482 233484 368510 238433
rect 369430 238417 369482 238423
rect 369430 238359 369482 238365
rect 369046 237381 369098 237387
rect 369046 237323 369098 237329
rect 368950 236271 369002 236277
rect 368950 236213 369002 236219
rect 368962 233484 368990 236213
rect 368352 233456 368510 233484
rect 368736 233456 368990 233484
rect 369058 233470 369086 237323
rect 369442 233470 369470 238359
rect 369634 236055 369662 246494
rect 369826 246480 370080 246508
rect 369826 240315 369854 246480
rect 370210 245749 370238 246776
rect 370292 246753 370348 246762
rect 370676 246818 370732 246827
rect 370676 246753 370732 246762
rect 373460 246818 373516 246827
rect 373460 246753 373516 246762
rect 389012 246818 389068 246827
rect 389012 246753 389068 246762
rect 389300 246818 389356 246827
rect 389300 246753 389356 246762
rect 390260 246818 390316 246827
rect 405908 246818 405964 246827
rect 390260 246753 390316 246762
rect 397270 246779 397322 246785
rect 370306 246480 370560 246508
rect 370198 245743 370250 245749
rect 370198 245685 370250 245691
rect 370102 245373 370154 245379
rect 370102 245315 370154 245321
rect 369910 245299 369962 245305
rect 370114 245287 370142 245315
rect 370198 245299 370250 245305
rect 370114 245259 370198 245287
rect 369910 245241 369962 245247
rect 370198 245241 370250 245247
rect 369922 245157 369950 245241
rect 369910 245151 369962 245157
rect 369910 245093 369962 245099
rect 370306 243899 370334 246480
rect 370690 246415 370718 246753
rect 370678 246409 370730 246415
rect 370678 246351 370730 246357
rect 370978 245601 371006 246494
rect 370966 245595 371018 245601
rect 370966 245537 371018 245543
rect 370294 243893 370346 243899
rect 370294 243835 370346 243841
rect 369812 240306 369868 240315
rect 369812 240241 369868 240250
rect 371362 240199 371390 246494
rect 371842 240347 371870 246494
rect 372034 246480 372288 246508
rect 372418 246480 372672 246508
rect 372898 246480 373152 246508
rect 372034 245083 372062 246480
rect 372022 245077 372074 245083
rect 372022 245019 372074 245025
rect 371830 240341 371882 240347
rect 371830 240283 371882 240289
rect 371350 240193 371402 240199
rect 371350 240135 371402 240141
rect 372418 240125 372446 246480
rect 372898 241499 372926 246480
rect 372982 246409 373034 246415
rect 372982 246351 373034 246357
rect 372994 245897 373022 246351
rect 372982 245891 373034 245897
rect 372982 245833 373034 245839
rect 373474 245823 373502 246753
rect 373462 245817 373514 245823
rect 373462 245759 373514 245765
rect 372884 241490 372940 241499
rect 372884 241425 372940 241434
rect 373570 240273 373598 246494
rect 374050 245009 374078 246494
rect 374038 245003 374090 245009
rect 374038 244945 374090 244951
rect 374434 241901 374462 246494
rect 374626 246480 374880 246508
rect 375106 246480 375360 246508
rect 374626 244861 374654 246480
rect 374614 244855 374666 244861
rect 374614 244797 374666 244803
rect 374422 241895 374474 241901
rect 374422 241837 374474 241843
rect 375106 240421 375134 246480
rect 375778 240791 375806 246494
rect 376054 241895 376106 241901
rect 376054 241837 376106 241843
rect 375766 240785 375818 240791
rect 375766 240727 375818 240733
rect 375094 240415 375146 240421
rect 375094 240357 375146 240363
rect 373558 240267 373610 240273
rect 373558 240209 373610 240215
rect 372406 240119 372458 240125
rect 372406 240061 372458 240067
rect 374806 239749 374858 239755
rect 374806 239691 374858 239697
rect 373846 239675 373898 239681
rect 373846 239617 373898 239623
rect 373366 239083 373418 239089
rect 373366 239025 373418 239031
rect 370390 238639 370442 238645
rect 370390 238581 370442 238587
rect 369814 238195 369866 238201
rect 369814 238137 369866 238143
rect 369622 236049 369674 236055
rect 369622 235991 369674 235997
rect 369826 233470 369854 238137
rect 370006 238121 370058 238127
rect 370004 238086 370006 238095
rect 370058 238086 370060 238095
rect 370004 238021 370060 238030
rect 370402 233484 370430 238581
rect 371638 238269 371690 238275
rect 371638 238211 371690 238217
rect 371158 238121 371210 238127
rect 371158 238063 371210 238069
rect 370774 236863 370826 236869
rect 370774 236805 370826 236811
rect 370786 233484 370814 236805
rect 371170 233484 371198 238063
rect 371254 237973 371306 237979
rect 371254 237915 371306 237921
rect 370176 233456 370430 233484
rect 370560 233456 370814 233484
rect 370944 233456 371198 233484
rect 371266 233470 371294 237915
rect 371650 233470 371678 238211
rect 372022 238047 372074 238053
rect 372022 237989 372074 237995
rect 372034 233470 372062 237989
rect 372598 237455 372650 237461
rect 372598 237397 372650 237403
rect 372610 233484 372638 237397
rect 372982 237159 373034 237165
rect 372982 237101 373034 237107
rect 372994 233484 373022 237101
rect 373378 233484 373406 239025
rect 373462 237677 373514 237683
rect 373462 237619 373514 237625
rect 372384 233456 372638 233484
rect 372768 233456 373022 233484
rect 373152 233456 373406 233484
rect 373474 233470 373502 237619
rect 373858 233470 373886 239617
rect 374230 237603 374282 237609
rect 374230 237545 374282 237551
rect 374242 233470 374270 237545
rect 374818 233484 374846 239691
rect 375670 239231 375722 239237
rect 375670 239173 375722 239179
rect 375190 239157 375242 239163
rect 375190 239099 375242 239105
rect 375202 233484 375230 239099
rect 375574 237825 375626 237831
rect 375574 237767 375626 237773
rect 375586 233484 375614 237767
rect 374592 233456 374846 233484
rect 374976 233456 375230 233484
rect 375360 233456 375614 233484
rect 375682 233470 375710 239173
rect 376066 233470 376094 241837
rect 376162 241087 376190 246494
rect 376150 241081 376202 241087
rect 376150 241023 376202 241029
rect 376438 240193 376490 240199
rect 376438 240135 376490 240141
rect 376450 233470 376478 240135
rect 376642 237535 376670 246494
rect 376834 246480 377088 246508
rect 377314 246480 377568 246508
rect 376834 241351 376862 246480
rect 376820 241342 376876 241351
rect 376820 241277 376876 241286
rect 377206 240267 377258 240273
rect 377206 240209 377258 240215
rect 377014 240119 377066 240125
rect 377014 240061 377066 240067
rect 376630 237529 376682 237535
rect 376630 237471 376682 237477
rect 376726 237529 376778 237535
rect 376726 237471 376778 237477
rect 376738 233761 376766 237471
rect 376726 233755 376778 233761
rect 376726 233697 376778 233703
rect 377026 233484 377054 240061
rect 377218 233780 377246 240209
rect 377314 238941 377342 246480
rect 377890 240907 377918 246494
rect 377876 240898 377932 240907
rect 377876 240833 377932 240842
rect 378262 240415 378314 240421
rect 378262 240357 378314 240363
rect 377782 240341 377834 240347
rect 377782 240283 377834 240289
rect 377302 238935 377354 238941
rect 377302 238877 377354 238883
rect 376800 233456 377054 233484
rect 377170 233752 377246 233780
rect 377170 233470 377198 233752
rect 377794 233484 377822 240283
rect 377878 239971 377930 239977
rect 377878 239913 377930 239919
rect 377568 233456 377822 233484
rect 377890 233470 377918 239913
rect 378274 233470 378302 240357
rect 378370 238571 378398 246494
rect 378646 241821 378698 241827
rect 378646 241763 378698 241769
rect 378742 241821 378794 241827
rect 378742 241763 378794 241769
rect 378658 241679 378686 241763
rect 378646 241673 378698 241679
rect 378646 241615 378698 241621
rect 378754 241605 378782 241763
rect 378742 241599 378794 241605
rect 378742 241541 378794 241547
rect 378646 239897 378698 239903
rect 378646 239839 378698 239845
rect 378358 238565 378410 238571
rect 378358 238507 378410 238513
rect 378658 233470 378686 239839
rect 378850 238391 378878 246494
rect 379042 246480 379296 246508
rect 379426 246480 379680 246508
rect 379042 239015 379070 246480
rect 379222 241081 379274 241087
rect 379222 241023 379274 241029
rect 379030 239009 379082 239015
rect 379030 238951 379082 238957
rect 378836 238382 378892 238391
rect 378836 238317 378892 238326
rect 379234 233484 379262 241023
rect 379426 234839 379454 246480
rect 379606 240785 379658 240791
rect 379606 240727 379658 240733
rect 379412 234830 379468 234839
rect 379412 234765 379468 234774
rect 379618 233484 379646 240727
rect 380098 239607 380126 246494
rect 380182 245299 380234 245305
rect 380182 245241 380234 245247
rect 380194 245083 380222 245241
rect 380182 245077 380234 245083
rect 380182 245019 380234 245025
rect 380578 239829 380606 246494
rect 380566 239823 380618 239829
rect 380566 239765 380618 239771
rect 380086 239601 380138 239607
rect 380086 239543 380138 239549
rect 380854 239527 380906 239533
rect 380854 239469 380906 239475
rect 380086 239453 380138 239459
rect 380086 239395 380138 239401
rect 379990 237307 380042 237313
rect 379990 237249 380042 237255
rect 380002 233484 380030 237249
rect 379008 233456 379262 233484
rect 379392 233456 379646 233484
rect 379776 233456 380030 233484
rect 380098 233470 380126 239395
rect 380470 239009 380522 239015
rect 380470 238951 380522 238957
rect 380180 236865 380236 236874
rect 380180 236800 380236 236809
rect 380194 236721 380222 236800
rect 380182 236715 380234 236721
rect 380182 236657 380234 236663
rect 380482 233470 380510 238951
rect 380866 233470 380894 239469
rect 380962 237905 380990 246494
rect 381154 246480 381408 246508
rect 381888 246480 382142 246508
rect 380950 237899 381002 237905
rect 380950 237841 381002 237847
rect 381154 236869 381182 246480
rect 381814 240045 381866 240051
rect 381814 239987 381866 239993
rect 381430 238787 381482 238793
rect 381430 238729 381482 238735
rect 381142 236863 381194 236869
rect 381142 236805 381194 236811
rect 381442 233484 381470 238729
rect 381826 233484 381854 239987
rect 381910 235975 381962 235981
rect 381910 235917 381962 235923
rect 381216 233456 381470 233484
rect 381600 233456 381854 233484
rect 381922 233336 381950 235917
rect 382114 233484 382142 246480
rect 382306 237239 382334 246494
rect 382690 239755 382718 246494
rect 382870 246483 382922 246489
rect 382870 246425 382922 246431
rect 382966 246483 383018 246489
rect 382966 246425 383018 246431
rect 383074 246480 383184 246508
rect 383362 246480 383616 246508
rect 383842 246480 384096 246508
rect 382882 245749 382910 246425
rect 382978 246193 383006 246425
rect 382966 246187 383018 246193
rect 382966 246129 383018 246135
rect 382870 245743 382922 245749
rect 382870 245685 382922 245691
rect 382678 239749 382730 239755
rect 383074 239723 383102 246480
rect 382678 239691 382730 239697
rect 383060 239714 383116 239723
rect 383060 239649 383116 239658
rect 383158 239675 383210 239681
rect 383158 239617 383210 239623
rect 383170 239589 383198 239617
rect 383074 239561 383198 239589
rect 383074 239533 383102 239561
rect 383062 239527 383114 239533
rect 383362 239515 383390 246480
rect 383540 240750 383596 240759
rect 383540 240685 383596 240694
rect 383554 239755 383582 240685
rect 383842 239903 383870 246480
rect 383830 239897 383882 239903
rect 383830 239839 383882 239845
rect 383542 239749 383594 239755
rect 383542 239691 383594 239697
rect 383638 239749 383690 239755
rect 383638 239691 383690 239697
rect 383362 239487 383582 239515
rect 383062 239469 383114 239475
rect 383060 239122 383116 239131
rect 382978 239080 383060 239108
rect 382294 237233 382346 237239
rect 382294 237175 382346 237181
rect 382978 233484 383006 239080
rect 383060 239057 383116 239066
rect 383158 239009 383210 239015
rect 383158 238951 383210 238957
rect 383170 238719 383198 238951
rect 383350 238861 383402 238867
rect 383554 238849 383582 239487
rect 383402 238821 383582 238849
rect 383350 238803 383402 238809
rect 383158 238713 383210 238719
rect 383158 238655 383210 238661
rect 383062 238565 383114 238571
rect 383062 238507 383114 238513
rect 383074 238095 383102 238507
rect 383060 238086 383116 238095
rect 383060 238021 383116 238030
rect 383062 237899 383114 237905
rect 383062 237841 383114 237847
rect 382114 233456 382320 233484
rect 382704 233456 383006 233484
rect 383074 233470 383102 237841
rect 383650 233484 383678 239691
rect 383734 239601 383786 239607
rect 383734 239543 383786 239549
rect 383746 233780 383774 239543
rect 384418 237905 384446 246494
rect 384610 246480 384912 246508
rect 384406 237899 384458 237905
rect 384406 237841 384458 237847
rect 384502 237899 384554 237905
rect 384502 237841 384554 237847
rect 384406 237751 384458 237757
rect 384406 237693 384458 237699
rect 383746 233752 383822 233780
rect 383424 233456 383678 233484
rect 383794 233470 383822 233752
rect 384418 233484 384446 237693
rect 384192 233456 384446 233484
rect 384514 233470 384542 237841
rect 384610 237535 384638 246480
rect 384886 239823 384938 239829
rect 384886 239765 384938 239771
rect 384598 237529 384650 237535
rect 384598 237471 384650 237477
rect 384898 233470 384926 239765
rect 385270 238343 385322 238349
rect 385270 238285 385322 238291
rect 385282 233470 385310 238285
rect 385378 237313 385406 246494
rect 385570 246480 385824 246508
rect 385954 246480 386208 246508
rect 385570 239755 385598 246480
rect 385558 239749 385610 239755
rect 385558 239691 385610 239697
rect 385954 238497 385982 246480
rect 386626 239533 386654 246494
rect 386614 239527 386666 239533
rect 386614 239469 386666 239475
rect 385942 238491 385994 238497
rect 385942 238433 385994 238439
rect 385366 237307 385418 237313
rect 385366 237249 385418 237255
rect 387106 236277 387134 246494
rect 387586 238719 387614 246494
rect 387682 246480 387936 246508
rect 388162 246480 388416 246508
rect 387574 238713 387626 238719
rect 387574 238655 387626 238661
rect 387682 237387 387710 246480
rect 388162 239681 388190 246480
rect 388150 239675 388202 239681
rect 388150 239617 388202 239623
rect 388834 238423 388862 246494
rect 388918 246335 388970 246341
rect 388918 246277 388970 246283
rect 388930 245823 388958 246277
rect 388918 245817 388970 245823
rect 388918 245759 388970 245765
rect 389026 245675 389054 246753
rect 389014 245669 389066 245675
rect 389014 245611 389066 245617
rect 388916 243414 388972 243423
rect 388916 243349 388972 243358
rect 388930 243127 388958 243349
rect 388916 243118 388972 243127
rect 388916 243053 388972 243062
rect 389218 238793 389246 246494
rect 389314 244787 389342 246753
rect 389398 246483 389450 246489
rect 389398 246425 389450 246431
rect 389410 245897 389438 246425
rect 389398 245891 389450 245897
rect 389398 245833 389450 245839
rect 389302 244781 389354 244787
rect 389302 244723 389354 244729
rect 389206 238787 389258 238793
rect 389206 238729 389258 238735
rect 388822 238417 388874 238423
rect 388822 238359 388874 238365
rect 389698 238201 389726 246494
rect 389890 246480 390144 246508
rect 389890 240051 389918 246480
rect 390274 245527 390302 246753
rect 397270 246721 397322 246727
rect 397750 246779 397802 246785
rect 397750 246721 397802 246727
rect 398230 246779 398282 246785
rect 398230 246721 398282 246727
rect 403030 246779 403082 246785
rect 405908 246753 405964 246762
rect 406100 246818 406156 246827
rect 406100 246753 406102 246762
rect 403030 246721 403082 246727
rect 390370 246480 390624 246508
rect 390262 245521 390314 245527
rect 390262 245463 390314 245469
rect 389878 240045 389930 240051
rect 389878 239987 389930 239993
rect 390370 238645 390398 246480
rect 390358 238639 390410 238645
rect 390358 238581 390410 238587
rect 389686 238195 389738 238201
rect 389686 238137 389738 238143
rect 387670 237381 387722 237387
rect 387670 237323 387722 237329
rect 390164 236754 390220 236763
rect 390164 236689 390166 236698
rect 390218 236689 390220 236698
rect 390166 236657 390218 236663
rect 387094 236271 387146 236277
rect 387094 236213 387146 236219
rect 390946 235981 390974 246494
rect 391222 246261 391274 246267
rect 391222 246203 391274 246209
rect 391234 246045 391262 246203
rect 391222 246039 391274 246045
rect 391222 245981 391274 245987
rect 391426 238571 391454 246494
rect 391414 238565 391466 238571
rect 391414 238507 391466 238513
rect 391906 238127 391934 246494
rect 392098 246480 392352 246508
rect 392482 246480 392736 246508
rect 392098 239311 392126 246480
rect 392086 239305 392138 239311
rect 392086 239247 392138 239253
rect 391894 238121 391946 238127
rect 391894 238063 391946 238069
rect 392482 237979 392510 246480
rect 392470 237973 392522 237979
rect 393154 237947 393182 246494
rect 393634 238275 393662 246494
rect 394114 241679 394142 246494
rect 394210 246480 394464 246508
rect 394690 246480 394944 246508
rect 394102 241673 394154 241679
rect 394102 241615 394154 241621
rect 393622 238269 393674 238275
rect 393622 238211 393674 238217
rect 394210 238053 394238 246480
rect 394198 238047 394250 238053
rect 394198 237989 394250 237995
rect 392470 237915 392522 237921
rect 393140 237938 393196 237947
rect 393140 237873 393196 237882
rect 394690 237799 394718 246480
rect 394676 237790 394732 237799
rect 394676 237725 394732 237734
rect 395362 237461 395390 246494
rect 395842 239385 395870 246494
rect 395830 239379 395882 239385
rect 395830 239321 395882 239327
rect 395350 237455 395402 237461
rect 395350 237397 395402 237403
rect 396226 237165 396254 246494
rect 396418 246480 396672 246508
rect 396898 246480 397152 246508
rect 396418 241827 396446 246480
rect 396406 241821 396458 241827
rect 396406 241763 396458 241769
rect 396898 239089 396926 246480
rect 397282 246267 397310 246721
rect 397366 246705 397418 246711
rect 397366 246647 397418 246653
rect 397270 246261 397322 246267
rect 397270 246203 397322 246209
rect 397378 246193 397406 246647
rect 397654 246557 397706 246563
rect 397654 246499 397706 246505
rect 397366 246187 397418 246193
rect 397366 246129 397418 246135
rect 397474 241309 397502 246494
rect 397666 246323 397694 246499
rect 397762 246489 397790 246721
rect 397750 246483 397802 246489
rect 397750 246425 397802 246431
rect 397846 246335 397898 246341
rect 397666 246295 397846 246323
rect 397846 246277 397898 246283
rect 397462 241303 397514 241309
rect 397462 241245 397514 241251
rect 396886 239083 396938 239089
rect 396886 239025 396938 239031
rect 397954 237683 397982 246494
rect 398242 245971 398270 246721
rect 398230 245965 398282 245971
rect 398230 245907 398282 245913
rect 398434 241457 398462 246494
rect 398626 246480 398880 246508
rect 399010 246480 399264 246508
rect 398422 241451 398474 241457
rect 398422 241393 398474 241399
rect 398626 240759 398654 246480
rect 398710 245151 398762 245157
rect 398710 245093 398762 245099
rect 398722 243571 398750 245093
rect 398708 243562 398764 243571
rect 398708 243497 398764 243506
rect 399010 241235 399038 246480
rect 398998 241229 399050 241235
rect 398998 241171 399050 241177
rect 398612 240750 398668 240759
rect 398612 240685 398668 240694
rect 397942 237677 397994 237683
rect 397942 237619 397994 237625
rect 399682 237609 399710 246494
rect 400162 241753 400190 246494
rect 400150 241747 400202 241753
rect 400150 241689 400202 241695
rect 400642 239163 400670 246494
rect 400738 246480 400992 246508
rect 401218 246480 401472 246508
rect 400738 241531 400766 246480
rect 400726 241525 400778 241531
rect 400726 241467 400778 241473
rect 400630 239157 400682 239163
rect 400630 239099 400682 239105
rect 401218 237831 401246 246480
rect 401890 241383 401918 246494
rect 401878 241377 401930 241383
rect 401878 241319 401930 241325
rect 402370 239237 402398 246494
rect 402754 241161 402782 246494
rect 403042 245601 403070 246721
rect 403200 246480 403262 246508
rect 403030 245595 403082 245601
rect 403030 245537 403082 245543
rect 403234 241901 403262 246480
rect 403426 246480 403680 246508
rect 403222 241895 403274 241901
rect 403222 241837 403274 241843
rect 402742 241155 402794 241161
rect 402742 241097 402794 241103
rect 403426 240717 403454 246480
rect 403414 240711 403466 240717
rect 403414 240653 403466 240659
rect 404098 240199 404126 246494
rect 404482 240939 404510 246494
rect 404470 240933 404522 240939
rect 404470 240875 404522 240881
rect 404086 240193 404138 240199
rect 404086 240135 404138 240141
rect 404962 240125 404990 246494
rect 405154 246480 405408 246508
rect 405538 246480 405792 246508
rect 405154 240643 405182 246480
rect 405142 240637 405194 240643
rect 405142 240579 405194 240585
rect 405538 240273 405566 246480
rect 405922 245527 405950 246753
rect 406154 246753 406156 246762
rect 406388 246818 406444 246827
rect 406772 246818 406828 246827
rect 406388 246753 406444 246762
rect 406580 246781 406636 246790
rect 406102 246721 406154 246727
rect 406402 246563 406430 246753
rect 406772 246753 406828 246762
rect 406964 246818 407020 246827
rect 406964 246753 406966 246762
rect 406580 246716 406636 246725
rect 406594 246637 406622 246716
rect 406582 246631 406634 246637
rect 406582 246573 406634 246579
rect 406390 246557 406442 246563
rect 406114 246480 406272 246508
rect 406390 246499 406442 246505
rect 406006 245817 406058 245823
rect 406006 245759 406058 245765
rect 405910 245521 405962 245527
rect 405910 245463 405962 245469
rect 406018 243571 406046 245759
rect 406004 243562 406060 243571
rect 406004 243497 406060 243506
rect 406114 240569 406142 246480
rect 406102 240563 406154 240569
rect 406102 240505 406154 240511
rect 406690 240347 406718 246494
rect 406786 245675 406814 246753
rect 407018 246753 407020 246762
rect 407348 246818 407404 246827
rect 407348 246753 407404 246762
rect 407732 246818 407788 246827
rect 407732 246753 407788 246762
rect 408116 246818 408172 246827
rect 408308 246818 408364 246827
rect 408172 246776 408254 246804
rect 408116 246753 408172 246762
rect 406966 246721 407018 246727
rect 406774 245669 406826 245675
rect 406774 245611 406826 245617
rect 407170 241013 407198 246494
rect 407362 246341 407390 246753
rect 407350 246335 407402 246341
rect 407350 246277 407402 246283
rect 407158 241007 407210 241013
rect 407158 240949 407210 240955
rect 406678 240341 406730 240347
rect 406678 240283 406730 240289
rect 405526 240267 405578 240273
rect 405526 240209 405578 240215
rect 404950 240119 405002 240125
rect 404950 240061 405002 240067
rect 407554 239977 407582 246494
rect 407746 246415 407774 246753
rect 407842 246480 408000 246508
rect 407734 246409 407786 246415
rect 407734 246351 407786 246357
rect 407842 240495 407870 246480
rect 408118 246409 408170 246415
rect 408118 246351 408170 246357
rect 408130 245971 408158 246351
rect 408118 245965 408170 245971
rect 408118 245907 408170 245913
rect 408226 245749 408254 246776
rect 408308 246753 408364 246762
rect 408980 246818 409036 246827
rect 408980 246753 408982 246762
rect 408322 246711 408350 246753
rect 409034 246753 409036 246762
rect 410324 246818 410380 246827
rect 410324 246753 410380 246762
rect 410516 246818 410572 246827
rect 410516 246753 410572 246762
rect 410804 246818 410860 246827
rect 410804 246753 410860 246762
rect 411188 246818 411244 246827
rect 411188 246753 411244 246762
rect 411380 246818 411436 246827
rect 411380 246753 411436 246762
rect 411764 246818 411820 246827
rect 411764 246753 411820 246762
rect 408982 246721 409034 246727
rect 408310 246705 408362 246711
rect 408310 246647 408362 246653
rect 408322 246480 408480 246508
rect 408214 245743 408266 245749
rect 408214 245685 408266 245691
rect 407830 240489 407882 240495
rect 407830 240431 407882 240437
rect 408322 240421 408350 246480
rect 408898 240865 408926 246494
rect 409282 241087 409310 246494
rect 409270 241081 409322 241087
rect 409270 241023 409322 241029
rect 408886 240859 408938 240865
rect 408886 240801 408938 240807
rect 409762 240463 409790 246494
rect 409954 246480 410208 246508
rect 409954 240791 409982 246480
rect 410338 245601 410366 246753
rect 410530 246415 410558 246753
rect 410626 246480 410688 246508
rect 410518 246409 410570 246415
rect 410518 246351 410570 246357
rect 410326 245595 410378 245601
rect 410326 245537 410378 245543
rect 409942 240785 409994 240791
rect 409942 240727 409994 240733
rect 409748 240454 409804 240463
rect 408310 240415 408362 240421
rect 409748 240389 409804 240398
rect 408310 240357 408362 240363
rect 407542 239971 407594 239977
rect 407542 239913 407594 239919
rect 402358 239231 402410 239237
rect 402358 239173 402410 239179
rect 401206 237825 401258 237831
rect 401206 237767 401258 237773
rect 410626 237757 410654 246480
rect 410818 246341 410846 246753
rect 410806 246335 410858 246341
rect 410806 246277 410858 246283
rect 411010 237905 411038 246494
rect 411202 246267 411230 246753
rect 411190 246261 411242 246267
rect 411190 246203 411242 246209
rect 411394 245897 411422 246753
rect 411382 245891 411434 245897
rect 411382 245833 411434 245839
rect 411490 245231 411518 246494
rect 411778 246193 411806 246753
rect 411766 246187 411818 246193
rect 411766 246129 411818 246135
rect 411478 245225 411530 245231
rect 411478 245167 411530 245173
rect 410998 237899 411050 237905
rect 410998 237841 411050 237847
rect 410614 237751 410666 237757
rect 410614 237693 410666 237699
rect 411970 237651 411998 246494
rect 412162 245527 412190 247197
rect 412150 245521 412202 245527
rect 412150 245463 412202 245469
rect 412258 241975 412286 272769
rect 413206 271347 413258 271353
rect 413206 271289 413258 271295
rect 413218 270909 413246 271289
rect 413206 270903 413258 270909
rect 413206 270845 413258 270851
rect 413398 267943 413450 267949
rect 413398 267885 413450 267891
rect 413302 267869 413354 267875
rect 413108 267834 413164 267843
rect 413108 267769 413164 267778
rect 413300 267834 413302 267843
rect 413354 267834 413356 267843
rect 413300 267769 413356 267778
rect 412918 266833 412970 266839
rect 412918 266775 412970 266781
rect 412822 265501 412874 265507
rect 412820 265466 412822 265475
rect 412874 265466 412876 265475
rect 412820 265401 412876 265410
rect 412930 265327 412958 266775
rect 413122 265623 413150 267769
rect 413302 266759 413354 266765
rect 413302 266701 413354 266707
rect 413108 265614 413164 265623
rect 413108 265549 413164 265558
rect 412916 265318 412972 265327
rect 412916 265253 412972 265262
rect 412724 265170 412780 265179
rect 412724 265105 412780 265114
rect 412738 265063 412766 265105
rect 412726 265057 412778 265063
rect 412628 265022 412684 265031
rect 412726 264999 412778 265005
rect 412628 264957 412630 264966
rect 412682 264957 412684 264966
rect 412630 264925 412682 264931
rect 413314 264883 413342 266701
rect 413410 265919 413438 267885
rect 414370 267727 414398 277870
rect 416674 269059 416702 277870
rect 417922 277569 417950 277870
rect 417910 277563 417962 277569
rect 417910 277505 417962 277511
rect 417334 273789 417386 273795
rect 417334 273731 417386 273737
rect 417346 273652 417374 273731
rect 417332 273643 417388 273652
rect 417332 273578 417388 273587
rect 416662 269053 416714 269059
rect 416662 268995 416714 269001
rect 414358 267721 414410 267727
rect 414358 267663 414410 267669
rect 419074 267579 419102 277870
rect 420226 274831 420254 277870
rect 420214 274825 420266 274831
rect 420214 274767 420266 274773
rect 419062 267573 419114 267579
rect 419062 267515 419114 267521
rect 421474 267505 421502 277870
rect 423874 269133 423902 277870
rect 425026 277347 425054 277870
rect 425014 277341 425066 277347
rect 425014 277283 425066 277289
rect 423862 269127 423914 269133
rect 423862 269069 423914 269075
rect 426274 268245 426302 277870
rect 427426 274979 427454 277870
rect 427414 274973 427466 274979
rect 427414 274915 427466 274921
rect 426262 268239 426314 268245
rect 426262 268181 426314 268187
rect 421462 267499 421514 267505
rect 421462 267441 421514 267447
rect 419350 267203 419402 267209
rect 419350 267145 419402 267151
rect 413396 265910 413452 265919
rect 413396 265845 413452 265854
rect 419362 265729 419390 267145
rect 428674 266691 428702 277870
rect 429826 273721 429854 277870
rect 429814 273715 429866 273721
rect 429814 273657 429866 273663
rect 429140 270794 429196 270803
rect 429140 270729 429196 270738
rect 429154 270336 429182 270729
rect 429058 270308 429182 270336
rect 428948 270054 429004 270063
rect 428948 269989 429004 269998
rect 428962 269059 428990 269989
rect 429058 269915 429086 270308
rect 429236 270054 429292 270063
rect 429236 269989 429292 269998
rect 429044 269906 429100 269915
rect 429044 269841 429100 269850
rect 429250 269059 429278 269989
rect 431074 269207 431102 277870
rect 432226 277273 432254 277870
rect 432214 277267 432266 277273
rect 432214 277209 432266 277215
rect 431062 269201 431114 269207
rect 431062 269143 431114 269149
rect 428950 269053 429002 269059
rect 428950 268995 429002 269001
rect 429238 269053 429290 269059
rect 429238 268995 429290 269001
rect 433378 267431 433406 277870
rect 434530 276385 434558 277870
rect 434518 276379 434570 276385
rect 434518 276321 434570 276327
rect 433462 271939 433514 271945
rect 433462 271881 433514 271887
rect 433474 271279 433502 271881
rect 433462 271273 433514 271279
rect 433462 271215 433514 271221
rect 433366 267425 433418 267431
rect 433366 267367 433418 267373
rect 428662 266685 428714 266691
rect 428662 266627 428714 266633
rect 435682 266469 435710 277870
rect 436642 277856 436944 277875
rect 438082 270465 438110 277870
rect 439330 277125 439358 277870
rect 439318 277119 439370 277125
rect 439318 277061 439370 277067
rect 438070 270459 438122 270465
rect 438070 270401 438122 270407
rect 440482 268023 440510 277870
rect 441730 276163 441758 277870
rect 441718 276157 441770 276163
rect 441718 276099 441770 276105
rect 440756 273902 440812 273911
rect 440578 273860 440756 273888
rect 440578 273763 440606 273860
rect 440756 273837 440812 273846
rect 440564 273754 440620 273763
rect 440564 273689 440620 273698
rect 440660 270498 440716 270507
rect 440660 270433 440662 270442
rect 440714 270433 440716 270442
rect 440662 270401 440714 270407
rect 440470 268017 440522 268023
rect 440470 267959 440522 267965
rect 435670 266463 435722 266469
rect 435670 266405 435722 266411
rect 442882 266395 442910 277870
rect 444130 273869 444158 277870
rect 444118 273863 444170 273869
rect 444118 273805 444170 273811
rect 445282 270317 445310 277870
rect 446530 276977 446558 277870
rect 446518 276971 446570 276977
rect 446518 276913 446570 276919
rect 445270 270311 445322 270317
rect 445270 270253 445322 270259
rect 447682 267283 447710 277870
rect 448834 276089 448862 277870
rect 448822 276083 448874 276089
rect 448822 276025 448874 276031
rect 449302 274381 449354 274387
rect 449302 274323 449354 274329
rect 449314 274239 449342 274323
rect 449302 274233 449354 274239
rect 449302 274175 449354 274181
rect 449204 270794 449260 270803
rect 449204 270729 449260 270738
rect 449218 269915 449246 270729
rect 449204 269906 449260 269915
rect 449204 269841 449260 269850
rect 447670 267277 447722 267283
rect 447670 267219 447722 267225
rect 442870 266389 442922 266395
rect 442870 266331 442922 266337
rect 449986 266321 450014 277870
rect 450850 277865 451152 277884
rect 450838 277859 451152 277865
rect 450890 277856 451152 277859
rect 450838 277801 450890 277807
rect 452386 270169 452414 277870
rect 453538 276829 453566 277870
rect 453526 276823 453578 276829
rect 453526 276765 453578 276771
rect 452374 270163 452426 270169
rect 452374 270105 452426 270111
rect 454786 268097 454814 277870
rect 455938 276015 455966 277870
rect 455926 276009 455978 276015
rect 455926 275951 455978 275957
rect 454774 268091 454826 268097
rect 454774 268033 454826 268039
rect 449974 266315 450026 266321
rect 449974 266257 450026 266263
rect 457186 266173 457214 277870
rect 457954 273971 458078 273999
rect 457954 273911 457982 273971
rect 457940 273902 457996 273911
rect 457940 273837 457996 273846
rect 458050 273467 458078 273971
rect 458036 273458 458092 273467
rect 458036 273393 458092 273402
rect 458338 267135 458366 277870
rect 459286 271569 459338 271575
rect 459286 271511 459338 271517
rect 459298 271279 459326 271511
rect 459286 271273 459338 271279
rect 459286 271215 459338 271221
rect 459586 269947 459614 277870
rect 460738 277199 460766 277870
rect 460726 277193 460778 277199
rect 460726 277135 460778 277141
rect 461986 274017 462014 277870
rect 463138 275867 463166 277870
rect 463126 275861 463178 275867
rect 463126 275803 463178 275809
rect 461974 274011 462026 274017
rect 461974 273953 462026 273959
rect 460724 270498 460780 270507
rect 460724 270433 460726 270442
rect 460778 270433 460780 270442
rect 460726 270401 460778 270407
rect 459574 269941 459626 269947
rect 459574 269883 459626 269889
rect 458326 267129 458378 267135
rect 458326 267071 458378 267077
rect 457174 266167 457226 266173
rect 457174 266109 457226 266115
rect 464290 266099 464318 277870
rect 465250 277856 465552 277884
rect 465250 277791 465278 277856
rect 465238 277785 465290 277791
rect 465238 277727 465290 277733
rect 466594 269725 466622 277870
rect 466582 269719 466634 269725
rect 466582 269661 466634 269667
rect 468994 268171 469022 277870
rect 470242 275719 470270 277870
rect 470230 275713 470282 275719
rect 470230 275655 470282 275661
rect 469462 274233 469514 274239
rect 469462 274175 469514 274181
rect 469474 274017 469502 274175
rect 469462 274011 469514 274017
rect 469462 273953 469514 273959
rect 469174 270459 469226 270465
rect 469174 270401 469226 270407
rect 469654 270459 469706 270465
rect 469654 270401 469706 270407
rect 469076 270350 469132 270359
rect 469076 270285 469078 270294
rect 469130 270285 469132 270294
rect 469078 270253 469130 270259
rect 469186 270063 469214 270401
rect 469556 270350 469612 270359
rect 469378 270308 469502 270336
rect 469378 270299 469406 270308
rect 469282 270271 469406 270299
rect 469172 270054 469228 270063
rect 469172 269989 469228 269998
rect 469282 269915 469310 270271
rect 469364 270202 469420 270211
rect 469364 270137 469366 270146
rect 469418 270137 469420 270146
rect 469366 270105 469418 270111
rect 469474 269947 469502 270308
rect 469556 270285 469558 270294
rect 469610 270285 469612 270294
rect 469558 270253 469610 270259
rect 469556 270202 469612 270211
rect 469556 270137 469558 270146
rect 469610 270137 469612 270146
rect 469558 270105 469610 270111
rect 469666 270063 469694 270401
rect 469652 270054 469708 270063
rect 469652 269989 469708 269998
rect 469462 269941 469514 269947
rect 469268 269906 469324 269915
rect 469462 269883 469514 269889
rect 469268 269841 469324 269850
rect 468982 268165 469034 268171
rect 468982 268107 469034 268113
rect 464278 266093 464330 266099
rect 464278 266035 464330 266041
rect 471394 266025 471422 277870
rect 472642 266913 472670 277870
rect 473794 269651 473822 277870
rect 476194 274091 476222 277870
rect 477442 275571 477470 277870
rect 477430 275565 477482 275571
rect 477430 275507 477482 275513
rect 476182 274085 476234 274091
rect 476182 274027 476234 274033
rect 473782 269645 473834 269651
rect 473782 269587 473834 269593
rect 472630 266907 472682 266913
rect 472630 266849 472682 266855
rect 471382 266019 471434 266025
rect 471382 265961 471434 265967
rect 478594 265877 478622 277870
rect 479746 274165 479774 277870
rect 479734 274159 479786 274165
rect 479734 274101 479786 274107
rect 479446 271569 479498 271575
rect 479446 271511 479498 271517
rect 479458 271279 479486 271511
rect 479446 271273 479498 271279
rect 479446 271215 479498 271221
rect 480994 269429 481022 277870
rect 480982 269423 481034 269429
rect 480982 269365 481034 269371
rect 483298 268319 483326 277870
rect 484450 274059 484478 277870
rect 484436 274050 484492 274059
rect 484436 273985 484492 273994
rect 483286 268313 483338 268319
rect 483286 268255 483338 268261
rect 478582 265871 478634 265877
rect 478582 265813 478634 265819
rect 485698 265803 485726 277870
rect 486850 277421 486878 277870
rect 486838 277415 486890 277421
rect 486838 277357 486890 277363
rect 488098 268139 488126 277870
rect 489004 277856 489264 277884
rect 488948 277833 489004 277842
rect 491650 274207 491678 277870
rect 491636 274198 491692 274207
rect 491636 274133 491692 274142
rect 489620 273754 489676 273763
rect 489620 273689 489676 273698
rect 489634 273467 489662 273689
rect 489620 273458 489676 273467
rect 489620 273393 489676 273402
rect 488278 269941 488330 269947
rect 488278 269883 488330 269889
rect 488290 268139 488318 269883
rect 488084 268130 488140 268139
rect 488084 268065 488140 268074
rect 488276 268130 488332 268139
rect 488276 268065 488332 268074
rect 485686 265797 485738 265803
rect 485686 265739 485738 265745
rect 419254 265723 419306 265729
rect 419254 265665 419306 265671
rect 419350 265723 419402 265729
rect 419350 265665 419402 265671
rect 419062 265427 419114 265433
rect 419062 265369 419114 265375
rect 419074 265285 419102 265369
rect 419062 265279 419114 265285
rect 419062 265221 419114 265227
rect 419158 265279 419210 265285
rect 419158 265221 419210 265227
rect 419170 265137 419198 265221
rect 419266 265137 419294 265665
rect 492898 265655 492926 277870
rect 494050 266617 494078 277870
rect 495202 269281 495230 277870
rect 496162 277856 496464 277884
rect 496162 277759 496190 277856
rect 496148 277750 496204 277759
rect 496148 277685 496204 277694
rect 495190 269275 495242 269281
rect 495190 269217 495242 269223
rect 494038 266611 494090 266617
rect 494038 266553 494090 266559
rect 497602 266543 497630 277870
rect 498850 274355 498878 277870
rect 498836 274346 498892 274355
rect 498836 274281 498892 274290
rect 499606 271569 499658 271575
rect 499606 271511 499658 271517
rect 499618 271279 499646 271511
rect 499606 271273 499658 271279
rect 499606 271215 499658 271221
rect 499508 270350 499564 270359
rect 499508 270285 499564 270294
rect 499414 268461 499466 268467
rect 499412 268426 499414 268435
rect 499466 268426 499468 268435
rect 499412 268361 499468 268370
rect 499318 268239 499370 268245
rect 499318 268181 499370 268187
rect 499330 268139 499358 268181
rect 499522 268139 499550 270285
rect 499700 270202 499756 270211
rect 499700 270137 499756 270146
rect 499604 270054 499660 270063
rect 499604 269989 499660 269998
rect 499618 268731 499646 269989
rect 499604 268722 499660 268731
rect 499604 268657 499660 268666
rect 499714 268435 499742 270137
rect 499796 270054 499852 270063
rect 499796 269989 499852 269998
rect 499700 268426 499756 268435
rect 499700 268361 499756 268370
rect 499810 268245 499838 269989
rect 499798 268239 499850 268245
rect 499798 268181 499850 268187
rect 499316 268130 499372 268139
rect 499316 268065 499372 268074
rect 499508 268130 499564 268139
rect 499508 268065 499564 268074
rect 497590 266537 497642 266543
rect 497590 266479 497642 266485
rect 492886 265649 492938 265655
rect 492886 265591 492938 265597
rect 499906 265581 499934 277870
rect 501154 268393 501182 277870
rect 502018 277856 502320 277884
rect 502018 268467 502046 277856
rect 503554 270539 503582 277870
rect 504706 277051 504734 277870
rect 504694 277045 504746 277051
rect 504694 276987 504746 276993
rect 505954 274503 505982 277870
rect 507106 277611 507134 277870
rect 507092 277602 507148 277611
rect 507092 277537 507148 277546
rect 505940 274494 505996 274503
rect 505940 274429 505996 274438
rect 508354 274017 508382 277870
rect 508342 274011 508394 274017
rect 508342 273953 508394 273959
rect 504020 273902 504076 273911
rect 504020 273837 504076 273846
rect 503924 273754 503980 273763
rect 504034 273740 504062 273837
rect 503980 273712 504062 273740
rect 503924 273689 503980 273698
rect 503542 270533 503594 270539
rect 503542 270475 503594 270481
rect 509506 270359 509534 277870
rect 510658 271057 510686 277870
rect 511906 274313 511934 277870
rect 511894 274307 511946 274313
rect 511894 274249 511946 274255
rect 510646 271051 510698 271057
rect 510646 270993 510698 270999
rect 509492 270350 509548 270359
rect 509492 270285 509548 270294
rect 513058 269175 513086 277870
rect 513044 269166 513100 269175
rect 513044 269101 513100 269110
rect 502006 268461 502058 268467
rect 502006 268403 502058 268409
rect 501142 268387 501194 268393
rect 501142 268329 501194 268335
rect 499894 265575 499946 265581
rect 499894 265517 499946 265523
rect 514306 265507 514334 277870
rect 515458 276903 515486 277870
rect 515446 276897 515498 276903
rect 515446 276839 515498 276845
rect 516610 274651 516638 277870
rect 517762 277463 517790 277870
rect 517748 277454 517804 277463
rect 517748 277389 517804 277398
rect 519010 276755 519038 277870
rect 518998 276749 519050 276755
rect 518998 276691 519050 276697
rect 520162 274799 520190 277870
rect 520148 274790 520204 274799
rect 520148 274725 520204 274734
rect 516596 274642 516652 274651
rect 516596 274577 516652 274586
rect 518326 271569 518378 271575
rect 518326 271511 518378 271517
rect 518338 271279 518366 271511
rect 518326 271273 518378 271279
rect 518326 271215 518378 271221
rect 519476 270350 519532 270359
rect 519476 270285 519532 270294
rect 519668 270350 519724 270359
rect 519668 270285 519724 270294
rect 519490 269175 519518 270285
rect 519476 269166 519532 269175
rect 519476 269101 519532 269110
rect 519682 268139 519710 270285
rect 519860 270202 519916 270211
rect 519860 270137 519916 270146
rect 519764 270054 519820 270063
rect 519764 269989 519820 269998
rect 519778 268731 519806 269989
rect 519764 268722 519820 268731
rect 519764 268657 519820 268666
rect 519874 268435 519902 270137
rect 519860 268426 519916 268435
rect 519860 268361 519916 268370
rect 519668 268130 519724 268139
rect 519668 268065 519724 268074
rect 514294 265501 514346 265507
rect 514294 265443 514346 265449
rect 521410 265433 521438 277870
rect 521590 266389 521642 266395
rect 521590 266331 521642 266337
rect 521398 265427 521450 265433
rect 521398 265369 521450 265375
rect 419158 265131 419210 265137
rect 419158 265073 419210 265079
rect 419254 265131 419306 265137
rect 419254 265073 419306 265079
rect 413300 264874 413356 264883
rect 413300 264809 413356 264818
rect 412340 246818 412396 246827
rect 412340 246753 412396 246762
rect 412354 246045 412382 246753
rect 505846 246113 505898 246119
rect 505846 246055 505898 246061
rect 412342 246039 412394 246045
rect 412342 245981 412394 245987
rect 443540 243710 443596 243719
rect 443540 243645 443542 243654
rect 443594 243645 443596 243654
rect 463604 243710 463660 243719
rect 463604 243645 463606 243654
rect 443542 243613 443594 243619
rect 463658 243645 463660 243654
rect 483860 243710 483916 243719
rect 483860 243645 483862 243654
rect 463606 243613 463658 243619
rect 483914 243645 483916 243654
rect 503924 243710 503980 243719
rect 503924 243645 503926 243654
rect 483862 243613 483914 243619
rect 503978 243645 503980 243654
rect 503926 243613 503978 243619
rect 443542 242561 443594 242567
rect 443540 242526 443542 242535
rect 463606 242561 463658 242567
rect 443594 242526 443596 242535
rect 443540 242461 443596 242470
rect 463604 242526 463606 242535
rect 483862 242561 483914 242567
rect 463658 242526 463660 242535
rect 463604 242461 463660 242470
rect 483860 242526 483862 242535
rect 503926 242561 503978 242567
rect 483914 242526 483916 242535
rect 483860 242461 483916 242470
rect 503924 242526 503926 242535
rect 503978 242526 503980 242535
rect 503924 242461 503980 242470
rect 412054 241969 412106 241975
rect 412054 241911 412106 241917
rect 412246 241969 412298 241975
rect 412246 241911 412298 241917
rect 412066 238835 412094 241911
rect 412052 238826 412108 238835
rect 412052 238761 412108 238770
rect 497494 237677 497546 237683
rect 411956 237642 412012 237651
rect 399670 237603 399722 237609
rect 505858 237651 505886 246055
rect 511124 242526 511180 242535
rect 511124 242461 511180 242470
rect 511138 237799 511166 242461
rect 521602 241943 521630 266331
rect 522562 266247 522590 277870
rect 523522 277856 523824 277884
rect 523522 266395 523550 277856
rect 524962 269873 524990 277870
rect 524950 269867 525002 269873
rect 524950 269809 525002 269815
rect 526114 268689 526142 277870
rect 526102 268683 526154 268689
rect 526102 268625 526154 268631
rect 523510 266389 523562 266395
rect 523510 266331 523562 266337
rect 522550 266241 522602 266247
rect 522550 266183 522602 266189
rect 527362 265327 527390 277870
rect 528514 277315 528542 277870
rect 528500 277306 528556 277315
rect 528500 277241 528556 277250
rect 529762 268837 529790 277870
rect 529844 273754 529900 273763
rect 529844 273689 529900 273698
rect 529858 273467 529886 273689
rect 529844 273458 529900 273467
rect 529844 273393 529900 273402
rect 529844 269906 529900 269915
rect 529844 269841 529900 269850
rect 529858 269175 529886 269841
rect 529844 269166 529900 269175
rect 529844 269101 529900 269110
rect 529750 268831 529802 268837
rect 529750 268773 529802 268779
rect 527348 265318 527404 265327
rect 527348 265253 527404 265262
rect 530914 265179 530942 277870
rect 532162 275793 532190 277870
rect 532150 275787 532202 275793
rect 532150 275729 532202 275735
rect 533218 265951 533246 277870
rect 534466 271205 534494 277870
rect 534454 271199 534506 271205
rect 534454 271141 534506 271147
rect 533206 265945 533258 265951
rect 533206 265887 533258 265893
rect 535618 265359 535646 277870
rect 536866 268985 536894 277870
rect 536854 268979 536906 268985
rect 536854 268921 536906 268927
rect 535606 265353 535658 265359
rect 535606 265295 535658 265301
rect 530900 265170 530956 265179
rect 530900 265105 530956 265114
rect 538018 265031 538046 277870
rect 539266 277167 539294 277870
rect 539252 277158 539308 277167
rect 539252 277093 539308 277102
rect 540418 274683 540446 277870
rect 540406 274677 540458 274683
rect 540406 274619 540458 274625
rect 541570 272241 541598 277870
rect 541558 272235 541610 272241
rect 541558 272177 541610 272183
rect 542818 269503 542846 277870
rect 543970 271279 543998 277870
rect 543958 271273 544010 271279
rect 543958 271215 544010 271221
rect 545218 270983 545246 277870
rect 545206 270977 545258 270983
rect 545206 270919 545258 270925
rect 544438 270533 544490 270539
rect 544436 270498 544438 270507
rect 544490 270498 544492 270507
rect 544436 270433 544492 270442
rect 542806 269497 542858 269503
rect 542806 269439 542858 269445
rect 546370 265285 546398 277870
rect 547618 265729 547646 277870
rect 548770 273763 548798 277870
rect 548756 273754 548812 273763
rect 548756 273689 548812 273698
rect 549922 270687 549950 277870
rect 551074 274905 551102 277870
rect 551062 274899 551114 274905
rect 551062 274841 551114 274847
rect 552322 272167 552350 277870
rect 552310 272161 552362 272167
rect 552310 272103 552362 272109
rect 549910 270681 549962 270687
rect 549910 270623 549962 270629
rect 553474 269355 553502 277870
rect 554722 276681 554750 277870
rect 554710 276675 554762 276681
rect 554710 276617 554762 276623
rect 553462 269349 553514 269355
rect 553462 269291 553514 269297
rect 547606 265723 547658 265729
rect 547606 265665 547658 265671
rect 546358 265279 546410 265285
rect 546358 265221 546410 265227
rect 538004 265022 538060 265031
rect 538004 264957 538060 264966
rect 555874 264883 555902 277870
rect 557026 273499 557054 277870
rect 558274 273943 558302 277870
rect 558262 273937 558314 273943
rect 558262 273879 558314 273885
rect 557014 273493 557066 273499
rect 557014 273435 557066 273441
rect 559426 271353 559454 277870
rect 559414 271347 559466 271353
rect 559414 271289 559466 271295
rect 560674 267991 560702 277870
rect 561826 270613 561854 277870
rect 563074 273319 563102 277870
rect 564226 275497 564254 277870
rect 565474 276311 565502 277870
rect 565462 276305 565514 276311
rect 565462 276247 565514 276253
rect 564214 275491 564266 275497
rect 564214 275433 564266 275439
rect 563060 273310 563116 273319
rect 563060 273245 563116 273254
rect 566530 271395 566558 277870
rect 566516 271386 566572 271395
rect 566516 271321 566572 271330
rect 561814 270607 561866 270613
rect 561814 270549 561866 270555
rect 564406 270533 564458 270539
rect 564404 270498 564406 270507
rect 564458 270498 564460 270507
rect 564404 270433 564460 270442
rect 567778 268583 567806 277870
rect 568930 270391 568958 277870
rect 570178 270761 570206 277870
rect 571330 275275 571358 277870
rect 572482 276237 572510 277870
rect 572470 276231 572522 276237
rect 572470 276173 572522 276179
rect 571318 275269 571370 275275
rect 571318 275211 571370 275217
rect 573730 272315 573758 277870
rect 573718 272309 573770 272315
rect 573718 272251 573770 272257
rect 570166 270755 570218 270761
rect 570166 270697 570218 270703
rect 568918 270385 568970 270391
rect 568918 270327 568970 270333
rect 574882 268879 574910 277870
rect 576130 270243 576158 277870
rect 576118 270237 576170 270243
rect 576118 270179 576170 270185
rect 577282 269767 577310 277870
rect 578530 275201 578558 277870
rect 579682 275941 579710 277870
rect 579670 275935 579722 275941
rect 579670 275877 579722 275883
rect 578518 275195 578570 275201
rect 578518 275137 578570 275143
rect 580930 271131 580958 277870
rect 580918 271125 580970 271131
rect 580918 271067 580970 271073
rect 582082 270359 582110 277870
rect 582068 270350 582124 270359
rect 582068 270285 582124 270294
rect 583234 270095 583262 277870
rect 584386 272463 584414 277870
rect 585634 275053 585662 277870
rect 585622 275047 585674 275053
rect 585622 274989 585674 274995
rect 584374 272457 584426 272463
rect 584374 272399 584426 272405
rect 583222 270089 583274 270095
rect 583222 270031 583274 270037
rect 586786 270021 586814 277870
rect 587938 272389 587966 277870
rect 587926 272383 587978 272389
rect 587926 272325 587978 272331
rect 589186 270211 589214 277870
rect 590338 271427 590366 277870
rect 591586 272611 591614 277870
rect 592738 276279 592766 277870
rect 592724 276270 592780 276279
rect 592724 276205 592780 276214
rect 591574 272605 591626 272611
rect 591574 272547 591626 272553
rect 593986 271501 594014 277870
rect 595138 273573 595166 277870
rect 595126 273567 595178 273573
rect 595126 273509 595178 273515
rect 596182 272827 596234 272833
rect 596182 272769 596234 272775
rect 593974 271495 594026 271501
rect 593974 271437 594026 271443
rect 590326 271421 590378 271427
rect 590326 271363 590378 271369
rect 589172 270202 589228 270211
rect 589172 270137 589228 270146
rect 586774 270015 586826 270021
rect 586774 269957 586826 269963
rect 577268 269758 577324 269767
rect 577268 269693 577324 269702
rect 574868 268870 574924 268879
rect 574868 268805 574924 268814
rect 567764 268574 567820 268583
rect 567764 268509 567820 268518
rect 560660 267982 560716 267991
rect 560660 267917 560716 267926
rect 555860 264874 555916 264883
rect 555860 264809 555916 264818
rect 524180 243710 524236 243719
rect 524180 243645 524182 243654
rect 524234 243645 524236 243654
rect 544244 243710 544300 243719
rect 544244 243645 544246 243654
rect 524182 243613 524234 243619
rect 544298 243645 544300 243654
rect 564500 243710 564556 243719
rect 564500 243645 564502 243654
rect 544246 243613 544298 243619
rect 564554 243645 564556 243654
rect 584564 243710 584620 243719
rect 584564 243645 584566 243654
rect 564502 243613 564554 243619
rect 584618 243645 584620 243654
rect 584566 243613 584618 243619
rect 521588 241934 521644 241943
rect 521588 241869 521644 241878
rect 596194 238983 596222 272769
rect 596386 270063 596414 277870
rect 596372 270054 596428 270063
rect 596372 269989 596428 269998
rect 597538 269799 597566 277870
rect 598498 277856 598800 277884
rect 598498 272833 598526 277856
rect 599842 275983 599870 277870
rect 599828 275974 599884 275983
rect 599828 275909 599884 275918
rect 601090 275645 601118 277870
rect 601078 275639 601130 275645
rect 601078 275581 601130 275587
rect 602242 275539 602270 277870
rect 602228 275530 602284 275539
rect 602228 275465 602284 275474
rect 598486 272827 598538 272833
rect 598486 272769 598538 272775
rect 603394 269915 603422 277870
rect 603380 269906 603436 269915
rect 603380 269841 603436 269850
rect 597526 269793 597578 269799
rect 597526 269735 597578 269741
rect 604642 269577 604670 277870
rect 605794 269619 605822 277870
rect 607042 276131 607070 277870
rect 607028 276122 607084 276131
rect 607028 276057 607084 276066
rect 605780 269610 605836 269619
rect 604630 269571 604682 269577
rect 605780 269545 605836 269554
rect 604630 269513 604682 269519
rect 608194 265211 608222 277870
rect 609442 265919 609470 277870
rect 610594 275835 610622 277870
rect 611842 276607 611870 277870
rect 611830 276601 611882 276607
rect 611830 276543 611882 276549
rect 610580 275826 610636 275835
rect 610580 275761 610636 275770
rect 612994 272685 613022 277870
rect 612982 272679 613034 272685
rect 612982 272621 613034 272627
rect 614242 267843 614270 277870
rect 614228 267834 614284 267843
rect 614228 267769 614284 267778
rect 609428 265910 609484 265919
rect 609428 265845 609484 265854
rect 608182 265205 608234 265211
rect 608182 265147 608234 265153
rect 615394 265137 615422 277870
rect 616546 275391 616574 277870
rect 617698 276871 617726 277870
rect 617684 276862 617740 276871
rect 617684 276797 617740 276806
rect 616532 275382 616588 275391
rect 616532 275317 616588 275326
rect 618850 272019 618878 277870
rect 618838 272013 618890 272019
rect 618838 271955 618890 271961
rect 620098 269471 620126 277870
rect 620084 269462 620140 269471
rect 620084 269397 620140 269406
rect 621250 267801 621278 277870
rect 622498 275423 622526 277870
rect 622486 275417 622538 275423
rect 622486 275359 622538 275365
rect 623650 275243 623678 277870
rect 624898 275687 624926 277870
rect 624884 275678 624940 275687
rect 624884 275613 624940 275622
rect 623636 275234 623692 275243
rect 623636 275169 623692 275178
rect 623062 270607 623114 270613
rect 623062 270549 623114 270555
rect 623074 270507 623102 270549
rect 623060 270498 623116 270507
rect 623060 270433 623116 270442
rect 626050 268287 626078 277870
rect 627298 275095 627326 277870
rect 627284 275086 627340 275095
rect 627284 275021 627340 275030
rect 626036 268278 626092 268287
rect 626036 268213 626092 268222
rect 621238 267795 621290 267801
rect 621238 267737 621290 267743
rect 628450 265623 628478 277870
rect 629698 267357 629726 277870
rect 630850 269323 630878 277870
rect 630836 269314 630892 269323
rect 630836 269249 630892 269258
rect 629686 267351 629738 267357
rect 629686 267293 629738 267299
rect 628436 265614 628492 265623
rect 628436 265549 628492 265558
rect 632098 265475 632126 277870
rect 633154 275349 633182 277870
rect 633142 275343 633194 275349
rect 633142 275285 633194 275291
rect 633622 271939 633674 271945
rect 633622 271881 633674 271887
rect 632084 265466 632140 265475
rect 632084 265401 632140 265410
rect 615382 265131 615434 265137
rect 615382 265073 615434 265079
rect 633634 262177 633662 271881
rect 634306 270655 634334 277870
rect 635554 276723 635582 277870
rect 635540 276714 635596 276723
rect 635540 276649 635596 276658
rect 637954 276427 637982 277870
rect 637940 276418 637996 276427
rect 637940 276353 637996 276362
rect 634292 270646 634348 270655
rect 634292 270581 634348 270590
rect 639106 267695 639134 277870
rect 640354 269027 640382 277870
rect 641506 270613 641534 277870
rect 642754 276575 642782 277870
rect 642740 276566 642796 276575
rect 642262 276527 642314 276533
rect 642740 276501 642796 276510
rect 642262 276469 642314 276475
rect 642274 271945 642302 276469
rect 643906 272907 643934 277870
rect 645154 274947 645182 277870
rect 647554 275127 647582 277870
rect 648034 277856 648720 277884
rect 647542 275121 647594 275127
rect 647542 275063 647594 275069
rect 645140 274938 645196 274947
rect 645140 274873 645196 274882
rect 645718 274307 645770 274313
rect 645718 274249 645770 274255
rect 643894 272901 643946 272907
rect 643894 272843 643946 272849
rect 642262 271939 642314 271945
rect 642262 271881 642314 271887
rect 641494 270607 641546 270613
rect 641494 270549 641546 270555
rect 640340 269018 640396 269027
rect 640340 268953 640396 268962
rect 639092 267686 639148 267695
rect 639092 267621 639148 267630
rect 633622 262171 633674 262177
rect 633622 262113 633674 262119
rect 625846 262097 625898 262103
rect 625846 262039 625898 262045
rect 625858 257811 625886 262039
rect 645730 260549 645758 274249
rect 642262 260543 642314 260549
rect 642262 260485 642314 260491
rect 645718 260543 645770 260549
rect 645718 260485 645770 260491
rect 616342 257805 616394 257811
rect 616342 257747 616394 257753
rect 625846 257805 625898 257811
rect 625846 257747 625898 257753
rect 616354 250633 616382 257747
rect 639286 256399 639338 256405
rect 639286 256341 639338 256347
rect 607702 250627 607754 250633
rect 607702 250569 607754 250575
rect 616342 250627 616394 250633
rect 616342 250569 616394 250575
rect 636502 250627 636554 250633
rect 636502 250569 636554 250575
rect 604822 243745 604874 243751
rect 604820 243710 604822 243719
rect 604874 243710 604876 243719
rect 604820 243645 604876 243654
rect 607714 241975 607742 250569
rect 636514 247747 636542 250569
rect 627862 247741 627914 247747
rect 627862 247683 627914 247689
rect 636502 247741 636554 247747
rect 636502 247683 636554 247689
rect 624886 243745 624938 243751
rect 624884 243710 624886 243719
rect 624938 243710 624940 243719
rect 624884 243645 624940 243654
rect 627874 242068 627902 247683
rect 627778 242040 627902 242068
rect 607702 241969 607754 241975
rect 607702 241911 607754 241917
rect 602902 241895 602954 241901
rect 602902 241837 602954 241843
rect 596180 238974 596236 238983
rect 596180 238909 596236 238918
rect 511124 237790 511180 237799
rect 511124 237725 511180 237734
rect 549238 237751 549290 237757
rect 497494 237619 497546 237625
rect 505844 237642 505900 237651
rect 411956 237577 412012 237586
rect 420598 237603 420650 237609
rect 399670 237545 399722 237551
rect 420598 237545 420650 237551
rect 396214 237159 396266 237165
rect 396214 237101 396266 237107
rect 420500 236754 420556 236763
rect 420500 236689 420502 236698
rect 420554 236689 420556 236698
rect 420502 236657 420554 236663
rect 420610 236467 420638 237545
rect 497506 236763 497534 237619
rect 505844 237577 505900 237586
rect 440564 236754 440620 236763
rect 440564 236689 440566 236698
rect 440618 236689 440620 236698
rect 460820 236754 460876 236763
rect 460820 236689 460822 236698
rect 440566 236657 440618 236663
rect 460874 236689 460876 236698
rect 480884 236754 480940 236763
rect 480884 236689 480886 236698
rect 460822 236657 460874 236663
rect 480938 236689 480940 236698
rect 497492 236754 497548 236763
rect 497492 236689 497548 236698
rect 480886 236657 480938 236663
rect 420596 236458 420652 236467
rect 420596 236393 420652 236402
rect 390934 235975 390986 235981
rect 390934 235917 390986 235923
rect 420610 233470 420638 236393
rect 497506 233470 497534 236689
rect 505858 233484 505886 237577
rect 511138 233484 511166 237725
rect 549238 237693 549290 237699
rect 549250 236203 549278 237693
rect 602914 237683 602942 241837
rect 627778 240495 627806 242040
rect 607606 240489 607658 240495
rect 607606 240431 607658 240437
rect 627766 240489 627818 240495
rect 627766 240431 627818 240437
rect 602902 237677 602954 237683
rect 602902 237619 602954 237625
rect 607618 237609 607646 240431
rect 607606 237603 607658 237609
rect 607606 237545 607658 237551
rect 638038 236567 638090 236573
rect 638038 236509 638090 236515
rect 637558 236493 637610 236499
rect 637558 236435 637610 236441
rect 547126 236197 547178 236203
rect 547126 236139 547178 236145
rect 549238 236197 549290 236203
rect 549238 236139 549290 236145
rect 547138 234691 547166 236139
rect 547124 234682 547180 234691
rect 547124 234617 547180 234626
rect 549250 233484 549278 236139
rect 637172 233646 637228 233655
rect 637172 233581 637228 233590
rect 505632 233456 505886 233484
rect 510384 233456 511166 233484
rect 549024 233456 549278 233484
rect 637186 233484 637214 233581
rect 637570 233484 637598 236435
rect 637942 236419 637994 236425
rect 637942 236361 637994 236367
rect 637954 233951 637982 236361
rect 638050 234099 638078 236509
rect 639190 236345 639242 236351
rect 638420 236310 638476 236319
rect 639298 236319 639326 256341
rect 642274 250633 642302 260485
rect 642262 250627 642314 250633
rect 642262 250569 642314 250575
rect 645140 243710 645196 243719
rect 648034 243677 648062 277856
rect 645140 243645 645142 243654
rect 645194 243645 645196 243654
rect 648022 243671 648074 243677
rect 645142 243613 645194 243619
rect 648022 243613 648074 243619
rect 649378 237757 649406 995157
rect 649750 995141 649802 995147
rect 649750 995083 649802 995089
rect 649654 995067 649706 995073
rect 649654 995009 649706 995015
rect 649558 983597 649610 983603
rect 649558 983539 649610 983545
rect 649462 983523 649514 983529
rect 649462 983465 649514 983471
rect 649474 274313 649502 983465
rect 649570 276533 649598 983539
rect 649666 964807 649694 995009
rect 649654 964801 649706 964807
rect 649654 964743 649706 964749
rect 649654 927431 649706 927437
rect 649654 927373 649706 927379
rect 649558 276527 649610 276533
rect 649558 276469 649610 276475
rect 649462 274307 649514 274313
rect 649462 274249 649514 274255
rect 649366 237751 649418 237757
rect 649366 237693 649418 237699
rect 639190 236287 639242 236293
rect 639284 236310 639340 236319
rect 638420 236245 638476 236254
rect 638806 236271 638858 236277
rect 638036 234090 638092 234099
rect 638036 234025 638092 234034
rect 637940 233942 637996 233951
rect 637940 233877 637996 233886
rect 637954 233484 637982 233877
rect 637186 233456 637598 233484
rect 637728 233456 637982 233484
rect 638050 233336 638078 234025
rect 638228 233498 638284 233507
rect 638434 233484 638462 236245
rect 638806 236213 638858 236219
rect 638818 233803 638846 236213
rect 638804 233794 638860 233803
rect 638804 233729 638860 233738
rect 638284 233470 638462 233484
rect 638818 233470 638846 233729
rect 638900 233646 638956 233655
rect 638900 233581 638956 233590
rect 638914 233484 638942 233581
rect 639202 233484 639230 236287
rect 649666 236277 649694 927373
rect 649762 754467 649790 995083
rect 649846 989961 649898 989967
rect 649846 989903 649898 989909
rect 649748 754458 649804 754467
rect 649748 754393 649804 754402
rect 649750 748869 649802 748875
rect 649750 748811 649802 748817
rect 639284 236245 639340 236254
rect 649654 236271 649706 236277
rect 649654 236213 649706 236219
rect 639766 236197 639818 236203
rect 639766 236139 639818 236145
rect 639778 233484 639806 236139
rect 638914 233470 639230 233484
rect 638284 233456 638448 233470
rect 638914 233456 639216 233470
rect 639552 233456 639806 233484
rect 638228 233433 638284 233442
rect 214114 233308 214176 233336
rect 227362 233308 227424 233336
rect 359842 233308 359904 233336
rect 381922 233308 381984 233336
rect 638050 233308 638112 233336
rect 210274 106176 210398 106204
rect 210274 86987 210302 106176
rect 210260 86978 210316 86987
rect 210260 86913 210316 86922
rect 210166 86791 210218 86797
rect 210166 86733 210218 86739
rect 210262 86495 210314 86501
rect 210262 86437 210314 86443
rect 210164 77802 210220 77811
rect 210164 77737 210220 77746
rect 210178 66096 210206 77737
rect 210274 66225 210302 86437
rect 210262 66219 210314 66225
rect 210262 66161 210314 66167
rect 210178 66068 210398 66096
rect 210262 65997 210314 66003
rect 210262 65939 210314 65945
rect 210164 56046 210220 56055
rect 210164 55981 210220 55990
rect 210178 55273 210206 55981
rect 210166 55267 210218 55273
rect 210166 55209 210218 55215
rect 210274 55144 210302 65939
rect 210178 55116 210302 55144
rect 210178 52905 210206 55116
rect 210260 55010 210316 55019
rect 210260 54945 210316 54954
rect 210274 53867 210302 54945
rect 210262 53861 210314 53867
rect 210262 53803 210314 53809
rect 210370 53571 210398 66068
rect 217174 54305 217226 54311
rect 210836 54270 210892 54279
rect 210836 54205 210892 54214
rect 214772 54270 214828 54279
rect 214828 54228 214896 54256
rect 228502 54305 228554 54311
rect 217174 54247 217226 54253
rect 214772 54205 214828 54214
rect 210740 54122 210796 54131
rect 210740 54057 210796 54066
rect 210358 53565 210410 53571
rect 210358 53507 210410 53513
rect 210754 53127 210782 54057
rect 210850 54015 210878 54205
rect 216980 54122 217036 54131
rect 217036 54080 217104 54108
rect 216980 54057 217036 54066
rect 210838 54009 210890 54015
rect 210838 53951 210890 53957
rect 216982 54009 217034 54015
rect 216982 53951 217034 53957
rect 213408 53784 213470 53812
rect 210742 53121 210794 53127
rect 210742 53063 210794 53069
rect 210166 52899 210218 52905
rect 210166 52841 210218 52847
rect 210070 48977 210122 48983
rect 210070 48919 210122 48925
rect 209014 48829 209066 48835
rect 209014 48771 209066 48777
rect 208918 48237 208970 48243
rect 208918 48179 208970 48185
rect 208822 48163 208874 48169
rect 208822 48105 208874 48111
rect 208726 46757 208778 46763
rect 208726 46699 208778 46705
rect 208630 46535 208682 46541
rect 208630 46477 208682 46483
rect 208534 46387 208586 46393
rect 208534 46329 208586 46335
rect 208438 46313 208490 46319
rect 208438 46255 208490 46261
rect 208342 46239 208394 46245
rect 208342 46181 208394 46187
rect 206902 42169 206954 42175
rect 206902 42111 206954 42117
rect 187604 41838 187660 41847
rect 187344 41796 187604 41824
rect 194324 41838 194380 41847
rect 194064 41796 194324 41824
rect 187604 41773 187660 41782
rect 194324 41773 194380 41782
rect 211042 40811 211070 53650
rect 211200 53636 211262 53664
rect 211392 53636 211454 53664
rect 211234 51795 211262 53636
rect 211222 51789 211274 51795
rect 211222 51731 211274 51737
rect 211426 45357 211454 53636
rect 211570 53368 211598 53650
rect 211714 53636 211776 53664
rect 211570 53340 211646 53368
rect 211618 49723 211646 53340
rect 211606 49717 211658 49723
rect 211606 49659 211658 49665
rect 211414 45351 211466 45357
rect 211414 45293 211466 45299
rect 211714 45103 211742 53636
rect 211954 53368 211982 53650
rect 211954 53340 212030 53368
rect 211894 52529 211946 52535
rect 211894 52471 211946 52477
rect 211906 52091 211934 52471
rect 211894 52085 211946 52091
rect 211894 52027 211946 52033
rect 212002 51911 212030 53340
rect 211988 51902 212044 51911
rect 211988 51837 212044 51846
rect 212098 45251 212126 53650
rect 212304 53636 212414 53664
rect 212182 52381 212234 52387
rect 212182 52323 212234 52329
rect 212194 52165 212222 52323
rect 212182 52159 212234 52165
rect 212182 52101 212234 52107
rect 212386 52091 212414 53636
rect 212374 52085 212426 52091
rect 212374 52027 212426 52033
rect 212084 45242 212140 45251
rect 212084 45177 212140 45186
rect 211700 45094 211756 45103
rect 211700 45029 211756 45038
rect 212482 42397 212510 53650
rect 212674 52059 212702 53650
rect 212660 52050 212716 52059
rect 212660 51985 212716 51994
rect 212866 45209 212894 53650
rect 213058 53539 213086 53650
rect 213044 53530 213100 53539
rect 213044 53465 213100 53474
rect 213250 45283 213278 53650
rect 213442 53349 213470 53784
rect 216994 53719 217022 53951
rect 216982 53713 217034 53719
rect 213600 53636 213662 53664
rect 213430 53343 213482 53349
rect 213430 53285 213482 53291
rect 213430 52085 213482 52091
rect 213430 52027 213482 52033
rect 213442 51869 213470 52027
rect 213430 51863 213482 51869
rect 213430 51805 213482 51811
rect 213238 45277 213290 45283
rect 213238 45219 213290 45225
rect 212854 45203 212906 45209
rect 212854 45145 212906 45151
rect 212470 42391 212522 42397
rect 212470 42333 212522 42339
rect 213634 42101 213662 53636
rect 213778 53627 213806 53650
rect 213730 53599 213806 53627
rect 213922 53636 213984 53664
rect 214114 53636 214176 53664
rect 213730 53275 213758 53599
rect 213718 53269 213770 53275
rect 213718 53211 213770 53217
rect 213922 45135 213950 53636
rect 214114 51721 214142 53636
rect 214102 51715 214154 51721
rect 214102 51657 214154 51663
rect 213910 45129 213962 45135
rect 213910 45071 213962 45077
rect 213622 42095 213674 42101
rect 213622 42037 213674 42043
rect 214306 42027 214334 53650
rect 214498 51647 214526 53650
rect 214486 51641 214538 51647
rect 214486 51583 214538 51589
rect 214690 44987 214718 53650
rect 215074 45061 215102 53650
rect 215266 53571 215294 53650
rect 215254 53565 215306 53571
rect 215254 53507 215306 53513
rect 215062 45055 215114 45061
rect 215062 44997 215114 45003
rect 214678 44981 214730 44987
rect 215458 44955 215486 53650
rect 215602 53571 215630 53650
rect 215794 53571 215822 53650
rect 215590 53565 215642 53571
rect 215590 53507 215642 53513
rect 215782 53565 215834 53571
rect 215986 53539 216014 53650
rect 216130 53636 216192 53664
rect 216982 53655 217034 53661
rect 215782 53507 215834 53513
rect 215972 53530 216028 53539
rect 215972 53465 216028 53474
rect 216130 50389 216158 53636
rect 216370 53497 216398 53650
rect 216358 53491 216410 53497
rect 216358 53433 216410 53439
rect 216118 50383 216170 50389
rect 216118 50325 216170 50331
rect 215830 49495 215882 49501
rect 215830 49437 215882 49443
rect 215926 49495 215978 49501
rect 215926 49437 215978 49443
rect 215842 49372 215870 49437
rect 215938 49372 215966 49437
rect 215842 49344 215966 49372
rect 216514 47725 216542 53650
rect 216706 53391 216734 53650
rect 216692 53382 216748 53391
rect 216692 53317 216748 53326
rect 216898 50315 216926 53650
rect 217186 53571 217214 54247
rect 219202 54237 219312 54256
rect 228502 54247 228554 54253
rect 219190 54231 219312 54237
rect 219242 54228 219312 54231
rect 219190 54173 219242 54179
rect 221410 54089 221520 54108
rect 221398 54083 221520 54089
rect 221450 54080 221520 54083
rect 221398 54025 221450 54031
rect 221396 53974 221452 53983
rect 221396 53909 221452 53918
rect 218194 53793 218222 53798
rect 218182 53787 218234 53793
rect 218182 53729 218234 53735
rect 217174 53565 217226 53571
rect 217174 53507 217226 53513
rect 217282 52757 217310 53650
rect 217474 53571 217502 53650
rect 217462 53565 217514 53571
rect 217462 53507 217514 53513
rect 217270 52751 217322 52757
rect 217270 52693 217322 52699
rect 216886 50309 216938 50315
rect 216886 50251 216938 50257
rect 217666 50241 217694 53650
rect 217824 53636 217886 53664
rect 218016 53636 218078 53664
rect 217858 53243 217886 53636
rect 217844 53234 217900 53243
rect 217844 53169 217900 53178
rect 217654 50235 217706 50241
rect 217654 50177 217706 50183
rect 216502 47719 216554 47725
rect 216502 47661 216554 47667
rect 218050 47651 218078 53636
rect 218338 53636 218400 53664
rect 218530 53636 218592 53664
rect 218038 47645 218090 47651
rect 218038 47587 218090 47593
rect 218338 47503 218366 53636
rect 218530 47651 218558 53636
rect 218518 47645 218570 47651
rect 218518 47587 218570 47593
rect 218722 47577 218750 53650
rect 218914 52905 218942 53650
rect 218902 52899 218954 52905
rect 218902 52841 218954 52847
rect 218806 49495 218858 49501
rect 218806 49437 218858 49443
rect 218818 49353 218846 49437
rect 218806 49347 218858 49353
rect 218806 49289 218858 49295
rect 219106 48021 219134 53650
rect 219490 48095 219518 53650
rect 219682 53497 219710 53650
rect 219670 53491 219722 53497
rect 219670 53433 219722 53439
rect 219874 52239 219902 53650
rect 220032 53636 220094 53664
rect 220224 53636 220286 53664
rect 220066 52979 220094 53636
rect 220054 52973 220106 52979
rect 220054 52915 220106 52921
rect 219862 52233 219914 52239
rect 219862 52175 219914 52181
rect 219478 48089 219530 48095
rect 219478 48031 219530 48037
rect 219094 48015 219146 48021
rect 219094 47957 219146 47963
rect 220258 47799 220286 53636
rect 220402 53368 220430 53650
rect 220354 53340 220430 53368
rect 220546 53636 220608 53664
rect 220738 53636 220800 53664
rect 220354 53053 220382 53340
rect 220342 53047 220394 53053
rect 220342 52989 220394 52995
rect 220546 47873 220574 53636
rect 220738 48983 220766 53636
rect 220930 52535 220958 53650
rect 221122 53539 221150 53650
rect 221108 53530 221164 53539
rect 221108 53465 221164 53474
rect 220918 52529 220970 52535
rect 220918 52471 220970 52477
rect 220726 48977 220778 48983
rect 220726 48919 220778 48925
rect 221314 47947 221342 53650
rect 221410 53053 221438 53909
rect 221398 53047 221450 53053
rect 221398 52989 221450 52995
rect 221698 48761 221726 53650
rect 221890 52355 221918 53650
rect 221876 52346 221932 52355
rect 221876 52281 221932 52290
rect 222082 48835 222110 53650
rect 222240 53636 222302 53664
rect 222432 53636 222494 53664
rect 222274 48909 222302 53636
rect 222262 48903 222314 48909
rect 222262 48845 222314 48851
rect 222070 48829 222122 48835
rect 222070 48771 222122 48777
rect 221686 48755 221738 48761
rect 221686 48697 221738 48703
rect 222466 48243 222494 53636
rect 222610 53368 222638 53650
rect 222754 53636 222816 53664
rect 222946 53636 223008 53664
rect 222610 53340 222686 53368
rect 222658 51763 222686 53340
rect 222644 51754 222700 51763
rect 222644 51689 222700 51698
rect 222454 48237 222506 48243
rect 222454 48179 222506 48185
rect 222754 48169 222782 53636
rect 222946 48835 222974 53636
rect 222934 48829 222986 48835
rect 222934 48771 222986 48777
rect 222742 48163 222794 48169
rect 222742 48105 222794 48111
rect 221302 47941 221354 47947
rect 221302 47883 221354 47889
rect 220534 47867 220586 47873
rect 220534 47809 220586 47815
rect 220246 47793 220298 47799
rect 220246 47735 220298 47741
rect 218710 47571 218762 47577
rect 218710 47513 218762 47519
rect 218326 47497 218378 47503
rect 218326 47439 218378 47445
rect 223138 46541 223166 53650
rect 223330 52207 223358 53650
rect 223316 52198 223372 52207
rect 223316 52133 223372 52142
rect 223522 46763 223550 53650
rect 223714 48983 223742 53650
rect 223702 48977 223754 48983
rect 223702 48919 223754 48925
rect 223510 46757 223562 46763
rect 223510 46699 223562 46705
rect 223906 46615 223934 53650
rect 224098 48761 224126 53650
rect 224290 49871 224318 53650
rect 224640 53636 224702 53664
rect 224278 49865 224330 49871
rect 224278 49807 224330 49813
rect 224086 48755 224138 48761
rect 224086 48697 224138 48703
rect 223894 46609 223946 46615
rect 223894 46551 223946 46557
rect 223126 46535 223178 46541
rect 223126 46477 223178 46483
rect 224674 46393 224702 53636
rect 224962 53636 225024 53664
rect 224962 49945 224990 53636
rect 224950 49939 225002 49945
rect 224950 49881 225002 49887
rect 225346 49797 225374 53650
rect 225730 52165 225758 53650
rect 225718 52159 225770 52165
rect 225718 52101 225770 52107
rect 225334 49791 225386 49797
rect 225334 49733 225386 49739
rect 224662 46387 224714 46393
rect 224662 46329 224714 46335
rect 226114 46319 226142 53650
rect 226102 46313 226154 46319
rect 226102 46255 226154 46261
rect 226498 46245 226526 53650
rect 226594 53636 226848 53664
rect 226978 53636 227232 53664
rect 226594 49649 226622 53636
rect 226978 52387 227006 53636
rect 226966 52381 227018 52387
rect 226966 52323 227018 52329
rect 227554 51943 227582 53650
rect 227542 51937 227594 51943
rect 227542 51879 227594 51885
rect 226582 49643 226634 49649
rect 226582 49585 226634 49591
rect 227938 46911 227966 53650
rect 228322 50759 228350 53650
rect 228514 53571 228542 54247
rect 256054 54157 256106 54163
rect 256054 54099 256106 54105
rect 228502 53565 228554 53571
rect 228502 53507 228554 53513
rect 228310 50753 228362 50759
rect 228310 50695 228362 50701
rect 228706 50685 228734 53650
rect 228802 53636 229056 53664
rect 229186 53636 229440 53664
rect 228694 50679 228746 50685
rect 228694 50621 228746 50627
rect 228802 50537 228830 53636
rect 228790 50531 228842 50537
rect 228790 50473 228842 50479
rect 227926 46905 227978 46911
rect 227926 46847 227978 46853
rect 229186 46467 229214 53636
rect 229762 50611 229790 53650
rect 229750 50605 229802 50611
rect 229750 50547 229802 50553
rect 229652 50422 229708 50431
rect 229652 50357 229708 50366
rect 229666 48983 229694 50357
rect 229654 48977 229706 48983
rect 229654 48919 229706 48925
rect 230146 46689 230174 53650
rect 230530 50833 230558 53650
rect 230518 50827 230570 50833
rect 230518 50769 230570 50775
rect 230914 47059 230942 53650
rect 231010 53636 231264 53664
rect 231394 53636 231648 53664
rect 231010 50981 231038 53636
rect 230998 50975 231050 50981
rect 230998 50917 231050 50923
rect 231394 50907 231422 53636
rect 231970 51055 231998 53650
rect 232354 51129 232382 53650
rect 232342 51123 232394 51129
rect 232342 51065 232394 51071
rect 231958 51049 232010 51055
rect 231958 50991 232010 50997
rect 231382 50901 231434 50907
rect 231382 50843 231434 50849
rect 232738 50019 232766 53650
rect 232726 50013 232778 50019
rect 232726 49955 232778 49961
rect 230902 47053 230954 47059
rect 230902 46995 230954 47001
rect 233122 46837 233150 53650
rect 233314 53636 233472 53664
rect 233602 53636 233856 53664
rect 233314 47207 233342 53636
rect 233602 51425 233630 53636
rect 233590 51419 233642 51425
rect 233590 51361 233642 51367
rect 234178 48613 234206 53650
rect 234562 51351 234590 53650
rect 234550 51345 234602 51351
rect 234550 51287 234602 51293
rect 234946 51203 234974 53650
rect 235330 51277 235358 53650
rect 235426 53636 235680 53664
rect 235810 53636 236064 53664
rect 235318 51271 235370 51277
rect 235318 51213 235370 51219
rect 234934 51197 234986 51203
rect 234934 51139 234986 51145
rect 235426 50093 235454 53636
rect 235810 50167 235838 53636
rect 235798 50161 235850 50167
rect 235798 50103 235850 50109
rect 235414 50087 235466 50093
rect 235414 50029 235466 50035
rect 236386 48687 236414 53650
rect 236770 51573 236798 53650
rect 236758 51567 236810 51573
rect 236758 51509 236810 51515
rect 237154 51499 237182 53650
rect 237430 51863 237482 51869
rect 237430 51805 237482 51811
rect 237442 51573 237470 51805
rect 237430 51567 237482 51573
rect 237430 51509 237482 51515
rect 237142 51493 237194 51499
rect 237142 51435 237194 51441
rect 237538 51319 237566 53650
rect 237634 53636 237888 53664
rect 238018 53636 238272 53664
rect 237634 51467 237662 53636
rect 237620 51458 237676 51467
rect 237620 51393 237676 51402
rect 237524 51310 237580 51319
rect 237524 51245 237580 51254
rect 236374 48681 236426 48687
rect 236374 48623 236426 48629
rect 234166 48607 234218 48613
rect 234166 48549 234218 48555
rect 238018 47429 238046 53636
rect 238006 47423 238058 47429
rect 238006 47365 238058 47371
rect 238594 47355 238622 53650
rect 238582 47349 238634 47355
rect 238582 47291 238634 47297
rect 238978 47281 239006 53650
rect 239062 52307 239114 52313
rect 239062 52249 239114 52255
rect 239074 51869 239102 52249
rect 239062 51863 239114 51869
rect 239062 51805 239114 51811
rect 238966 47275 239018 47281
rect 238966 47217 239018 47223
rect 233302 47201 233354 47207
rect 233302 47143 233354 47149
rect 239362 47133 239390 53650
rect 239746 48391 239774 53650
rect 239842 53636 240096 53664
rect 240226 53636 240480 53664
rect 239842 48465 239870 53636
rect 240226 48539 240254 53636
rect 240214 48533 240266 48539
rect 240214 48475 240266 48481
rect 239830 48459 239882 48465
rect 239830 48401 239882 48407
rect 239734 48385 239786 48391
rect 239734 48327 239786 48333
rect 239350 47127 239402 47133
rect 239350 47069 239402 47075
rect 240802 46985 240830 53650
rect 241186 49353 241214 53650
rect 241174 49347 241226 49353
rect 241174 49289 241226 49295
rect 241570 48317 241598 53650
rect 241558 48311 241610 48317
rect 241558 48253 241610 48259
rect 241954 48211 241982 53650
rect 242050 53636 242304 53664
rect 242434 53636 242688 53664
rect 242050 48655 242078 53636
rect 242434 48803 242462 53636
rect 242420 48794 242476 48803
rect 242420 48729 242476 48738
rect 242036 48646 242092 48655
rect 242036 48581 242092 48590
rect 243010 48507 243038 53650
rect 243394 51615 243422 53650
rect 243380 51606 243436 51615
rect 243380 51541 243436 51550
rect 242996 48498 243052 48507
rect 242996 48433 243052 48442
rect 243778 48359 243806 53650
rect 244162 51869 244190 53650
rect 256066 53516 256094 54099
rect 282166 53935 282218 53941
rect 282166 53877 282218 53883
rect 282178 53775 282206 53877
rect 282178 53747 282398 53775
rect 256066 53497 256286 53516
rect 256066 53491 256298 53497
rect 256066 53488 256246 53491
rect 256246 53433 256298 53439
rect 255958 53417 256010 53423
rect 256150 53417 256202 53423
rect 256010 53365 256150 53368
rect 255958 53359 256202 53365
rect 255970 53340 256190 53359
rect 273620 53271 273676 53280
rect 273620 53206 273676 53215
rect 276406 53121 276458 53127
rect 276598 53121 276650 53127
rect 276458 53081 276598 53109
rect 276406 53063 276458 53069
rect 276598 53063 276650 53069
rect 244150 51863 244202 51869
rect 244150 51805 244202 51811
rect 254422 51863 254474 51869
rect 254422 51805 254474 51811
rect 251926 51715 251978 51721
rect 251926 51657 251978 51663
rect 251938 51499 251966 51657
rect 253558 51641 253610 51647
rect 253558 51583 253610 51589
rect 251926 51493 251978 51499
rect 251926 51435 251978 51441
rect 253462 51493 253514 51499
rect 253570 51444 253598 51583
rect 253514 51441 253598 51444
rect 253462 51435 253598 51441
rect 253474 51416 253598 51435
rect 254434 51425 254462 51805
rect 254422 51419 254474 51425
rect 254422 51361 254474 51367
rect 282370 48983 282398 53747
rect 357430 53639 357482 53645
rect 357430 53581 357482 53587
rect 383158 53639 383210 53645
rect 383158 53581 383210 53587
rect 403126 53639 403178 53645
rect 403126 53581 403178 53587
rect 443362 53636 443678 53664
rect 293686 53343 293738 53349
rect 293686 53285 293738 53291
rect 293698 53243 293726 53285
rect 321046 53269 321098 53275
rect 293684 53234 293740 53243
rect 321046 53211 321098 53217
rect 293684 53169 293740 53178
rect 321058 53053 321086 53211
rect 331126 53195 331178 53201
rect 331126 53137 331178 53143
rect 331138 53053 331166 53137
rect 321046 53047 321098 53053
rect 321046 52989 321098 52995
rect 331126 53047 331178 53053
rect 331126 52989 331178 52995
rect 331126 52011 331178 52017
rect 331126 51953 331178 51959
rect 342550 52011 342602 52017
rect 342550 51953 342602 51959
rect 331138 51869 331166 51953
rect 322582 51863 322634 51869
rect 322498 51823 322582 51851
rect 322498 51795 322526 51823
rect 322582 51805 322634 51811
rect 331126 51863 331178 51869
rect 331126 51805 331178 51811
rect 308086 51789 308138 51795
rect 308182 51789 308234 51795
rect 308138 51737 308182 51740
rect 308086 51731 308234 51737
rect 322486 51789 322538 51795
rect 322486 51731 322538 51737
rect 342562 51740 342590 51953
rect 342742 51863 342794 51869
rect 342742 51805 342794 51811
rect 342754 51740 342782 51805
rect 308098 51712 308222 51731
rect 322390 51715 322442 51721
rect 342562 51712 342782 51740
rect 322390 51657 322442 51663
rect 308086 51641 308138 51647
rect 308182 51641 308234 51647
rect 308138 51601 308182 51629
rect 308086 51583 308138 51589
rect 308182 51583 308234 51589
rect 322402 51573 322430 51657
rect 342742 51641 342794 51647
rect 342658 51589 342742 51592
rect 342658 51583 342794 51589
rect 342658 51573 342782 51583
rect 322390 51567 322442 51573
rect 322390 51509 322442 51515
rect 342646 51567 342782 51573
rect 342698 51564 342782 51567
rect 342646 51509 342698 51515
rect 282358 48977 282410 48983
rect 282358 48919 282410 48925
rect 302422 48977 302474 48983
rect 302422 48919 302474 48925
rect 243764 48350 243820 48359
rect 243764 48285 243820 48294
rect 241940 48202 241996 48211
rect 241940 48137 241996 48146
rect 240790 46979 240842 46985
rect 240790 46921 240842 46927
rect 233110 46831 233162 46837
rect 233110 46773 233162 46779
rect 230134 46683 230186 46689
rect 230134 46625 230186 46631
rect 229174 46461 229226 46467
rect 229174 46403 229226 46409
rect 226486 46239 226538 46245
rect 226486 46181 226538 46187
rect 214678 44923 214730 44929
rect 215444 44946 215500 44955
rect 215444 44881 215500 44890
rect 302434 42143 302462 48919
rect 302516 43318 302572 43327
rect 302516 43253 302572 43262
rect 302420 42134 302476 42143
rect 302530 42120 302558 43253
rect 310102 42391 310154 42397
rect 310102 42333 310154 42339
rect 306740 42134 306796 42143
rect 302530 42092 302688 42120
rect 302420 42069 302476 42078
rect 306796 42092 307008 42120
rect 310114 42106 310142 42333
rect 357442 42106 357470 53581
rect 362722 53340 363038 53368
rect 362722 53201 362750 53340
rect 363010 53201 363038 53340
rect 383062 53269 383114 53275
rect 383170 53257 383198 53581
rect 398326 53565 398378 53571
rect 398326 53507 398378 53513
rect 403138 53516 403166 53581
rect 443362 53571 443390 53636
rect 423574 53565 423626 53571
rect 383114 53229 383198 53257
rect 383062 53211 383114 53217
rect 362710 53195 362762 53201
rect 362710 53137 362762 53143
rect 362998 53195 363050 53201
rect 362998 53137 363050 53143
rect 368482 51869 368606 51888
rect 368470 51863 368618 51869
rect 368522 51860 368566 51863
rect 368470 51805 368522 51811
rect 368566 51805 368618 51811
rect 394306 51712 394526 51740
rect 362998 51641 363050 51647
rect 362818 51589 362998 51592
rect 374422 51641 374474 51647
rect 362818 51583 363050 51589
rect 374420 51606 374422 51615
rect 394306 51615 394334 51712
rect 394498 51647 394526 51712
rect 394486 51641 394538 51647
rect 374474 51606 374476 51615
rect 362818 51573 363038 51583
rect 362806 51567 363038 51573
rect 362858 51564 363038 51567
rect 374420 51541 374476 51550
rect 394292 51606 394348 51615
rect 394486 51583 394538 51589
rect 394292 51541 394348 51550
rect 362806 51509 362858 51515
rect 398338 46171 398366 53507
rect 403138 53488 403454 53516
rect 423574 53507 423626 53513
rect 443350 53565 443402 53571
rect 443350 53507 443402 53513
rect 403138 53340 403358 53368
rect 403426 53349 403454 53488
rect 403138 53201 403166 53340
rect 403330 53201 403358 53340
rect 403414 53343 403466 53349
rect 403414 53285 403466 53291
rect 423382 53343 423434 53349
rect 423382 53285 423434 53291
rect 423394 53257 423422 53285
rect 423586 53257 423614 53507
rect 443446 53491 443498 53497
rect 443446 53433 443498 53439
rect 443350 53417 443402 53423
rect 443350 53359 443402 53365
rect 423394 53229 423614 53257
rect 440660 53234 440716 53243
rect 403126 53195 403178 53201
rect 403126 53137 403178 53143
rect 403318 53195 403370 53201
rect 440660 53169 440662 53178
rect 403318 53137 403370 53143
rect 440714 53169 440716 53178
rect 440662 53137 440714 53143
rect 443362 52609 443390 53359
rect 443350 52603 443402 52609
rect 443350 52545 443402 52551
rect 408898 51869 409022 51888
rect 408886 51863 409034 51869
rect 408938 51860 408982 51863
rect 408886 51805 408938 51811
rect 408982 51805 409034 51811
rect 414646 51715 414698 51721
rect 414646 51657 414698 51663
rect 414658 51425 414686 51657
rect 423286 51641 423338 51647
rect 423382 51641 423434 51647
rect 423338 51589 423382 51592
rect 423286 51583 423434 51589
rect 417526 51567 417578 51573
rect 423298 51564 423422 51583
rect 417526 51509 417578 51515
rect 417538 51425 417566 51509
rect 414646 51419 414698 51425
rect 414646 51361 414698 51367
rect 417526 51419 417578 51425
rect 417526 51361 417578 51367
rect 443458 49057 443486 53433
rect 443650 53349 443678 53636
rect 490966 53639 491018 53645
rect 490966 53581 491018 53587
rect 460822 53565 460874 53571
rect 460822 53507 460874 53513
rect 460834 53423 460862 53507
rect 460822 53417 460874 53423
rect 460822 53359 460874 53365
rect 490978 53349 491006 53581
rect 443638 53343 443690 53349
rect 443638 53285 443690 53291
rect 490966 53343 491018 53349
rect 490966 53285 491018 53291
rect 512278 53343 512330 53349
rect 512278 53285 512330 53291
rect 443734 53269 443786 53275
rect 443732 53234 443734 53243
rect 443786 53234 443788 53243
rect 443732 53169 443788 53178
rect 460726 52603 460778 52609
rect 460726 52545 460778 52551
rect 449218 51869 449342 51888
rect 449206 51863 449354 51869
rect 449258 51860 449302 51863
rect 449206 51805 449258 51811
rect 449302 51805 449354 51811
rect 460738 51740 460766 52545
rect 460822 52011 460874 52017
rect 460822 51953 460874 51959
rect 470806 52011 470858 52017
rect 470806 51953 470858 51959
rect 460834 51869 460862 51953
rect 460822 51863 460874 51869
rect 460822 51805 460874 51811
rect 460738 51712 460862 51740
rect 470818 51721 470846 51953
rect 509782 51863 509834 51869
rect 509782 51805 509834 51811
rect 457942 51641 457994 51647
rect 457940 51606 457942 51615
rect 457994 51606 457996 51615
rect 457940 51541 457996 51550
rect 443446 49051 443498 49057
rect 443446 48993 443498 48999
rect 398326 46165 398378 46171
rect 460834 46139 460862 51712
rect 470806 51715 470858 51721
rect 470806 51657 470858 51663
rect 509686 51715 509738 51721
rect 509794 51703 509822 51805
rect 509738 51675 509822 51703
rect 509686 51657 509738 51663
rect 480886 51641 480938 51647
rect 478004 51606 478060 51615
rect 498262 51641 498314 51647
rect 480886 51583 480938 51589
rect 498260 51606 498262 51615
rect 498314 51606 498316 51615
rect 478004 51541 478060 51550
rect 478018 51499 478046 51541
rect 480898 51499 480926 51583
rect 498260 51541 498316 51550
rect 478006 51493 478058 51499
rect 478006 51435 478058 51441
rect 480886 51493 480938 51499
rect 480886 51435 480938 51441
rect 512290 49099 512318 53285
rect 525910 53269 525962 53275
rect 525910 53211 525962 53217
rect 518326 51715 518378 51721
rect 518326 51657 518378 51663
rect 518338 51615 518366 51657
rect 518324 51606 518380 51615
rect 518324 51541 518380 51550
rect 512276 49090 512332 49099
rect 512276 49025 512332 49034
rect 471382 48977 471434 48983
rect 471382 48919 471434 48925
rect 398326 46107 398378 46113
rect 460820 46130 460876 46139
rect 408886 46091 408938 46097
rect 460820 46065 460876 46074
rect 465812 46130 465868 46139
rect 465812 46065 465868 46074
rect 408886 46033 408938 46039
rect 361750 45351 361802 45357
rect 361750 45293 361802 45299
rect 361762 42106 361790 45293
rect 406102 45277 406154 45283
rect 406102 45219 406154 45225
rect 364916 43318 364972 43327
rect 364916 43253 364972 43262
rect 364930 42106 364958 43253
rect 406114 43211 406142 45219
rect 406102 43205 406154 43211
rect 406102 43147 406154 43153
rect 405238 42169 405290 42175
rect 405290 42117 405552 42120
rect 405238 42111 405552 42117
rect 405250 42092 405552 42111
rect 306740 42069 306796 42078
rect 214294 42021 214346 42027
rect 214294 41963 214346 41969
rect 408898 41824 408926 46033
rect 411574 45203 411626 45209
rect 411574 45145 411626 45151
rect 410998 43205 411050 43211
rect 411050 43153 411102 43156
rect 410998 43147 411102 43153
rect 411010 43128 411102 43147
rect 411586 42143 411614 45145
rect 443926 45129 443978 45135
rect 443926 45071 443978 45077
rect 411572 42134 411628 42143
rect 411572 42069 411628 42078
rect 416276 42134 416332 42143
rect 416332 42092 416592 42120
rect 416276 42069 416332 42078
rect 408898 41796 409296 41824
rect 211028 40802 211084 40811
rect 211028 40737 211084 40746
rect 136532 40210 136588 40219
rect 136532 40145 136588 40154
rect 443938 37439 443966 45071
rect 465826 44340 465854 46065
rect 465826 44312 465856 44340
rect 465828 44178 465856 44312
rect 460066 42101 460368 42120
rect 471394 42106 471422 48919
rect 509686 45055 509738 45061
rect 509686 44997 509738 45003
rect 508246 44981 508298 44987
rect 508246 44923 508298 44929
rect 508258 43285 508286 44923
rect 508246 43279 508298 43285
rect 508246 43221 508298 43227
rect 460054 42095 460368 42101
rect 460106 42092 460368 42095
rect 460054 42037 460106 42043
rect 509698 41847 509726 44997
rect 521494 43205 521546 43211
rect 521494 43147 521546 43153
rect 520436 42134 520492 42143
rect 521506 42120 521534 43147
rect 525922 42120 525950 53211
rect 639682 52017 639710 233456
rect 649762 233243 649790 748811
rect 649858 707551 649886 989903
rect 649844 707542 649900 707551
rect 649844 707477 649900 707486
rect 649846 702767 649898 702773
rect 649846 702709 649898 702715
rect 649858 236351 649886 702709
rect 649954 660635 649982 995749
rect 650228 994070 650284 994079
rect 650228 994005 650284 994014
rect 650038 992107 650090 992113
rect 650038 992049 650090 992055
rect 650050 801383 650078 992049
rect 650134 989369 650186 989375
rect 650134 989311 650186 989317
rect 650146 848299 650174 989311
rect 650242 907161 650270 994005
rect 658102 989295 658154 989301
rect 658102 989237 658154 989243
rect 658006 986483 658058 986489
rect 658006 986425 658058 986431
rect 655124 976754 655180 976763
rect 655124 976689 655180 976698
rect 653782 964801 653834 964807
rect 653782 964743 653834 964749
rect 653794 941539 653822 964743
rect 653780 941530 653836 941539
rect 653780 941465 653836 941474
rect 655138 939129 655166 976689
rect 655220 965062 655276 965071
rect 655220 964997 655276 965006
rect 655234 939277 655262 964997
rect 655316 953370 655372 953379
rect 655316 953305 655372 953314
rect 655330 939425 655358 953305
rect 655318 939419 655370 939425
rect 655318 939361 655370 939367
rect 655222 939271 655274 939277
rect 655222 939213 655274 939219
rect 655126 939123 655178 939129
rect 655126 939065 655178 939071
rect 658018 936317 658046 986425
rect 658114 939573 658142 989237
rect 660886 986409 660938 986415
rect 660886 986351 660938 986357
rect 658102 939567 658154 939573
rect 658102 939509 658154 939515
rect 660898 938019 660926 986351
rect 674518 983745 674570 983751
rect 674518 983687 674570 983693
rect 674134 983671 674186 983677
rect 674134 983613 674186 983619
rect 674146 959299 674174 983613
rect 674530 966551 674558 983687
rect 675106 966722 675408 966750
rect 674516 966542 674572 966551
rect 674516 966477 674572 966486
rect 675106 960756 675134 966722
rect 675284 966542 675340 966551
rect 675284 966477 675340 966486
rect 675298 961348 675326 966477
rect 675778 965811 675806 966070
rect 675764 965802 675820 965811
rect 675764 965737 675820 965746
rect 675394 965071 675422 965435
rect 675380 965062 675436 965071
rect 675380 964997 675436 965006
rect 675778 963443 675806 963595
rect 675764 963434 675820 963443
rect 675764 963369 675820 963378
rect 675682 962555 675710 963036
rect 675668 962546 675724 962555
rect 675668 962481 675724 962490
rect 675394 962259 675422 962399
rect 675380 962250 675436 962259
rect 675380 962185 675436 962194
rect 675778 961519 675806 961778
rect 675764 961510 675820 961519
rect 675764 961445 675820 961454
rect 675298 961320 675422 961348
rect 675394 961200 675422 961320
rect 675394 961186 675504 961200
rect 675408 961172 675518 961186
rect 675490 960779 675518 961172
rect 674914 960728 675134 960756
rect 675476 960770 675532 960779
rect 674132 959290 674188 959299
rect 674132 959225 674188 959234
rect 669526 954737 669578 954743
rect 669526 954679 669578 954685
rect 660886 938013 660938 938019
rect 660886 937955 660938 937961
rect 658006 936311 658058 936317
rect 658006 936253 658058 936259
rect 654452 929838 654508 929847
rect 654452 929773 654508 929782
rect 654466 927511 654494 929773
rect 654454 927505 654506 927511
rect 654454 927447 654506 927453
rect 666742 927505 666794 927511
rect 666742 927447 666794 927453
rect 653972 918146 654028 918155
rect 653972 918081 654028 918090
rect 653986 915893 654014 918081
rect 653974 915887 654026 915893
rect 653974 915829 654026 915835
rect 660982 915887 661034 915893
rect 660982 915829 661034 915835
rect 650230 907155 650282 907161
rect 650230 907097 650282 907103
rect 653782 907155 653834 907161
rect 653782 907097 653834 907103
rect 653794 894623 653822 907097
rect 654452 906454 654508 906463
rect 654452 906389 654508 906398
rect 654466 904423 654494 906389
rect 654454 904417 654506 904423
rect 654454 904359 654506 904365
rect 653780 894614 653836 894623
rect 653780 894549 653836 894558
rect 653972 882922 654028 882931
rect 653972 882857 654028 882866
rect 653986 881335 654014 882857
rect 653974 881329 654026 881335
rect 653974 881271 654026 881277
rect 660886 881329 660938 881335
rect 660886 881271 660938 881277
rect 654452 871230 654508 871239
rect 654452 871165 654508 871174
rect 654466 869865 654494 871165
rect 654454 869859 654506 869865
rect 654454 869801 654506 869807
rect 654164 859538 654220 859547
rect 654164 859473 654220 859482
rect 654178 858321 654206 859473
rect 654166 858315 654218 858321
rect 654166 858257 654218 858263
rect 650132 848290 650188 848299
rect 650132 848225 650188 848234
rect 653972 836006 654028 836015
rect 653972 835941 654028 835950
rect 653986 835233 654014 835941
rect 653974 835227 654026 835233
rect 653974 835169 654026 835175
rect 653972 824314 654028 824323
rect 653972 824249 654028 824258
rect 653986 823763 654014 824249
rect 653974 823757 654026 823763
rect 653974 823699 654026 823705
rect 654452 812622 654508 812631
rect 654452 812557 654508 812566
rect 654466 812219 654494 812557
rect 654454 812213 654506 812219
rect 654454 812155 654506 812161
rect 650036 801374 650092 801383
rect 650036 801309 650092 801318
rect 654068 789090 654124 789099
rect 654068 789025 654124 789034
rect 654082 786319 654110 789025
rect 654070 786313 654122 786319
rect 654070 786255 654122 786261
rect 654068 777398 654124 777407
rect 654068 777333 654124 777342
rect 654082 774775 654110 777333
rect 654070 774769 654122 774775
rect 654070 774711 654122 774717
rect 653972 765558 654028 765567
rect 653972 765493 654028 765502
rect 653986 763305 654014 765493
rect 653974 763299 654026 763305
rect 653974 763241 654026 763247
rect 653972 742174 654028 742183
rect 653972 742109 654028 742118
rect 653986 740217 654014 742109
rect 653974 740211 654026 740217
rect 653974 740153 654026 740159
rect 655220 730482 655276 730491
rect 655220 730417 655276 730426
rect 654260 718642 654316 718651
rect 654260 718577 654316 718586
rect 654274 717203 654302 718577
rect 654262 717197 654314 717203
rect 654262 717139 654314 717145
rect 654452 695258 654508 695267
rect 654452 695193 654508 695202
rect 654466 694115 654494 695193
rect 654454 694109 654506 694115
rect 654454 694051 654506 694057
rect 655124 683566 655180 683575
rect 655124 683501 655180 683510
rect 654452 671726 654508 671735
rect 654452 671661 654508 671670
rect 654466 671101 654494 671661
rect 654454 671095 654506 671101
rect 654454 671037 654506 671043
rect 649940 660626 649996 660635
rect 649940 660561 649996 660570
rect 650038 659551 650090 659557
rect 650038 659493 650090 659499
rect 649942 613523 649994 613529
rect 649942 613465 649994 613471
rect 649846 236345 649898 236351
rect 649846 236287 649898 236293
rect 649954 236203 649982 613465
rect 649942 236197 649994 236203
rect 649942 236139 649994 236145
rect 645526 233237 645578 233243
rect 645526 233179 645578 233185
rect 649750 233237 649802 233243
rect 649750 233179 649802 233185
rect 645238 233163 645290 233169
rect 645238 233105 645290 233111
rect 645142 232941 645194 232947
rect 645142 232883 645194 232889
rect 645154 231583 645182 232883
rect 645140 231574 645196 231583
rect 645140 231509 645196 231518
rect 640726 73471 640778 73477
rect 640726 73413 640778 73419
rect 625942 52011 625994 52017
rect 625942 51953 625994 51959
rect 639670 52011 639722 52017
rect 639670 51953 639722 51959
rect 541366 51937 541418 51943
rect 558742 51937 558794 51943
rect 541418 51897 541502 51925
rect 541366 51879 541418 51885
rect 541474 51869 541502 51897
rect 558794 51897 558878 51925
rect 558742 51879 558794 51885
rect 541462 51863 541514 51869
rect 541462 51805 541514 51811
rect 558850 51795 558878 51897
rect 590338 51869 590462 51888
rect 590326 51863 590474 51869
rect 590378 51860 590422 51863
rect 590326 51805 590378 51811
rect 590422 51805 590474 51811
rect 558838 51789 558890 51795
rect 558838 51731 558890 51737
rect 604726 51715 604778 51721
rect 604726 51657 604778 51663
rect 538582 51641 538634 51647
rect 538580 51606 538582 51615
rect 541462 51641 541514 51647
rect 538634 51606 538636 51615
rect 538580 51541 538636 51550
rect 541460 51606 541462 51615
rect 584662 51641 584714 51647
rect 541514 51606 541516 51615
rect 541460 51541 541516 51550
rect 584660 51606 584662 51615
rect 604738 51615 604766 51657
rect 625954 51647 625982 51953
rect 625942 51641 625994 51647
rect 584714 51606 584716 51615
rect 584660 51541 584716 51550
rect 604724 51606 604780 51615
rect 625942 51583 625994 51589
rect 604724 51541 604780 51550
rect 529268 43318 529324 43327
rect 529268 43253 529324 43262
rect 520492 42092 520656 42120
rect 521506 42092 521856 42120
rect 525922 42092 526176 42120
rect 529282 42106 529310 43253
rect 520436 42069 520492 42078
rect 514870 42021 514922 42027
rect 514922 41969 515136 41972
rect 514870 41963 515136 41969
rect 514882 41944 515136 41963
rect 509684 41838 509740 41847
rect 509684 41773 509740 41782
rect 518516 41838 518572 41847
rect 518572 41796 518832 41824
rect 518516 41773 518572 41782
rect 459190 41577 459242 41583
rect 459190 41519 459242 41525
rect 459202 37439 459230 41519
rect 640738 40663 640766 73413
rect 645154 48909 645182 231509
rect 645250 231139 645278 233105
rect 645334 233015 645386 233021
rect 645334 232957 645386 232963
rect 645236 231130 645292 231139
rect 645236 231065 645292 231074
rect 645142 48903 645194 48909
rect 645142 48845 645194 48851
rect 645250 48835 645278 231065
rect 645346 230695 645374 232957
rect 645538 232027 645566 233179
rect 650050 232619 650078 659493
rect 654260 648342 654316 648351
rect 654260 648277 654316 648286
rect 654274 648087 654302 648277
rect 654262 648081 654314 648087
rect 654262 648023 654314 648029
rect 654356 624810 654412 624819
rect 654356 624745 654412 624754
rect 654370 622261 654398 624745
rect 654358 622255 654410 622261
rect 654358 622197 654410 622203
rect 654358 613449 654410 613455
rect 654358 613391 654410 613397
rect 654370 613127 654398 613391
rect 654356 613118 654412 613127
rect 654356 613053 654412 613062
rect 654452 601426 654508 601435
rect 654452 601361 654508 601370
rect 654466 599099 654494 601361
rect 654454 599093 654506 599099
rect 654454 599035 654506 599041
rect 654452 589586 654508 589595
rect 654452 589521 654508 589530
rect 654466 587555 654494 589521
rect 654454 587549 654506 587555
rect 654454 587491 654506 587497
rect 654452 577894 654508 577903
rect 654452 577829 654508 577838
rect 654466 576085 654494 577829
rect 654454 576079 654506 576085
rect 654454 576021 654506 576027
rect 650134 567421 650186 567427
rect 650134 567363 650186 567369
rect 650146 233021 650174 567363
rect 654454 567347 654506 567353
rect 654454 567289 654506 567295
rect 654466 566211 654494 567289
rect 654452 566202 654508 566211
rect 654452 566137 654508 566146
rect 654452 554510 654508 554519
rect 654452 554445 654508 554454
rect 654466 552997 654494 554445
rect 654454 552991 654506 552997
rect 654454 552933 654506 552939
rect 654452 542670 654508 542679
rect 654452 542605 654508 542614
rect 654466 541527 654494 542605
rect 654454 541521 654506 541527
rect 654454 541463 654506 541469
rect 655138 535829 655166 683501
rect 655234 582005 655262 730417
rect 660898 717647 660926 881271
rect 660994 762935 661022 915829
rect 663958 904417 664010 904423
rect 663958 904359 664010 904365
rect 663766 869859 663818 869865
rect 663766 869801 663818 869807
rect 661078 858315 661130 858321
rect 661078 858257 661130 858263
rect 660982 762929 661034 762935
rect 660982 762871 661034 762877
rect 660982 737325 661034 737331
rect 660982 737267 661034 737273
rect 660886 717641 660938 717647
rect 660886 717583 660938 717589
rect 655316 636650 655372 636659
rect 655316 636585 655372 636594
rect 655222 581999 655274 582005
rect 655222 581941 655274 581947
rect 655126 535823 655178 535829
rect 655126 535765 655178 535771
rect 654068 530978 654124 530987
rect 654068 530913 654124 530922
rect 654082 529983 654110 530913
rect 654070 529977 654122 529983
rect 654070 529919 654122 529925
rect 650230 524353 650282 524359
rect 650230 524295 650282 524301
rect 650242 236499 650270 524295
rect 654454 519321 654506 519327
rect 654452 519286 654454 519295
rect 654506 519286 654508 519295
rect 654452 519221 654508 519230
rect 654452 507446 654508 507455
rect 654452 507381 654508 507390
rect 654466 506969 654494 507381
rect 654454 506963 654506 506969
rect 654454 506905 654506 506911
rect 654356 495754 654412 495763
rect 654356 495689 654412 495698
rect 654370 495425 654398 495689
rect 654358 495419 654410 495425
rect 654358 495361 654410 495367
rect 655330 492539 655358 636585
rect 660886 555877 660938 555883
rect 660886 555819 660938 555825
rect 655318 492533 655370 492539
rect 655318 492475 655370 492481
rect 654260 484062 654316 484071
rect 654260 483997 654316 484006
rect 654274 483881 654302 483997
rect 654262 483875 654314 483881
rect 654262 483817 654314 483823
rect 650326 479509 650378 479515
rect 650326 479451 650378 479457
rect 650230 236493 650282 236499
rect 650230 236435 650282 236441
rect 650338 236425 650366 479451
rect 654454 472257 654506 472263
rect 654452 472222 654454 472231
rect 654506 472222 654508 472231
rect 654452 472157 654508 472166
rect 654452 460530 654508 460539
rect 654452 460465 654508 460474
rect 654466 457981 654494 460465
rect 654454 457975 654506 457981
rect 654454 457917 654506 457923
rect 654356 448838 654412 448847
rect 654356 448773 654412 448782
rect 654370 446437 654398 448773
rect 654358 446431 654410 446437
rect 654358 446373 654410 446379
rect 654452 436998 654508 437007
rect 654452 436933 654508 436942
rect 654466 434967 654494 436933
rect 654454 434961 654506 434967
rect 654454 434903 654506 434909
rect 654454 426229 654506 426235
rect 654454 426171 654506 426177
rect 654466 425463 654494 426171
rect 654452 425454 654508 425463
rect 654452 425389 654508 425398
rect 653876 413614 653932 413623
rect 653876 413549 653932 413558
rect 653890 411879 653918 413549
rect 653878 411873 653930 411879
rect 653878 411815 653930 411821
rect 654452 401774 654508 401783
rect 654452 401709 654508 401718
rect 654466 400409 654494 401709
rect 654454 400403 654506 400409
rect 654454 400345 654506 400351
rect 650422 391819 650474 391825
rect 650422 391761 650474 391767
rect 650326 236419 650378 236425
rect 650326 236361 650378 236367
rect 650434 233169 650462 391761
rect 654452 390082 654508 390091
rect 654452 390017 654508 390026
rect 654466 388865 654494 390017
rect 654454 388859 654506 388865
rect 654454 388801 654506 388807
rect 654454 380127 654506 380133
rect 654454 380069 654506 380075
rect 654466 378547 654494 380069
rect 654452 378538 654508 378547
rect 654452 378473 654508 378482
rect 654452 366550 654508 366559
rect 654452 366485 654508 366494
rect 654466 365851 654494 366485
rect 654454 365845 654506 365851
rect 654454 365787 654506 365793
rect 655220 354858 655276 354867
rect 655220 354793 655276 354802
rect 650518 345643 650570 345649
rect 650518 345585 650570 345591
rect 650530 236573 650558 345585
rect 654452 343166 654508 343175
rect 654452 343101 654508 343110
rect 654466 342763 654494 343101
rect 654454 342757 654506 342763
rect 654454 342699 654506 342705
rect 654454 332323 654506 332329
rect 654454 332265 654506 332271
rect 654466 331631 654494 332265
rect 654452 331622 654508 331631
rect 654452 331557 654508 331566
rect 655124 319782 655180 319791
rect 655124 319717 655180 319726
rect 650614 302649 650666 302655
rect 650614 302591 650666 302597
rect 650518 236567 650570 236573
rect 650518 236509 650570 236515
rect 650422 233163 650474 233169
rect 650422 233105 650474 233111
rect 650134 233015 650186 233021
rect 650134 232957 650186 232963
rect 650626 232947 650654 302591
rect 654548 296250 654604 296259
rect 654548 296185 654604 296194
rect 654562 293849 654590 296185
rect 654550 293843 654602 293849
rect 654550 293785 654602 293791
rect 654070 284815 654122 284821
rect 654070 284757 654122 284763
rect 654082 284715 654110 284757
rect 654068 284706 654124 284715
rect 654068 284641 654124 284650
rect 650614 232941 650666 232947
rect 650614 232883 650666 232889
rect 646292 232610 646348 232619
rect 646292 232545 646348 232554
rect 650036 232610 650092 232619
rect 650036 232545 650092 232554
rect 645524 232018 645580 232027
rect 645524 231953 645580 231962
rect 645332 230686 645388 230695
rect 645332 230621 645388 230630
rect 645238 48829 645290 48835
rect 645238 48771 645290 48777
rect 645346 48761 645374 230621
rect 645430 121201 645482 121207
rect 645428 121166 645430 121175
rect 645482 121166 645484 121175
rect 645428 121101 645484 121110
rect 645430 104551 645482 104557
rect 645430 104493 645482 104499
rect 645442 104303 645470 104493
rect 645428 104294 645484 104303
rect 645428 104229 645484 104238
rect 645428 87718 645484 87727
rect 645428 87653 645484 87662
rect 645442 87093 645470 87653
rect 645430 87087 645482 87093
rect 645430 87029 645482 87035
rect 645428 86682 645484 86691
rect 645428 86617 645484 86626
rect 645442 86501 645470 86617
rect 645430 86495 645482 86501
rect 645430 86437 645482 86443
rect 645538 51795 645566 231953
rect 646306 221815 646334 232545
rect 646100 221806 646156 221815
rect 646100 221741 646156 221750
rect 646292 221806 646348 221815
rect 646292 221741 646348 221750
rect 645620 210410 645676 210419
rect 645620 210345 645676 210354
rect 645634 210303 645662 210345
rect 645622 210297 645674 210303
rect 645622 210239 645674 210245
rect 645526 51789 645578 51795
rect 645526 51731 645578 51737
rect 645334 48755 645386 48761
rect 645334 48697 645386 48703
rect 645634 47651 645662 210239
rect 646114 201645 646142 221741
rect 645910 201639 645962 201645
rect 645910 201581 645962 201587
rect 646102 201639 646154 201645
rect 646102 201581 646154 201587
rect 645922 198727 645950 201581
rect 645908 198718 645964 198727
rect 645908 198653 645964 198662
rect 646100 198718 646156 198727
rect 646100 198653 646156 198662
rect 646114 187141 646142 198653
rect 645718 187135 645770 187141
rect 645718 187077 645770 187083
rect 646102 187135 646154 187141
rect 646102 187077 646154 187083
rect 645730 161315 645758 187077
rect 647062 167303 647114 167309
rect 647062 167245 647114 167251
rect 647074 166315 647102 167245
rect 647830 167229 647882 167235
rect 647830 167171 647882 167177
rect 647060 166306 647116 166315
rect 647060 166241 647116 166250
rect 647842 166019 647870 167171
rect 647926 167155 647978 167161
rect 647926 167097 647978 167103
rect 647938 167055 647966 167097
rect 647924 167046 647980 167055
rect 647924 166981 647980 166990
rect 647828 166010 647884 166019
rect 647828 165945 647884 165954
rect 645718 161309 645770 161315
rect 645716 161274 645718 161283
rect 645910 161309 645962 161315
rect 645770 161274 645772 161283
rect 645716 161209 645772 161218
rect 645908 161274 645910 161283
rect 645962 161274 645964 161283
rect 645908 161209 645964 161218
rect 645730 146959 645758 161209
rect 645718 146953 645770 146959
rect 645718 146895 645770 146901
rect 645814 146879 645866 146885
rect 645814 146821 645866 146827
rect 645826 126776 645854 146821
rect 655138 132677 655166 319717
rect 655234 178705 655262 354793
rect 655316 307942 655372 307951
rect 655316 307877 655372 307886
rect 655222 178699 655274 178705
rect 655222 178641 655274 178647
rect 655330 132825 655358 307877
rect 660898 284821 660926 555819
rect 660994 472263 661022 737267
rect 661090 717055 661118 858257
rect 661174 763299 661226 763305
rect 661174 763241 661226 763247
rect 661078 717049 661130 717055
rect 661078 716991 661130 716997
rect 661078 671095 661130 671101
rect 661078 671037 661130 671043
rect 661090 536643 661118 671037
rect 661186 626627 661214 763241
rect 663778 718091 663806 869801
rect 663862 780541 663914 780547
rect 663862 780483 663914 780489
rect 663766 718085 663818 718091
rect 663766 718027 663818 718033
rect 661174 626621 661226 626627
rect 661174 626563 661226 626569
rect 663766 601979 663818 601985
rect 663766 601921 663818 601927
rect 661078 536637 661130 536643
rect 661078 536579 661130 536585
rect 661174 495419 661226 495425
rect 661174 495361 661226 495367
rect 660982 472257 661034 472263
rect 660982 472199 661034 472205
rect 660982 457975 661034 457981
rect 660982 457917 661034 457923
rect 660886 284815 660938 284821
rect 660886 284757 660938 284763
rect 660994 269799 661022 457917
rect 661078 365845 661130 365851
rect 661078 365787 661130 365793
rect 660982 269793 661034 269799
rect 660982 269735 661034 269741
rect 661090 179371 661118 365787
rect 661186 315087 661214 495361
rect 663778 332329 663806 601921
rect 663874 519327 663902 780483
rect 663970 762047 663998 904359
rect 666646 865345 666698 865351
rect 666646 865287 666698 865293
rect 664054 812213 664106 812219
rect 664054 812155 664106 812161
rect 663958 762041 664010 762047
rect 663958 761983 664010 761989
rect 663958 740211 664010 740217
rect 663958 740153 664010 740159
rect 663970 582079 663998 740153
rect 664066 671915 664094 812155
rect 664054 671909 664106 671915
rect 664054 671851 664106 671857
rect 664054 648081 664106 648087
rect 664054 648023 664106 648029
rect 663958 582073 664010 582079
rect 663958 582015 664010 582021
rect 663862 519321 663914 519327
rect 663862 519263 663914 519269
rect 663862 506963 663914 506969
rect 663862 506905 663914 506911
rect 663766 332323 663818 332329
rect 663766 332265 663818 332271
rect 661174 315081 661226 315087
rect 661174 315023 661226 315029
rect 663874 314791 663902 506905
rect 664066 493279 664094 648023
rect 666658 567353 666686 865287
rect 666754 762343 666782 927447
rect 666838 835227 666890 835233
rect 666838 835169 666890 835175
rect 666742 762337 666794 762343
rect 666742 762279 666794 762285
rect 666850 672359 666878 835169
rect 666934 717197 666986 717203
rect 666934 717139 666986 717145
rect 666838 672353 666890 672359
rect 666838 672295 666890 672301
rect 666742 641125 666794 641131
rect 666742 641067 666794 641073
rect 666646 567347 666698 567353
rect 666646 567289 666698 567295
rect 666646 552991 666698 552997
rect 666646 552933 666698 552939
rect 664054 493273 664106 493279
rect 664054 493215 664106 493221
rect 663958 434961 664010 434967
rect 663958 434903 664010 434909
rect 663862 314785 663914 314791
rect 663862 314727 663914 314733
rect 663766 293843 663818 293849
rect 663766 293785 663818 293791
rect 661078 179365 661130 179371
rect 661078 179307 661130 179313
rect 663778 133639 663806 293785
rect 663970 269207 663998 434903
rect 666658 359783 666686 552933
rect 666754 380133 666782 641067
rect 666838 587549 666890 587555
rect 666838 587491 666890 587497
rect 666850 405515 666878 587491
rect 666946 581635 666974 717139
rect 669538 613455 669566 954679
rect 674134 953997 674186 954003
rect 674134 953939 674186 953945
rect 674038 952073 674090 952079
rect 674038 952015 674090 952021
rect 673844 939162 673900 939171
rect 673844 939097 673900 939106
rect 673366 872153 673418 872159
rect 673366 872095 673418 872101
rect 673270 869193 673322 869199
rect 673270 869135 673322 869141
rect 673174 867861 673226 867867
rect 673174 867803 673226 867809
rect 669910 823757 669962 823763
rect 669910 823699 669962 823705
rect 669718 786313 669770 786319
rect 669718 786255 669770 786261
rect 669622 686265 669674 686271
rect 669622 686207 669674 686213
rect 669526 613449 669578 613455
rect 669526 613391 669578 613397
rect 666934 581629 666986 581635
rect 666934 581571 666986 581577
rect 666934 483875 666986 483881
rect 666934 483817 666986 483823
rect 666838 405509 666890 405515
rect 666838 405451 666890 405457
rect 666838 400403 666890 400409
rect 666838 400345 666890 400351
rect 666742 380127 666794 380133
rect 666742 380069 666794 380075
rect 666646 359777 666698 359783
rect 666646 359719 666698 359725
rect 666646 342757 666698 342763
rect 666646 342699 666698 342705
rect 663958 269201 664010 269207
rect 663958 269143 664010 269149
rect 666658 178853 666686 342699
rect 666850 225103 666878 400345
rect 666946 314051 666974 483817
rect 669634 426235 669662 686207
rect 669730 627367 669758 786255
rect 669814 694109 669866 694115
rect 669814 694051 669866 694057
rect 669718 627361 669770 627367
rect 669718 627303 669770 627309
rect 669718 541521 669770 541527
rect 669718 541463 669770 541469
rect 669622 426229 669674 426235
rect 669622 426171 669674 426177
rect 669526 411873 669578 411879
rect 669526 411815 669578 411821
rect 666934 314045 666986 314051
rect 666934 313987 666986 313993
rect 666838 225097 666890 225103
rect 666838 225039 666890 225045
rect 669538 224363 669566 411815
rect 669622 388859 669674 388865
rect 669622 388801 669674 388807
rect 669526 224357 669578 224363
rect 669526 224299 669578 224305
rect 669634 224067 669662 388801
rect 669730 360079 669758 541463
rect 669826 537235 669854 694051
rect 669922 672951 669950 823699
rect 672310 783501 672362 783507
rect 672310 783443 672362 783449
rect 672214 779357 672266 779363
rect 672214 779299 672266 779305
rect 672226 708693 672254 779299
rect 672322 709951 672350 783443
rect 672886 783131 672938 783137
rect 672886 783073 672938 783079
rect 672502 782539 672554 782545
rect 672502 782481 672554 782487
rect 672406 774769 672458 774775
rect 672406 774711 672458 774717
rect 672310 709945 672362 709951
rect 672310 709887 672362 709893
rect 672214 708687 672266 708693
rect 672214 708629 672266 708635
rect 672310 692925 672362 692931
rect 672310 692867 672362 692873
rect 669910 672945 669962 672951
rect 669910 672887 669962 672893
rect 670966 625511 671018 625517
rect 670966 625453 671018 625459
rect 670978 580895 671006 625453
rect 671926 622181 671978 622187
rect 671926 622123 671978 622129
rect 671830 604125 671882 604131
rect 671830 604067 671882 604073
rect 670966 580889 671018 580895
rect 670966 580831 671018 580837
rect 669910 576079 669962 576085
rect 669910 576021 669962 576027
rect 669814 537229 669866 537235
rect 669814 537171 669866 537177
rect 669814 446431 669866 446437
rect 669814 446373 669866 446379
rect 669718 360073 669770 360079
rect 669718 360015 669770 360021
rect 669826 270095 669854 446373
rect 669922 404479 669950 576021
rect 671842 529909 671870 604067
rect 671938 587555 671966 622123
rect 672022 622107 672074 622113
rect 672022 622049 672074 622055
rect 671926 587549 671978 587555
rect 671926 587491 671978 587497
rect 672034 579827 672062 622049
rect 672322 617895 672350 692867
rect 672418 627737 672446 774711
rect 672514 740217 672542 782481
rect 672694 777655 672746 777661
rect 672694 777597 672746 777603
rect 672502 740211 672554 740217
rect 672502 740153 672554 740159
rect 672598 732367 672650 732373
rect 672598 732309 672650 732315
rect 672610 664219 672638 732309
rect 672706 709211 672734 777597
rect 672898 745989 672926 783073
rect 673078 779801 673130 779807
rect 673078 779743 673130 779749
rect 672982 778617 673034 778623
rect 672982 778559 673034 778565
rect 672886 745983 672938 745989
rect 672886 745925 672938 745931
rect 672790 734439 672842 734445
rect 672790 734381 672842 734387
rect 672694 709205 672746 709211
rect 672694 709147 672746 709153
rect 672694 699881 672746 699887
rect 672694 699823 672746 699829
rect 672706 693005 672734 699823
rect 672694 692999 672746 693005
rect 672694 692941 672746 692947
rect 672598 664213 672650 664219
rect 672598 664155 672650 664161
rect 672706 653785 672734 692941
rect 672802 665255 672830 734381
rect 672886 733625 672938 733631
rect 672886 733567 672938 733573
rect 672790 665249 672842 665255
rect 672790 665191 672842 665197
rect 672898 662369 672926 733567
rect 672994 707065 673022 778559
rect 673090 707551 673118 779743
rect 673186 752099 673214 867803
rect 673282 752543 673310 869135
rect 673378 753135 673406 872095
rect 673462 782983 673514 782989
rect 673462 782925 673514 782931
rect 673364 753126 673420 753135
rect 673364 753061 673420 753070
rect 673268 752534 673324 752543
rect 673268 752469 673324 752478
rect 673172 752090 673228 752099
rect 673172 752025 673228 752034
rect 673174 738139 673226 738145
rect 673174 738081 673226 738087
rect 673076 707542 673132 707551
rect 673076 707477 673132 707486
rect 672982 707059 673034 707065
rect 672982 707001 673034 707007
rect 673186 699887 673214 738081
rect 673366 737917 673418 737923
rect 673366 737859 673418 737865
rect 673270 734809 673322 734815
rect 673270 734751 673322 734757
rect 673174 699881 673226 699887
rect 673174 699823 673226 699829
rect 673078 689817 673130 689823
rect 673078 689759 673130 689765
rect 672982 689373 673034 689379
rect 672982 689315 673034 689321
rect 672886 662363 672938 662369
rect 672886 662305 672938 662311
rect 672694 653779 672746 653785
rect 672694 653721 672746 653727
rect 672790 644603 672842 644609
rect 672790 644545 672842 644551
rect 672502 644085 672554 644091
rect 672502 644027 672554 644033
rect 672406 627731 672458 627737
rect 672406 627673 672458 627679
rect 672310 617889 672362 617895
rect 672310 617831 672362 617837
rect 672118 602867 672170 602873
rect 672118 602809 672170 602815
rect 672020 579818 672076 579827
rect 672020 579753 672076 579762
rect 671926 579187 671978 579193
rect 671926 579129 671978 579135
rect 671938 536199 671966 579129
rect 672130 564393 672158 602809
rect 672310 602497 672362 602503
rect 672310 602439 672362 602445
rect 672214 597169 672266 597175
rect 672214 597111 672266 597117
rect 672118 564387 672170 564393
rect 672118 564329 672170 564335
rect 671926 536193 671978 536199
rect 671926 536135 671978 536141
rect 671830 529903 671882 529909
rect 671830 529845 671882 529851
rect 672226 529095 672254 597111
rect 672322 564467 672350 602439
rect 672406 599093 672458 599099
rect 672406 599035 672458 599041
rect 672310 564461 672362 564467
rect 672310 564403 672362 564409
rect 672214 529089 672266 529095
rect 672214 529031 672266 529037
rect 672418 406107 672446 599035
rect 672514 573643 672542 644027
rect 672694 642309 672746 642315
rect 672694 642251 672746 642257
rect 672598 622255 672650 622261
rect 672598 622197 672650 622203
rect 672502 573637 672554 573643
rect 672502 573579 672554 573585
rect 672502 529977 672554 529983
rect 672502 529919 672554 529925
rect 672406 406101 672458 406107
rect 672406 406043 672458 406049
rect 669910 404473 669962 404479
rect 669910 404415 669962 404421
rect 672514 359043 672542 529919
rect 672610 492465 672638 622197
rect 672706 576011 672734 642251
rect 672694 576005 672746 576011
rect 672694 575947 672746 575953
rect 672802 573125 672830 644545
rect 672886 643419 672938 643425
rect 672886 643361 672938 643367
rect 672790 573119 672842 573125
rect 672790 573061 672842 573067
rect 672898 571645 672926 643361
rect 672994 618487 673022 689315
rect 672982 618481 673034 618487
rect 672982 618423 673034 618429
rect 673090 617599 673118 689759
rect 673174 688633 673226 688639
rect 673174 688575 673226 688581
rect 673078 617593 673130 617599
rect 673078 617535 673130 617541
rect 673186 616827 673214 688575
rect 673282 662411 673310 734751
rect 673378 662855 673406 737859
rect 673474 708143 673502 782925
rect 673858 761275 673886 939097
rect 674050 934731 674078 952015
rect 674146 938981 674174 953939
rect 674914 953527 674942 960728
rect 675476 960705 675532 960714
rect 675106 960545 675408 960573
rect 675106 959299 675134 960545
rect 675092 959290 675148 959299
rect 675092 959225 675148 959234
rect 675490 959151 675518 959262
rect 675476 959142 675532 959151
rect 675476 959077 675532 959086
rect 675778 958411 675806 958744
rect 675764 958402 675820 958411
rect 675764 958337 675820 958346
rect 675394 957671 675422 958078
rect 675380 957662 675436 957671
rect 675380 957597 675436 957606
rect 675490 957037 675518 957412
rect 675190 957031 675242 957037
rect 675190 956973 675242 956979
rect 675478 957031 675530 957037
rect 675478 956973 675530 956979
rect 674900 953518 674956 953527
rect 674900 953453 674956 953462
rect 675202 953379 675230 956973
rect 675490 956043 675518 956228
rect 675476 956034 675532 956043
rect 675476 955969 675532 955978
rect 675394 954743 675422 955044
rect 675382 954737 675434 954743
rect 675382 954679 675434 954685
rect 675490 954003 675518 954378
rect 675478 953997 675530 954003
rect 675478 953939 675530 953945
rect 675188 953370 675244 953379
rect 675188 953305 675244 953314
rect 675490 952079 675518 952528
rect 675478 952073 675530 952079
rect 675478 952015 675530 952021
rect 676820 940938 676876 940947
rect 676820 940873 676876 940882
rect 674516 939902 674572 939911
rect 674516 939837 674572 939846
rect 674420 939606 674476 939615
rect 674420 939541 674422 939550
rect 674474 939541 674476 939550
rect 674422 939509 674474 939515
rect 674530 939425 674558 939837
rect 674518 939419 674570 939425
rect 674518 939361 674570 939367
rect 676834 939277 676862 940873
rect 676916 940494 676972 940503
rect 676916 940429 676972 940438
rect 676822 939271 676874 939277
rect 676822 939213 676874 939219
rect 676930 939129 676958 940429
rect 676918 939123 676970 939129
rect 676918 939065 676970 939071
rect 674134 938975 674186 938981
rect 674134 938917 674186 938923
rect 676918 938975 676970 938981
rect 676918 938917 676970 938923
rect 676820 938274 676876 938283
rect 676820 938209 676876 938218
rect 674422 938013 674474 938019
rect 674420 937978 674422 937987
rect 674474 937978 674476 937987
rect 674420 937913 674476 937922
rect 676834 936317 676862 938209
rect 676930 937247 676958 938917
rect 676916 937238 676972 937247
rect 676916 937173 676972 937182
rect 676822 936311 676874 936317
rect 676822 936253 676874 936259
rect 674036 934722 674092 934731
rect 674036 934657 674092 934666
rect 677012 929542 677068 929551
rect 677012 929477 677068 929486
rect 676820 928950 676876 928959
rect 676820 928885 676876 928894
rect 676834 928515 676862 928885
rect 677026 928515 677054 929477
rect 676820 928506 676876 928515
rect 676820 928441 676876 928450
rect 677012 928506 677068 928515
rect 677012 928441 677068 928450
rect 677026 927437 677054 928441
rect 677014 927431 677066 927437
rect 677014 927373 677066 927379
rect 675394 877011 675422 877523
rect 675380 877002 675436 877011
rect 675380 876937 675436 876946
rect 675778 876567 675806 876900
rect 675764 876558 675820 876567
rect 675764 876493 675820 876502
rect 675490 875827 675518 876234
rect 675092 875818 675148 875827
rect 675092 875753 675148 875762
rect 675476 875818 675532 875827
rect 675476 875753 675532 875762
rect 674614 872671 674666 872677
rect 674614 872613 674666 872619
rect 674230 871709 674282 871715
rect 674230 871651 674282 871657
rect 674242 789205 674270 871651
rect 674326 868379 674378 868385
rect 674326 868321 674378 868327
rect 674230 789199 674282 789205
rect 674230 789141 674282 789147
rect 674338 772967 674366 868321
rect 674518 862977 674570 862983
rect 674518 862919 674570 862925
rect 674530 775631 674558 862919
rect 674516 775622 674572 775631
rect 674516 775557 674572 775566
rect 674324 772958 674380 772967
rect 674324 772893 674380 772902
rect 674626 772671 674654 872613
rect 675106 871715 675134 875753
rect 675188 875670 675244 875679
rect 675188 875605 675244 875614
rect 675094 871709 675146 871715
rect 675094 871651 675146 871657
rect 675202 871493 675230 875605
rect 675490 874051 675518 874384
rect 675476 874042 675532 874051
rect 675476 873977 675532 873986
rect 675394 873607 675422 873866
rect 675380 873598 675436 873607
rect 675380 873533 675436 873542
rect 675394 872677 675422 873200
rect 675382 872671 675434 872677
rect 675382 872613 675434 872619
rect 675490 872159 675518 872534
rect 675478 872153 675530 872159
rect 675478 872095 675530 872101
rect 675394 871715 675422 872016
rect 675382 871709 675434 871715
rect 675382 871651 675434 871657
rect 674902 871487 674954 871493
rect 674902 871429 674954 871435
rect 675190 871487 675242 871493
rect 675190 871429 675242 871435
rect 675382 871487 675434 871493
rect 675382 871429 675434 871435
rect 674914 855657 674942 871429
rect 675394 871350 675422 871429
rect 675394 869907 675422 870092
rect 675380 869898 675436 869907
rect 675380 869833 675436 869842
rect 675490 869199 675518 869500
rect 675478 869193 675530 869199
rect 675478 869135 675530 869141
rect 675394 868385 675422 868875
rect 675382 868379 675434 868385
rect 675382 868321 675434 868327
rect 675394 867867 675422 868242
rect 675382 867861 675434 867867
rect 675382 867803 675434 867809
rect 675394 866535 675422 867058
rect 675094 866529 675146 866535
rect 675094 866471 675146 866477
rect 675382 866529 675434 866535
rect 675382 866471 675434 866477
rect 675106 855805 675134 866471
rect 675394 865351 675422 865839
rect 675382 865345 675434 865351
rect 675382 865287 675434 865293
rect 675490 864727 675518 865208
rect 675476 864718 675532 864727
rect 675476 864653 675532 864662
rect 675394 862983 675422 863358
rect 675382 862977 675434 862983
rect 675382 862919 675434 862925
rect 675094 855799 675146 855805
rect 675094 855741 675146 855747
rect 675478 855799 675530 855805
rect 675478 855741 675530 855747
rect 674902 855651 674954 855657
rect 674902 855593 674954 855599
rect 675490 790611 675518 855741
rect 675574 855651 675626 855657
rect 675574 855593 675626 855599
rect 674710 790605 674762 790611
rect 674710 790547 674762 790553
rect 675478 790605 675530 790611
rect 675478 790547 675530 790553
rect 674722 775039 674750 790547
rect 675586 789279 675614 855593
rect 674998 789273 675050 789279
rect 674998 789215 675050 789221
rect 675574 789273 675626 789279
rect 675574 789215 675626 789221
rect 675010 782545 675038 789215
rect 675094 789199 675146 789205
rect 675094 789141 675146 789147
rect 675106 783137 675134 789141
rect 675394 788063 675422 788322
rect 675380 788054 675436 788063
rect 675380 787989 675436 787998
rect 675490 787175 675518 787656
rect 675476 787166 675532 787175
rect 675476 787101 675532 787110
rect 675778 786731 675806 787035
rect 675764 786722 675820 786731
rect 675764 786657 675820 786666
rect 675778 784955 675806 785214
rect 675764 784946 675820 784955
rect 675764 784881 675820 784890
rect 675682 784215 675710 784622
rect 675668 784206 675724 784215
rect 675668 784141 675724 784150
rect 675394 783507 675422 783999
rect 675382 783501 675434 783507
rect 675382 783443 675434 783449
rect 675094 783131 675146 783137
rect 675094 783073 675146 783079
rect 675394 782989 675422 783364
rect 675478 783131 675530 783137
rect 675478 783073 675530 783079
rect 675382 782983 675434 782989
rect 675382 782925 675434 782931
rect 675490 782803 675518 783073
rect 674998 782539 675050 782545
rect 674998 782481 675050 782487
rect 675478 782539 675530 782545
rect 675478 782481 675530 782487
rect 675490 782180 675518 782481
rect 675778 780663 675806 780848
rect 675764 780654 675820 780663
rect 675764 780589 675820 780598
rect 675094 780541 675146 780547
rect 675094 780483 675146 780489
rect 675106 777069 675134 780483
rect 675394 779807 675422 780330
rect 675382 779801 675434 779807
rect 675382 779743 675434 779749
rect 675490 779363 675518 779664
rect 675478 779357 675530 779363
rect 675478 779299 675530 779305
rect 675394 778623 675422 779031
rect 675382 778617 675434 778623
rect 675382 778559 675434 778565
rect 675490 777661 675518 777814
rect 675478 777655 675530 777661
rect 675478 777597 675530 777603
rect 675094 777063 675146 777069
rect 675094 777005 675146 777011
rect 675382 777063 675434 777069
rect 675382 777005 675434 777011
rect 675394 776630 675422 777005
rect 675394 775483 675422 775995
rect 675380 775474 675436 775483
rect 675380 775409 675436 775418
rect 674708 775030 674764 775039
rect 674708 774965 674764 774974
rect 675778 773707 675806 774155
rect 675764 773698 675820 773707
rect 675764 773633 675820 773642
rect 676628 773106 676684 773115
rect 676628 773041 676684 773050
rect 674612 772662 674668 772671
rect 674612 772597 674668 772606
rect 674422 762929 674474 762935
rect 674420 762894 674422 762903
rect 674474 762894 674476 762903
rect 674420 762829 674476 762838
rect 674422 762337 674474 762343
rect 674420 762302 674422 762311
rect 674474 762302 674476 762311
rect 674420 762237 674476 762246
rect 674614 762041 674666 762047
rect 674612 762006 674614 762015
rect 674666 762006 674668 762015
rect 674612 761941 674668 761950
rect 673844 761266 673900 761275
rect 673844 761201 673900 761210
rect 673844 760674 673900 760683
rect 673844 760609 673900 760618
rect 673858 716283 673886 760609
rect 676642 758315 676670 773041
rect 677780 764670 677836 764679
rect 677780 764605 677836 764614
rect 676628 758306 676684 758315
rect 676628 758241 676684 758250
rect 677794 754467 677822 764605
rect 677780 754458 677836 754467
rect 677780 754393 677836 754402
rect 677012 751202 677068 751211
rect 677012 751137 677068 751146
rect 677026 750619 677054 751137
rect 676820 750610 676876 750619
rect 676820 750545 676876 750554
rect 677012 750610 677068 750619
rect 677012 750545 677068 750554
rect 676834 750175 676862 750545
rect 676820 750166 676876 750175
rect 676820 750101 676876 750110
rect 677026 748875 677054 750545
rect 677014 748869 677066 748875
rect 677014 748811 677066 748817
rect 675094 745983 675146 745989
rect 675094 745925 675146 745931
rect 674710 740211 674762 740217
rect 674710 740153 674762 740159
rect 674722 737701 674750 740153
rect 675106 738145 675134 745925
rect 675394 743219 675422 743330
rect 675380 743210 675436 743219
rect 675380 743145 675436 743154
rect 675490 742183 675518 742664
rect 675476 742174 675532 742183
rect 675476 742109 675532 742118
rect 675778 741739 675806 742035
rect 675764 741730 675820 741739
rect 675764 741665 675820 741674
rect 675394 740111 675422 740222
rect 675380 740102 675436 740111
rect 675380 740037 675436 740046
rect 675490 739223 675518 739630
rect 675476 739214 675532 739223
rect 675476 739149 675532 739158
rect 675394 738631 675422 738999
rect 675380 738622 675436 738631
rect 675380 738557 675436 738566
rect 675094 738139 675146 738145
rect 675094 738081 675146 738087
rect 675394 737923 675422 738372
rect 675478 738139 675530 738145
rect 675478 738081 675530 738087
rect 675382 737917 675434 737923
rect 675382 737859 675434 737865
rect 675490 737780 675518 738081
rect 674710 737695 674762 737701
rect 674710 737637 674762 737643
rect 675382 737695 675434 737701
rect 675382 737637 675434 737643
rect 674722 737572 674750 737637
rect 674434 737544 674750 737572
rect 674038 728667 674090 728673
rect 674038 728609 674090 728615
rect 673844 716274 673900 716283
rect 673844 716209 673900 716218
rect 673844 715682 673900 715691
rect 673844 715617 673900 715626
rect 673460 708134 673516 708143
rect 673460 708069 673516 708078
rect 673858 671143 673886 715617
rect 674050 685624 674078 728609
rect 674326 711351 674378 711357
rect 674326 711293 674378 711299
rect 674050 685596 674270 685624
rect 673942 685525 673994 685531
rect 673942 685467 673994 685473
rect 673844 671134 673900 671143
rect 673844 671069 673900 671078
rect 673846 665249 673898 665255
rect 673846 665191 673898 665197
rect 673858 663447 673886 665191
rect 673844 663438 673900 663447
rect 673844 663373 673900 663382
rect 673364 662846 673420 662855
rect 673364 662781 673420 662790
rect 673268 662402 673324 662411
rect 673268 662337 673324 662346
rect 673846 662363 673898 662369
rect 673846 662305 673898 662311
rect 673858 661819 673886 662305
rect 673844 661810 673900 661819
rect 673844 661745 673900 661754
rect 673270 648303 673322 648309
rect 673270 648245 673322 648251
rect 673172 616818 673228 616827
rect 673172 616753 673228 616762
rect 673078 599833 673130 599839
rect 673078 599775 673130 599781
rect 672982 599315 673034 599321
rect 672982 599257 673034 599263
rect 672886 571639 672938 571645
rect 672886 571581 672938 571587
rect 672886 553213 672938 553219
rect 672886 553155 672938 553161
rect 672598 492459 672650 492465
rect 672598 492401 672650 492407
rect 672898 483807 672926 553155
rect 672994 528503 673022 599257
rect 672982 528497 673034 528503
rect 672982 528439 673034 528445
rect 673090 527139 673118 599775
rect 673174 598427 673226 598433
rect 673174 598369 673226 598375
rect 673076 527130 673132 527139
rect 673076 527065 673132 527074
rect 673186 526695 673214 598369
rect 673282 574351 673310 648245
rect 673750 648081 673802 648087
rect 673750 648023 673802 648029
rect 673366 647119 673418 647125
rect 673366 647061 673418 647067
rect 673378 613455 673406 647061
rect 673366 613449 673418 613455
rect 673366 613391 673418 613397
rect 673558 603311 673610 603317
rect 673558 603253 673610 603259
rect 673366 602719 673418 602725
rect 673366 602661 673418 602667
rect 673268 574342 673324 574351
rect 673268 574277 673324 574286
rect 673270 553805 673322 553811
rect 673270 553747 673322 553753
rect 673172 526686 673228 526695
rect 673172 526621 673228 526630
rect 673282 484219 673310 553747
rect 673378 527731 673406 602661
rect 673570 529359 673598 603253
rect 673762 572723 673790 648023
rect 673954 642283 673982 685467
rect 674242 666185 674270 685596
rect 674338 671027 674366 711293
rect 674434 709359 674462 737544
rect 675094 737325 675146 737331
rect 675094 737267 675146 737273
rect 674614 735475 674666 735481
rect 674614 735417 674666 735423
rect 674626 731559 674654 735417
rect 675106 732077 675134 737267
rect 675394 737159 675422 737637
rect 675490 735481 675518 735856
rect 675478 735475 675530 735481
rect 675478 735417 675530 735423
rect 675394 734815 675422 735338
rect 675382 734809 675434 734815
rect 675382 734751 675434 734757
rect 675394 734445 675422 734672
rect 675382 734439 675434 734445
rect 675382 734381 675434 734387
rect 675490 733631 675518 734006
rect 675478 733625 675530 733631
rect 675478 733567 675530 733573
rect 675490 732373 675518 732822
rect 675478 732367 675530 732373
rect 675478 732309 675530 732315
rect 675094 732071 675146 732077
rect 675094 732013 675146 732019
rect 675382 732071 675434 732077
rect 675382 732013 675434 732019
rect 675394 731638 675422 732013
rect 674614 731553 674666 731559
rect 674614 731495 674666 731501
rect 674806 731553 674858 731559
rect 674806 731495 674858 731501
rect 674518 730517 674570 730523
rect 674518 730459 674570 730465
rect 674530 711357 674558 730459
rect 674614 718085 674666 718091
rect 674612 718050 674614 718059
rect 674666 718050 674668 718059
rect 674612 717985 674668 717994
rect 674614 717641 674666 717647
rect 674612 717606 674614 717615
rect 674666 717606 674668 717615
rect 674612 717541 674668 717550
rect 674614 717049 674666 717055
rect 674612 717014 674614 717023
rect 674666 717014 674668 717023
rect 674612 716949 674668 716958
rect 674818 715723 674846 731495
rect 675490 730523 675518 730972
rect 675478 730517 675530 730523
rect 675478 730459 675530 730465
rect 675490 728673 675518 729155
rect 675478 728667 675530 728673
rect 675478 728609 675530 728615
rect 674614 715717 674666 715723
rect 674614 715659 674666 715665
rect 674806 715717 674858 715723
rect 674806 715659 674858 715665
rect 674518 711351 674570 711357
rect 674626 711339 674654 715659
rect 677108 714794 677164 714803
rect 677108 714729 677164 714738
rect 674626 711311 674750 711339
rect 674518 711293 674570 711299
rect 674614 709945 674666 709951
rect 674612 709910 674614 709919
rect 674666 709910 674668 709919
rect 674612 709845 674668 709854
rect 674422 709353 674474 709359
rect 674422 709295 674474 709301
rect 674614 709353 674666 709359
rect 674614 709295 674666 709301
rect 674422 709205 674474 709211
rect 674420 709170 674422 709179
rect 674474 709170 674476 709179
rect 674420 709105 674476 709114
rect 674422 708687 674474 708693
rect 674420 708652 674422 708661
rect 674474 708652 674476 708661
rect 674420 708587 674476 708596
rect 674422 707059 674474 707065
rect 674420 707024 674422 707033
rect 674474 707024 674476 707033
rect 674420 706959 674476 706968
rect 674626 692709 674654 709295
rect 674722 705659 674750 711311
rect 677012 706210 677068 706219
rect 677012 706145 677068 706154
rect 674710 705653 674762 705659
rect 674710 705595 674762 705601
rect 674998 705653 675050 705659
rect 677026 705627 677054 706145
rect 677122 705775 677150 714729
rect 677108 705766 677164 705775
rect 677108 705701 677164 705710
rect 674998 705595 675050 705601
rect 676820 705618 676876 705627
rect 674614 692703 674666 692709
rect 674614 692645 674666 692651
rect 675010 692580 675038 705595
rect 676820 705553 676876 705562
rect 677012 705618 677068 705627
rect 677012 705553 677068 705562
rect 676834 705183 676862 705553
rect 676820 705174 676876 705183
rect 676820 705109 676876 705118
rect 677026 702773 677054 705553
rect 677014 702767 677066 702773
rect 677014 702709 677066 702715
rect 675394 697931 675422 698338
rect 675380 697922 675436 697931
rect 675380 697857 675436 697866
rect 675778 697339 675806 697672
rect 675764 697330 675820 697339
rect 675764 697265 675820 697274
rect 675394 696895 675422 697035
rect 675380 696886 675436 696895
rect 675380 696821 675436 696830
rect 675778 694823 675806 695195
rect 675764 694814 675820 694823
rect 675764 694749 675820 694758
rect 675490 694379 675518 694638
rect 675476 694370 675532 694379
rect 675476 694305 675532 694314
rect 675778 693491 675806 693972
rect 675764 693482 675820 693491
rect 675764 693417 675820 693426
rect 675394 692931 675422 693380
rect 675478 692999 675530 693005
rect 675478 692941 675530 692947
rect 675382 692925 675434 692931
rect 675382 692867 675434 692873
rect 675490 692788 675518 692941
rect 675382 692703 675434 692709
rect 675382 692645 675434 692651
rect 674626 692552 675038 692580
rect 674626 681184 674654 692552
rect 675394 692173 675422 692645
rect 675394 692159 675792 692173
rect 675408 692145 675806 692159
rect 675778 692011 675806 692145
rect 675764 692002 675820 692011
rect 675764 691937 675820 691946
rect 675490 690711 675518 690864
rect 674806 690705 674858 690711
rect 674806 690647 674858 690653
rect 675478 690705 675530 690711
rect 675478 690647 675530 690653
rect 674710 687375 674762 687381
rect 674710 687317 674762 687323
rect 674434 681156 674654 681184
rect 674326 671021 674378 671027
rect 674326 670963 674378 670969
rect 674434 666703 674462 681156
rect 674722 679408 674750 687317
rect 674626 679380 674750 679408
rect 674420 666694 674476 666703
rect 674420 666629 674476 666638
rect 674228 666176 674284 666185
rect 674228 666111 674284 666120
rect 674422 658515 674474 658521
rect 674422 658457 674474 658463
rect 674132 642311 674188 642320
rect 673940 642274 673996 642283
rect 674132 642246 674188 642255
rect 673940 642209 673996 642218
rect 674146 642167 674174 642246
rect 673942 642161 673994 642167
rect 673942 642103 673994 642109
rect 674134 642161 674186 642167
rect 674134 642103 674186 642109
rect 673954 623339 673982 642103
rect 674434 627885 674462 658457
rect 674518 653779 674570 653785
rect 674518 653721 674570 653727
rect 674530 647125 674558 653721
rect 674518 647119 674570 647125
rect 674518 647061 674570 647067
rect 674518 645935 674570 645941
rect 674518 645877 674570 645883
rect 674422 627879 674474 627885
rect 674422 627821 674474 627827
rect 674422 627731 674474 627737
rect 674420 627696 674422 627705
rect 674474 627696 674476 627705
rect 674420 627631 674476 627640
rect 674422 626621 674474 626627
rect 674420 626586 674422 626595
rect 674474 626586 674476 626595
rect 674420 626521 674476 626530
rect 674420 625550 674476 625559
rect 674420 625485 674422 625494
rect 674474 625485 674476 625494
rect 674422 625453 674474 625459
rect 673940 623330 673996 623339
rect 673940 623265 673996 623274
rect 674530 622007 674558 645877
rect 674516 621998 674572 622007
rect 674516 621933 674572 621942
rect 674626 619195 674654 679380
rect 674818 676300 674846 690647
rect 675394 689823 675422 690346
rect 675382 689817 675434 689823
rect 675382 689759 675434 689765
rect 675394 689379 675422 689680
rect 675382 689373 675434 689379
rect 675382 689315 675434 689321
rect 675490 688639 675518 689014
rect 675478 688633 675530 688639
rect 675478 688575 675530 688581
rect 675490 687381 675518 687830
rect 675478 687375 675530 687381
rect 675478 687317 675530 687323
rect 675394 686271 675422 686646
rect 675382 686265 675434 686271
rect 675382 686207 675434 686213
rect 675490 685531 675518 685980
rect 675478 685525 675530 685531
rect 675478 685467 675530 685473
rect 675490 683681 675518 684130
rect 675478 683675 675530 683681
rect 675478 683617 675530 683623
rect 675478 683379 675530 683385
rect 675478 683321 675530 683327
rect 674722 676272 674846 676300
rect 674722 673099 674750 676272
rect 674710 673093 674762 673099
rect 674710 673035 674762 673041
rect 674998 673093 675050 673099
rect 674998 673035 675050 673041
rect 674710 672945 674762 672951
rect 674708 672910 674710 672919
rect 674762 672910 674764 672919
rect 674708 672845 674764 672854
rect 674710 672353 674762 672359
rect 674708 672318 674710 672327
rect 674762 672318 674764 672327
rect 674708 672253 674764 672262
rect 674710 671909 674762 671915
rect 674708 671874 674710 671883
rect 674762 671874 674764 671883
rect 674708 671809 674764 671818
rect 674710 671021 674762 671027
rect 674710 670963 674762 670969
rect 674722 668627 674750 670963
rect 674708 668618 674764 668627
rect 674708 668553 674764 668562
rect 674710 664213 674762 664219
rect 674708 664178 674710 664187
rect 674762 664178 674764 664187
rect 674708 664113 674764 664122
rect 674708 660922 674764 660931
rect 674708 660857 674764 660866
rect 674722 660487 674750 660857
rect 674708 660478 674764 660487
rect 674708 660413 674764 660422
rect 674722 659557 674750 660413
rect 674710 659551 674762 659557
rect 674710 659493 674762 659499
rect 674708 653670 674764 653679
rect 674708 653605 674764 653614
rect 674722 646404 674750 653605
rect 674722 646385 674846 646404
rect 674722 646379 674858 646385
rect 674722 646376 674806 646379
rect 674806 646321 674858 646327
rect 674818 638245 674846 646321
rect 675010 645941 675038 673035
rect 675092 660478 675148 660487
rect 675092 660413 675148 660422
rect 675106 659895 675134 660413
rect 675092 659886 675148 659895
rect 675092 659821 675148 659830
rect 675490 658521 675518 683321
rect 675478 658515 675530 658521
rect 675478 658457 675530 658463
rect 675394 652643 675422 653124
rect 675380 652634 675436 652643
rect 675380 652569 675436 652578
rect 675490 652199 675518 652458
rect 675476 652190 675532 652199
rect 675476 652125 675532 652134
rect 675490 651459 675518 651835
rect 675476 651450 675532 651459
rect 675476 651385 675532 651394
rect 675682 649831 675710 650016
rect 675668 649822 675724 649831
rect 675668 649757 675724 649766
rect 675490 648943 675518 649424
rect 675476 648934 675532 648943
rect 675476 648869 675532 648878
rect 675394 648309 675422 648799
rect 675382 648303 675434 648309
rect 675382 648245 675434 648251
rect 675394 648087 675422 648166
rect 675382 648081 675434 648087
rect 675382 648023 675434 648029
rect 675394 647125 675422 647603
rect 675382 647119 675434 647125
rect 675382 647061 675434 647067
rect 675394 646459 675422 646982
rect 675382 646453 675434 646459
rect 675382 646395 675434 646401
rect 674998 645935 675050 645941
rect 674998 645877 675050 645883
rect 675490 645391 675518 645650
rect 675476 645382 675532 645391
rect 675476 645317 675532 645326
rect 675490 644609 675518 645132
rect 675478 644603 675530 644609
rect 675478 644545 675530 644551
rect 675490 644091 675518 644466
rect 675478 644085 675530 644091
rect 675478 644027 675530 644033
rect 675394 643425 675422 643831
rect 675382 643419 675434 643425
rect 675382 643361 675434 643367
rect 675490 642315 675518 642616
rect 675478 642309 675530 642315
rect 675478 642251 675530 642257
rect 675490 641131 675518 641432
rect 675478 641125 675530 641131
rect 675478 641067 675530 641073
rect 675778 640359 675806 640795
rect 675764 640350 675820 640359
rect 675764 640285 675820 640294
rect 675778 638583 675806 638955
rect 675764 638574 675820 638583
rect 675764 638509 675820 638518
rect 674806 638239 674858 638245
rect 674806 638181 674858 638187
rect 675478 638239 675530 638245
rect 675478 638181 675530 638187
rect 675094 627879 675146 627885
rect 675094 627821 675146 627827
rect 674902 627361 674954 627367
rect 674900 627326 674902 627335
rect 674954 627326 674956 627335
rect 674900 627261 674956 627270
rect 675106 621415 675134 627821
rect 675092 621406 675148 621415
rect 675092 621341 675148 621350
rect 674612 619186 674668 619195
rect 674612 619121 674668 619130
rect 674422 618481 674474 618487
rect 674420 618446 674422 618455
rect 674474 618446 674476 618455
rect 674420 618381 674476 618390
rect 674422 617889 674474 617895
rect 674420 617854 674422 617863
rect 674474 617854 674476 617863
rect 674420 617789 674476 617798
rect 674710 617593 674762 617599
rect 674708 617558 674710 617567
rect 674762 617558 674764 617567
rect 674708 617493 674764 617502
rect 674998 613449 675050 613455
rect 674998 613391 675050 613397
rect 675010 602873 675038 613391
rect 675490 612197 675518 638181
rect 676820 624810 676876 624819
rect 676820 624745 676876 624754
rect 676834 622113 676862 624745
rect 676916 624070 676972 624079
rect 676916 624005 676972 624014
rect 676930 622187 676958 624005
rect 676918 622181 676970 622187
rect 676918 622123 676970 622129
rect 676822 622107 676874 622113
rect 676822 622049 676874 622055
rect 677108 615930 677164 615939
rect 677108 615865 677164 615874
rect 677122 615347 677150 615865
rect 676916 615338 676972 615347
rect 676916 615273 676972 615282
rect 677108 615338 677164 615347
rect 677108 615273 677164 615282
rect 676930 614903 676958 615273
rect 676916 614894 676972 614903
rect 676916 614829 676972 614838
rect 677122 613529 677150 615273
rect 677110 613523 677162 613529
rect 677110 613465 677162 613471
rect 675094 612191 675146 612197
rect 675094 612133 675146 612139
rect 675478 612191 675530 612197
rect 675478 612133 675530 612139
rect 674998 602867 675050 602873
rect 674998 602809 675050 602815
rect 675106 602503 675134 612133
rect 675394 607799 675422 608132
rect 675380 607790 675436 607799
rect 675380 607725 675436 607734
rect 675490 607207 675518 607466
rect 675476 607198 675532 607207
rect 675476 607133 675532 607142
rect 675490 606467 675518 606835
rect 675476 606458 675532 606467
rect 675476 606393 675532 606402
rect 675394 604839 675422 604995
rect 675380 604830 675436 604839
rect 675380 604765 675436 604774
rect 675490 604131 675518 604432
rect 675478 604125 675530 604131
rect 675478 604067 675530 604073
rect 675394 603317 675422 603799
rect 675382 603311 675434 603317
rect 675382 603253 675434 603259
rect 675394 602725 675422 603174
rect 675478 602867 675530 602873
rect 675478 602809 675530 602815
rect 675382 602719 675434 602725
rect 675382 602661 675434 602667
rect 675490 602582 675518 602809
rect 675094 602497 675146 602503
rect 675094 602439 675146 602445
rect 675382 602497 675434 602503
rect 675382 602439 675434 602445
rect 674422 601979 674474 601985
rect 675394 601959 675422 602439
rect 674422 601921 674474 601927
rect 674434 596879 674462 601921
rect 675778 600251 675806 600658
rect 675764 600242 675820 600251
rect 675764 600177 675820 600186
rect 675394 599839 675422 600140
rect 675382 599833 675434 599839
rect 675382 599775 675434 599781
rect 675394 599321 675422 599474
rect 675382 599315 675434 599321
rect 675382 599257 675434 599263
rect 675490 598433 675518 598808
rect 675478 598427 675530 598433
rect 675478 598369 675530 598375
rect 675490 597175 675518 597624
rect 675478 597169 675530 597175
rect 675478 597111 675530 597117
rect 674422 596873 674474 596879
rect 674422 596815 674474 596821
rect 675382 596873 675434 596879
rect 675382 596815 675434 596821
rect 675394 596440 675422 596815
rect 675778 595367 675806 595774
rect 675764 595358 675820 595367
rect 675764 595293 675820 595302
rect 675778 593443 675806 593955
rect 675764 593434 675820 593443
rect 675764 593369 675820 593378
rect 676822 587549 676874 587555
rect 676822 587491 676874 587497
rect 674612 582186 674668 582195
rect 674612 582121 674668 582130
rect 674422 582073 674474 582079
rect 674422 582015 674474 582021
rect 674434 581973 674462 582015
rect 674626 582005 674654 582121
rect 674614 581999 674666 582005
rect 674420 581964 674476 581973
rect 674614 581941 674666 581947
rect 674420 581899 674476 581908
rect 674614 581629 674666 581635
rect 674612 581594 674614 581603
rect 674666 581594 674668 581603
rect 674612 581529 674668 581538
rect 674422 580889 674474 580895
rect 674420 580854 674422 580863
rect 674474 580854 674476 580863
rect 674420 580789 674476 580798
rect 673844 580262 673900 580271
rect 673844 580197 673900 580206
rect 673858 579193 673886 580197
rect 676834 579531 676862 587491
rect 676820 579522 676876 579531
rect 676820 579457 676876 579466
rect 673846 579187 673898 579193
rect 673846 579129 673898 579135
rect 673846 576005 673898 576011
rect 673846 575947 673898 575953
rect 673858 573759 673886 575947
rect 673844 573750 673900 573759
rect 673844 573685 673900 573694
rect 673846 573637 673898 573643
rect 673846 573579 673898 573585
rect 673858 573315 673886 573579
rect 673844 573306 673900 573315
rect 673844 573241 673900 573250
rect 673846 573119 673898 573125
rect 673846 573061 673898 573067
rect 673748 572714 673804 572723
rect 673748 572649 673804 572658
rect 673858 572131 673886 573061
rect 673844 572122 673900 572131
rect 673844 572057 673900 572066
rect 674422 571639 674474 571645
rect 674420 571604 674422 571613
rect 674474 571604 674476 571613
rect 674420 571539 674476 571548
rect 677012 570790 677068 570799
rect 677012 570725 677068 570734
rect 676820 570198 676876 570207
rect 676820 570133 676876 570142
rect 676834 569763 676862 570133
rect 676820 569754 676876 569763
rect 676820 569689 676876 569698
rect 677026 569615 677054 570725
rect 677012 569606 677068 569615
rect 677012 569541 677068 569550
rect 677026 567427 677054 569541
rect 677014 567421 677066 567427
rect 677014 567363 677066 567369
rect 675094 564461 675146 564467
rect 675094 564403 675146 564409
rect 674998 564387 675050 564393
rect 674998 564329 675050 564335
rect 674230 559577 674282 559583
rect 674230 559519 674282 559525
rect 673750 557653 673802 557659
rect 673750 557595 673802 557601
rect 673652 529942 673708 529951
rect 673652 529877 673654 529886
rect 673706 529877 673708 529886
rect 673654 529845 673706 529851
rect 673556 529350 673612 529359
rect 673556 529285 673612 529294
rect 673364 527722 673420 527731
rect 673364 527657 673420 527666
rect 673268 484210 673324 484219
rect 673268 484145 673324 484154
rect 672886 483801 672938 483807
rect 673762 483775 673790 557595
rect 673846 492459 673898 492465
rect 673846 492401 673898 492407
rect 673858 492359 673886 492401
rect 673844 492350 673900 492359
rect 673844 492285 673900 492294
rect 674242 488067 674270 559519
rect 674710 558097 674762 558103
rect 674710 558039 674762 558045
rect 674422 555285 674474 555291
rect 674422 555227 674474 555233
rect 674326 551955 674378 551961
rect 674326 551897 674378 551903
rect 674228 488058 674284 488067
rect 674228 487993 674284 488002
rect 674338 484811 674366 551897
rect 674434 487475 674462 555227
rect 674518 550105 674570 550111
rect 674518 550047 674570 550053
rect 674530 489399 674558 550047
rect 674614 548255 674666 548261
rect 674614 548197 674666 548203
rect 674516 489390 674572 489399
rect 674516 489325 674572 489334
rect 674420 487466 674476 487475
rect 674420 487401 674476 487410
rect 674626 487179 674654 548197
rect 674722 509652 674750 558039
rect 675010 557881 675038 564329
rect 674998 557875 675050 557881
rect 674998 557817 675050 557823
rect 675106 557141 675134 564403
rect 675490 562659 675518 562918
rect 675476 562650 675532 562659
rect 675476 562585 675532 562594
rect 675490 561771 675518 562252
rect 675476 561762 675532 561771
rect 675476 561697 675532 561706
rect 675394 561475 675422 561660
rect 675380 561466 675436 561475
rect 675380 561401 675436 561410
rect 675394 559583 675422 559810
rect 675382 559577 675434 559583
rect 675382 559519 675434 559525
rect 675490 558959 675518 559218
rect 675476 558950 675532 558959
rect 675476 558885 675532 558894
rect 675394 558103 675422 558626
rect 675382 558097 675434 558103
rect 675382 558039 675434 558045
rect 675382 557875 675434 557881
rect 675382 557817 675434 557823
rect 675394 557403 675422 557817
rect 675490 557659 675518 557960
rect 675478 557653 675530 557659
rect 675478 557595 675530 557601
rect 675094 557135 675146 557141
rect 675094 557077 675146 557083
rect 675478 557135 675530 557141
rect 675478 557077 675530 557083
rect 675490 556776 675518 557077
rect 674998 555877 675050 555883
rect 674998 555819 675050 555825
rect 675010 551665 675038 555819
rect 675490 555291 675518 555444
rect 675478 555285 675530 555291
rect 675478 555227 675530 555233
rect 675778 554519 675806 554926
rect 675764 554510 675820 554519
rect 675764 554445 675820 554454
rect 675490 553811 675518 554260
rect 675478 553805 675530 553811
rect 675478 553747 675530 553753
rect 675394 553219 675422 553631
rect 675382 553213 675434 553219
rect 675382 553155 675434 553161
rect 675490 551961 675518 552410
rect 675478 551955 675530 551961
rect 675478 551897 675530 551903
rect 674998 551659 675050 551665
rect 674998 551601 675050 551607
rect 675382 551659 675434 551665
rect 675382 551601 675434 551607
rect 675394 551226 675422 551601
rect 675490 550111 675518 550595
rect 675478 550105 675530 550111
rect 675478 550047 675530 550053
rect 675490 548261 675518 548755
rect 675478 548255 675530 548261
rect 675478 548197 675530 548203
rect 674806 537229 674858 537235
rect 674804 537194 674806 537203
rect 674858 537194 674860 537203
rect 674804 537129 674860 537138
rect 676820 537194 676876 537203
rect 676820 537129 676876 537138
rect 674806 536637 674858 536643
rect 674804 536602 674806 536611
rect 674858 536602 674860 536611
rect 674804 536537 674860 536546
rect 674806 536193 674858 536199
rect 674804 536158 674806 536167
rect 674858 536158 674860 536167
rect 674804 536093 674860 536102
rect 676834 535829 676862 537129
rect 676822 535823 676874 535829
rect 676822 535765 676874 535771
rect 677300 535122 677356 535131
rect 677300 535057 677356 535066
rect 676916 533938 676972 533947
rect 676916 533873 676972 533882
rect 674806 529089 674858 529095
rect 674804 529054 674806 529063
rect 674858 529054 674860 529063
rect 674804 528989 674860 528998
rect 674806 528497 674858 528503
rect 674804 528462 674806 528471
rect 674858 528462 674860 528471
rect 674804 528397 674860 528406
rect 676820 525206 676876 525215
rect 676820 525141 676876 525150
rect 676834 524771 676862 525141
rect 676820 524762 676876 524771
rect 676820 524697 676876 524706
rect 674722 509624 674846 509652
rect 674612 487170 674668 487179
rect 674612 487105 674668 487114
rect 674818 485551 674846 509624
rect 675094 493273 675146 493279
rect 674900 493238 674956 493247
rect 674900 493173 674956 493182
rect 675092 493238 675094 493247
rect 675146 493238 675148 493247
rect 675092 493173 675148 493182
rect 674914 492539 674942 493173
rect 674902 492533 674954 492539
rect 674902 492475 674954 492481
rect 676930 489991 676958 533873
rect 677206 525981 677258 525987
rect 677206 525923 677258 525929
rect 677012 525798 677068 525807
rect 677012 525733 677068 525742
rect 677026 525215 677054 525733
rect 677012 525206 677068 525215
rect 677012 525141 677068 525150
rect 677026 524359 677054 525141
rect 677014 524353 677066 524359
rect 677014 524295 677066 524301
rect 677218 490583 677246 525923
rect 677314 492211 677342 535057
rect 677396 534530 677452 534539
rect 677396 534465 677452 534474
rect 677410 525987 677438 534465
rect 677398 525981 677450 525987
rect 677398 525923 677450 525929
rect 677300 492202 677356 492211
rect 677300 492137 677356 492146
rect 677396 491018 677452 491027
rect 677396 490953 677452 490962
rect 677204 490574 677260 490583
rect 677204 490509 677260 490518
rect 676916 489982 676972 489991
rect 676916 489917 676972 489926
rect 674804 485542 674860 485551
rect 674804 485477 674860 485486
rect 674324 484802 674380 484811
rect 674324 484737 674380 484746
rect 673846 483801 673898 483807
rect 672886 483743 672938 483749
rect 673748 483766 673804 483775
rect 673846 483743 673898 483749
rect 673748 483701 673804 483710
rect 673858 482591 673886 483743
rect 673844 482582 673900 482591
rect 673844 482517 673900 482526
rect 676820 481250 676876 481259
rect 676820 481185 676876 481194
rect 676834 480815 676862 481185
rect 676820 480806 676876 480815
rect 676820 480741 676876 480750
rect 673846 406101 673898 406107
rect 673846 406043 673898 406049
rect 673858 404743 673886 406043
rect 674710 405509 674762 405515
rect 674708 405474 674710 405483
rect 674762 405474 674764 405483
rect 674708 405409 674764 405418
rect 673844 404734 673900 404743
rect 673844 404669 673900 404678
rect 674710 404473 674762 404479
rect 674708 404438 674710 404447
rect 674762 404438 674764 404447
rect 674708 404373 674764 404382
rect 673844 403106 673900 403115
rect 673844 403041 673900 403050
rect 673366 400477 673418 400483
rect 673366 400419 673418 400425
rect 673378 373367 673406 400419
rect 673750 400403 673802 400409
rect 673750 400345 673802 400351
rect 673762 374403 673790 400345
rect 673748 374394 673804 374403
rect 673748 374329 673804 374338
rect 673364 373358 673420 373367
rect 673364 373293 673420 373302
rect 672502 359037 672554 359043
rect 672502 358979 672554 358985
rect 673858 358419 673886 403041
rect 676930 402227 676958 489917
rect 677012 481694 677068 481703
rect 677012 481629 677068 481638
rect 677026 480815 677054 481629
rect 677012 480806 677068 480815
rect 677012 480741 677068 480750
rect 677026 479515 677054 480741
rect 677014 479509 677066 479515
rect 677014 479451 677066 479457
rect 677218 402819 677246 490509
rect 677410 404003 677438 490953
rect 677396 403994 677452 404003
rect 677396 403929 677452 403938
rect 677204 402810 677260 402819
rect 677204 402745 677260 402754
rect 676916 402218 676972 402227
rect 676916 402153 676972 402162
rect 675092 401330 675148 401339
rect 675092 401265 675148 401274
rect 674132 399850 674188 399859
rect 674132 399785 674188 399794
rect 673940 396594 673996 396603
rect 673940 396529 673996 396538
rect 673954 375767 673982 396529
rect 674146 383167 674174 399785
rect 674228 397630 674284 397639
rect 674228 397565 674284 397574
rect 674134 383161 674186 383167
rect 674134 383103 674186 383109
rect 674242 382501 674270 397565
rect 674900 396890 674956 396899
rect 674900 396825 674956 396834
rect 674516 395854 674572 395863
rect 674516 395789 674572 395798
rect 674230 382495 674282 382501
rect 674230 382437 674282 382443
rect 674530 377617 674558 395789
rect 674804 394670 674860 394679
rect 674804 394605 674860 394614
rect 674612 394226 674668 394235
rect 674612 394161 674668 394170
rect 674518 377611 674570 377617
rect 674518 377553 674570 377559
rect 674626 376951 674654 394161
rect 674818 378209 674846 394605
rect 674914 384721 674942 396825
rect 674996 395262 675052 395271
rect 674996 395197 675052 395206
rect 674902 384715 674954 384721
rect 674902 384657 674954 384663
rect 675010 381336 675038 395197
rect 675106 384869 675134 401265
rect 676930 400483 676958 402153
rect 676918 400477 676970 400483
rect 676918 400419 676970 400425
rect 677218 400409 677246 402745
rect 677206 400403 677258 400409
rect 677206 400345 677258 400351
rect 675380 400146 675436 400155
rect 675380 400081 675436 400090
rect 675188 397926 675244 397935
rect 675188 397861 675244 397870
rect 675202 385461 675230 397861
rect 675394 386423 675422 400081
rect 677108 393486 677164 393495
rect 677108 393421 677164 393430
rect 677122 393051 677150 393421
rect 676916 393042 676972 393051
rect 676916 392977 676972 392986
rect 677108 393042 677164 393051
rect 677108 392977 677164 392986
rect 676930 392607 676958 392977
rect 676916 392598 676972 392607
rect 676916 392533 676972 392542
rect 677122 391825 677150 392977
rect 677110 391819 677162 391825
rect 677110 391761 677162 391767
rect 675382 386417 675434 386423
rect 675382 386359 675434 386365
rect 675382 386195 675434 386201
rect 675382 386137 675434 386143
rect 675394 385723 675422 386137
rect 675190 385455 675242 385461
rect 675190 385397 675242 385403
rect 675478 385455 675530 385461
rect 675478 385397 675530 385403
rect 675490 385096 675518 385397
rect 675094 384863 675146 384869
rect 675094 384805 675146 384811
rect 675382 384863 675434 384869
rect 675382 384805 675434 384811
rect 675094 384715 675146 384721
rect 675094 384657 675146 384663
rect 675106 381410 675134 384657
rect 675394 384430 675422 384805
rect 675286 383161 675338 383167
rect 675286 383103 675338 383109
rect 675298 382668 675326 383103
rect 675298 382640 675422 382668
rect 675394 382580 675422 382640
rect 675478 382495 675530 382501
rect 675478 382437 675530 382443
rect 675490 382062 675518 382437
rect 675106 381382 675408 381410
rect 675010 381308 675422 381336
rect 675394 380730 675422 381308
rect 675106 380198 675408 380226
rect 674806 378203 674858 378209
rect 674806 378145 674858 378151
rect 674614 376945 674666 376951
rect 674614 376887 674666 376893
rect 673942 375761 673994 375767
rect 673942 375703 673994 375709
rect 675106 374551 675134 380198
rect 675202 379532 675408 379560
rect 675092 374542 675148 374551
rect 675092 374477 675148 374486
rect 675202 374107 675230 379532
rect 675476 378834 675532 378843
rect 675476 378769 675532 378778
rect 675490 378288 675518 378769
rect 675382 378203 675434 378209
rect 675382 378145 675434 378151
rect 675394 377696 675422 378145
rect 675382 377611 675434 377617
rect 675382 377553 675434 377559
rect 675394 377075 675422 377553
rect 675478 376945 675530 376951
rect 675478 376887 675530 376893
rect 675490 376438 675518 376887
rect 675478 375761 675530 375767
rect 675478 375703 675530 375709
rect 675490 375254 675518 375703
rect 675188 374098 675244 374107
rect 675188 374033 675244 374042
rect 675476 373950 675532 373959
rect 675476 373885 675532 373894
rect 675490 373404 675518 373885
rect 675380 372026 675436 372035
rect 675380 371961 675436 371970
rect 675394 371554 675422 371961
rect 674422 360073 674474 360079
rect 674420 360038 674422 360047
rect 674474 360038 674476 360047
rect 674420 359973 674476 359982
rect 674710 359777 674762 359783
rect 674708 359742 674710 359751
rect 674762 359742 674764 359751
rect 674708 359677 674764 359686
rect 674422 359037 674474 359043
rect 674420 359002 674422 359011
rect 674474 359002 674476 359011
rect 674420 358937 674476 358946
rect 673844 358410 673900 358419
rect 673844 358345 673900 358354
rect 674900 356042 674956 356051
rect 674900 355977 674956 355986
rect 673940 354118 673996 354127
rect 673940 354053 673996 354062
rect 673954 333587 673982 354053
rect 674324 351898 674380 351907
rect 674324 351833 674380 351842
rect 674132 350862 674188 350871
rect 674132 350797 674188 350806
rect 674036 349678 674092 349687
rect 674036 349613 674092 349622
rect 673942 333581 673994 333587
rect 673942 333523 673994 333529
rect 674050 332773 674078 349613
rect 674038 332767 674090 332773
rect 674038 332709 674090 332715
rect 674146 332255 674174 350797
rect 674338 336621 674366 351833
rect 674708 350122 674764 350131
rect 674708 350057 674764 350066
rect 674516 348938 674572 348947
rect 674516 348873 674572 348882
rect 674326 336615 674378 336621
rect 674326 336557 674378 336563
rect 674134 332249 674186 332255
rect 674134 332191 674186 332197
rect 674530 331811 674558 348873
rect 674722 335569 674750 350057
rect 674914 339581 674942 355977
rect 675188 355006 675244 355015
rect 675188 354941 675244 354950
rect 674996 354414 675052 354423
rect 674996 354349 675052 354358
rect 675010 340839 675038 354349
rect 675092 352194 675148 352203
rect 675092 352129 675148 352138
rect 674998 340833 675050 340839
rect 674998 340775 675050 340781
rect 674902 339575 674954 339581
rect 674902 339517 674954 339523
rect 675106 336862 675134 352129
rect 675202 340987 675230 354941
rect 677108 353230 677164 353239
rect 677108 353165 677164 353174
rect 675284 352786 675340 352795
rect 675284 352721 675340 352730
rect 675190 340981 675242 340987
rect 675190 340923 675242 340929
rect 675190 340833 675242 340839
rect 675190 340775 675242 340781
rect 675202 337409 675230 340775
rect 675298 339896 675326 352721
rect 676916 351158 676972 351167
rect 676916 351093 676972 351102
rect 676820 347754 676876 347763
rect 676820 347689 676876 347698
rect 676834 347319 676862 347689
rect 676820 347310 676876 347319
rect 676820 347245 676876 347254
rect 676930 344211 676958 351093
rect 677012 348346 677068 348355
rect 677012 348281 677068 348290
rect 677026 347319 677054 348281
rect 677012 347310 677068 347319
rect 677012 347245 677068 347254
rect 677026 345649 677054 347245
rect 677014 345643 677066 345649
rect 677014 345585 677066 345591
rect 677122 345247 677150 353165
rect 677108 345238 677164 345247
rect 677108 345173 677164 345182
rect 676916 344202 676972 344211
rect 676916 344137 676972 344146
rect 675478 340981 675530 340987
rect 675478 340923 675530 340929
rect 675490 340548 675518 340923
rect 675298 339868 675408 339896
rect 675382 339575 675434 339581
rect 675382 339517 675434 339523
rect 675394 339216 675422 339517
rect 675202 337381 675408 337409
rect 675106 336834 675408 336862
rect 675382 336615 675434 336621
rect 675382 336557 675434 336563
rect 675394 336182 675422 336557
rect 674722 335541 675408 335569
rect 675284 335026 675340 335035
rect 675010 334984 675284 335012
rect 674518 331805 674570 331811
rect 674518 331747 674570 331753
rect 675010 329559 675038 334984
rect 675340 334984 675408 335012
rect 675284 334961 675340 334970
rect 675298 334901 675326 334961
rect 675476 334582 675532 334591
rect 675476 334517 675532 334526
rect 675298 334392 675422 334420
rect 675298 334346 675326 334392
rect 675106 334318 675326 334346
rect 675394 334346 675422 334392
rect 675490 334346 675518 334517
rect 675394 334332 675518 334346
rect 675408 334318 675504 334332
rect 675106 331187 675134 334318
rect 675382 333581 675434 333587
rect 675382 333523 675434 333529
rect 675394 333074 675422 333523
rect 675382 332767 675434 332773
rect 675382 332709 675434 332715
rect 675394 332519 675422 332709
rect 675478 332249 675530 332255
rect 675478 332191 675530 332197
rect 675490 331890 675518 332191
rect 675382 331805 675434 331811
rect 675382 331747 675434 331753
rect 675394 331224 675422 331747
rect 675092 331178 675148 331187
rect 675092 331113 675148 331122
rect 675764 330586 675820 330595
rect 675764 330521 675820 330530
rect 675778 330040 675806 330521
rect 674996 329550 675052 329559
rect 674996 329485 675052 329494
rect 675380 328366 675436 328375
rect 675380 328301 675436 328310
rect 675394 328190 675422 328301
rect 675764 326886 675820 326895
rect 675764 326821 675820 326830
rect 675778 326340 675806 326821
rect 674422 315081 674474 315087
rect 674420 315046 674422 315055
rect 674474 315046 674476 315055
rect 674420 314981 674476 314990
rect 674710 314785 674762 314791
rect 674708 314750 674710 314759
rect 674762 314750 674764 314759
rect 674708 314685 674764 314694
rect 674422 314045 674474 314051
rect 674420 314010 674422 314019
rect 674474 314010 674476 314019
rect 674420 313945 674476 313954
rect 674036 311346 674092 311355
rect 674036 311281 674092 311290
rect 674050 294811 674078 311281
rect 675092 310014 675148 310023
rect 675092 309949 675148 309958
rect 674324 309644 674380 309653
rect 674324 309579 674380 309588
rect 674132 305870 674188 305879
rect 674132 305805 674188 305814
rect 674038 294805 674090 294811
rect 674038 294747 674090 294753
rect 673940 289590 673996 289599
rect 673940 289525 673996 289534
rect 673954 289483 673982 289525
rect 673942 289477 673994 289483
rect 673994 289425 674038 289428
rect 673942 289419 674038 289425
rect 673954 289400 674038 289419
rect 673954 284715 673982 289400
rect 674146 287263 674174 305805
rect 674228 304242 674284 304251
rect 674228 304177 674284 304186
rect 674134 287257 674186 287263
rect 674134 287199 674186 287205
rect 674242 286819 674270 304177
rect 674338 292961 674366 309579
rect 674996 308830 675052 308839
rect 674996 308765 675052 308774
rect 674900 307794 674956 307803
rect 674900 307729 674956 307738
rect 674804 307202 674860 307211
rect 674804 307137 674860 307146
rect 674612 306758 674668 306767
rect 674612 306693 674668 306702
rect 674516 304538 674572 304547
rect 674516 304473 674572 304482
rect 674420 303650 674476 303659
rect 674420 303585 674476 303594
rect 674434 302655 674462 303585
rect 674422 302649 674474 302655
rect 674420 302614 674422 302623
rect 674474 302614 674476 302623
rect 674420 302549 674476 302558
rect 674530 300676 674558 304473
rect 674434 300648 674558 300676
rect 674326 292955 674378 292961
rect 674326 292897 674378 292903
rect 674434 287781 674462 300648
rect 674626 300528 674654 306693
rect 674708 305130 674764 305139
rect 674708 305065 674764 305074
rect 674530 300500 674654 300528
rect 674530 291703 674558 300500
rect 674722 291777 674750 305065
rect 674818 293553 674846 307137
rect 674914 295477 674942 307729
rect 674902 295471 674954 295477
rect 674902 295413 674954 295419
rect 674806 293547 674858 293553
rect 674806 293489 674858 293495
rect 674710 291771 674762 291777
rect 674710 291713 674762 291719
rect 674518 291697 674570 291703
rect 674518 291639 674570 291645
rect 675010 288595 675038 308765
rect 675106 295537 675134 309949
rect 677012 308238 677068 308247
rect 677012 308173 677068 308182
rect 676916 306018 676972 306027
rect 676916 305953 676972 305962
rect 676820 302762 676876 302771
rect 676820 302697 676876 302706
rect 676834 302327 676862 302697
rect 676820 302318 676876 302327
rect 676820 302253 676876 302262
rect 676930 299515 676958 305953
rect 676916 299506 676972 299515
rect 676916 299441 676972 299450
rect 677026 299367 677054 308173
rect 677012 299358 677068 299367
rect 677012 299293 677068 299302
rect 675106 295509 675408 295537
rect 675094 295471 675146 295477
rect 675094 295413 675146 295419
rect 675106 294904 675134 295413
rect 675106 294876 675408 294904
rect 675094 294805 675146 294811
rect 675094 294747 675146 294753
rect 675106 294238 675134 294747
rect 675106 294210 675408 294238
rect 675094 293547 675146 293553
rect 675094 293489 675146 293495
rect 675106 291870 675134 293489
rect 675382 292955 675434 292961
rect 675382 292897 675434 292903
rect 675394 292374 675422 292897
rect 675106 291842 675408 291870
rect 675094 291771 675146 291777
rect 675094 291713 675146 291719
rect 675106 290569 675134 291713
rect 675190 291697 675242 291703
rect 675190 291639 675242 291645
rect 675202 291204 675230 291639
rect 675202 291176 675408 291204
rect 675106 290541 675408 290569
rect 675284 290034 675340 290043
rect 675106 289992 675284 290020
rect 674998 288589 675050 288595
rect 674998 288531 675050 288537
rect 674422 287775 674474 287781
rect 674422 287717 674474 287723
rect 674230 286813 674282 286819
rect 674230 286755 674282 286761
rect 675106 285011 675134 289992
rect 675340 289992 675408 290020
rect 675284 289969 675340 289978
rect 675298 289909 675326 289969
rect 675382 289477 675434 289483
rect 675382 289419 675434 289425
rect 675394 289340 675422 289419
rect 675478 288589 675530 288595
rect 675478 288531 675530 288537
rect 675490 288082 675518 288531
rect 675382 287775 675434 287781
rect 675382 287717 675434 287723
rect 675394 287519 675422 287717
rect 675478 287257 675530 287263
rect 675478 287199 675530 287205
rect 675490 286898 675518 287199
rect 675382 286813 675434 286819
rect 675382 286755 675434 286761
rect 675394 286232 675422 286755
rect 675092 285002 675148 285011
rect 675092 284937 675148 284946
rect 675778 284863 675806 285048
rect 675764 284854 675820 284863
rect 675764 284789 675820 284798
rect 673940 284706 673996 284715
rect 673940 284641 673996 284650
rect 675380 283670 675436 283679
rect 675380 283605 675436 283614
rect 675394 283198 675422 283605
rect 675764 281894 675820 281903
rect 675764 281829 675820 281838
rect 675778 281348 675806 281829
rect 669814 270089 669866 270095
rect 674422 270089 674474 270095
rect 669814 270031 669866 270037
rect 674420 270054 674422 270063
rect 674474 270054 674476 270063
rect 674420 269989 674476 269998
rect 674710 269793 674762 269799
rect 674708 269758 674710 269767
rect 674762 269758 674764 269767
rect 674708 269693 674764 269702
rect 674710 269201 674762 269207
rect 674708 269166 674710 269175
rect 674762 269166 674764 269175
rect 674708 269101 674764 269110
rect 674516 266058 674572 266067
rect 674516 265993 674572 266002
rect 674324 262506 674380 262515
rect 674324 262441 674380 262450
rect 674132 260878 674188 260887
rect 674132 260813 674188 260822
rect 674146 242419 674174 260813
rect 674338 247303 674366 262441
rect 674530 250411 674558 265993
rect 677108 265466 677164 265475
rect 677108 265401 677164 265410
rect 675188 265022 675244 265031
rect 675188 264957 675244 264966
rect 675092 264430 675148 264439
rect 675092 264365 675148 264374
rect 674804 261766 674860 261775
rect 674804 261701 674860 261710
rect 674708 261174 674764 261183
rect 674708 261109 674764 261118
rect 674612 259546 674668 259555
rect 674612 259481 674668 259490
rect 674518 250405 674570 250411
rect 674518 250347 674570 250353
rect 674326 247297 674378 247303
rect 674326 247239 674378 247245
rect 674626 243011 674654 259481
rect 674614 243005 674666 243011
rect 674614 242947 674666 242953
rect 674134 242413 674186 242419
rect 674134 242355 674186 242361
rect 674722 240569 674750 261109
rect 674818 247229 674846 261701
rect 674900 260138 674956 260147
rect 674900 260073 674956 260082
rect 674806 247223 674858 247229
rect 674806 247165 674858 247171
rect 674914 246341 674942 260073
rect 674996 258954 675052 258963
rect 674996 258889 675052 258898
rect 674902 246335 674954 246341
rect 674902 246277 674954 246283
rect 675010 241605 675038 258889
rect 675106 247396 675134 264365
rect 675202 251003 675230 264957
rect 676916 263246 676972 263255
rect 676916 263181 676972 263190
rect 675284 262802 675340 262811
rect 675284 262737 675340 262746
rect 675190 250997 675242 251003
rect 675190 250939 675242 250945
rect 675190 250405 675242 250411
rect 675190 250347 675242 250353
rect 675202 249246 675230 250347
rect 675298 250208 675326 262737
rect 676820 257770 676876 257779
rect 676820 257705 676876 257714
rect 676834 257335 676862 257705
rect 676820 257326 676876 257335
rect 676820 257261 676876 257270
rect 676930 253339 676958 263181
rect 677012 258362 677068 258371
rect 677012 258297 677068 258306
rect 677026 257779 677054 258297
rect 677012 257770 677068 257779
rect 677012 257705 677068 257714
rect 677026 256405 677054 257705
rect 677014 256399 677066 256405
rect 677014 256341 677066 256347
rect 676916 253330 676972 253339
rect 676916 253265 676972 253274
rect 677122 253191 677150 265401
rect 677108 253182 677164 253191
rect 677108 253117 677164 253126
rect 675382 250997 675434 251003
rect 675382 250939 675434 250945
rect 675394 250523 675422 250939
rect 675298 250180 675518 250208
rect 675490 249898 675518 250180
rect 675202 249218 675408 249246
rect 675106 247368 675408 247396
rect 675190 247297 675242 247303
rect 675190 247239 675242 247245
rect 675094 247223 675146 247229
rect 675094 247165 675146 247171
rect 675106 246212 675134 247165
rect 675202 246878 675230 247239
rect 675202 246850 675326 246878
rect 675298 246804 675326 246850
rect 675394 246804 675422 246864
rect 675298 246776 675422 246804
rect 675106 246184 675408 246212
rect 675286 246113 675338 246119
rect 675286 246055 675338 246061
rect 675298 245916 675326 246055
rect 675298 245888 675422 245916
rect 675394 245532 675422 245888
rect 675188 245338 675244 245347
rect 675188 245273 675244 245282
rect 675202 244362 675230 245273
rect 675394 244755 675422 245014
rect 675380 244746 675436 244755
rect 675380 244681 675436 244690
rect 675202 244334 675408 244362
rect 674998 241599 675050 241605
rect 674998 241541 675050 241547
rect 674710 240563 674762 240569
rect 674710 240505 674762 240511
rect 675202 238983 675230 244334
rect 675476 243562 675532 243571
rect 675476 243497 675532 243506
rect 675490 243090 675518 243497
rect 675382 243005 675434 243011
rect 675382 242947 675434 242953
rect 675394 242498 675422 242947
rect 675382 242413 675434 242419
rect 675382 242355 675434 242361
rect 675394 241875 675422 242355
rect 675478 241599 675530 241605
rect 675478 241541 675530 241547
rect 675490 241240 675518 241541
rect 675478 240563 675530 240569
rect 675478 240505 675530 240511
rect 675490 240056 675518 240505
rect 675188 238974 675244 238983
rect 675188 238909 675244 238918
rect 675764 238678 675820 238687
rect 675764 238613 675820 238622
rect 675778 238206 675806 238613
rect 675764 236902 675820 236911
rect 675764 236837 675820 236846
rect 675778 236356 675806 236837
rect 674710 225097 674762 225103
rect 674708 225062 674710 225071
rect 674762 225062 674764 225071
rect 674708 224997 674764 225006
rect 674422 224357 674474 224363
rect 674420 224322 674422 224331
rect 674474 224322 674476 224331
rect 674420 224257 674476 224266
rect 669622 224061 669674 224067
rect 674710 224061 674762 224067
rect 669622 224003 669674 224009
rect 674708 224026 674710 224035
rect 674762 224026 674764 224035
rect 674708 223961 674764 223970
rect 674900 220918 674956 220927
rect 674900 220853 674956 220862
rect 674228 216774 674284 216783
rect 674228 216709 674284 216718
rect 674242 201349 674270 216709
rect 674516 215442 674572 215451
rect 674516 215377 674572 215386
rect 674230 201343 674282 201349
rect 674230 201285 674282 201291
rect 674530 197057 674558 215377
rect 674804 214850 674860 214859
rect 674804 214785 674860 214794
rect 674708 214406 674764 214415
rect 674708 214341 674764 214350
rect 674612 213814 674668 213823
rect 674612 213749 674668 213758
rect 674518 197051 674570 197057
rect 674518 196993 674570 196999
rect 674626 196613 674654 213749
rect 674722 197797 674750 214341
rect 674818 200387 674846 214785
rect 674914 204457 674942 220853
rect 675476 219734 675532 219743
rect 675476 219669 675532 219678
rect 674996 219290 675052 219299
rect 674996 219225 675052 219234
rect 674902 204451 674954 204457
rect 674902 204393 674954 204399
rect 675010 202237 675038 219225
rect 675188 217662 675244 217671
rect 675188 217597 675244 217606
rect 675092 216922 675148 216931
rect 675092 216857 675148 216866
rect 674998 202231 675050 202237
rect 674998 202173 675050 202179
rect 675106 202089 675134 216857
rect 675202 205049 675230 217597
rect 675490 206011 675518 219669
rect 677108 218106 677164 218115
rect 677108 218041 677164 218050
rect 676916 216034 676972 216043
rect 676916 215969 676972 215978
rect 676820 212630 676876 212639
rect 676820 212565 676876 212574
rect 676834 212195 676862 212565
rect 676820 212186 676876 212195
rect 676820 212121 676876 212130
rect 676930 210271 676958 215969
rect 677012 213222 677068 213231
rect 677012 213157 677068 213166
rect 677026 212639 677054 213157
rect 677012 212630 677068 212639
rect 677012 212565 677068 212574
rect 677026 210303 677054 212565
rect 677014 210297 677066 210303
rect 676916 210262 676972 210271
rect 677014 210239 677066 210245
rect 676916 210197 676972 210206
rect 677122 210123 677150 218041
rect 677108 210114 677164 210123
rect 677108 210049 677164 210058
rect 675478 206005 675530 206011
rect 675478 205947 675530 205953
rect 675478 205783 675530 205789
rect 675478 205725 675530 205731
rect 675490 205350 675518 205725
rect 675190 205043 675242 205049
rect 675190 204985 675242 204991
rect 675478 205043 675530 205049
rect 675478 204985 675530 204991
rect 675490 204684 675518 204985
rect 675382 204451 675434 204457
rect 675382 204393 675434 204399
rect 675394 204018 675422 204393
rect 675298 202237 675422 202256
rect 675286 202231 675422 202237
rect 675338 202228 675422 202231
rect 675286 202173 675338 202179
rect 675394 202168 675422 202228
rect 675094 202083 675146 202089
rect 675094 202025 675146 202031
rect 675286 202083 675338 202089
rect 675286 202025 675338 202031
rect 675298 201664 675326 202025
rect 675298 201636 675408 201664
rect 675382 201343 675434 201349
rect 675382 201285 675434 201291
rect 675394 200984 675422 201285
rect 674806 200381 674858 200387
rect 674806 200323 674858 200329
rect 675286 200381 675338 200387
rect 675338 200341 675408 200369
rect 675286 200323 675338 200329
rect 675394 199319 675422 199800
rect 675380 199310 675436 199319
rect 675380 199245 675436 199254
rect 675490 198727 675518 199134
rect 675476 198718 675532 198727
rect 675476 198653 675532 198662
rect 675476 198422 675532 198431
rect 675476 198357 675532 198366
rect 675490 197876 675518 198357
rect 674710 197791 674762 197797
rect 674710 197733 674762 197739
rect 675382 197791 675434 197797
rect 675382 197733 675434 197739
rect 675394 197319 675422 197733
rect 675478 197051 675530 197057
rect 675478 196993 675530 196999
rect 675490 196692 675518 196993
rect 674614 196607 674666 196613
rect 674614 196549 674666 196555
rect 675382 196607 675434 196613
rect 675382 196549 675434 196555
rect 675394 196026 675422 196549
rect 675764 195314 675820 195323
rect 675764 195249 675820 195258
rect 675778 194842 675806 195249
rect 675380 193538 675436 193547
rect 675380 193473 675436 193482
rect 675394 192992 675422 193473
rect 675764 191614 675820 191623
rect 675764 191549 675820 191558
rect 675778 191142 675806 191549
rect 674708 179626 674764 179635
rect 674708 179561 674764 179570
rect 674422 179365 674474 179371
rect 674420 179330 674422 179339
rect 674474 179330 674476 179339
rect 674420 179265 674476 179274
rect 666646 178847 666698 178853
rect 674422 178847 674474 178853
rect 666646 178789 666698 178795
rect 674420 178812 674422 178821
rect 674474 178812 674476 178821
rect 674420 178747 674476 178756
rect 674722 178705 674750 179561
rect 674710 178699 674762 178705
rect 674710 178641 674762 178647
rect 674036 176074 674092 176083
rect 674036 176009 674092 176018
rect 674050 159465 674078 176009
rect 676916 175186 676972 175195
rect 676916 175121 676972 175130
rect 675572 174742 675628 174751
rect 675572 174677 675628 174686
rect 674804 174298 674860 174307
rect 674804 174233 674860 174242
rect 674324 169562 674380 169571
rect 674324 169497 674380 169506
rect 674038 159459 674090 159465
rect 674038 159401 674090 159407
rect 674338 152657 674366 169497
rect 674516 168822 674572 168831
rect 674516 168757 674572 168766
rect 674420 167342 674476 167351
rect 674420 167277 674422 167286
rect 674474 167277 674476 167286
rect 674422 167245 674474 167251
rect 674326 152651 674378 152657
rect 674326 152593 674378 152599
rect 674530 151547 674558 168757
rect 674612 168230 674668 168239
rect 674612 168165 674668 168174
rect 674626 167235 674654 168165
rect 674708 167638 674764 167647
rect 674708 167573 674764 167582
rect 674614 167229 674666 167235
rect 674614 167171 674666 167177
rect 674722 167161 674750 167573
rect 674710 167155 674762 167161
rect 674710 167097 674762 167103
rect 674818 157763 674846 174233
rect 675092 172078 675148 172087
rect 675092 172013 675148 172022
rect 674996 171486 675052 171495
rect 674996 171421 675052 171430
rect 674900 169858 674956 169867
rect 674900 169793 674956 169802
rect 674806 157757 674858 157763
rect 674806 157699 674858 157705
rect 674914 155369 674942 169793
rect 675010 156006 675038 171421
rect 675106 156672 675134 172013
rect 675586 161019 675614 174677
rect 676820 173114 676876 173123
rect 676820 173049 676876 173058
rect 675764 172670 675820 172679
rect 675764 172605 675820 172614
rect 675778 161019 675806 172605
rect 676834 161431 676862 173049
rect 676930 161579 676958 175121
rect 676916 161570 676972 161579
rect 676916 161505 676972 161514
rect 676820 161422 676876 161431
rect 676820 161357 676876 161366
rect 675574 161013 675626 161019
rect 675574 160955 675626 160961
rect 675766 161013 675818 161019
rect 675766 160955 675818 160961
rect 675574 160791 675626 160797
rect 675574 160733 675626 160739
rect 675586 160323 675614 160733
rect 675766 160051 675818 160057
rect 675766 159993 675818 159999
rect 675778 159692 675806 159993
rect 675382 159459 675434 159465
rect 675382 159401 675434 159407
rect 675394 159026 675422 159401
rect 675478 157757 675530 157763
rect 675478 157699 675530 157705
rect 675490 157176 675518 157699
rect 675106 156644 675326 156672
rect 675298 156524 675326 156644
rect 675394 156524 675422 156658
rect 675298 156496 675422 156524
rect 675010 155978 675408 156006
rect 674914 155341 675408 155369
rect 675284 155206 675340 155215
rect 675284 155141 675340 155150
rect 675298 154822 675326 155141
rect 675298 154794 675408 154822
rect 675476 154466 675532 154475
rect 675476 154401 675532 154410
rect 675490 154142 675518 154401
rect 675476 153430 675532 153439
rect 675476 153365 675532 153374
rect 675490 152884 675518 153365
rect 675382 152651 675434 152657
rect 675382 152593 675434 152599
rect 675394 152292 675422 152593
rect 675476 151950 675532 151959
rect 675476 151885 675532 151894
rect 675490 151700 675518 151885
rect 674518 151541 674570 151547
rect 674518 151483 674570 151489
rect 675382 151541 675434 151547
rect 675382 151483 675434 151489
rect 675394 151034 675422 151483
rect 675476 150322 675532 150331
rect 675476 150257 675532 150266
rect 675490 149850 675518 150257
rect 675764 148546 675820 148555
rect 675764 148481 675820 148490
rect 675778 148000 675806 148481
rect 675764 146622 675820 146631
rect 675764 146557 675820 146566
rect 675778 146150 675806 146557
rect 676916 134338 676972 134347
rect 676916 134273 676972 134282
rect 676820 133894 676876 133903
rect 676820 133829 676876 133838
rect 663766 133633 663818 133639
rect 674422 133633 674474 133639
rect 663766 133575 663818 133581
rect 674420 133598 674422 133607
rect 674474 133598 674476 133607
rect 674420 133533 674476 133542
rect 655318 132819 655370 132825
rect 655318 132761 655370 132767
rect 676834 132677 676862 133829
rect 676930 132825 676958 134273
rect 676918 132819 676970 132825
rect 676918 132761 676970 132767
rect 655126 132671 655178 132677
rect 655126 132613 655178 132619
rect 676822 132671 676874 132677
rect 676822 132613 676874 132619
rect 674420 132562 674476 132571
rect 647734 132523 647786 132529
rect 674420 132497 674422 132506
rect 647734 132465 647786 132471
rect 674474 132497 674476 132506
rect 674422 132465 674474 132471
rect 645826 126748 645950 126776
rect 645716 121462 645772 121471
rect 645716 121397 645772 121406
rect 645730 121281 645758 121397
rect 645718 121275 645770 121281
rect 645718 121217 645770 121223
rect 645718 121127 645770 121133
rect 645718 121069 645770 121075
rect 645730 120879 645758 121069
rect 645922 120985 645950 126748
rect 645910 120979 645962 120985
rect 645910 120921 645962 120927
rect 646102 120979 646154 120985
rect 646102 120921 646154 120927
rect 645716 120870 645772 120879
rect 645716 120805 645772 120814
rect 646114 100857 646142 120921
rect 647746 120435 647774 132465
rect 674516 130638 674572 130647
rect 674516 130573 674572 130582
rect 674324 127086 674380 127095
rect 674324 127021 674380 127030
rect 673940 125458 673996 125467
rect 673940 125393 673996 125402
rect 647732 120426 647788 120435
rect 647732 120361 647788 120370
rect 673954 106925 673982 125393
rect 674228 123830 674284 123839
rect 674228 123765 674284 123774
rect 673942 106919 673994 106925
rect 673942 106861 673994 106867
rect 668182 106549 668234 106555
rect 668180 106514 668182 106523
rect 668234 106514 668236 106523
rect 668180 106449 668236 106458
rect 674242 106407 674270 123765
rect 674338 111883 674366 127021
rect 674530 114177 674558 130573
rect 677108 130046 677164 130055
rect 677108 129981 677164 129990
rect 675188 129602 675244 129611
rect 675188 129537 675244 129546
rect 675092 129010 675148 129019
rect 675092 128945 675148 128954
rect 674900 127382 674956 127391
rect 674900 127317 674956 127326
rect 674804 126346 674860 126355
rect 674804 126281 674860 126290
rect 674612 124718 674668 124727
rect 674612 124653 674668 124662
rect 674518 114171 674570 114177
rect 674518 114113 674570 114119
rect 674326 111877 674378 111883
rect 674326 111819 674378 111825
rect 674626 111365 674654 124653
rect 674708 121906 674764 121915
rect 674708 121841 674764 121850
rect 674722 121281 674750 121841
rect 674710 121275 674762 121281
rect 674710 121217 674762 121223
rect 674818 120856 674846 126281
rect 674722 120828 674846 120856
rect 674614 111359 674666 111365
rect 674614 111301 674666 111307
rect 674722 111217 674750 120828
rect 674914 120708 674942 127317
rect 674996 124126 675052 124135
rect 674996 124061 675052 124070
rect 674818 120680 674942 120708
rect 674818 114843 674846 120680
rect 674806 114837 674858 114843
rect 674806 114779 674858 114785
rect 674710 111211 674762 111217
rect 674710 111153 674762 111159
rect 675010 107591 675038 124061
rect 675106 112009 675134 128945
rect 675202 115435 675230 129537
rect 677012 127826 677068 127835
rect 677012 127761 677068 127770
rect 676916 122942 676972 122951
rect 676916 122877 676972 122886
rect 676820 122350 676876 122359
rect 676820 122285 676876 122294
rect 676834 121133 676862 122285
rect 676930 121207 676958 122877
rect 676918 121201 676970 121207
rect 676918 121143 676970 121149
rect 676822 121127 676874 121133
rect 676822 121069 676874 121075
rect 677026 118067 677054 127761
rect 677012 118058 677068 118067
rect 677012 117993 677068 118002
rect 677122 117919 677150 129981
rect 677108 117910 677164 117919
rect 677108 117845 677164 117854
rect 675190 115429 675242 115435
rect 675190 115371 675242 115377
rect 675478 115429 675530 115435
rect 675478 115371 675530 115377
rect 675490 115144 675518 115371
rect 675382 114837 675434 114843
rect 675382 114779 675434 114785
rect 675394 114478 675422 114779
rect 675382 114171 675434 114177
rect 675382 114113 675434 114119
rect 675394 113812 675422 114113
rect 675106 111981 675408 112009
rect 675094 111877 675146 111883
rect 675094 111819 675146 111825
rect 675106 111458 675134 111819
rect 675106 111430 675408 111458
rect 675094 111359 675146 111365
rect 675094 111301 675146 111307
rect 675106 110169 675134 111301
rect 675382 111211 675434 111217
rect 675382 111153 675434 111159
rect 675394 110778 675422 111153
rect 675106 110141 675408 110169
rect 675380 110066 675436 110075
rect 675380 110001 675436 110010
rect 675394 109594 675422 110001
rect 675476 109326 675532 109335
rect 675476 109261 675532 109270
rect 675490 108973 675518 109261
rect 675106 108959 675518 108973
rect 675106 108945 675504 108959
rect 674998 107585 675050 107591
rect 674998 107527 675050 107533
rect 675106 106555 675134 108945
rect 675380 108142 675436 108151
rect 675380 108077 675436 108086
rect 675394 107670 675422 108077
rect 675382 107585 675434 107591
rect 675382 107527 675434 107533
rect 675394 107119 675422 107527
rect 675478 106919 675530 106925
rect 675478 106861 675530 106867
rect 675094 106549 675146 106555
rect 675094 106491 675146 106497
rect 675490 106486 675518 106861
rect 674230 106401 674282 106407
rect 674230 106343 674282 106349
rect 675382 106401 675434 106407
rect 675382 106343 675434 106349
rect 675394 105820 675422 106343
rect 665204 105182 665260 105191
rect 665122 105140 665204 105168
rect 665122 103743 665150 105140
rect 665204 105117 665260 105126
rect 675380 105182 675436 105191
rect 675380 105117 675436 105126
rect 675394 104636 675422 105117
rect 665204 104590 665260 104599
rect 665204 104525 665206 104534
rect 665258 104525 665260 104534
rect 665206 104493 665258 104499
rect 663190 103737 663242 103743
rect 663190 103679 663242 103685
rect 665110 103737 665162 103743
rect 665110 103679 665162 103685
rect 645814 100851 645866 100857
rect 645814 100793 645866 100799
rect 646102 100851 646154 100857
rect 646102 100793 646154 100799
rect 645826 100728 645854 100793
rect 645826 100700 645950 100728
rect 645716 88162 645772 88171
rect 645716 88097 645772 88106
rect 645730 87019 645758 88097
rect 645718 87013 645770 87019
rect 645718 86955 645770 86961
rect 645922 86871 645950 100700
rect 646390 92711 646442 92717
rect 646390 92653 646442 92659
rect 659830 92711 659882 92717
rect 659830 92653 659882 92659
rect 646102 92267 646154 92273
rect 646102 92209 646154 92215
rect 645718 86865 645770 86871
rect 645718 86807 645770 86813
rect 645910 86865 645962 86871
rect 645910 86807 645962 86813
rect 645730 80803 645758 86807
rect 646114 85803 646142 92209
rect 646100 85794 646156 85803
rect 646100 85729 646156 85738
rect 646294 85237 646346 85243
rect 646294 85179 646346 85185
rect 646306 85063 646334 85179
rect 646292 85054 646348 85063
rect 646292 84989 646348 84998
rect 645908 84166 645964 84175
rect 645908 84101 645964 84110
rect 645922 81839 645950 84101
rect 645910 81833 645962 81839
rect 645910 81775 645962 81781
rect 645718 80797 645770 80803
rect 645718 80739 645770 80745
rect 645814 80723 645866 80729
rect 645814 80665 645866 80671
rect 645826 49797 645854 80665
rect 646102 79169 646154 79175
rect 646102 79111 646154 79117
rect 646114 78699 646142 79111
rect 646100 78690 646156 78699
rect 646100 78625 646156 78634
rect 646402 74902 646430 92653
rect 647542 92637 647594 92643
rect 647542 92579 647594 92585
rect 647158 92563 647210 92569
rect 647158 92505 647210 92511
rect 646678 92193 646730 92199
rect 646678 92135 646730 92141
rect 646486 76949 646538 76955
rect 646484 76914 646486 76923
rect 646538 76914 646540 76923
rect 646484 76849 646540 76858
rect 646486 76801 646538 76807
rect 646486 76743 646538 76749
rect 646498 76035 646526 76743
rect 646484 76026 646540 76035
rect 646484 75961 646540 75970
rect 646402 74874 646526 74902
rect 646498 72779 646526 74874
rect 646484 72770 646540 72779
rect 646484 72705 646540 72714
rect 646690 72187 646718 92135
rect 647170 80919 647198 92505
rect 647348 87422 647404 87431
rect 647348 87357 647404 87366
rect 647156 80910 647212 80919
rect 647156 80845 647212 80854
rect 646870 78651 646922 78657
rect 646870 78593 646922 78599
rect 646882 78551 646910 78593
rect 646868 78542 646924 78551
rect 646868 78477 646924 78486
rect 647362 77769 647390 87357
rect 647554 82251 647582 92579
rect 647830 92489 647882 92495
rect 647830 92431 647882 92437
rect 647734 92341 647786 92347
rect 647734 92283 647786 92289
rect 647636 89050 647692 89059
rect 647636 88985 647692 88994
rect 647540 82242 647596 82251
rect 647540 82177 647596 82186
rect 647650 81691 647678 88985
rect 647746 85507 647774 92283
rect 647842 86247 647870 92431
rect 658870 92193 658922 92199
rect 658870 92135 658922 92141
rect 658882 87986 658910 92135
rect 659842 88000 659870 92653
rect 661750 92637 661802 92643
rect 661750 92579 661802 92585
rect 660694 92563 660746 92569
rect 660694 92505 660746 92511
rect 659842 87972 660144 88000
rect 660706 87986 660734 92505
rect 661174 92267 661226 92273
rect 661174 92209 661226 92215
rect 661186 88000 661214 92209
rect 661762 88000 661790 92579
rect 663094 92489 663146 92495
rect 663094 92431 663146 92437
rect 662518 92341 662570 92347
rect 662518 92283 662570 92289
rect 661186 87972 661440 88000
rect 661762 87972 662016 88000
rect 662530 87986 662558 92283
rect 663106 87986 663134 92431
rect 659362 87389 659616 87408
rect 651382 87383 651434 87389
rect 651382 87325 651434 87331
rect 659350 87383 659616 87389
rect 659402 87380 659616 87383
rect 659350 87325 659402 87331
rect 650998 87013 651050 87019
rect 650900 86978 650956 86987
rect 650998 86955 651050 86961
rect 650900 86913 650956 86922
rect 647828 86238 647884 86247
rect 647828 86173 647884 86182
rect 647732 85498 647788 85507
rect 647732 85433 647788 85442
rect 650914 85243 650942 86913
rect 651010 85359 651038 86955
rect 651094 86495 651146 86501
rect 651094 86437 651146 86443
rect 650996 85350 651052 85359
rect 650996 85285 651052 85294
rect 650902 85237 650954 85243
rect 650902 85179 650954 85185
rect 650996 84314 651052 84323
rect 650996 84249 651052 84258
rect 647926 83461 647978 83467
rect 647924 83426 647926 83435
rect 647978 83426 647980 83435
rect 647924 83361 647980 83370
rect 650900 82686 650956 82695
rect 650900 82621 650956 82630
rect 647924 82538 647980 82547
rect 647924 82473 647980 82482
rect 647938 81913 647966 82473
rect 647926 81907 647978 81913
rect 647926 81849 647978 81855
rect 647638 81685 647690 81691
rect 647638 81627 647690 81633
rect 647924 81354 647980 81363
rect 647924 81289 647926 81298
rect 647978 81289 647980 81298
rect 647926 81257 647978 81263
rect 647828 80466 647884 80475
rect 647828 80401 647884 80410
rect 647842 78731 647870 80401
rect 647926 80205 647978 80211
rect 647924 80170 647926 80179
rect 647978 80170 647980 80179
rect 647924 80105 647980 80114
rect 647924 79282 647980 79291
rect 647924 79217 647980 79226
rect 647830 78725 647882 78731
rect 647830 78667 647882 78673
rect 647938 78361 647966 79217
rect 647926 78355 647978 78361
rect 647926 78297 647978 78303
rect 647350 77763 647402 77769
rect 647350 77705 647402 77711
rect 647926 77689 647978 77695
rect 647924 77654 647926 77663
rect 647978 77654 647980 77663
rect 647924 77589 647980 77598
rect 647926 77319 647978 77325
rect 647926 77261 647978 77267
rect 647938 77071 647966 77261
rect 647924 77062 647980 77071
rect 647924 76997 647980 77006
rect 650914 76807 650942 82621
rect 651010 77695 651038 84249
rect 651106 83435 651134 86437
rect 651188 86238 651244 86247
rect 651188 86173 651244 86182
rect 651092 83426 651148 83435
rect 651092 83361 651148 83370
rect 651202 78657 651230 86173
rect 651394 83879 651422 87325
rect 658006 87309 658058 87315
rect 656866 87232 657792 87260
rect 658058 87257 658320 87260
rect 658006 87251 658320 87257
rect 658018 87232 658320 87251
rect 651380 83870 651436 83879
rect 651380 83805 651436 83814
rect 651190 78651 651242 78657
rect 651190 78593 651242 78599
rect 650998 77689 651050 77695
rect 650998 77631 651050 77637
rect 650902 76801 650954 76807
rect 650902 76743 650954 76749
rect 656866 75623 656894 87232
rect 657046 87161 657098 87167
rect 657046 87103 657098 87109
rect 657058 83467 657086 87103
rect 657046 83461 657098 83467
rect 657046 83403 657098 83409
rect 661078 81685 661130 81691
rect 661130 81633 661440 81636
rect 661078 81627 661440 81633
rect 661090 81608 661440 81627
rect 657538 81321 657792 81340
rect 657526 81315 657792 81321
rect 657578 81312 657792 81315
rect 657526 81257 657578 81263
rect 662900 81206 662956 81215
rect 662900 81141 662956 81150
rect 656962 81016 657216 81044
rect 656962 80211 656990 81016
rect 656950 80205 657002 80211
rect 656950 80147 657002 80153
rect 658306 76955 658334 81030
rect 658882 79175 658910 81030
rect 659602 80748 659630 81030
rect 659554 80729 659630 80748
rect 659446 80723 659498 80729
rect 659446 80665 659498 80671
rect 659542 80723 659630 80729
rect 659594 80720 659630 80723
rect 659542 80665 659594 80671
rect 658870 79169 658922 79175
rect 658870 79111 658922 79117
rect 659458 77769 659486 80665
rect 659446 77763 659498 77769
rect 659446 77705 659498 77711
rect 658294 76949 658346 76955
rect 658294 76891 658346 76897
rect 646870 75617 646922 75623
rect 646870 75559 646922 75565
rect 656854 75617 656906 75623
rect 656854 75559 656906 75565
rect 646882 75443 646910 75559
rect 646868 75434 646924 75443
rect 646868 75369 646924 75378
rect 647926 75321 647978 75327
rect 647926 75263 647978 75269
rect 647938 75147 647966 75263
rect 647924 75138 647980 75147
rect 647924 75073 647980 75082
rect 646964 74398 647020 74407
rect 646964 74333 647020 74342
rect 646978 72663 647006 74333
rect 647828 73806 647884 73815
rect 647828 73741 647884 73750
rect 646966 72657 647018 72663
rect 646966 72599 647018 72605
rect 647842 72293 647870 73741
rect 647924 73066 647980 73075
rect 647924 73001 647980 73010
rect 647938 72737 647966 73001
rect 647926 72731 647978 72737
rect 647926 72673 647978 72679
rect 660130 72293 660158 81030
rect 660706 78731 660734 81030
rect 661762 81016 662016 81044
rect 660694 78725 660746 78731
rect 660694 78667 660746 78673
rect 661762 75327 661790 81016
rect 662530 78361 662558 81030
rect 662518 78355 662570 78361
rect 662518 78297 662570 78303
rect 662914 77325 662942 81141
rect 662902 77319 662954 77325
rect 662902 77261 662954 77267
rect 661750 75321 661802 75327
rect 661750 75263 661802 75269
rect 663202 73477 663230 103679
rect 675764 103258 675820 103267
rect 675764 103193 675820 103202
rect 675778 102786 675806 103193
rect 675764 101482 675820 101491
rect 675764 101417 675820 101426
rect 675778 100936 675806 101417
rect 663286 87087 663338 87093
rect 663286 87029 663338 87035
rect 663298 85211 663326 87029
rect 663572 85646 663628 85655
rect 663572 85581 663628 85590
rect 663284 85202 663340 85211
rect 663284 85137 663340 85146
rect 663476 84758 663532 84767
rect 663476 84693 663532 84702
rect 663380 82834 663436 82843
rect 663380 82769 663436 82778
rect 663284 82094 663340 82103
rect 663284 82029 663340 82038
rect 663298 81913 663326 82029
rect 663286 81907 663338 81913
rect 663286 81849 663338 81855
rect 663394 81839 663422 82769
rect 663382 81833 663434 81839
rect 663382 81775 663434 81781
rect 663490 80156 663518 84693
rect 663298 80128 663518 80156
rect 663190 73471 663242 73477
rect 663190 73413 663242 73419
rect 663298 72737 663326 80128
rect 663586 80008 663614 85581
rect 663490 79980 663614 80008
rect 663286 72731 663338 72737
rect 663286 72673 663338 72679
rect 663490 72663 663518 79980
rect 663478 72657 663530 72663
rect 663478 72599 663530 72605
rect 647830 72287 647882 72293
rect 647830 72229 647882 72235
rect 660118 72287 660170 72293
rect 660118 72229 660170 72235
rect 646676 72178 646732 72187
rect 646676 72113 646732 72122
rect 645814 49791 645866 49797
rect 645814 49733 645866 49739
rect 645622 47645 645674 47651
rect 645622 47587 645674 47593
rect 640724 40654 640780 40663
rect 640724 40589 640780 40598
rect 443926 37433 443978 37439
rect 443926 37375 443978 37381
rect 459190 37433 459242 37439
rect 459190 37375 459242 37381
<< via2 >>
rect 148532 1015918 148588 1015974
rect 251348 1015918 251404 1015974
rect 353396 1015918 353452 1015974
rect 145364 1007926 145420 1007982
rect 148532 1007926 148588 1007982
rect 81044 995790 81100 995846
rect 81620 995642 81676 995698
rect 42164 968706 42220 968762
rect 41780 967078 41836 967134
rect 41780 965006 41836 965062
rect 42164 963970 42220 964026
rect 41780 963378 41836 963434
rect 41780 962638 41836 962694
rect 42164 962342 42220 962398
rect 41876 962194 41932 962250
rect 42452 962046 42508 962102
rect 41780 959678 41836 959734
rect 41876 959086 41932 959142
rect 41780 958494 41836 958550
rect 42164 957754 42220 957810
rect 42068 956126 42124 956182
rect 40436 942954 40492 943010
rect 40052 941918 40108 941974
rect 39956 941770 40012 941826
rect 40052 940290 40108 940346
rect 39956 939106 40012 939162
rect 35252 932594 35308 932650
rect 35252 932150 35308 932206
rect 42548 944621 42550 944638
rect 42550 944621 42602 944638
rect 42602 944621 42604 944638
rect 42548 944582 42604 944621
rect 42548 944177 42550 944194
rect 42550 944177 42602 944194
rect 42602 944177 42604 944194
rect 42548 944138 42604 944177
rect 42548 944029 42550 944046
rect 42550 944029 42602 944046
rect 42602 944029 42604 944046
rect 42548 943990 42604 944029
rect 42548 942993 42550 943010
rect 42550 942993 42602 943010
rect 42602 942993 42604 943010
rect 42548 942954 42604 942993
rect 42548 942379 42604 942418
rect 42548 942362 42550 942379
rect 42550 942362 42602 942379
rect 42602 942362 42604 942379
rect 41780 941918 41836 941974
rect 42836 937774 42892 937830
rect 42548 933186 42604 933242
rect 42548 932167 42604 932206
rect 42548 932150 42550 932167
rect 42550 932150 42602 932167
rect 42602 932150 42604 932167
rect 42548 819265 42550 819282
rect 42550 819265 42602 819282
rect 42602 819265 42604 819282
rect 42548 819226 42604 819265
rect 42836 818525 42838 818542
rect 42838 818525 42890 818542
rect 42890 818525 42892 818542
rect 42836 818486 42892 818525
rect 42548 818229 42550 818246
rect 42550 818229 42602 818246
rect 42602 818229 42604 818246
rect 42548 818190 42604 818229
rect 43220 817450 43276 817506
rect 40436 817154 40492 817210
rect 40340 816710 40396 816766
rect 41684 814934 41740 814990
rect 40244 813898 40300 813954
rect 40148 811678 40204 811734
rect 35156 806794 35212 806850
rect 35156 806350 35212 806406
rect 41492 810494 41548 810550
rect 40244 802058 40300 802114
rect 40148 801910 40204 801966
rect 41588 808866 41644 808922
rect 41492 800726 41548 800782
rect 41588 800578 41644 800634
rect 42548 814342 42604 814398
rect 41972 813306 42028 813362
rect 41876 812270 41932 812326
rect 41780 808422 41836 808478
rect 41684 800430 41740 800486
rect 41780 800282 41836 800338
rect 42068 812714 42124 812770
rect 42164 809458 42220 809514
rect 43124 811382 43180 811438
rect 42932 810346 42988 810402
rect 42164 800282 42220 800338
rect 42068 794214 42124 794270
rect 41780 793770 41836 793826
rect 42452 792142 42508 792198
rect 43028 808126 43084 808182
rect 42740 796138 42796 796194
rect 42452 791846 42508 791902
rect 42068 791106 42124 791162
rect 41780 790514 41836 790570
rect 42836 791846 42892 791902
rect 42932 791698 42988 791754
rect 42836 789330 42892 789386
rect 42740 789182 42796 789238
rect 42740 775901 42742 775918
rect 42742 775901 42794 775918
rect 42794 775901 42796 775918
rect 42740 775862 42796 775901
rect 42740 775309 42742 775326
rect 42742 775309 42794 775326
rect 42794 775309 42796 775326
rect 42740 775270 42796 775309
rect 42740 774791 42742 774808
rect 42742 774791 42794 774808
rect 42794 774791 42796 774808
rect 42740 774752 42796 774791
rect 44660 806498 44716 806554
rect 43220 774234 43276 774290
rect 42932 772014 42988 772070
rect 41972 771126 42028 771182
rect 40244 770682 40300 770738
rect 35156 763578 35212 763634
rect 35156 763134 35212 763190
rect 41492 770090 41548 770146
rect 40244 757658 40300 757714
rect 41780 769498 41836 769554
rect 41588 767426 41644 767482
rect 41492 757362 41548 757418
rect 41684 766242 41740 766298
rect 41876 769054 41932 769110
rect 41780 757214 41836 757270
rect 42068 766242 42124 766298
rect 41972 757066 42028 757122
rect 41876 754846 41932 754902
rect 43124 767130 43180 767186
rect 43028 765502 43084 765558
rect 43412 773642 43468 773698
rect 42932 751886 42988 751942
rect 42068 751738 42124 751794
rect 42932 750998 42988 751054
rect 42068 749814 42124 749870
rect 42452 749222 42508 749278
rect 41972 747742 42028 747798
rect 41780 747150 41836 747206
rect 42068 746262 42124 746318
rect 43124 747002 43180 747058
rect 43028 746854 43084 746910
rect 42836 732685 42838 732702
rect 42838 732685 42890 732702
rect 42890 732685 42892 732702
rect 42836 732646 42892 732685
rect 42836 732093 42838 732110
rect 42838 732093 42890 732110
rect 42890 732093 42892 732110
rect 42836 732054 42892 732093
rect 42836 731797 42838 731814
rect 42838 731797 42890 731814
rect 42890 731797 42892 731814
rect 42836 731758 42892 731797
rect 43700 731018 43756 731074
rect 43412 730426 43468 730482
rect 41492 728650 41548 728706
rect 35156 720362 35212 720418
rect 35156 719918 35212 719974
rect 42452 727910 42508 727966
rect 41588 726874 41644 726930
rect 41876 725838 41932 725894
rect 41684 724654 41740 724710
rect 41780 724210 41836 724266
rect 41780 713850 41836 713906
rect 41972 723618 42028 723674
rect 42068 722582 42124 722638
rect 42164 721990 42220 722046
rect 42452 721990 42508 722046
rect 43124 726282 43180 726338
rect 42068 713998 42124 714054
rect 42452 721546 42508 721602
rect 42164 713850 42220 713906
rect 43316 721990 43372 722046
rect 42452 713258 42508 713314
rect 43028 711038 43084 711094
rect 42068 708522 42124 708578
rect 41780 707930 41836 707986
rect 42740 707782 42796 707838
rect 42164 707338 42220 707394
rect 42452 705414 42508 705470
rect 41876 704674 41932 704730
rect 41780 704082 41836 704138
rect 43220 711334 43276 711390
rect 43028 703490 43084 703546
rect 42836 689469 42838 689486
rect 42838 689469 42890 689486
rect 42890 689469 42892 689486
rect 42836 689430 42892 689469
rect 42452 689134 42508 689190
rect 42452 688581 42454 688598
rect 42454 688581 42506 688598
rect 42506 688581 42508 688598
rect 42452 688542 42508 688581
rect 43700 711334 43756 711390
rect 43220 687654 43276 687710
rect 43220 687506 43276 687562
rect 41876 685434 41932 685490
rect 40244 684250 40300 684306
rect 35252 677146 35308 677202
rect 35252 676702 35308 676758
rect 41684 683658 41740 683714
rect 41588 683066 41644 683122
rect 40532 680994 40588 681050
rect 40244 673298 40300 673354
rect 40628 679810 40684 679866
rect 41492 679810 41548 679866
rect 40532 671078 40588 671134
rect 40628 670930 40684 670986
rect 41588 670930 41644 670986
rect 42452 684842 42508 684898
rect 41972 682622 42028 682678
rect 41780 670634 41836 670690
rect 42164 681438 42220 681494
rect 42068 678330 42124 678386
rect 43028 680698 43084 680754
rect 43124 679070 43180 679126
rect 43124 670782 43180 670838
rect 42740 668562 42796 668618
rect 41780 664566 41836 664622
rect 42164 664122 42220 664178
rect 42452 662790 42508 662846
rect 41780 661458 41836 661514
rect 41876 661310 41932 661366
rect 41780 660274 41836 660330
rect 43124 659090 43180 659146
rect 42164 656130 42220 656186
rect 42932 646214 42988 646270
rect 42452 645474 42508 645530
rect 42932 645217 42934 645234
rect 42934 645217 42986 645234
rect 42986 645217 42988 645234
rect 42932 645178 42988 645217
rect 43796 647102 43852 647158
rect 43604 646954 43660 647010
rect 43412 644586 43468 644642
rect 43220 644438 43276 644494
rect 41492 642218 41548 642274
rect 39860 641034 39916 641090
rect 35156 633930 35212 633986
rect 35156 633486 35212 633542
rect 40244 638814 40300 638870
rect 41300 638370 41356 638426
rect 40244 628010 40300 628066
rect 39860 627862 39916 627918
rect 42932 641922 42988 641978
rect 41588 640442 41644 640498
rect 41492 627862 41548 627918
rect 41684 639998 41740 640054
rect 41300 627714 41356 627770
rect 41588 627714 41644 627770
rect 41876 639406 41932 639462
rect 42068 636742 42124 636798
rect 41972 636150 42028 636206
rect 41972 627418 42028 627474
rect 42164 635558 42220 635614
rect 43124 638074 43180 638130
rect 43028 635558 43084 635614
rect 43796 643550 43852 643606
rect 43604 642958 43660 643014
rect 42164 623422 42220 623478
rect 43124 621498 43180 621554
rect 42452 619574 42508 619630
rect 41780 618390 41836 618446
rect 41780 618242 41836 618298
rect 41972 617798 42028 617854
rect 41780 616614 41836 616670
rect 42164 613506 42220 613562
rect 41780 612766 41836 612822
rect 42836 602998 42892 603054
rect 42740 602275 42796 602314
rect 42740 602258 42742 602275
rect 42742 602258 42794 602275
rect 42794 602258 42796 602275
rect 42164 602110 42220 602166
rect 43316 601222 43372 601278
rect 43988 601370 44044 601426
rect 43796 600334 43852 600390
rect 43604 599742 43660 599798
rect 43124 599150 43180 599206
rect 41972 598410 42028 598466
rect 41588 597226 41644 597282
rect 41492 596782 41548 596838
rect 41876 596190 41932 596246
rect 41780 595154 41836 595210
rect 41684 594562 41740 594618
rect 41588 584646 41644 584702
rect 41684 584498 41740 584554
rect 42164 593526 42220 593582
rect 42068 592934 42124 592990
rect 42068 584350 42124 584406
rect 42836 592712 42892 592768
rect 42740 588346 42796 588402
rect 42836 584498 42892 584554
rect 41972 584202 42028 584258
rect 42164 584202 42220 584258
rect 41876 581982 41932 582038
rect 41780 580206 41836 580262
rect 42068 578430 42124 578486
rect 42932 578282 42988 578338
rect 42164 577542 42220 577598
rect 42068 574878 42124 574934
rect 42068 574582 42124 574638
rect 41780 574434 41836 574490
rect 41780 573990 41836 574046
rect 43220 573102 43276 573158
rect 41780 570438 41836 570494
rect 42836 559634 42892 559690
rect 43028 559355 43084 559394
rect 43028 559338 43030 559355
rect 43030 559338 43082 559355
rect 43082 559338 43084 559355
rect 43508 559042 43564 559098
rect 42932 558746 42988 558802
rect 43412 557118 43468 557174
rect 41588 555786 41644 555842
rect 41492 554010 41548 554066
rect 41396 549718 41452 549774
rect 35156 547498 35212 547554
rect 35156 547054 35212 547110
rect 41492 541430 41548 541486
rect 41396 541282 41452 541338
rect 41876 555194 41932 555250
rect 41780 551346 41836 551402
rect 41684 549126 41740 549182
rect 41684 541282 41740 541338
rect 42164 553566 42220 553622
rect 41972 551938 42028 551994
rect 41780 540986 41836 541042
rect 42068 550310 42124 550366
rect 42452 552974 42508 553030
rect 42164 541134 42220 541190
rect 43124 550754 43180 550810
rect 42068 536990 42124 537046
rect 41780 534326 41836 534382
rect 41972 533734 42028 533790
rect 43124 548978 43180 549034
rect 43028 541578 43084 541634
rect 43028 538026 43084 538082
rect 42068 532698 42124 532754
rect 41780 531810 41836 531866
rect 41780 531218 41836 531274
rect 42932 532550 42988 532606
rect 42164 529442 42220 529498
rect 43028 530034 43084 530090
rect 43124 524114 43180 524170
rect 43316 524114 43372 524170
rect 42164 509906 42220 509962
rect 42164 503986 42220 504042
rect 42068 483710 42124 483766
rect 42068 463878 42124 463934
rect 42836 432245 42838 432262
rect 42838 432245 42890 432262
rect 42890 432245 42892 432262
rect 42836 432206 42892 432245
rect 42548 431949 42550 431966
rect 42550 431949 42602 431966
rect 42602 431949 42604 431966
rect 42548 431910 42604 431949
rect 41876 431318 41932 431374
rect 42932 430578 42988 430634
rect 42548 427618 42604 427674
rect 40244 425398 40300 425454
rect 39956 422734 40012 422790
rect 35156 419922 35212 419978
rect 35156 419478 35212 419534
rect 40148 422142 40204 422198
rect 40052 421550 40108 421606
rect 42356 423326 42412 423382
rect 42452 419478 42508 419534
rect 43220 430134 43276 430190
rect 43124 429690 43180 429746
rect 43700 558450 43756 558506
rect 43988 558006 44044 558062
rect 43796 557118 43852 557174
rect 44564 547350 44620 547406
rect 43508 428950 43564 429006
rect 43124 424066 43180 424122
rect 42932 421402 42988 421458
rect 42356 408082 42412 408138
rect 42068 406010 42124 406066
rect 42068 404234 42124 404290
rect 41780 403790 41836 403846
rect 43028 409266 43084 409322
rect 41780 402606 41836 402662
rect 41780 401866 41836 401922
rect 41780 400090 41836 400146
rect 41780 399498 41836 399554
rect 41780 398758 41836 398814
rect 42356 389325 42358 389342
rect 42358 389325 42410 389342
rect 42410 389325 42412 389342
rect 42356 389286 42412 389325
rect 42644 388733 42646 388750
rect 42646 388733 42698 388750
rect 42698 388733 42700 388750
rect 42644 388694 42700 388733
rect 42644 387993 42646 388010
rect 42646 387993 42698 388010
rect 42698 387993 42700 388010
rect 42644 387954 42700 387993
rect 43412 387214 43468 387270
rect 42932 387066 42988 387122
rect 42740 384698 42796 384754
rect 42356 382182 42412 382238
rect 39956 380554 40012 380610
rect 35156 376706 35212 376762
rect 35156 376262 35212 376318
rect 40052 380110 40108 380166
rect 40244 378334 40300 378390
rect 42644 377594 42700 377650
rect 42644 376575 42700 376614
rect 42644 376558 42646 376575
rect 42646 376558 42698 376575
rect 42698 376558 42700 376575
rect 43028 379814 43084 379870
rect 42932 378186 42988 378242
rect 41780 362794 41836 362850
rect 42164 361906 42220 361962
rect 42260 361166 42316 361222
rect 42164 360574 42220 360630
rect 42068 359390 42124 359446
rect 41780 358650 41836 358706
rect 41780 356874 41836 356930
rect 41780 356430 41836 356486
rect 41780 355542 41836 355598
rect 42836 345887 42838 345904
rect 42838 345887 42890 345904
rect 42890 345887 42892 345904
rect 42836 345848 42892 345887
rect 42836 345369 42838 345386
rect 42838 345369 42890 345386
rect 42890 345369 42892 345386
rect 42836 345330 42892 345369
rect 42836 344777 42838 344794
rect 42838 344777 42890 344794
rect 42890 344777 42892 344794
rect 42836 344738 42892 344777
rect 43412 344146 43468 344202
rect 43220 343702 43276 343758
rect 42836 341482 42892 341538
rect 41780 338966 41836 339022
rect 40052 336894 40108 336950
rect 35156 333490 35212 333546
rect 35156 333046 35212 333102
rect 40148 336302 40204 336358
rect 42260 337486 42316 337542
rect 42548 334674 42604 334730
rect 43220 333342 43276 333398
rect 42836 324758 42892 324814
rect 41780 320466 41836 320522
rect 42068 319726 42124 319782
rect 42164 318394 42220 318450
rect 42068 317950 42124 318006
rect 41780 316174 41836 316230
rect 41780 315434 41836 315490
rect 41876 313658 41932 313714
rect 41780 313214 41836 313270
rect 41780 312326 41836 312382
rect 42836 302671 42838 302688
rect 42838 302671 42890 302688
rect 42890 302671 42892 302688
rect 42836 302632 42892 302671
rect 42452 302301 42454 302318
rect 42454 302301 42506 302318
rect 42506 302301 42508 302318
rect 42452 302262 42508 302301
rect 42836 301522 42892 301578
rect 43124 300930 43180 300986
rect 43220 300486 43276 300542
rect 41780 297970 41836 298026
rect 40244 293678 40300 293734
rect 40052 293086 40108 293142
rect 39956 292494 40012 292550
rect 35156 290422 35212 290478
rect 35156 289830 35212 289886
rect 40148 292050 40204 292106
rect 42260 295750 42316 295806
rect 42356 294270 42412 294326
rect 42836 290143 42892 290182
rect 42836 290126 42838 290143
rect 42838 290126 42890 290143
rect 42890 290126 42892 290143
rect 42356 284798 42412 284854
rect 42356 281542 42412 281598
rect 42164 278582 42220 278638
rect 42068 276510 42124 276566
rect 41972 274734 42028 274790
rect 42164 274586 42220 274642
rect 41780 272958 41836 273014
rect 41780 272218 41836 272274
rect 41780 270590 41836 270646
rect 43124 270590 43180 270646
rect 41780 269998 41836 270054
rect 41780 269110 41836 269166
rect 42548 259677 42550 259694
rect 42550 259677 42602 259694
rect 42602 259677 42604 259694
rect 42548 259638 42604 259677
rect 42644 258937 42646 258954
rect 42646 258937 42698 258954
rect 42698 258937 42700 258954
rect 42644 258898 42700 258937
rect 42548 258197 42550 258214
rect 42550 258197 42602 258214
rect 42602 258197 42604 258214
rect 42548 258158 42604 258197
rect 41780 252534 41836 252590
rect 40244 250462 40300 250518
rect 39956 249870 40012 249926
rect 35252 247206 35308 247262
rect 35252 246762 35308 246818
rect 40052 249278 40108 249334
rect 40148 248834 40204 248890
rect 42548 257566 42604 257622
rect 43220 257270 43276 257326
rect 43028 255050 43084 255106
rect 42548 247798 42604 247854
rect 42548 247206 42604 247262
rect 42260 243802 42316 243858
rect 42260 240694 42316 240750
rect 42356 236550 42412 236606
rect 41780 233294 41836 233350
rect 41972 231666 42028 231722
rect 41780 231074 41836 231130
rect 43124 248538 43180 248594
rect 41780 230334 41836 230390
rect 41780 229594 41836 229650
rect 41780 229002 41836 229058
rect 41780 227374 41836 227430
rect 41780 226782 41836 226838
rect 41780 225894 41836 225950
rect 42740 216313 42742 216330
rect 42742 216313 42794 216330
rect 42794 216313 42796 216330
rect 42740 216274 42796 216313
rect 42740 215721 42742 215738
rect 42742 215721 42794 215738
rect 42794 215721 42796 215738
rect 42740 215682 42796 215721
rect 42740 215203 42742 215220
rect 42742 215203 42794 215220
rect 42794 215203 42796 215220
rect 42740 215164 42796 215203
rect 43412 256678 43468 256734
rect 43316 255790 43372 255846
rect 47444 941622 47500 941678
rect 44660 246170 44716 246226
rect 43316 242766 43372 242822
rect 43220 214054 43276 214110
rect 59444 975366 59500 975422
rect 43412 213610 43468 213666
rect 43316 213018 43372 213074
rect 41972 211538 42028 211594
rect 40244 209466 40300 209522
rect 40148 206654 40204 206710
rect 40052 206062 40108 206118
rect 35156 203990 35212 204046
rect 35156 203546 35212 203602
rect 40244 205618 40300 205674
rect 42356 209910 42412 209966
rect 42740 207690 42796 207746
rect 42932 207246 42988 207302
rect 42740 204804 42796 204860
rect 42740 203694 42796 203750
rect 42356 201178 42412 201234
rect 42164 197478 42220 197534
rect 42356 195110 42412 195166
rect 42068 190226 42124 190282
rect 41972 189042 42028 189098
rect 41780 188302 41836 188358
rect 41780 186674 41836 186730
rect 41780 185786 41836 185842
rect 43028 205322 43084 205378
rect 62036 992090 62092 992146
rect 78356 993718 78412 993774
rect 85364 995494 85420 995550
rect 84788 995346 84844 995402
rect 87764 995198 87820 995254
rect 89396 994902 89452 994958
rect 88724 993866 88780 993922
rect 104660 996547 104716 996586
rect 104660 996530 104662 996547
rect 104662 996530 104714 996547
rect 104714 996530 104716 996547
rect 94964 995790 95020 995846
rect 94964 995681 94966 995698
rect 94966 995681 95018 995698
rect 95018 995681 95020 995698
rect 94964 995642 95020 995681
rect 83444 993570 83500 993626
rect 92660 993570 92716 993626
rect 83444 992090 83500 992146
rect 62036 962342 62092 962398
rect 61844 962046 61900 962102
rect 59540 960862 59596 960918
rect 59540 946654 59596 946710
rect 59540 932150 59596 932206
rect 59540 917794 59596 917850
rect 53300 763282 53356 763338
rect 59540 903438 59596 903494
rect 59540 889082 59596 889138
rect 59540 874726 59596 874782
rect 58580 860370 58636 860426
rect 59540 846014 59596 846070
rect 59540 831658 59596 831714
rect 59540 817302 59596 817358
rect 59540 802798 59596 802854
rect 59540 788590 59596 788646
rect 59540 774086 59596 774142
rect 59540 759730 59596 759786
rect 53492 720066 53548 720122
rect 59540 745522 59596 745578
rect 59540 731018 59596 731074
rect 59540 716662 59596 716718
rect 59540 702306 59596 702362
rect 59540 687950 59596 688006
rect 53684 676850 53740 676906
rect 59540 673594 59596 673650
rect 59540 659238 59596 659294
rect 59540 644882 59596 644938
rect 56084 633930 56140 633986
rect 53780 590566 53836 590622
rect 59540 630526 59596 630582
rect 59540 616170 59596 616226
rect 59540 601853 59542 601870
rect 59542 601853 59594 601870
rect 59594 601853 59596 601870
rect 59540 601814 59596 601853
rect 59540 587458 59596 587514
rect 59540 572954 59596 573010
rect 59540 558911 59596 558950
rect 59540 558894 59542 558911
rect 59542 558894 59594 558911
rect 59594 558894 59596 558911
rect 59540 544390 59596 544446
rect 59540 530034 59596 530090
rect 59540 515678 59596 515734
rect 59540 501191 59596 501230
rect 59540 501174 59542 501191
rect 59542 501174 59594 501191
rect 59594 501174 59596 501191
rect 58580 486818 58636 486874
rect 59540 472462 59596 472518
rect 59540 458106 59596 458162
rect 59540 443750 59596 443806
rect 59540 429394 59596 429450
rect 58388 415038 58444 415094
rect 57620 400682 57676 400738
rect 59252 386326 59308 386382
rect 59540 371822 59596 371878
rect 59540 357614 59596 357670
rect 58388 343110 58444 343166
rect 57812 328754 57868 328810
rect 58004 314546 58060 314602
rect 59444 300042 59500 300098
rect 58100 285834 58156 285890
rect 53684 246466 53740 246522
rect 53300 246318 53356 246374
rect 99764 995938 99820 995994
rect 102836 995955 102892 995994
rect 102836 995938 102838 995955
rect 102838 995938 102890 995955
rect 102890 995938 102892 995955
rect 98036 995790 98092 995846
rect 100724 995790 100780 995846
rect 101204 995829 101206 995846
rect 101206 995829 101258 995846
rect 101258 995829 101260 995846
rect 101204 995790 101260 995829
rect 102452 995790 102508 995846
rect 103988 995807 104044 995846
rect 103988 995790 103990 995807
rect 103990 995790 104042 995807
rect 104042 995790 104044 995807
rect 102356 995659 102412 995698
rect 108980 995977 108982 995994
rect 108982 995977 109034 995994
rect 109034 995977 109036 995994
rect 108980 995938 109036 995977
rect 109556 995938 109612 995994
rect 107924 995790 107980 995846
rect 102356 995642 102358 995659
rect 102358 995642 102410 995659
rect 102410 995642 102412 995659
rect 105332 995642 105388 995698
rect 105908 995642 105964 995698
rect 107540 995642 107596 995698
rect 97940 995050 97996 995106
rect 106772 995198 106828 995254
rect 106772 993718 106828 993774
rect 109172 995642 109228 995698
rect 109364 995494 109420 995550
rect 110132 995642 110188 995698
rect 129716 994014 129772 994070
rect 133652 995494 133708 995550
rect 132788 994458 132844 994514
rect 126644 993570 126700 993626
rect 136148 994162 136204 994218
rect 140756 994310 140812 994366
rect 134324 993718 134380 993774
rect 140372 993718 140428 993774
rect 160436 1003207 160492 1003246
rect 160436 1003190 160438 1003207
rect 160438 1003190 160490 1003207
rect 160490 1003190 160492 1003207
rect 161492 1003153 161548 1003209
rect 153332 1002615 153388 1002654
rect 153332 1002598 153334 1002615
rect 153334 1002598 153386 1002615
rect 153386 1002598 153388 1002615
rect 151604 1002467 151660 1002506
rect 151604 1002450 151606 1002467
rect 151606 1002450 151658 1002467
rect 151658 1002450 151660 1002467
rect 152660 1002489 152662 1002506
rect 152662 1002489 152714 1002506
rect 152714 1002489 152716 1002506
rect 152660 1002450 152716 1002489
rect 151028 1002341 151030 1002358
rect 151030 1002341 151082 1002358
rect 151082 1002341 151084 1002358
rect 151028 1002302 151084 1002341
rect 155540 999381 155542 999398
rect 155542 999381 155594 999398
rect 155594 999381 155596 999398
rect 155540 999342 155596 999381
rect 159188 996251 159244 996290
rect 159188 996234 159190 996251
rect 159190 996234 159242 996251
rect 159242 996234 159244 996251
rect 159764 996103 159820 996142
rect 159764 996086 159766 996103
rect 159766 996086 159818 996103
rect 159818 996086 159820 996103
rect 156596 995938 156652 995994
rect 160436 995977 160438 995994
rect 160438 995977 160490 995994
rect 160490 995977 160492 995994
rect 160436 995938 160492 995977
rect 154868 995807 154924 995846
rect 154868 995790 154870 995807
rect 154870 995790 154922 995807
rect 154922 995790 154924 995807
rect 146804 995237 146806 995254
rect 146806 995237 146858 995254
rect 146858 995237 146860 995254
rect 146804 995198 146860 995237
rect 149684 995346 149740 995402
rect 149684 994458 149740 994514
rect 156404 995198 156460 995254
rect 156116 994310 156172 994366
rect 161492 995790 161548 995846
rect 157268 995346 157324 995402
rect 161684 995198 161740 995254
rect 213812 1005114 213868 1005170
rect 218804 1005153 218806 1005170
rect 218806 1005153 218858 1005170
rect 218858 1005153 218860 1005170
rect 218804 1005114 218860 1005153
rect 183764 995790 183820 995846
rect 192500 995790 192556 995846
rect 209108 1003207 209164 1003246
rect 209108 1003190 209110 1003207
rect 209110 1003190 209162 1003207
rect 209162 1003190 209164 1003207
rect 211796 1003207 211852 1003246
rect 211796 1003190 211798 1003207
rect 211798 1003190 211850 1003207
rect 211850 1003190 211852 1003207
rect 195284 995790 195340 995846
rect 189428 995494 189484 995550
rect 187316 994014 187372 994070
rect 206900 999381 206902 999398
rect 206902 999381 206954 999398
rect 206954 999381 206956 999398
rect 206900 999342 206956 999381
rect 205172 996547 205228 996586
rect 205172 996530 205174 996547
rect 205174 996530 205226 996547
rect 205226 996530 205228 996547
rect 207956 996547 208012 996586
rect 207956 996530 207958 996547
rect 207958 996530 208010 996547
rect 208010 996530 208012 996547
rect 210164 996103 210220 996142
rect 210164 996086 210166 996103
rect 210166 996086 210218 996103
rect 210218 996086 210220 996103
rect 204020 995938 204076 995994
rect 210644 995977 210646 995994
rect 210646 995977 210698 995994
rect 210698 995977 210700 995994
rect 210644 995938 210700 995977
rect 211796 995955 211852 995994
rect 211796 995938 211798 995955
rect 211798 995938 211850 995955
rect 211850 995938 211852 995955
rect 219092 995938 219148 995994
rect 203060 995790 203116 995846
rect 203636 995790 203692 995846
rect 204692 995807 204748 995846
rect 204692 995790 204694 995807
rect 204694 995790 204746 995807
rect 204746 995790 204748 995807
rect 197204 995642 197260 995698
rect 186164 993570 186220 993626
rect 195476 993570 195532 993626
rect 213332 995790 213388 995846
rect 208724 995346 208780 995402
rect 198644 995198 198700 995254
rect 209780 995198 209836 995254
rect 216020 995642 216076 995698
rect 239540 995790 239596 995846
rect 240788 995642 240844 995698
rect 232148 994458 232204 994514
rect 234356 994162 234412 994218
rect 235796 994606 235852 994662
rect 240212 995346 240268 995402
rect 241748 995198 241804 995254
rect 243860 995494 243916 995550
rect 250484 995790 250540 995846
rect 250100 995494 250156 995550
rect 250100 995050 250156 995106
rect 247604 994606 247660 994662
rect 247508 994458 247564 994514
rect 243188 994014 243244 994070
rect 348884 1007778 348940 1007834
rect 353300 1007778 353356 1007834
rect 316436 1003190 316492 1003246
rect 258356 999381 258358 999398
rect 258358 999381 258410 999398
rect 258410 999381 258412 999398
rect 258356 999342 258412 999381
rect 270644 997122 270700 997178
rect 298100 997139 298156 997178
rect 298100 997122 298102 997139
rect 298102 997122 298154 997139
rect 298154 997122 298156 997139
rect 262484 996399 262540 996438
rect 262484 996382 262486 996399
rect 262486 996382 262538 996399
rect 262538 996382 262540 996399
rect 257780 996103 257836 996142
rect 257780 996086 257782 996103
rect 257782 996086 257834 996103
rect 257834 996086 257836 996103
rect 262004 996103 262060 996142
rect 262004 996086 262006 996103
rect 262006 996086 262058 996103
rect 262058 996086 262060 996103
rect 263060 996125 263062 996142
rect 263062 996125 263114 996142
rect 263114 996125 263116 996142
rect 263060 996086 263116 996125
rect 254516 995955 254572 995994
rect 254516 995938 254518 995955
rect 254518 995938 254570 995955
rect 254570 995938 254572 995955
rect 254900 995938 254956 995994
rect 261044 995938 261100 995994
rect 263252 995977 263254 995994
rect 263254 995977 263306 995994
rect 263306 995977 263308 995994
rect 263252 995938 263308 995977
rect 256148 995790 256204 995846
rect 257108 995790 257164 995846
rect 259220 995790 259276 995846
rect 255956 995659 256012 995698
rect 255956 995642 255958 995659
rect 255958 995642 256010 995659
rect 256010 995642 256012 995659
rect 259028 995494 259084 995550
rect 256148 995198 256204 995254
rect 260084 995198 260140 995254
rect 259220 994162 259276 994218
rect 270740 995790 270796 995846
rect 267860 995642 267916 995698
rect 267956 995494 268012 995550
rect 287924 995790 287980 995846
rect 286772 995642 286828 995698
rect 308852 1002911 308908 1002950
rect 308852 1002894 308854 1002911
rect 308854 1002894 308906 1002911
rect 308906 1002894 308908 1002911
rect 312116 1002933 312118 1002950
rect 312118 1002933 312170 1002950
rect 312170 1002933 312172 1002950
rect 312116 1002894 312172 1002933
rect 287444 995494 287500 995550
rect 286004 994458 286060 994514
rect 291476 995198 291532 995254
rect 298964 995642 299020 995698
rect 296660 994310 296716 994366
rect 294548 994162 294604 994218
rect 308276 1002763 308332 1002802
rect 308276 1002746 308278 1002763
rect 308278 1002746 308330 1002763
rect 308330 1002746 308332 1002763
rect 309332 1002785 309334 1002802
rect 309334 1002785 309386 1002802
rect 309386 1002785 309388 1002802
rect 309332 1002746 309388 1002785
rect 309908 999381 309910 999398
rect 309910 999381 309962 999398
rect 309962 999381 309964 999398
rect 309908 999342 309964 999381
rect 314804 997879 314860 997918
rect 314804 997862 314806 997879
rect 314806 997862 314858 997879
rect 314858 997862 314860 997879
rect 313748 997139 313804 997178
rect 313748 997122 313750 997139
rect 313750 997122 313802 997139
rect 313802 997122 313804 997139
rect 311540 996547 311596 996586
rect 311540 996530 311542 996547
rect 311542 996530 311594 996547
rect 311594 996530 311596 996547
rect 299540 996086 299596 996142
rect 299348 995790 299404 995846
rect 303956 995938 304012 995994
rect 304340 995938 304396 995994
rect 305492 995938 305548 995994
rect 305972 995790 306028 995846
rect 307604 995790 307660 995846
rect 299252 995494 299308 995550
rect 299540 995494 299596 995550
rect 313172 996103 313228 996142
rect 313172 996086 313174 996103
rect 313174 996086 313226 996103
rect 313226 996086 313228 996103
rect 314804 996125 314806 996142
rect 314806 996125 314858 996142
rect 314858 996125 314860 996142
rect 314804 996086 314860 996125
rect 310292 995938 310348 995994
rect 319604 995938 319660 995994
rect 312788 995346 312844 995402
rect 319700 995642 319756 995698
rect 357428 1003207 357484 1003246
rect 357428 1003190 357430 1003207
rect 357430 1003190 357482 1003207
rect 357482 1003190 357484 1003207
rect 362516 1003207 362572 1003246
rect 362516 1003190 362518 1003207
rect 362518 1003190 362570 1003207
rect 362570 1003190 362572 1003207
rect 358580 1002763 358636 1002802
rect 358580 1002746 358582 1002763
rect 358582 1002746 358634 1002763
rect 358634 1002746 358636 1002763
rect 358004 1002637 358006 1002654
rect 358006 1002637 358058 1002654
rect 358058 1002637 358060 1002654
rect 358004 1002598 358060 1002637
rect 361844 1002489 361846 1002506
rect 361846 1002489 361898 1002506
rect 361898 1002489 361900 1002506
rect 361844 1002450 361900 1002489
rect 359060 1002319 359116 1002358
rect 359060 1002302 359062 1002319
rect 359062 1002302 359114 1002319
rect 359114 1002302 359116 1002319
rect 362900 1002341 362902 1002358
rect 362902 1002341 362954 1002358
rect 362954 1002341 362956 1002358
rect 362900 1002302 362956 1002341
rect 361364 1002193 361366 1002210
rect 361366 1002193 361418 1002210
rect 361418 1002193 361420 1002210
rect 361364 1002154 361420 1002193
rect 356372 1001283 356428 1001322
rect 356372 1001266 356374 1001283
rect 356374 1001266 356426 1001283
rect 356426 1001266 356428 1001283
rect 357044 1001118 357100 1001174
rect 359636 1000839 359692 1000878
rect 359636 1000822 359638 1000839
rect 359638 1000822 359690 1000839
rect 359690 1000822 359692 1000839
rect 360212 1000861 360214 1000878
rect 360214 1000861 360266 1000878
rect 360266 1000861 360268 1000878
rect 360212 1000822 360268 1000861
rect 364532 999359 364588 999398
rect 364532 999342 364534 999359
rect 364534 999342 364586 999359
rect 364586 999342 364588 999359
rect 365204 997879 365260 997918
rect 365204 997862 365206 997879
rect 365206 997862 365258 997879
rect 365258 997862 365260 997879
rect 363956 995977 363958 995994
rect 363958 995977 364010 995994
rect 364010 995977 364012 995994
rect 363956 995938 364012 995977
rect 360884 995807 360940 995846
rect 360884 995790 360886 995807
rect 360886 995790 360938 995807
rect 360938 995790 360940 995807
rect 366164 995790 366220 995846
rect 366740 995807 366796 995846
rect 366740 995790 366742 995807
rect 366742 995790 366794 995807
rect 366794 995790 366796 995807
rect 371540 995790 371596 995846
rect 368660 995642 368716 995698
rect 383060 995642 383116 995698
rect 383540 995790 383596 995846
rect 428660 1003207 428716 1003246
rect 428660 1003190 428662 1003207
rect 428662 1003190 428714 1003207
rect 428714 1003190 428716 1003207
rect 425396 1003081 425398 1003098
rect 425398 1003081 425450 1003098
rect 425450 1003081 425452 1003098
rect 425396 1003042 425452 1003081
rect 428276 1003059 428332 1003098
rect 428276 1003042 428278 1003059
rect 428278 1003042 428330 1003059
rect 428330 1003042 428332 1003059
rect 423860 1002911 423916 1002950
rect 423860 1002894 423862 1002911
rect 423862 1002894 423914 1002911
rect 423914 1002894 423916 1002911
rect 426068 1002933 426070 1002950
rect 426070 1002933 426122 1002950
rect 426122 1002933 426124 1002950
rect 426068 1002894 426124 1002933
rect 424340 1002785 424342 1002802
rect 424342 1002785 424394 1002802
rect 424394 1002785 424396 1002802
rect 424340 1002746 424396 1002785
rect 424820 1002763 424876 1002802
rect 424820 1002746 424822 1002763
rect 424822 1002746 424874 1002763
rect 424874 1002746 424876 1002763
rect 427604 1002637 427606 1002654
rect 427606 1002637 427658 1002654
rect 427658 1002637 427660 1002654
rect 427604 1002598 427660 1002637
rect 426644 1002489 426646 1002506
rect 426646 1002489 426698 1002506
rect 426698 1002489 426700 1002506
rect 426644 1002450 426700 1002489
rect 427124 1002467 427180 1002506
rect 427124 1002450 427126 1002467
rect 427126 1002450 427178 1002467
rect 427178 1002450 427180 1002467
rect 430292 1003059 430348 1003098
rect 430292 1003042 430294 1003059
rect 430294 1003042 430346 1003059
rect 430346 1003042 430348 1003059
rect 432020 1002785 432022 1002802
rect 432022 1002785 432074 1002802
rect 432074 1002785 432076 1002802
rect 432020 1002746 432076 1002785
rect 429236 1002615 429292 1002654
rect 435284 1006298 435340 1006354
rect 465620 1006298 465676 1006354
rect 435188 1006002 435244 1006058
rect 435092 1005854 435148 1005910
rect 429236 1002598 429238 1002615
rect 429238 1002598 429290 1002615
rect 429290 1002598 429292 1002615
rect 429908 1000839 429964 1000878
rect 429908 1000822 429910 1000839
rect 429910 1000822 429962 1000839
rect 429962 1000822 429964 1000839
rect 430964 1000861 430966 1000878
rect 430966 1000861 431018 1000878
rect 431018 1000861 431020 1000878
rect 430964 1000822 431020 1000861
rect 432500 996234 432556 996290
rect 432500 996125 432502 996142
rect 432502 996125 432554 996142
rect 432554 996125 432556 996142
rect 432500 996086 432556 996125
rect 465236 1005854 465292 1005910
rect 421556 995938 421612 995994
rect 430964 995977 430966 995994
rect 430966 995977 431018 995994
rect 431018 995977 431020 995994
rect 430964 995938 431020 995977
rect 437876 995938 437932 995994
rect 387476 995790 387532 995846
rect 391796 995642 391852 995698
rect 385940 995198 385996 995254
rect 377300 994754 377356 994810
rect 373364 994458 373420 994514
rect 377300 994310 377356 994366
rect 390836 994754 390892 994810
rect 396308 995198 396364 995254
rect 395156 994458 395212 994514
rect 403124 993587 403180 993626
rect 403124 993570 403126 993587
rect 403126 993570 403178 993587
rect 403178 993570 403180 993587
rect 437780 995642 437836 995698
rect 437972 995494 438028 995550
rect 466100 1006002 466156 1006058
rect 465620 995494 465676 995550
rect 466100 995346 466156 995402
rect 472052 995642 472108 995698
rect 502388 1003207 502444 1003246
rect 502388 1003190 502390 1003207
rect 502390 1003190 502442 1003207
rect 502442 1003190 502444 1003207
rect 501332 1003059 501388 1003098
rect 501332 1003042 501334 1003059
rect 501334 1003042 501386 1003059
rect 501386 1003042 501388 1003059
rect 502964 1003059 503020 1003098
rect 502964 1003042 502966 1003059
rect 502966 1003042 503018 1003059
rect 503018 1003042 503020 1003059
rect 472244 995790 472300 995846
rect 478388 995790 478444 995846
rect 482036 995642 482092 995698
rect 477044 995494 477100 995550
rect 477716 995346 477772 995402
rect 479828 994458 479884 994514
rect 479156 993570 479212 993626
rect 506324 1000987 506380 1001026
rect 506324 1000970 506326 1000987
rect 506326 1000970 506378 1000987
rect 506378 1000970 506380 1000987
rect 507860 1000839 507916 1000878
rect 507860 1000822 507862 1000839
rect 507862 1000822 507914 1000839
rect 507914 1000822 507916 1000839
rect 506900 1000691 506956 1000730
rect 506900 1000674 506902 1000691
rect 506902 1000674 506954 1000691
rect 506954 1000674 506956 1000691
rect 504692 999825 504694 999842
rect 504694 999825 504746 999842
rect 504746 999825 504748 999842
rect 504692 999786 504748 999825
rect 512084 999825 512086 999842
rect 512086 999825 512138 999842
rect 512138 999825 512140 999842
rect 512084 999786 512140 999825
rect 500756 999655 500812 999694
rect 500756 999638 500758 999655
rect 500758 999638 500810 999655
rect 500810 999638 500812 999655
rect 503636 999677 503638 999694
rect 503638 999677 503690 999694
rect 503690 999677 503692 999694
rect 503636 999638 503692 999677
rect 502004 999507 502060 999546
rect 502004 999490 502006 999507
rect 502006 999490 502058 999507
rect 502058 999490 502060 999507
rect 503636 999529 503638 999546
rect 503638 999529 503690 999546
rect 503690 999529 503692 999546
rect 503636 999490 503692 999529
rect 512084 999655 512140 999694
rect 512084 999638 512086 999655
rect 512086 999638 512138 999655
rect 512138 999638 512140 999655
rect 515540 1000230 515596 1000286
rect 512660 1000082 512716 1000138
rect 512276 999934 512332 999990
rect 512180 999490 512236 999546
rect 512084 999342 512140 999398
rect 505748 996547 505804 996586
rect 505748 996530 505750 996547
rect 505750 996530 505802 996547
rect 505802 996530 505804 996547
rect 507476 996569 507478 996586
rect 507478 996569 507530 996586
rect 507530 996569 507532 996586
rect 507476 996530 507532 996569
rect 508916 996103 508972 996142
rect 508916 996086 508918 996103
rect 508918 996086 508970 996103
rect 508970 996086 508972 996103
rect 509588 996125 509590 996142
rect 509590 996125 509642 996142
rect 509642 996125 509644 996142
rect 509588 996086 509644 996125
rect 508340 995977 508342 995994
rect 508342 995977 508394 995994
rect 508394 995977 508396 995994
rect 508340 995938 508396 995977
rect 499316 995790 499372 995846
rect 515540 995938 515596 995994
rect 509972 995642 510028 995698
rect 499316 995494 499372 995550
rect 501812 995494 501868 995550
rect 510260 995533 510262 995550
rect 510262 995533 510314 995550
rect 510314 995533 510316 995550
rect 510260 995494 510316 995533
rect 489140 993570 489196 993626
rect 515636 995642 515692 995698
rect 515732 995494 515788 995550
rect 555380 1003059 555436 1003098
rect 555380 1003042 555382 1003059
rect 555382 1003042 555434 1003059
rect 555434 1003042 555436 1003059
rect 553748 1002911 553804 1002950
rect 553748 1002894 553750 1002911
rect 553750 1002894 553802 1002911
rect 553802 1002894 553804 1002911
rect 554324 1002933 554326 1002950
rect 554326 1002933 554378 1002950
rect 554378 1002933 554380 1002950
rect 554324 1002894 554380 1002933
rect 554900 1002763 554956 1002802
rect 554900 1002746 554902 1002763
rect 554902 1002746 554954 1002763
rect 554954 1002746 554956 1002763
rect 553268 1002615 553324 1002654
rect 553268 1002598 553270 1002615
rect 553270 1002598 553322 1002615
rect 553322 1002598 553324 1002615
rect 552308 1000839 552364 1000878
rect 552308 1000822 552310 1000839
rect 552310 1000822 552362 1000839
rect 552362 1000822 552364 1000839
rect 523508 1000230 523564 1000286
rect 519860 996086 519916 996142
rect 519764 995938 519820 995994
rect 519668 995494 519724 995550
rect 523604 1000082 523660 1000138
rect 523508 995642 523564 995698
rect 518324 994606 518380 994662
rect 523700 999934 523756 999990
rect 523988 999786 524044 999842
rect 523796 999638 523852 999694
rect 523700 995790 523756 995846
rect 523892 999490 523948 999546
rect 524084 999342 524140 999398
rect 552884 999342 552940 999398
rect 558836 999233 558838 999250
rect 558838 999233 558890 999250
rect 558890 999233 558892 999250
rect 558836 999194 558892 999233
rect 557204 998789 557206 998806
rect 557206 998789 557258 998806
rect 557258 998789 557260 998806
rect 557204 998750 557260 998789
rect 555956 997879 556012 997918
rect 555956 997862 555958 997879
rect 555958 997862 556010 997879
rect 556010 997862 556012 997879
rect 558164 997753 558166 997770
rect 558166 997753 558218 997770
rect 558218 997753 558220 997770
rect 558164 997714 558220 997753
rect 557780 997605 557782 997622
rect 557782 997605 557834 997622
rect 557834 997605 557836 997622
rect 557780 997566 557836 997605
rect 559412 997583 559468 997622
rect 559412 997566 559414 997583
rect 559414 997566 559466 997583
rect 559466 997566 559468 997583
rect 561044 996125 561046 996142
rect 561046 996125 561098 996142
rect 561098 996125 561100 996142
rect 561044 996086 561100 996125
rect 528404 995790 528460 995846
rect 532820 995790 532876 995846
rect 550484 995790 550540 995846
rect 556532 995807 556588 995846
rect 556532 995790 556534 995807
rect 556534 995790 556586 995807
rect 556586 995790 556588 995807
rect 527828 995642 527884 995698
rect 533396 995642 533452 995698
rect 558932 995642 558988 995698
rect 559604 995659 559660 995698
rect 559604 995642 559606 995659
rect 559606 995642 559658 995659
rect 559658 995642 559660 995659
rect 535316 995494 535372 995550
rect 534356 994606 534412 994662
rect 531188 994458 531244 994514
rect 533684 993866 533740 993922
rect 536756 993866 536812 993922
rect 550484 995494 550540 995550
rect 560180 995642 560236 995698
rect 567284 995346 567340 995402
rect 569972 995790 570028 995846
rect 569876 995642 569932 995698
rect 569780 995494 569836 995550
rect 625940 995790 625996 995846
rect 629588 995790 629644 995846
rect 627668 995198 627724 995254
rect 573908 994754 573964 994810
rect 573716 994606 573772 994662
rect 634292 994754 634348 994810
rect 633044 994458 633100 994514
rect 639188 994606 639244 994662
rect 640532 993866 640588 993922
rect 643316 994162 643372 994218
rect 641108 993718 641164 993774
rect 70580 272514 70636 272570
rect 71732 272366 71788 272422
rect 69428 272070 69484 272126
rect 74132 272218 74188 272274
rect 72980 271330 73036 271386
rect 76532 272662 76588 272718
rect 78932 272810 78988 272866
rect 77780 270886 77836 270942
rect 65108 246022 65164 246078
rect 80468 246614 80524 246670
rect 81332 272958 81388 273014
rect 83636 273402 83692 273458
rect 86036 273106 86092 273162
rect 82580 271182 82636 271238
rect 88436 273550 88492 273606
rect 90836 271922 90892 271978
rect 87188 271034 87244 271090
rect 86516 246614 86572 246670
rect 93236 271774 93292 271830
rect 96788 271626 96844 271682
rect 100340 271478 100396 271534
rect 54740 242766 54796 242822
rect 106580 242618 106636 242674
rect 126644 242618 126700 242674
rect 126836 242618 126892 242674
rect 138260 242618 138316 242674
rect 54836 242470 54892 242526
rect 95060 242487 95116 242526
rect 95060 242470 95062 242487
rect 95062 242470 95114 242487
rect 95114 242470 95116 242487
rect 144020 242322 144076 242378
rect 146036 240546 146092 240602
rect 144116 238622 144172 238678
rect 142484 237586 142540 237642
rect 144020 236271 144076 236310
rect 144020 236254 144022 236271
rect 144022 236254 144074 236271
rect 144074 236254 144076 236271
rect 144020 233590 144076 233646
rect 144116 232110 144172 232166
rect 144020 231370 144076 231426
rect 144212 230186 144268 230242
rect 144116 228410 144172 228466
rect 144020 227818 144076 227874
rect 144404 223674 144460 223730
rect 144404 220122 144460 220178
rect 149588 245726 149644 245782
rect 146228 236846 146284 236902
rect 146132 225006 146188 225062
rect 146516 235070 146572 235126
rect 144404 215238 144460 215294
rect 145364 214498 145420 214554
rect 145268 211686 145324 211742
rect 144020 203250 144076 203306
rect 144500 199550 144556 199606
rect 144020 198975 144076 199014
rect 144020 198958 144022 198975
rect 144022 198958 144074 198975
rect 144074 198958 144076 198975
rect 144692 197774 144748 197830
rect 144596 196590 144652 196646
rect 144404 194814 144460 194870
rect 144308 192890 144364 192946
rect 144020 191706 144076 191762
rect 144020 188154 144076 188210
rect 41780 184158 41836 184214
rect 41780 183566 41836 183622
rect 41780 182826 41836 182882
rect 144020 184454 144076 184510
rect 144212 183270 144268 183326
rect 144020 181790 144076 181846
rect 144116 180458 144172 180514
rect 144020 178573 144022 178590
rect 144022 178573 144074 178590
rect 144074 178573 144076 178590
rect 144020 178534 144076 178573
rect 144020 176758 144076 176814
rect 144116 174390 144172 174446
rect 144020 173354 144076 173410
rect 144020 171282 144076 171338
rect 144020 167582 144076 167638
rect 144020 157518 144076 157574
rect 144212 163586 144268 163642
rect 144116 146862 144172 146918
rect 144020 145974 144076 146030
rect 144020 143162 144076 143218
rect 144020 142422 144076 142478
rect 144020 140942 144076 140998
rect 144020 138574 144076 138630
rect 144020 134726 144076 134782
rect 144020 132802 144076 132858
rect 144116 131026 144172 131082
rect 144020 130138 144076 130194
rect 144020 129250 144076 129306
rect 39860 125293 39862 125310
rect 39862 125293 39914 125310
rect 39914 125293 39916 125310
rect 39860 125254 39916 125293
rect 144116 125106 144172 125162
rect 144020 124366 144076 124422
rect 144116 122738 144172 122794
rect 144020 121554 144076 121610
rect 141044 118594 141100 118650
rect 144116 120814 144172 120870
rect 141044 118298 141100 118354
rect 144020 118315 144076 118354
rect 144020 118298 144022 118315
rect 144022 118298 144074 118315
rect 144074 118298 144076 118315
rect 144020 114154 144076 114210
rect 144116 113118 144172 113174
rect 144020 112395 144076 112434
rect 144020 112378 144022 112395
rect 144022 112378 144074 112395
rect 144074 112378 144076 112395
rect 144116 111194 144172 111250
rect 144020 109714 144076 109770
rect 144020 107494 144076 107550
rect 143924 106902 143980 106958
rect 144020 105866 144076 105922
rect 144308 159886 144364 159942
rect 144308 139462 144364 139518
rect 144308 133986 144364 134042
rect 144116 104682 144172 104738
rect 144020 104255 144076 104294
rect 144020 104238 144022 104255
rect 144022 104238 144074 104255
rect 144074 104238 144076 104255
rect 144116 102758 144172 102814
rect 144020 101591 144076 101630
rect 144020 101574 144022 101591
rect 144022 101574 144074 101591
rect 144074 101574 144076 101591
rect 144212 99798 144268 99854
rect 144116 99058 144172 99114
rect 144020 98061 144022 98078
rect 144022 98061 144074 98078
rect 144074 98061 144076 98078
rect 144020 98022 144076 98061
rect 144116 96246 144172 96302
rect 144020 95506 144076 95562
rect 144116 94322 144172 94378
rect 144020 92842 144076 92898
rect 144212 91362 144268 91418
rect 144116 90770 144172 90826
rect 144020 89586 144076 89642
rect 144116 87070 144172 87126
rect 144020 85886 144076 85942
rect 144020 82334 144076 82390
rect 144116 79374 144172 79430
rect 144020 78634 144076 78690
rect 144116 77450 144172 77506
rect 144020 75674 144076 75730
rect 144020 73898 144076 73954
rect 144116 72714 144172 72770
rect 144020 71234 144076 71290
rect 144020 69754 144076 69810
rect 144020 67682 144076 67738
rect 144020 65462 144076 65518
rect 144020 62650 144076 62706
rect 144020 59581 144022 59598
rect 144022 59581 144074 59598
rect 144074 59581 144076 59598
rect 144020 59542 144076 59581
rect 144020 58654 144076 58710
rect 144020 57065 144022 57082
rect 144022 57065 144074 57082
rect 144074 57065 144076 57082
rect 144020 57026 144076 57065
rect 144020 56138 144076 56194
rect 144020 54675 144076 54714
rect 144020 54658 144022 54675
rect 144022 54658 144074 54675
rect 144074 54658 144076 54675
rect 144020 53770 144076 53826
rect 144212 66350 144268 66406
rect 144500 154410 144556 154466
rect 144500 151598 144556 151654
rect 144500 149674 144556 149730
rect 144500 126734 144556 126790
rect 144404 80706 144460 80762
rect 144884 179718 144940 179774
rect 144692 166546 144748 166602
rect 145268 176018 145324 176074
rect 145172 172022 145228 172078
rect 144980 170098 145036 170154
rect 144884 164770 144940 164826
rect 144692 162846 144748 162902
rect 144788 161366 144844 161422
rect 144692 159294 144748 159350
rect 144692 156334 144748 156390
rect 144692 108234 144748 108290
rect 144596 106606 144652 106662
rect 144692 83518 144748 83574
rect 145076 168322 145132 168378
rect 144884 64761 144886 64778
rect 144886 64761 144938 64778
rect 144938 64761 144940 64778
rect 144884 64722 144940 64761
rect 145460 210502 145516 210558
rect 145556 207986 145612 208042
rect 145652 205618 145708 205674
rect 145748 205026 145804 205082
rect 145844 202066 145900 202122
rect 145748 201326 145804 201382
rect 145940 193630 145996 193686
rect 146036 190078 146092 190134
rect 146228 189338 146284 189394
rect 146132 186378 146188 186434
rect 146420 185194 146476 185250
rect 146804 226634 146860 226690
rect 146804 222934 146860 222990
rect 146708 221750 146764 221806
rect 146804 218198 146860 218254
rect 146804 213314 146860 213370
rect 146612 209762 146668 209818
rect 146804 207411 146860 207450
rect 146804 207394 146806 207411
rect 146806 207394 146858 207411
rect 146858 207394 146860 207411
rect 146132 135170 146188 135226
rect 146132 126734 146188 126790
rect 146228 106754 146284 106810
rect 146228 106458 146284 106514
rect 146036 76414 146092 76470
rect 146420 87810 146476 87866
rect 146516 75970 146572 76026
rect 146516 69014 146572 69070
rect 146900 155633 146902 155650
rect 146902 155633 146954 155650
rect 146954 155633 146956 155650
rect 146900 155594 146956 155633
rect 146804 152930 146860 152986
rect 146804 150858 146860 150914
rect 146804 147898 146860 147954
rect 146708 144198 146764 144254
rect 146708 135614 146764 135670
rect 146996 136075 147052 136114
rect 146996 136058 146998 136075
rect 146998 136058 147050 136075
rect 147050 136058 147052 136075
rect 146708 127474 146764 127530
rect 146900 119055 146956 119094
rect 146900 119038 146902 119055
rect 146902 119038 146954 119055
rect 146954 119038 146956 119055
rect 146708 84110 146764 84166
rect 146900 116687 146956 116726
rect 146900 116670 146902 116687
rect 146902 116670 146954 116687
rect 146954 116670 146956 116687
rect 146900 115947 146956 115986
rect 146900 115930 146902 115947
rect 146902 115930 146954 115947
rect 146954 115930 146956 115947
rect 147092 126899 147148 126938
rect 147092 126882 147094 126899
rect 147094 126882 147146 126899
rect 147146 126882 147148 126899
rect 146900 75082 146956 75138
rect 146900 62354 146956 62410
rect 146900 60726 146956 60782
rect 152468 237734 152524 237790
rect 155348 245430 155404 245486
rect 158324 245134 158380 245190
rect 161108 244986 161164 245042
rect 163988 247650 164044 247706
rect 166868 246910 166924 246966
rect 161108 137538 161164 137594
rect 175508 247502 175564 247558
rect 172724 246614 172780 246670
rect 171380 242618 171436 242674
rect 168404 48738 168460 48794
rect 171284 48590 171340 48646
rect 178388 243506 178444 243562
rect 175700 242361 175702 242378
rect 175702 242361 175754 242378
rect 175754 242361 175756 242378
rect 175700 242322 175756 242361
rect 174164 48442 174220 48498
rect 165524 48146 165580 48202
rect 181268 247354 181324 247410
rect 181364 247058 181420 247114
rect 181364 245874 181420 245930
rect 187028 247206 187084 247262
rect 187220 247650 187276 247706
rect 187220 247058 187276 247114
rect 190004 245874 190060 245930
rect 191444 238770 191500 238826
rect 182804 48294 182860 48350
rect 201524 270590 201580 270646
rect 206036 276954 206092 277010
rect 196916 247650 196972 247706
rect 196916 247354 196972 247410
rect 196916 247206 196972 247262
rect 197396 247502 197452 247558
rect 197012 247058 197068 247114
rect 197300 246466 197356 246522
rect 196724 246318 196780 246374
rect 196916 246318 196972 246374
rect 197204 246170 197260 246226
rect 197204 245578 197260 245634
rect 197588 246318 197644 246374
rect 197588 245874 197644 245930
rect 197300 245282 197356 245338
rect 196724 244838 196780 244894
rect 195764 242470 195820 242526
rect 204596 232554 204652 232610
rect 204692 232110 204748 232166
rect 204500 231518 204556 231574
rect 204788 230926 204844 230982
rect 204980 227670 205036 227726
rect 211508 268222 211564 268278
rect 207188 261266 207244 261322
rect 207092 249278 207148 249334
rect 205268 232554 205324 232610
rect 206612 244542 206668 244598
rect 205460 230482 205516 230538
rect 205364 226634 205420 226690
rect 205556 226042 205612 226098
rect 205172 225598 205228 225654
rect 204500 223970 204556 224026
rect 204596 223378 204652 223434
rect 204692 222786 204748 222842
rect 204788 221750 204844 221806
rect 204500 221158 204556 221214
rect 204596 221010 204652 221066
rect 204692 220122 204748 220178
rect 204788 219530 204844 219586
rect 204884 219382 204940 219438
rect 204500 218494 204556 218550
rect 204596 217902 204652 217958
rect 204692 217754 204748 217810
rect 204788 216866 204844 216922
rect 204500 215830 204556 215886
rect 204596 215238 204652 215294
rect 201716 92250 201772 92306
rect 204500 102018 204556 102074
rect 204596 101574 204652 101630
rect 204692 100982 204748 101038
rect 204596 100390 204652 100446
rect 204500 100242 204556 100298
rect 204692 99354 204748 99410
rect 204788 98762 204844 98818
rect 204884 98614 204940 98670
rect 204500 97765 204502 97782
rect 204502 97765 204554 97782
rect 204554 97765 204556 97782
rect 204500 97726 204556 97765
rect 204500 97134 204556 97190
rect 204596 96986 204652 97042
rect 204788 96098 204844 96154
rect 204692 95506 204748 95562
rect 204596 94766 204652 94822
rect 204500 94470 204556 94526
rect 205268 93878 205324 93934
rect 204788 93730 204844 93786
rect 204692 92842 204748 92898
rect 204500 91954 204556 92010
rect 204500 90622 204556 90678
rect 204596 90030 204652 90086
rect 205364 91214 205420 91270
rect 204692 89586 204748 89642
rect 204500 88994 204556 89050
rect 204596 88402 204652 88458
rect 204692 87958 204748 88014
rect 204788 87366 204844 87422
rect 204884 86774 204940 86830
rect 204500 86330 204556 86386
rect 204500 85738 204556 85794
rect 204596 85146 204652 85202
rect 204692 84702 204748 84758
rect 204788 84110 204844 84166
rect 204884 83518 204940 83574
rect 204500 83074 204556 83130
rect 204596 82482 204652 82538
rect 204500 81890 204556 81946
rect 204692 81446 204748 81502
rect 204788 80854 204844 80910
rect 204500 78634 204556 78690
rect 205460 80114 205516 80170
rect 204692 79226 204748 79282
rect 204596 78486 204652 78542
rect 204596 77598 204652 77654
rect 204500 77006 204556 77062
rect 204692 76858 204748 76914
rect 204788 75970 204844 76026
rect 204884 75378 204940 75434
rect 204980 75230 205036 75286
rect 204500 74342 204556 74398
rect 204596 73750 204652 73806
rect 204692 73602 204748 73658
rect 204788 72714 204844 72770
rect 204884 72122 204940 72178
rect 204500 71695 204556 71734
rect 204500 71678 204502 71695
rect 204502 71678 204554 71695
rect 204554 71678 204556 71695
rect 204596 71086 204652 71142
rect 204692 70494 204748 70550
rect 204788 69902 204844 69958
rect 204884 69458 204940 69514
rect 204500 68866 204556 68922
rect 204596 68274 204652 68330
rect 204692 67830 204748 67886
rect 204788 67238 204844 67294
rect 204884 66646 204940 66702
rect 204596 66202 204652 66258
rect 204500 65610 204556 65666
rect 204692 65018 204748 65074
rect 204500 64574 204556 64630
rect 204596 63982 204652 64038
rect 204500 63407 204556 63446
rect 204500 63390 204502 63407
rect 204502 63390 204554 63407
rect 204554 63390 204556 63407
rect 204596 62946 204652 63002
rect 204692 62354 204748 62410
rect 204500 60726 204556 60782
rect 204884 61762 204940 61818
rect 204788 61318 204844 61374
rect 204596 60134 204652 60190
rect 204500 59986 204556 60042
rect 204692 59098 204748 59154
rect 205748 227226 205804 227282
rect 205940 228262 205996 228318
rect 206132 229298 206188 229354
rect 205748 211982 205804 212038
rect 206324 214646 206380 214702
rect 206228 214498 206284 214554
rect 206420 213610 206476 213666
rect 206900 244542 206956 244598
rect 206900 243358 206956 243414
rect 206900 227374 206956 227430
rect 206900 225006 206956 225062
rect 207284 255346 207340 255402
rect 208724 247650 208780 247706
rect 210356 247058 210412 247114
rect 210164 246762 210220 246818
rect 210260 246466 210316 246522
rect 210356 246318 210412 246374
rect 210356 246022 210412 246078
rect 210356 245765 210358 245782
rect 210358 245765 210410 245782
rect 210410 245765 210412 245782
rect 210356 245726 210412 245765
rect 210356 245578 210412 245634
rect 210260 245282 210316 245338
rect 210164 245134 210220 245190
rect 210068 244986 210124 245042
rect 209972 244838 210028 244894
rect 209972 243654 210028 243710
rect 210452 243654 210508 243710
rect 210356 243210 210412 243266
rect 210260 243062 210316 243118
rect 210644 242322 210700 242378
rect 208532 239066 208588 239122
rect 209876 239066 209932 239122
rect 209588 237586 209644 237642
rect 208052 230926 208108 230982
rect 207092 227374 207148 227430
rect 206996 224414 207052 224470
rect 206804 222342 206860 222398
rect 206708 216274 206764 216330
rect 206612 213018 206668 213074
rect 206516 212870 206572 212926
rect 205844 211390 205900 211446
rect 207092 202658 207148 202714
rect 206900 80262 206956 80318
rect 206900 55842 206956 55898
rect 207284 229890 207340 229946
rect 207284 57470 207340 57526
rect 209204 232110 209260 232166
rect 209492 231518 209548 231574
rect 209396 230482 209452 230538
rect 209300 56582 209356 56638
rect 209780 236994 209836 237050
rect 209684 236846 209740 236902
rect 210164 234774 210220 234830
rect 210164 228854 210220 228910
rect 211700 271034 211756 271090
rect 211988 271182 212044 271238
rect 212276 267926 212332 267982
rect 211508 242174 211564 242230
rect 211412 241878 211468 241934
rect 249812 273994 249868 274050
rect 250676 274142 250732 274198
rect 250292 268074 250348 268130
rect 252404 274438 252460 274494
rect 251828 274290 251884 274346
rect 252020 268370 252076 268426
rect 254132 274734 254188 274790
rect 253940 274586 253996 274642
rect 253364 269110 253420 269166
rect 252884 268666 252940 268722
rect 255860 268518 255916 268574
rect 254612 268222 254668 268278
rect 255092 267778 255148 267834
rect 256820 273698 256876 273754
rect 256628 267778 256684 267834
rect 257588 278434 257644 278490
rect 368564 278582 368620 278638
rect 259412 273254 259468 273310
rect 258932 270442 258988 270498
rect 261620 274882 261676 274938
rect 260660 270738 260716 270794
rect 260564 268962 260620 269018
rect 261140 269702 261196 269758
rect 262004 269850 262060 269906
rect 262868 276362 262924 276418
rect 264404 275474 264460 275530
rect 263348 273846 263404 273902
rect 263732 267926 263788 267982
rect 265940 275326 265996 275382
rect 265460 271034 265516 271090
rect 264884 269554 264940 269610
rect 265076 268222 265132 268278
rect 266612 269406 266668 269462
rect 267092 275178 267148 275234
rect 267188 275030 267244 275086
rect 269396 276066 269452 276122
rect 268148 269998 268204 270054
rect 267668 269258 267724 269314
rect 267764 267778 267820 267834
rect 269204 267926 269260 267982
rect 276212 267778 276268 267834
rect 293972 278434 294028 278490
rect 299540 278434 299596 278490
rect 299732 278451 299788 278490
rect 299732 278434 299734 278451
rect 299734 278434 299786 278451
rect 299786 278434 299788 278451
rect 300404 278451 300460 278490
rect 300404 278434 300406 278451
rect 300406 278434 300458 278451
rect 300458 278434 300460 278451
rect 315284 278434 315340 278490
rect 299540 278325 299542 278342
rect 299542 278325 299594 278342
rect 299594 278325 299596 278342
rect 299540 278286 299596 278325
rect 300308 278325 300310 278342
rect 300310 278325 300362 278342
rect 300362 278325 300364 278342
rect 300308 278286 300364 278325
rect 303380 278286 303436 278342
rect 298004 268518 298060 268574
rect 299636 277842 299692 277898
rect 299540 277694 299596 277750
rect 298004 267926 298060 267982
rect 297812 267778 297868 267834
rect 298196 267926 298252 267982
rect 298388 267778 298444 267834
rect 300404 277842 300460 277898
rect 300308 277694 300364 277750
rect 304532 278138 304588 278194
rect 305204 277990 305260 278046
rect 306356 277842 306412 277898
rect 307124 277694 307180 277750
rect 308372 277546 308428 277602
rect 309524 277398 309580 277454
rect 310964 277250 311020 277306
rect 312308 277102 312364 277158
rect 314420 270015 314476 270054
rect 314420 269998 314422 270015
rect 314422 269998 314474 270015
rect 314474 269998 314476 270015
rect 315284 270886 315340 270942
rect 315860 267926 315916 267982
rect 316724 268814 316780 268870
rect 317492 270590 317548 270646
rect 317684 270590 317740 270646
rect 317684 268518 317740 268574
rect 318644 276214 318700 276270
rect 317876 268518 317932 268574
rect 317876 267926 317932 267982
rect 318164 270294 318220 270350
rect 318068 269850 318124 269906
rect 318068 267926 318124 267982
rect 319796 275918 319852 275974
rect 318932 270146 318988 270202
rect 319700 269850 319756 269906
rect 320852 275770 320908 275826
rect 320180 269998 320236 270054
rect 321908 276806 321964 276862
rect 322868 275622 322924 275678
rect 324692 276510 324748 276566
rect 324500 271182 324556 271238
rect 325556 276658 325612 276714
rect 325460 276066 325516 276122
rect 325652 276066 325708 276122
rect 325268 270886 325324 270942
rect 325268 270590 325324 270646
rect 325460 270590 325516 270646
rect 267860 264818 267916 264874
rect 276500 264818 276556 264874
rect 308084 264818 308140 264874
rect 325748 267926 325804 267982
rect 327188 269850 327244 269906
rect 327092 267926 327148 267982
rect 328628 271182 328684 271238
rect 328436 270886 328492 270942
rect 329012 270886 329068 270942
rect 328436 269850 328492 269906
rect 332564 270886 332620 270942
rect 336884 271051 336940 271090
rect 336884 271034 336886 271051
rect 336886 271034 336938 271051
rect 336938 271034 336940 271051
rect 336212 267965 336214 267982
rect 336214 267965 336266 267982
rect 336266 267965 336268 267982
rect 336212 267926 336268 267965
rect 336404 267926 336460 267982
rect 338708 270294 338764 270350
rect 338036 269850 338092 269906
rect 339188 270886 339244 270942
rect 348692 272514 348748 272570
rect 348692 271182 348748 271238
rect 358676 272366 358732 272422
rect 358676 272070 358732 272126
rect 383828 278582 383884 278638
rect 368852 278434 368908 278490
rect 369044 271922 369100 271978
rect 369044 271034 369100 271090
rect 370388 271626 370444 271682
rect 370484 270442 370540 270498
rect 370676 270442 370732 270498
rect 370868 270442 370924 270498
rect 371444 270442 371500 270498
rect 371732 270442 371788 270498
rect 371252 268962 371308 269018
rect 371444 268962 371500 269018
rect 372788 272070 372844 272126
rect 373364 274882 373420 274938
rect 372980 273550 373036 273606
rect 373172 273550 373228 273606
rect 373172 272958 373228 273014
rect 373364 272958 373420 273014
rect 372980 270886 373036 270942
rect 374132 276362 374188 276418
rect 374324 276362 374380 276418
rect 373844 271330 373900 271386
rect 375668 273402 375724 273458
rect 375860 273402 375916 273458
rect 375860 272810 375916 272866
rect 376148 272662 376204 272718
rect 376340 272070 376396 272126
rect 378260 276954 378316 277010
rect 377300 273106 377356 273162
rect 377300 272070 377356 272126
rect 377108 268222 377164 268278
rect 377396 267778 377452 267834
rect 378068 274882 378124 274938
rect 378452 276954 378508 277010
rect 378068 273698 378124 273754
rect 378260 273698 378316 273754
rect 378068 273106 378124 273162
rect 378356 270886 378412 270942
rect 378548 270886 378604 270942
rect 378548 270442 378604 270498
rect 378836 270442 378892 270498
rect 379220 270442 379276 270498
rect 379412 270442 379468 270498
rect 379988 272070 380044 272126
rect 380180 272070 380236 272126
rect 380564 271626 380620 271682
rect 379796 268962 379852 269018
rect 379988 268962 380044 269018
rect 380276 268962 380332 269018
rect 383060 276954 383116 277010
rect 383252 276954 383308 277010
rect 382676 274882 382732 274938
rect 383252 274882 383308 274938
rect 382196 273550 382252 273606
rect 381236 272366 381292 272422
rect 382004 272514 382060 272570
rect 382196 272514 382252 272570
rect 381428 272366 381484 272422
rect 381332 271626 381388 271682
rect 381620 271182 381676 271238
rect 381908 271221 381910 271238
rect 381910 271221 381962 271238
rect 381962 271221 381964 271238
rect 381908 271182 381964 271221
rect 382964 273846 383020 273902
rect 382964 273550 383020 273606
rect 382868 271626 382924 271682
rect 383060 271626 383116 271682
rect 383348 272810 383404 272866
rect 383252 272218 383308 272274
rect 383444 271182 383500 271238
rect 384404 273402 384460 273458
rect 384884 272514 384940 272570
rect 378932 264855 378988 264911
rect 385364 273402 385420 273458
rect 387668 272958 387724 273014
rect 387572 272810 387628 272866
rect 385940 272366 385996 272422
rect 385556 271182 385612 271238
rect 386420 271182 386476 271238
rect 386612 272218 386668 272274
rect 387476 271034 387532 271090
rect 387668 271034 387724 271090
rect 397460 278451 397516 278490
rect 397460 278434 397462 278451
rect 397462 278434 397514 278451
rect 397514 278434 397516 278451
rect 417428 278451 417484 278490
rect 417428 278434 417430 278451
rect 417430 278434 417482 278451
rect 417482 278434 417484 278451
rect 428852 278434 428908 278490
rect 429044 278434 429100 278490
rect 440660 278473 440662 278490
rect 440662 278473 440714 278490
rect 440714 278473 440716 278490
rect 440660 278434 440716 278473
rect 489620 278473 489622 278490
rect 489622 278473 489674 278490
rect 489674 278473 489676 278490
rect 489620 278434 489676 278473
rect 495380 278473 495382 278490
rect 495382 278473 495434 278490
rect 495434 278473 495436 278490
rect 495380 278434 495436 278473
rect 501332 278473 501334 278490
rect 501334 278473 501386 278490
rect 501386 278473 501388 278490
rect 501332 278434 501388 278473
rect 525524 278451 525580 278490
rect 525524 278434 525526 278451
rect 525526 278434 525578 278451
rect 525578 278434 525580 278451
rect 551252 278451 551308 278490
rect 551252 278434 551254 278451
rect 551254 278434 551306 278451
rect 551306 278434 551308 278451
rect 610484 278451 610540 278490
rect 610484 278434 610486 278451
rect 610486 278434 610538 278451
rect 610538 278434 610540 278451
rect 610772 278451 610828 278490
rect 610772 278434 610774 278451
rect 610774 278434 610826 278451
rect 610826 278434 610828 278451
rect 625076 278473 625078 278490
rect 625078 278473 625130 278490
rect 625130 278473 625132 278490
rect 625076 278434 625132 278473
rect 631028 278473 631030 278490
rect 631030 278473 631082 278490
rect 631082 278473 631084 278490
rect 631028 278434 631084 278473
rect 467540 278286 467596 278342
rect 389684 272366 389740 272422
rect 388148 271922 388204 271978
rect 389588 271922 389644 271978
rect 389396 271774 389452 271830
rect 388724 271182 388780 271238
rect 388628 270442 388684 270498
rect 388820 270442 388876 270498
rect 388724 268222 388780 268278
rect 388916 268222 388972 268278
rect 388820 267778 388876 267834
rect 389012 267778 389068 267834
rect 389300 267778 389356 267834
rect 390836 271774 390892 271830
rect 389876 271478 389932 271534
rect 392468 272070 392524 272126
rect 394100 272958 394156 273014
rect 393140 272810 393196 272866
rect 393812 270738 393868 270794
rect 394292 272514 394348 272570
rect 394484 271073 394486 271090
rect 394486 271073 394538 271090
rect 394538 271073 394540 271090
rect 394484 271034 394540 271073
rect 394484 270886 394540 270942
rect 395156 271478 395212 271534
rect 474740 278138 474796 278194
rect 481844 277990 481900 278046
rect 646004 277990 646060 278046
rect 396692 276954 396748 277010
rect 397364 273567 397420 273606
rect 397364 273550 397366 273567
rect 397366 273550 397418 273567
rect 397418 273550 397420 273567
rect 395828 272662 395884 272718
rect 395636 270738 395692 270794
rect 395924 270738 395980 270794
rect 397364 273106 397420 273162
rect 397556 273106 397612 273162
rect 396980 272514 397036 272570
rect 396884 271182 396940 271238
rect 397556 272366 397612 272422
rect 397268 271626 397324 271682
rect 397844 270886 397900 270942
rect 397556 267778 397612 267834
rect 398420 272514 398476 272570
rect 399476 271034 399532 271090
rect 379124 264818 379180 264874
rect 385076 264855 385132 264911
rect 400148 272366 400204 272422
rect 401876 271626 401932 271682
rect 401204 270738 401260 270794
rect 403124 273846 403180 273902
rect 402740 272070 402796 272126
rect 403700 268222 403756 268278
rect 403892 268222 403948 268278
rect 404852 268222 404908 268278
rect 405716 268222 405772 268278
rect 406100 268222 406156 268278
rect 407060 271626 407116 271682
rect 407060 271182 407116 271238
rect 408596 272662 408652 272718
rect 408500 272514 408556 272570
rect 408404 272366 408460 272422
rect 408596 272070 408652 272126
rect 408500 271774 408556 271830
rect 408404 271626 408460 271682
rect 406484 264855 406540 264911
rect 407252 264855 407308 264911
rect 407732 264855 407788 264911
rect 408116 264855 408172 264911
rect 408788 264855 408844 264911
rect 409556 264855 409612 264911
rect 410804 264855 410860 264911
rect 411188 264855 411244 264911
rect 412148 247206 412204 247262
rect 223124 246762 223180 246818
rect 224852 246762 224908 246818
rect 225332 246762 225388 246818
rect 212276 238918 212332 238974
rect 211892 236550 211948 236606
rect 211316 236402 211372 236458
rect 210164 161514 210220 161570
rect 210164 158406 210220 158462
rect 210164 141534 210220 141590
rect 210164 138426 210220 138482
rect 210164 129102 210220 129158
rect 210164 126142 210220 126198
rect 210164 121110 210220 121166
rect 210164 113710 210220 113766
rect 211796 233442 211852 233498
rect 212276 236254 212332 236310
rect 212180 233590 212236 233646
rect 212660 236698 212716 236754
rect 212372 235070 212428 235126
rect 212564 233442 212620 233498
rect 212852 233442 212908 233498
rect 213236 243654 213292 243710
rect 214100 234922 214156 234978
rect 214964 243210 215020 243266
rect 215828 238178 215884 238234
rect 215252 238030 215308 238086
rect 214868 237882 214924 237938
rect 214772 237586 214828 237642
rect 214772 236550 214828 236606
rect 214292 233442 214348 233498
rect 216212 237586 216268 237642
rect 217172 243062 217228 243118
rect 216692 237734 216748 237790
rect 218900 242914 218956 242970
rect 218228 235218 218284 235274
rect 219764 235662 219820 235718
rect 220820 242766 220876 242822
rect 221396 242026 221452 242082
rect 221972 242618 222028 242674
rect 221300 235514 221356 235570
rect 223988 242509 223990 242526
rect 223990 242509 224042 242526
rect 224042 242509 224044 242526
rect 223988 242470 224044 242509
rect 223508 242174 223564 242230
rect 223700 242174 223756 242230
rect 223028 235366 223084 235422
rect 228116 246762 228172 246818
rect 228308 246762 228364 246818
rect 228596 246762 228652 246818
rect 224468 235810 224524 235866
rect 227060 243671 227116 243710
rect 227060 243654 227062 243671
rect 227062 243654 227114 243671
rect 227114 243654 227116 243671
rect 227060 243062 227116 243118
rect 227348 243654 227404 243710
rect 227348 243210 227404 243266
rect 227348 242914 227404 242970
rect 227636 242783 227692 242822
rect 227636 242766 227638 242783
rect 227638 242766 227690 242783
rect 227690 242766 227692 242783
rect 227540 242618 227596 242674
rect 227732 242657 227734 242674
rect 227734 242657 227786 242674
rect 227786 242657 227788 242674
rect 227732 242618 227788 242657
rect 227252 242322 227308 242378
rect 227540 242322 227596 242378
rect 227636 242174 227692 242230
rect 225812 236106 225868 236162
rect 227444 238178 227500 238234
rect 227636 238030 227692 238086
rect 227444 236994 227500 237050
rect 227636 236698 227692 236754
rect 246164 246762 246220 246818
rect 246452 246762 246508 246818
rect 247316 246762 247372 246818
rect 247796 246762 247852 246818
rect 229556 235958 229612 236014
rect 231668 242914 231724 242970
rect 238196 234330 238252 234386
rect 238676 234478 238732 234534
rect 239060 238030 239116 238086
rect 239060 236737 239062 236754
rect 239062 236737 239114 236754
rect 239114 236737 239116 236754
rect 239060 236698 239116 236737
rect 240980 240398 241036 240454
rect 241364 238178 241420 238234
rect 241940 242339 241996 242378
rect 241940 242322 241942 242339
rect 241942 242322 241994 242339
rect 241994 242322 241996 242339
rect 241748 240546 241804 240602
rect 242324 242339 242380 242378
rect 242324 242322 242326 242339
rect 242326 242322 242378 242339
rect 242378 242322 242380 242339
rect 242324 238474 242380 238530
rect 243188 240990 243244 241046
rect 242708 240694 242764 240750
rect 243092 237290 243148 237346
rect 243572 238622 243628 238678
rect 244532 241138 244588 241194
rect 243956 237438 244012 237494
rect 245396 241730 245452 241786
rect 245300 237142 245356 237198
rect 246740 241582 246796 241638
rect 247316 242509 247318 242526
rect 247318 242509 247370 242526
rect 247370 242509 247372 242526
rect 247316 242470 247372 242509
rect 248180 246779 248236 246818
rect 248180 246762 248182 246779
rect 248182 246762 248234 246779
rect 248234 246762 248236 246779
rect 248372 246762 248428 246818
rect 247796 242470 247852 242526
rect 247700 240102 247756 240158
rect 260948 246762 261004 246818
rect 269204 246762 269260 246818
rect 247988 239954 248044 240010
rect 259028 240842 259084 240898
rect 258644 238326 258700 238382
rect 259124 238030 259180 238086
rect 259604 239806 259660 239862
rect 259124 236737 259126 236754
rect 259126 236737 259178 236754
rect 259178 236737 259180 236754
rect 259124 236698 259180 236737
rect 261236 241286 261292 241342
rect 262964 240250 263020 240306
rect 267956 243654 268012 243710
rect 268244 242914 268300 242970
rect 267764 242470 267820 242526
rect 267956 242470 268012 242526
rect 267956 241730 268012 241786
rect 267668 241434 267724 241490
rect 267572 241286 267628 241342
rect 267764 241286 267820 241342
rect 267764 239806 267820 239862
rect 267956 239658 268012 239714
rect 281300 246762 281356 246818
rect 284948 246779 285004 246818
rect 284948 246762 284950 246779
rect 284950 246762 285002 246779
rect 285002 246762 285004 246779
rect 277556 240398 277612 240454
rect 278132 241138 278188 241194
rect 277748 240990 277804 241046
rect 278036 240694 278092 240750
rect 277556 239806 277612 239862
rect 278132 239658 278188 239714
rect 278804 239510 278860 239566
rect 280244 239510 280300 239566
rect 285236 246762 285292 246818
rect 287540 246762 287596 246818
rect 283412 234182 283468 234238
rect 307412 246762 307468 246818
rect 307892 246762 307948 246818
rect 285044 239658 285100 239714
rect 284948 234034 285004 234090
rect 287636 242914 287692 242970
rect 287252 239510 287308 239566
rect 287828 242470 287884 242526
rect 288116 243654 288172 243710
rect 288308 243654 288364 243710
rect 288020 242470 288076 242526
rect 288116 239658 288172 239714
rect 289652 241730 289708 241786
rect 289652 241138 289708 241194
rect 289076 236994 289132 237050
rect 289844 241138 289900 241194
rect 289844 240694 289900 240750
rect 289940 233886 289996 233942
rect 289844 233442 289900 233498
rect 290708 236271 290764 236310
rect 290708 236254 290710 236271
rect 290710 236254 290762 236271
rect 290762 236254 290764 236271
rect 292244 239214 292300 239270
rect 293108 239362 293164 239418
rect 293780 239658 293836 239714
rect 293780 239510 293836 239566
rect 294068 236254 294124 236310
rect 295604 241138 295660 241194
rect 295892 240990 295948 241046
rect 295700 239214 295756 239270
rect 295796 233886 295852 233942
rect 296084 233442 296140 233498
rect 298196 243210 298252 243266
rect 297908 243062 297964 243118
rect 298004 240398 298060 240454
rect 298004 239806 298060 239862
rect 298388 234182 298444 234238
rect 299156 234034 299212 234090
rect 301076 239658 301132 239714
rect 305300 239362 305356 239418
rect 307700 242470 307756 242526
rect 308084 246762 308140 246818
rect 311156 246762 311212 246818
rect 307892 243210 307948 243266
rect 308084 243210 308140 243266
rect 308084 242766 308140 242822
rect 308276 242805 308278 242822
rect 308278 242805 308330 242822
rect 308330 242805 308332 242822
rect 308276 242766 308332 242805
rect 307892 242470 307948 242526
rect 328340 246762 328396 246818
rect 312788 236994 312844 237050
rect 319700 238030 319756 238086
rect 319700 236994 319756 237050
rect 319700 236698 319756 236754
rect 328532 246762 328588 246818
rect 328916 246762 328972 246818
rect 329300 246762 329356 246818
rect 342548 246762 342604 246818
rect 348596 246762 348652 246818
rect 349076 246762 349132 246818
rect 349652 246762 349708 246818
rect 366452 246762 366508 246818
rect 366836 246762 366892 246818
rect 367316 246762 367372 246818
rect 369524 246762 369580 246818
rect 328340 242914 328396 242970
rect 328532 242914 328588 242970
rect 328436 242766 328492 242822
rect 328724 242657 328726 242674
rect 328726 242657 328778 242674
rect 328778 242657 328780 242674
rect 328724 242618 328780 242657
rect 334964 235070 335020 235126
rect 338132 242914 338188 242970
rect 338516 243062 338572 243118
rect 338516 242026 338572 242082
rect 338804 242026 338860 242082
rect 338996 242618 339052 242674
rect 339188 242618 339244 242674
rect 339764 238030 339820 238086
rect 339764 236994 339820 237050
rect 339764 236698 339820 236754
rect 341204 242766 341260 242822
rect 341108 235218 341164 235274
rect 342068 242322 342124 242378
rect 341588 235662 341644 235718
rect 342932 242174 342988 242230
rect 342740 238069 342742 238086
rect 342742 238069 342794 238086
rect 342794 238069 342796 238086
rect 342740 238030 342796 238069
rect 342548 235514 342604 235570
rect 343412 242618 343468 242674
rect 343316 235366 343372 235422
rect 344276 242026 344332 242082
rect 343796 235810 343852 235866
rect 344756 236106 344812 236162
rect 346004 235958 346060 236014
rect 347732 234330 347788 234386
rect 348212 234922 348268 234978
rect 349172 234478 349228 234534
rect 351284 239954 351340 240010
rect 351380 239066 351436 239122
rect 352244 242766 352300 242822
rect 352820 240102 352876 240158
rect 354644 243062 354700 243118
rect 354452 241582 354508 241638
rect 356756 241730 356812 241786
rect 357812 237142 357868 237198
rect 358964 241138 359020 241194
rect 359252 236550 359308 236606
rect 360020 237438 360076 237494
rect 360692 238622 360748 238678
rect 361652 240990 361708 241046
rect 363092 240694 363148 240750
rect 362708 237290 362764 237346
rect 363860 238474 363916 238530
rect 364820 240546 364876 240602
rect 365780 238178 365836 238234
rect 366548 240398 366604 240454
rect 367604 240398 367660 240454
rect 370292 246762 370348 246818
rect 370676 246762 370732 246818
rect 373460 246762 373516 246818
rect 389012 246762 389068 246818
rect 389300 246762 389356 246818
rect 390260 246762 390316 246818
rect 369812 240250 369868 240306
rect 372884 241434 372940 241490
rect 370004 238069 370006 238086
rect 370006 238069 370058 238086
rect 370058 238069 370060 238086
rect 370004 238030 370060 238069
rect 376820 241286 376876 241342
rect 377876 240842 377932 240898
rect 378836 238326 378892 238382
rect 379412 234774 379468 234830
rect 380180 236809 380236 236865
rect 383060 239658 383116 239714
rect 383540 240694 383596 240750
rect 383060 239066 383116 239122
rect 383060 238030 383116 238086
rect 388916 243358 388972 243414
rect 388916 243062 388972 243118
rect 405908 246762 405964 246818
rect 406100 246779 406156 246818
rect 406100 246762 406102 246779
rect 406102 246762 406154 246779
rect 406154 246762 406156 246779
rect 390164 236715 390220 236754
rect 390164 236698 390166 236715
rect 390166 236698 390218 236715
rect 390218 236698 390220 236715
rect 393140 237882 393196 237938
rect 394676 237734 394732 237790
rect 398708 243506 398764 243562
rect 398612 240694 398668 240750
rect 406388 246762 406444 246818
rect 406580 246725 406636 246781
rect 406772 246762 406828 246818
rect 406964 246779 407020 246818
rect 406964 246762 406966 246779
rect 406966 246762 407018 246779
rect 407018 246762 407020 246779
rect 406004 243506 406060 243562
rect 407348 246762 407404 246818
rect 407732 246762 407788 246818
rect 408116 246762 408172 246818
rect 408308 246762 408364 246818
rect 408980 246779 409036 246818
rect 408980 246762 408982 246779
rect 408982 246762 409034 246779
rect 409034 246762 409036 246779
rect 410324 246762 410380 246818
rect 410516 246762 410572 246818
rect 410804 246762 410860 246818
rect 411188 246762 411244 246818
rect 411380 246762 411436 246818
rect 411764 246762 411820 246818
rect 409748 240398 409804 240454
rect 413108 267778 413164 267834
rect 413300 267817 413302 267834
rect 413302 267817 413354 267834
rect 413354 267817 413356 267834
rect 413300 267778 413356 267817
rect 412820 265449 412822 265466
rect 412822 265449 412874 265466
rect 412874 265449 412876 265466
rect 412820 265410 412876 265449
rect 413108 265558 413164 265614
rect 412916 265262 412972 265318
rect 412724 265114 412780 265170
rect 412628 264983 412684 265022
rect 412628 264966 412630 264983
rect 412630 264966 412682 264983
rect 412682 264966 412684 264983
rect 417332 273587 417388 273643
rect 413396 265854 413452 265910
rect 429140 270738 429196 270794
rect 428948 269998 429004 270054
rect 429236 269998 429292 270054
rect 429044 269850 429100 269906
rect 440756 273846 440812 273902
rect 440564 273698 440620 273754
rect 440660 270459 440716 270498
rect 440660 270442 440662 270459
rect 440662 270442 440714 270459
rect 440714 270442 440716 270459
rect 449204 270738 449260 270794
rect 449204 269850 449260 269906
rect 457940 273846 457996 273902
rect 458036 273402 458092 273458
rect 460724 270459 460780 270498
rect 460724 270442 460726 270459
rect 460726 270442 460778 270459
rect 460778 270442 460780 270459
rect 469076 270311 469132 270350
rect 469076 270294 469078 270311
rect 469078 270294 469130 270311
rect 469130 270294 469132 270311
rect 469172 269998 469228 270054
rect 469364 270163 469420 270202
rect 469364 270146 469366 270163
rect 469366 270146 469418 270163
rect 469418 270146 469420 270163
rect 469556 270311 469612 270350
rect 469556 270294 469558 270311
rect 469558 270294 469610 270311
rect 469610 270294 469612 270311
rect 469556 270163 469612 270202
rect 469556 270146 469558 270163
rect 469558 270146 469610 270163
rect 469610 270146 469612 270163
rect 469652 269998 469708 270054
rect 469268 269850 469324 269906
rect 484436 273994 484492 274050
rect 488948 277842 489004 277898
rect 491636 274142 491692 274198
rect 489620 273698 489676 273754
rect 489620 273402 489676 273458
rect 488084 268074 488140 268130
rect 488276 268074 488332 268130
rect 496148 277694 496204 277750
rect 498836 274290 498892 274346
rect 499508 270294 499564 270350
rect 499412 268409 499414 268426
rect 499414 268409 499466 268426
rect 499466 268409 499468 268426
rect 499412 268370 499468 268409
rect 499700 270146 499756 270202
rect 499604 269998 499660 270054
rect 499604 268666 499660 268722
rect 499796 269998 499852 270054
rect 499700 268370 499756 268426
rect 499316 268074 499372 268130
rect 499508 268074 499564 268130
rect 507092 277546 507148 277602
rect 505940 274438 505996 274494
rect 504020 273846 504076 273902
rect 503924 273698 503980 273754
rect 509492 270294 509548 270350
rect 513044 269110 513100 269166
rect 517748 277398 517804 277454
rect 520148 274734 520204 274790
rect 516596 274586 516652 274642
rect 519476 270294 519532 270350
rect 519668 270294 519724 270350
rect 519476 269110 519532 269166
rect 519860 270146 519916 270202
rect 519764 269998 519820 270054
rect 519764 268666 519820 268722
rect 519860 268370 519916 268426
rect 519668 268074 519724 268130
rect 413300 264818 413356 264874
rect 412340 246762 412396 246818
rect 443540 243671 443596 243710
rect 443540 243654 443542 243671
rect 443542 243654 443594 243671
rect 443594 243654 443596 243671
rect 463604 243671 463660 243710
rect 463604 243654 463606 243671
rect 463606 243654 463658 243671
rect 463658 243654 463660 243671
rect 483860 243671 483916 243710
rect 483860 243654 483862 243671
rect 483862 243654 483914 243671
rect 483914 243654 483916 243671
rect 503924 243671 503980 243710
rect 503924 243654 503926 243671
rect 503926 243654 503978 243671
rect 503978 243654 503980 243671
rect 443540 242509 443542 242526
rect 443542 242509 443594 242526
rect 443594 242509 443596 242526
rect 443540 242470 443596 242509
rect 463604 242509 463606 242526
rect 463606 242509 463658 242526
rect 463658 242509 463660 242526
rect 463604 242470 463660 242509
rect 483860 242509 483862 242526
rect 483862 242509 483914 242526
rect 483914 242509 483916 242526
rect 483860 242470 483916 242509
rect 503924 242509 503926 242526
rect 503926 242509 503978 242526
rect 503978 242509 503980 242526
rect 503924 242470 503980 242509
rect 412052 238770 412108 238826
rect 411956 237586 412012 237642
rect 511124 242470 511180 242526
rect 528500 277250 528556 277306
rect 529844 273698 529900 273754
rect 529844 273402 529900 273458
rect 529844 269850 529900 269906
rect 529844 269110 529900 269166
rect 527348 265262 527404 265318
rect 530900 265114 530956 265170
rect 539252 277102 539308 277158
rect 544436 270481 544438 270498
rect 544438 270481 544490 270498
rect 544490 270481 544492 270498
rect 544436 270442 544492 270481
rect 548756 273698 548812 273754
rect 538004 264966 538060 265022
rect 563060 273254 563116 273310
rect 566516 271330 566572 271386
rect 564404 270481 564406 270498
rect 564406 270481 564458 270498
rect 564458 270481 564460 270498
rect 564404 270442 564460 270481
rect 582068 270294 582124 270350
rect 592724 276214 592780 276270
rect 589172 270146 589228 270202
rect 577268 269702 577324 269758
rect 574868 268814 574924 268870
rect 567764 268518 567820 268574
rect 560660 267926 560716 267982
rect 555860 264818 555916 264874
rect 524180 243671 524236 243710
rect 524180 243654 524182 243671
rect 524182 243654 524234 243671
rect 524234 243654 524236 243671
rect 544244 243671 544300 243710
rect 544244 243654 544246 243671
rect 544246 243654 544298 243671
rect 544298 243654 544300 243671
rect 564500 243671 564556 243710
rect 564500 243654 564502 243671
rect 564502 243654 564554 243671
rect 564554 243654 564556 243671
rect 584564 243671 584620 243710
rect 584564 243654 584566 243671
rect 584566 243654 584618 243671
rect 584618 243654 584620 243671
rect 521588 241878 521644 241934
rect 596372 269998 596428 270054
rect 599828 275918 599884 275974
rect 602228 275474 602284 275530
rect 603380 269850 603436 269906
rect 607028 276066 607084 276122
rect 605780 269554 605836 269610
rect 610580 275770 610636 275826
rect 614228 267778 614284 267834
rect 609428 265854 609484 265910
rect 617684 276806 617740 276862
rect 616532 275326 616588 275382
rect 620084 269406 620140 269462
rect 624884 275622 624940 275678
rect 623636 275178 623692 275234
rect 623060 270442 623116 270498
rect 627284 275030 627340 275086
rect 626036 268222 626092 268278
rect 630836 269258 630892 269314
rect 628436 265558 628492 265614
rect 632084 265410 632140 265466
rect 635540 276658 635596 276714
rect 637940 276362 637996 276418
rect 634292 270590 634348 270646
rect 642740 276510 642796 276566
rect 645140 274882 645196 274938
rect 640340 268962 640396 269018
rect 639092 267630 639148 267686
rect 604820 243693 604822 243710
rect 604822 243693 604874 243710
rect 604874 243693 604876 243710
rect 604820 243654 604876 243693
rect 624884 243693 624886 243710
rect 624886 243693 624938 243710
rect 624938 243693 624940 243710
rect 624884 243654 624940 243693
rect 596180 238918 596236 238974
rect 511124 237734 511180 237790
rect 420500 236715 420556 236754
rect 420500 236698 420502 236715
rect 420502 236698 420554 236715
rect 420554 236698 420556 236715
rect 505844 237586 505900 237642
rect 440564 236715 440620 236754
rect 440564 236698 440566 236715
rect 440566 236698 440618 236715
rect 440618 236698 440620 236715
rect 460820 236715 460876 236754
rect 460820 236698 460822 236715
rect 460822 236698 460874 236715
rect 460874 236698 460876 236715
rect 480884 236715 480940 236754
rect 480884 236698 480886 236715
rect 480886 236698 480938 236715
rect 480938 236698 480940 236715
rect 497492 236698 497548 236754
rect 420596 236402 420652 236458
rect 547124 234626 547180 234682
rect 637172 233590 637228 233646
rect 638420 236254 638476 236310
rect 645140 243671 645196 243710
rect 645140 243654 645142 243671
rect 645142 243654 645194 243671
rect 645194 243654 645196 243671
rect 638036 234034 638092 234090
rect 637940 233886 637996 233942
rect 638228 233442 638284 233498
rect 638804 233738 638860 233794
rect 638900 233590 638956 233646
rect 639284 236254 639340 236310
rect 649748 754402 649804 754458
rect 210260 86922 210316 86978
rect 210164 77746 210220 77802
rect 210164 55990 210220 56046
rect 210260 54954 210316 55010
rect 210836 54214 210892 54270
rect 214772 54214 214828 54270
rect 210740 54066 210796 54122
rect 216980 54066 217036 54122
rect 187604 41782 187660 41838
rect 194324 41782 194380 41838
rect 211988 51846 212044 51902
rect 212084 45186 212140 45242
rect 211700 45038 211756 45094
rect 212660 51994 212716 52050
rect 213044 53474 213100 53530
rect 215972 53474 216028 53530
rect 216692 53326 216748 53382
rect 221396 53918 221452 53974
rect 217844 53178 217900 53234
rect 221108 53474 221164 53530
rect 221876 52290 221932 52346
rect 222644 51698 222700 51754
rect 223316 52142 223372 52198
rect 229652 50366 229708 50422
rect 237620 51402 237676 51458
rect 237524 51254 237580 51310
rect 242420 48738 242476 48794
rect 242036 48590 242092 48646
rect 243380 51550 243436 51606
rect 242996 48442 243052 48498
rect 273620 53269 273676 53271
rect 273620 53217 273622 53269
rect 273622 53217 273674 53269
rect 273674 53217 273676 53269
rect 273620 53215 273676 53217
rect 293684 53178 293740 53234
rect 243764 48294 243820 48350
rect 241940 48146 241996 48202
rect 215444 44890 215500 44946
rect 302516 43262 302572 43318
rect 302420 42078 302476 42134
rect 306740 42078 306796 42134
rect 374420 51589 374422 51606
rect 374422 51589 374474 51606
rect 374474 51589 374476 51606
rect 374420 51550 374476 51589
rect 394292 51550 394348 51606
rect 440660 53195 440716 53234
rect 440660 53178 440662 53195
rect 440662 53178 440714 53195
rect 440714 53178 440716 53195
rect 443732 53217 443734 53234
rect 443734 53217 443786 53234
rect 443786 53217 443788 53234
rect 443732 53178 443788 53217
rect 457940 51589 457942 51606
rect 457942 51589 457994 51606
rect 457994 51589 457996 51606
rect 457940 51550 457996 51589
rect 478004 51550 478060 51606
rect 498260 51589 498262 51606
rect 498262 51589 498314 51606
rect 498314 51589 498316 51606
rect 498260 51550 498316 51589
rect 518324 51550 518380 51606
rect 512276 49034 512332 49090
rect 460820 46074 460876 46130
rect 465812 46074 465868 46130
rect 364916 43262 364972 43318
rect 411572 42078 411628 42134
rect 416276 42078 416332 42134
rect 211028 40746 211084 40802
rect 136532 40154 136588 40210
rect 520436 42078 520492 42134
rect 649844 707486 649900 707542
rect 650228 994014 650284 994070
rect 655124 976698 655180 976754
rect 653780 941474 653836 941530
rect 655220 965006 655276 965062
rect 655316 953314 655372 953370
rect 674516 966486 674572 966542
rect 675284 966486 675340 966542
rect 675764 965746 675820 965802
rect 675380 965006 675436 965062
rect 675764 963378 675820 963434
rect 675668 962490 675724 962546
rect 675380 962194 675436 962250
rect 675764 961454 675820 961510
rect 674132 959234 674188 959290
rect 654452 929782 654508 929838
rect 653972 918090 654028 918146
rect 654452 906398 654508 906454
rect 653780 894558 653836 894614
rect 653972 882866 654028 882922
rect 654452 871174 654508 871230
rect 654164 859482 654220 859538
rect 650132 848234 650188 848290
rect 653972 835950 654028 836006
rect 653972 824258 654028 824314
rect 654452 812566 654508 812622
rect 650036 801318 650092 801374
rect 654068 789034 654124 789090
rect 654068 777342 654124 777398
rect 653972 765502 654028 765558
rect 653972 742118 654028 742174
rect 655220 730426 655276 730482
rect 654260 718586 654316 718642
rect 654452 695202 654508 695258
rect 655124 683510 655180 683566
rect 654452 671670 654508 671726
rect 649940 660570 649996 660626
rect 645140 231518 645196 231574
rect 538580 51589 538582 51606
rect 538582 51589 538634 51606
rect 538634 51589 538636 51606
rect 538580 51550 538636 51589
rect 541460 51589 541462 51606
rect 541462 51589 541514 51606
rect 541514 51589 541516 51606
rect 541460 51550 541516 51589
rect 584660 51589 584662 51606
rect 584662 51589 584714 51606
rect 584714 51589 584716 51606
rect 584660 51550 584716 51589
rect 604724 51550 604780 51606
rect 529268 43262 529324 43318
rect 509684 41782 509740 41838
rect 518516 41782 518572 41838
rect 645236 231074 645292 231130
rect 654260 648286 654316 648342
rect 654356 624754 654412 624810
rect 654356 613062 654412 613118
rect 654452 601370 654508 601426
rect 654452 589530 654508 589586
rect 654452 577838 654508 577894
rect 654452 566146 654508 566202
rect 654452 554454 654508 554510
rect 654452 542614 654508 542670
rect 655316 636594 655372 636650
rect 654068 530922 654124 530978
rect 654452 519269 654454 519286
rect 654454 519269 654506 519286
rect 654506 519269 654508 519286
rect 654452 519230 654508 519269
rect 654452 507390 654508 507446
rect 654356 495698 654412 495754
rect 654260 484006 654316 484062
rect 654452 472205 654454 472222
rect 654454 472205 654506 472222
rect 654506 472205 654508 472222
rect 654452 472166 654508 472205
rect 654452 460474 654508 460530
rect 654356 448782 654412 448838
rect 654452 436942 654508 436998
rect 654452 425398 654508 425454
rect 653876 413558 653932 413614
rect 654452 401718 654508 401774
rect 654452 390026 654508 390082
rect 654452 378482 654508 378538
rect 654452 366494 654508 366550
rect 655220 354802 655276 354858
rect 654452 343110 654508 343166
rect 654452 331566 654508 331622
rect 655124 319726 655180 319782
rect 654548 296194 654604 296250
rect 654068 284650 654124 284706
rect 646292 232554 646348 232610
rect 650036 232554 650092 232610
rect 645524 231962 645580 232018
rect 645332 230630 645388 230686
rect 645428 121149 645430 121166
rect 645430 121149 645482 121166
rect 645482 121149 645484 121166
rect 645428 121110 645484 121149
rect 645428 104238 645484 104294
rect 645428 87662 645484 87718
rect 645428 86626 645484 86682
rect 646100 221750 646156 221806
rect 646292 221750 646348 221806
rect 645620 210354 645676 210410
rect 645908 198662 645964 198718
rect 646100 198662 646156 198718
rect 647060 166250 647116 166306
rect 647924 166990 647980 167046
rect 647828 165954 647884 166010
rect 645716 161257 645718 161274
rect 645718 161257 645770 161274
rect 645770 161257 645772 161274
rect 645716 161218 645772 161257
rect 645908 161257 645910 161274
rect 645910 161257 645962 161274
rect 645962 161257 645964 161274
rect 645908 161218 645964 161257
rect 655316 307886 655372 307942
rect 673844 939106 673900 939162
rect 673364 753070 673420 753126
rect 673268 752478 673324 752534
rect 673172 752034 673228 752090
rect 673076 707486 673132 707542
rect 672020 579762 672076 579818
rect 675476 960714 675532 960770
rect 675092 959234 675148 959290
rect 675476 959086 675532 959142
rect 675764 958346 675820 958402
rect 675380 957606 675436 957662
rect 674900 953462 674956 953518
rect 675476 955978 675532 956034
rect 675188 953314 675244 953370
rect 676820 940882 676876 940938
rect 674516 939846 674572 939902
rect 674420 939567 674476 939606
rect 674420 939550 674422 939567
rect 674422 939550 674474 939567
rect 674474 939550 674476 939567
rect 676916 940438 676972 940494
rect 676820 938218 676876 938274
rect 674420 937961 674422 937978
rect 674422 937961 674474 937978
rect 674474 937961 674476 937978
rect 674420 937922 674476 937961
rect 676916 937182 676972 937238
rect 674036 934666 674092 934722
rect 677012 929486 677068 929542
rect 676820 928894 676876 928950
rect 676820 928450 676876 928506
rect 677012 928450 677068 928506
rect 675380 876946 675436 877002
rect 675764 876502 675820 876558
rect 675092 875762 675148 875818
rect 675476 875762 675532 875818
rect 674516 775566 674572 775622
rect 674324 772902 674380 772958
rect 675188 875614 675244 875670
rect 675476 873986 675532 874042
rect 675380 873542 675436 873598
rect 675380 869842 675436 869898
rect 675476 864662 675532 864718
rect 675380 787998 675436 788054
rect 675476 787110 675532 787166
rect 675764 786666 675820 786722
rect 675764 784890 675820 784946
rect 675668 784150 675724 784206
rect 675764 780598 675820 780654
rect 675380 775418 675436 775474
rect 674708 774974 674764 775030
rect 675764 773642 675820 773698
rect 676628 773050 676684 773106
rect 674612 772606 674668 772662
rect 674420 762877 674422 762894
rect 674422 762877 674474 762894
rect 674474 762877 674476 762894
rect 674420 762838 674476 762877
rect 674420 762285 674422 762302
rect 674422 762285 674474 762302
rect 674474 762285 674476 762302
rect 674420 762246 674476 762285
rect 674612 761989 674614 762006
rect 674614 761989 674666 762006
rect 674666 761989 674668 762006
rect 674612 761950 674668 761989
rect 673844 761210 673900 761266
rect 673844 760618 673900 760674
rect 677780 764614 677836 764670
rect 676628 758250 676684 758306
rect 677780 754402 677836 754458
rect 677012 751146 677068 751202
rect 676820 750554 676876 750610
rect 677012 750554 677068 750610
rect 676820 750110 676876 750166
rect 675380 743154 675436 743210
rect 675476 742118 675532 742174
rect 675764 741674 675820 741730
rect 675380 740046 675436 740102
rect 675476 739158 675532 739214
rect 675380 738566 675436 738622
rect 673844 716218 673900 716274
rect 673844 715626 673900 715682
rect 673460 708078 673516 708134
rect 673844 671078 673900 671134
rect 673844 663382 673900 663438
rect 673364 662790 673420 662846
rect 673268 662346 673324 662402
rect 673844 661754 673900 661810
rect 673172 616762 673228 616818
rect 673076 527074 673132 527130
rect 673268 574286 673324 574342
rect 673172 526630 673228 526686
rect 674612 718033 674614 718050
rect 674614 718033 674666 718050
rect 674666 718033 674668 718050
rect 674612 717994 674668 718033
rect 674612 717589 674614 717606
rect 674614 717589 674666 717606
rect 674666 717589 674668 717606
rect 674612 717550 674668 717589
rect 674612 716997 674614 717014
rect 674614 716997 674666 717014
rect 674666 716997 674668 717014
rect 674612 716958 674668 716997
rect 677108 714738 677164 714794
rect 674612 709893 674614 709910
rect 674614 709893 674666 709910
rect 674666 709893 674668 709910
rect 674612 709854 674668 709893
rect 674420 709153 674422 709170
rect 674422 709153 674474 709170
rect 674474 709153 674476 709170
rect 674420 709114 674476 709153
rect 674420 708635 674422 708652
rect 674422 708635 674474 708652
rect 674474 708635 674476 708652
rect 674420 708596 674476 708635
rect 674420 707007 674422 707024
rect 674422 707007 674474 707024
rect 674474 707007 674476 707024
rect 674420 706968 674476 707007
rect 677012 706154 677068 706210
rect 677108 705710 677164 705766
rect 676820 705562 676876 705618
rect 677012 705562 677068 705618
rect 676820 705118 676876 705174
rect 675380 697866 675436 697922
rect 675764 697274 675820 697330
rect 675380 696830 675436 696886
rect 675764 694758 675820 694814
rect 675476 694314 675532 694370
rect 675764 693426 675820 693482
rect 675764 691946 675820 692002
rect 674420 666638 674476 666694
rect 674228 666120 674284 666176
rect 673940 642218 673996 642274
rect 674132 642255 674188 642311
rect 674420 627679 674422 627696
rect 674422 627679 674474 627696
rect 674474 627679 674476 627696
rect 674420 627640 674476 627679
rect 674420 626569 674422 626586
rect 674422 626569 674474 626586
rect 674474 626569 674476 626586
rect 674420 626530 674476 626569
rect 674420 625511 674476 625550
rect 674420 625494 674422 625511
rect 674422 625494 674474 625511
rect 674474 625494 674476 625511
rect 673940 623274 673996 623330
rect 674516 621942 674572 621998
rect 674708 672893 674710 672910
rect 674710 672893 674762 672910
rect 674762 672893 674764 672910
rect 674708 672854 674764 672893
rect 674708 672301 674710 672318
rect 674710 672301 674762 672318
rect 674762 672301 674764 672318
rect 674708 672262 674764 672301
rect 674708 671857 674710 671874
rect 674710 671857 674762 671874
rect 674762 671857 674764 671874
rect 674708 671818 674764 671857
rect 674708 668562 674764 668618
rect 674708 664161 674710 664178
rect 674710 664161 674762 664178
rect 674762 664161 674764 664178
rect 674708 664122 674764 664161
rect 674708 660866 674764 660922
rect 674708 660422 674764 660478
rect 674708 653614 674764 653670
rect 675092 660422 675148 660478
rect 675092 659830 675148 659886
rect 675380 652578 675436 652634
rect 675476 652134 675532 652190
rect 675476 651394 675532 651450
rect 675668 649766 675724 649822
rect 675476 648878 675532 648934
rect 675476 645326 675532 645382
rect 675764 640294 675820 640350
rect 675764 638518 675820 638574
rect 674900 627309 674902 627326
rect 674902 627309 674954 627326
rect 674954 627309 674956 627326
rect 674900 627270 674956 627309
rect 675092 621350 675148 621406
rect 674612 619130 674668 619186
rect 674420 618429 674422 618446
rect 674422 618429 674474 618446
rect 674474 618429 674476 618446
rect 674420 618390 674476 618429
rect 674420 617837 674422 617854
rect 674422 617837 674474 617854
rect 674474 617837 674476 617854
rect 674420 617798 674476 617837
rect 674708 617541 674710 617558
rect 674710 617541 674762 617558
rect 674762 617541 674764 617558
rect 674708 617502 674764 617541
rect 676820 624754 676876 624810
rect 676916 624014 676972 624070
rect 677108 615874 677164 615930
rect 676916 615282 676972 615338
rect 677108 615282 677164 615338
rect 676916 614838 676972 614894
rect 675380 607734 675436 607790
rect 675476 607142 675532 607198
rect 675476 606402 675532 606458
rect 675380 604774 675436 604830
rect 675764 600186 675820 600242
rect 675764 595302 675820 595358
rect 675764 593378 675820 593434
rect 674612 582130 674668 582186
rect 674420 581908 674476 581964
rect 674612 581577 674614 581594
rect 674614 581577 674666 581594
rect 674666 581577 674668 581594
rect 674612 581538 674668 581577
rect 674420 580837 674422 580854
rect 674422 580837 674474 580854
rect 674474 580837 674476 580854
rect 674420 580798 674476 580837
rect 673844 580206 673900 580262
rect 676820 579466 676876 579522
rect 673844 573694 673900 573750
rect 673844 573250 673900 573306
rect 673748 572658 673804 572714
rect 673844 572066 673900 572122
rect 674420 571587 674422 571604
rect 674422 571587 674474 571604
rect 674474 571587 674476 571604
rect 674420 571548 674476 571587
rect 677012 570734 677068 570790
rect 676820 570142 676876 570198
rect 676820 569698 676876 569754
rect 677012 569550 677068 569606
rect 673652 529903 673708 529942
rect 673652 529886 673654 529903
rect 673654 529886 673706 529903
rect 673706 529886 673708 529903
rect 673556 529294 673612 529350
rect 673364 527666 673420 527722
rect 673268 484154 673324 484210
rect 673844 492294 673900 492350
rect 674228 488002 674284 488058
rect 674516 489334 674572 489390
rect 674420 487410 674476 487466
rect 675476 562594 675532 562650
rect 675476 561706 675532 561762
rect 675380 561410 675436 561466
rect 675476 558894 675532 558950
rect 675764 554454 675820 554510
rect 674804 537177 674806 537194
rect 674806 537177 674858 537194
rect 674858 537177 674860 537194
rect 674804 537138 674860 537177
rect 676820 537138 676876 537194
rect 674804 536585 674806 536602
rect 674806 536585 674858 536602
rect 674858 536585 674860 536602
rect 674804 536546 674860 536585
rect 674804 536141 674806 536158
rect 674806 536141 674858 536158
rect 674858 536141 674860 536158
rect 674804 536102 674860 536141
rect 677300 535066 677356 535122
rect 676916 533882 676972 533938
rect 674804 529037 674806 529054
rect 674806 529037 674858 529054
rect 674858 529037 674860 529054
rect 674804 528998 674860 529037
rect 674804 528445 674806 528462
rect 674806 528445 674858 528462
rect 674858 528445 674860 528462
rect 674804 528406 674860 528445
rect 676820 525150 676876 525206
rect 676820 524706 676876 524762
rect 674612 487114 674668 487170
rect 674900 493182 674956 493238
rect 675092 493221 675094 493238
rect 675094 493221 675146 493238
rect 675146 493221 675148 493238
rect 675092 493182 675148 493221
rect 677012 525742 677068 525798
rect 677012 525150 677068 525206
rect 677396 534474 677452 534530
rect 677300 492146 677356 492202
rect 677396 490962 677452 491018
rect 677204 490518 677260 490574
rect 676916 489926 676972 489982
rect 674804 485486 674860 485542
rect 674324 484746 674380 484802
rect 673748 483710 673804 483766
rect 673844 482526 673900 482582
rect 676820 481194 676876 481250
rect 676820 480750 676876 480806
rect 674708 405457 674710 405474
rect 674710 405457 674762 405474
rect 674762 405457 674764 405474
rect 674708 405418 674764 405457
rect 673844 404678 673900 404734
rect 674708 404421 674710 404438
rect 674710 404421 674762 404438
rect 674762 404421 674764 404438
rect 674708 404382 674764 404421
rect 673844 403050 673900 403106
rect 673748 374338 673804 374394
rect 673364 373302 673420 373358
rect 677012 481638 677068 481694
rect 677012 480750 677068 480806
rect 677396 403938 677452 403994
rect 677204 402754 677260 402810
rect 676916 402162 676972 402218
rect 675092 401274 675148 401330
rect 674132 399794 674188 399850
rect 673940 396538 673996 396594
rect 674228 397574 674284 397630
rect 674900 396834 674956 396890
rect 674516 395798 674572 395854
rect 674804 394614 674860 394670
rect 674612 394170 674668 394226
rect 674996 395206 675052 395262
rect 675380 400090 675436 400146
rect 675188 397870 675244 397926
rect 677108 393430 677164 393486
rect 676916 392986 676972 393042
rect 677108 392986 677164 393042
rect 676916 392542 676972 392598
rect 675092 374486 675148 374542
rect 675476 378778 675532 378834
rect 675188 374042 675244 374098
rect 675476 373894 675532 373950
rect 675380 371970 675436 372026
rect 674420 360021 674422 360038
rect 674422 360021 674474 360038
rect 674474 360021 674476 360038
rect 674420 359982 674476 360021
rect 674708 359725 674710 359742
rect 674710 359725 674762 359742
rect 674762 359725 674764 359742
rect 674708 359686 674764 359725
rect 674420 358985 674422 359002
rect 674422 358985 674474 359002
rect 674474 358985 674476 359002
rect 674420 358946 674476 358985
rect 673844 358354 673900 358410
rect 674900 355986 674956 356042
rect 673940 354062 673996 354118
rect 674324 351842 674380 351898
rect 674132 350806 674188 350862
rect 674036 349622 674092 349678
rect 674708 350066 674764 350122
rect 674516 348882 674572 348938
rect 675188 354950 675244 355006
rect 674996 354358 675052 354414
rect 675092 352138 675148 352194
rect 677108 353174 677164 353230
rect 675284 352730 675340 352786
rect 676916 351102 676972 351158
rect 676820 347698 676876 347754
rect 676820 347254 676876 347310
rect 677012 348290 677068 348346
rect 677012 347254 677068 347310
rect 677108 345182 677164 345238
rect 676916 344146 676972 344202
rect 675284 334970 675340 335026
rect 675476 334526 675532 334582
rect 675092 331122 675148 331178
rect 675764 330530 675820 330586
rect 674996 329494 675052 329550
rect 675380 328310 675436 328366
rect 675764 326830 675820 326886
rect 674420 315029 674422 315046
rect 674422 315029 674474 315046
rect 674474 315029 674476 315046
rect 674420 314990 674476 315029
rect 674708 314733 674710 314750
rect 674710 314733 674762 314750
rect 674762 314733 674764 314750
rect 674708 314694 674764 314733
rect 674420 313993 674422 314010
rect 674422 313993 674474 314010
rect 674474 313993 674476 314010
rect 674420 313954 674476 313993
rect 674036 311290 674092 311346
rect 675092 309958 675148 310014
rect 674324 309588 674380 309644
rect 674132 305814 674188 305870
rect 673940 289534 673996 289590
rect 674228 304186 674284 304242
rect 674996 308774 675052 308830
rect 674900 307738 674956 307794
rect 674804 307146 674860 307202
rect 674612 306702 674668 306758
rect 674516 304482 674572 304538
rect 674420 303594 674476 303650
rect 674420 302597 674422 302614
rect 674422 302597 674474 302614
rect 674474 302597 674476 302614
rect 674420 302558 674476 302597
rect 674708 305074 674764 305130
rect 677012 308182 677068 308238
rect 676916 305962 676972 306018
rect 676820 302706 676876 302762
rect 676820 302262 676876 302318
rect 676916 299450 676972 299506
rect 677012 299302 677068 299358
rect 675284 289978 675340 290034
rect 675092 284946 675148 285002
rect 675764 284798 675820 284854
rect 673940 284650 673996 284706
rect 675380 283614 675436 283670
rect 675764 281838 675820 281894
rect 674420 270037 674422 270054
rect 674422 270037 674474 270054
rect 674474 270037 674476 270054
rect 674420 269998 674476 270037
rect 674708 269741 674710 269758
rect 674710 269741 674762 269758
rect 674762 269741 674764 269758
rect 674708 269702 674764 269741
rect 674708 269149 674710 269166
rect 674710 269149 674762 269166
rect 674762 269149 674764 269166
rect 674708 269110 674764 269149
rect 674516 266002 674572 266058
rect 674324 262450 674380 262506
rect 674132 260822 674188 260878
rect 677108 265410 677164 265466
rect 675188 264966 675244 265022
rect 675092 264374 675148 264430
rect 674804 261710 674860 261766
rect 674708 261118 674764 261174
rect 674612 259490 674668 259546
rect 674900 260082 674956 260138
rect 674996 258898 675052 258954
rect 676916 263190 676972 263246
rect 675284 262746 675340 262802
rect 676820 257714 676876 257770
rect 676820 257270 676876 257326
rect 677012 258306 677068 258362
rect 677012 257714 677068 257770
rect 676916 253274 676972 253330
rect 677108 253126 677164 253182
rect 675188 245282 675244 245338
rect 675380 244690 675436 244746
rect 675476 243506 675532 243562
rect 675188 238918 675244 238974
rect 675764 238622 675820 238678
rect 675764 236846 675820 236902
rect 674708 225045 674710 225062
rect 674710 225045 674762 225062
rect 674762 225045 674764 225062
rect 674708 225006 674764 225045
rect 674420 224305 674422 224322
rect 674422 224305 674474 224322
rect 674474 224305 674476 224322
rect 674420 224266 674476 224305
rect 674708 224009 674710 224026
rect 674710 224009 674762 224026
rect 674762 224009 674764 224026
rect 674708 223970 674764 224009
rect 674900 220862 674956 220918
rect 674228 216718 674284 216774
rect 674516 215386 674572 215442
rect 674804 214794 674860 214850
rect 674708 214350 674764 214406
rect 674612 213758 674668 213814
rect 675476 219678 675532 219734
rect 674996 219234 675052 219290
rect 675188 217606 675244 217662
rect 675092 216866 675148 216922
rect 677108 218050 677164 218106
rect 676916 215978 676972 216034
rect 676820 212574 676876 212630
rect 676820 212130 676876 212186
rect 677012 213166 677068 213222
rect 677012 212574 677068 212630
rect 676916 210206 676972 210262
rect 677108 210058 677164 210114
rect 675380 199254 675436 199310
rect 675476 198662 675532 198718
rect 675476 198366 675532 198422
rect 675764 195258 675820 195314
rect 675380 193482 675436 193538
rect 675764 191558 675820 191614
rect 674708 179570 674764 179626
rect 674420 179313 674422 179330
rect 674422 179313 674474 179330
rect 674474 179313 674476 179330
rect 674420 179274 674476 179313
rect 674420 178795 674422 178812
rect 674422 178795 674474 178812
rect 674474 178795 674476 178812
rect 674420 178756 674476 178795
rect 674036 176018 674092 176074
rect 676916 175130 676972 175186
rect 675572 174686 675628 174742
rect 674804 174242 674860 174298
rect 674324 169506 674380 169562
rect 674516 168766 674572 168822
rect 674420 167303 674476 167342
rect 674420 167286 674422 167303
rect 674422 167286 674474 167303
rect 674474 167286 674476 167303
rect 674612 168174 674668 168230
rect 674708 167582 674764 167638
rect 675092 172022 675148 172078
rect 674996 171430 675052 171486
rect 674900 169802 674956 169858
rect 676820 173058 676876 173114
rect 675764 172614 675820 172670
rect 676916 161514 676972 161570
rect 676820 161366 676876 161422
rect 675284 155150 675340 155206
rect 675476 154410 675532 154466
rect 675476 153374 675532 153430
rect 675476 151894 675532 151950
rect 675476 150266 675532 150322
rect 675764 148490 675820 148546
rect 675764 146566 675820 146622
rect 676916 134282 676972 134338
rect 676820 133838 676876 133894
rect 674420 133581 674422 133598
rect 674422 133581 674474 133598
rect 674474 133581 674476 133598
rect 674420 133542 674476 133581
rect 674420 132523 674476 132562
rect 674420 132506 674422 132523
rect 674422 132506 674474 132523
rect 674474 132506 674476 132523
rect 645716 121406 645772 121462
rect 645716 120814 645772 120870
rect 674516 130582 674572 130638
rect 674324 127030 674380 127086
rect 673940 125402 673996 125458
rect 647732 120370 647788 120426
rect 674228 123774 674284 123830
rect 668180 106497 668182 106514
rect 668182 106497 668234 106514
rect 668234 106497 668236 106514
rect 668180 106458 668236 106497
rect 677108 129990 677164 130046
rect 675188 129546 675244 129602
rect 675092 128954 675148 129010
rect 674900 127326 674956 127382
rect 674804 126290 674860 126346
rect 674612 124662 674668 124718
rect 674708 121850 674764 121906
rect 674996 124070 675052 124126
rect 677012 127770 677068 127826
rect 676916 122886 676972 122942
rect 676820 122294 676876 122350
rect 677012 118002 677068 118058
rect 677108 117854 677164 117910
rect 675380 110010 675436 110066
rect 675476 109270 675532 109326
rect 675380 108086 675436 108142
rect 665204 105126 665260 105182
rect 675380 105126 675436 105182
rect 665204 104551 665260 104590
rect 665204 104534 665206 104551
rect 665206 104534 665258 104551
rect 665258 104534 665260 104551
rect 645716 88106 645772 88162
rect 646100 85738 646156 85794
rect 646292 84998 646348 85054
rect 645908 84110 645964 84166
rect 646100 78634 646156 78690
rect 646484 76897 646486 76914
rect 646486 76897 646538 76914
rect 646538 76897 646540 76914
rect 646484 76858 646540 76897
rect 646484 75970 646540 76026
rect 646484 72714 646540 72770
rect 647348 87366 647404 87422
rect 647156 80854 647212 80910
rect 646868 78486 646924 78542
rect 647636 88994 647692 89050
rect 647540 82186 647596 82242
rect 650900 86922 650956 86978
rect 647828 86182 647884 86238
rect 647732 85442 647788 85498
rect 650996 85294 651052 85350
rect 650996 84258 651052 84314
rect 647924 83409 647926 83426
rect 647926 83409 647978 83426
rect 647978 83409 647980 83426
rect 647924 83370 647980 83409
rect 650900 82630 650956 82686
rect 647924 82482 647980 82538
rect 647924 81315 647980 81354
rect 647924 81298 647926 81315
rect 647926 81298 647978 81315
rect 647978 81298 647980 81315
rect 647828 80410 647884 80466
rect 647924 80153 647926 80170
rect 647926 80153 647978 80170
rect 647978 80153 647980 80170
rect 647924 80114 647980 80153
rect 647924 79226 647980 79282
rect 647924 77637 647926 77654
rect 647926 77637 647978 77654
rect 647978 77637 647980 77654
rect 647924 77598 647980 77637
rect 647924 77006 647980 77062
rect 651188 86182 651244 86238
rect 651092 83370 651148 83426
rect 651380 83814 651436 83870
rect 662900 81150 662956 81206
rect 646868 75378 646924 75434
rect 647924 75082 647980 75138
rect 646964 74342 647020 74398
rect 647828 73750 647884 73806
rect 647924 73010 647980 73066
rect 675764 103202 675820 103258
rect 675764 101426 675820 101482
rect 663572 85590 663628 85646
rect 663284 85146 663340 85202
rect 663476 84702 663532 84758
rect 663380 82778 663436 82834
rect 663284 82038 663340 82094
rect 646676 72122 646732 72178
rect 640724 40598 640780 40654
<< metal3 >>
rect 148527 1015976 148593 1015979
rect 251343 1015976 251409 1015979
rect 353391 1015976 353457 1015979
rect 98562 1015916 99486 1015976
rect 98562 1015680 98622 1015916
rect 99426 1015798 99486 1015916
rect 148527 1015974 150846 1015976
rect 148527 1015918 148532 1015974
rect 148588 1015918 150846 1015974
rect 148527 1015916 150846 1015918
rect 148527 1015913 148593 1015916
rect 149730 1015798 149790 1015916
rect 150786 1015798 150846 1015916
rect 200610 1015916 201726 1015976
rect 200610 1015798 200670 1015916
rect 201666 1015798 201726 1015916
rect 251343 1015974 253662 1015976
rect 251343 1015918 251348 1015974
rect 251404 1015918 253662 1015974
rect 251343 1015916 253662 1015918
rect 251343 1015913 251409 1015916
rect 252546 1015798 252606 1015916
rect 253602 1015798 253662 1015916
rect 353391 1015974 355326 1015976
rect 353391 1015918 353396 1015974
rect 353452 1015918 355326 1015974
rect 353391 1015916 355326 1015918
rect 353391 1015913 353457 1015916
rect 354498 1015798 354558 1015916
rect 355266 1015828 355326 1015916
rect 422274 1015916 423102 1015976
rect 422274 1015828 422334 1015916
rect 355266 1015768 355680 1015828
rect 421920 1015798 422334 1015828
rect 423042 1015798 423102 1015916
rect 421890 1015768 422334 1015798
rect 98400 1015650 98622 1015680
rect 98370 1015620 98622 1015650
rect 81039 995848 81105 995851
rect 94959 995848 95025 995851
rect 81039 995846 95025 995848
rect 81039 995790 81044 995846
rect 81100 995790 94964 995846
rect 95020 995790 95025 995846
rect 98031 995848 98097 995851
rect 98370 995848 98430 1015620
rect 145359 1007984 145425 1007987
rect 148527 1007984 148593 1007987
rect 145359 1007982 148593 1007984
rect 145359 1007926 145364 1007982
rect 145420 1007926 148532 1007982
rect 148588 1007926 148593 1007982
rect 145359 1007924 148593 1007926
rect 145359 1007921 145425 1007924
rect 148527 1007921 148593 1007924
rect 348879 1007836 348945 1007839
rect 353295 1007836 353361 1007839
rect 348879 1007834 353361 1007836
rect 348879 1007778 348884 1007834
rect 348940 1007778 353300 1007834
rect 353356 1007778 353361 1007834
rect 348879 1007776 353361 1007778
rect 348879 1007773 348945 1007776
rect 353295 1007773 353361 1007776
rect 161184 1005408 161598 1005468
rect 160431 1003248 160497 1003251
rect 160032 1003246 160497 1003248
rect 160032 1003190 160436 1003246
rect 160492 1003190 160497 1003246
rect 161538 1003214 161598 1005408
rect 213807 1005172 213873 1005175
rect 218799 1005172 218865 1005175
rect 213807 1005170 218865 1005172
rect 213807 1005114 213812 1005170
rect 213868 1005114 218804 1005170
rect 218860 1005114 218865 1005170
rect 213807 1005112 218865 1005114
rect 213807 1005109 213873 1005112
rect 218799 1005109 218865 1005112
rect 160032 1003188 160497 1003190
rect 160431 1003185 160497 1003188
rect 161487 1003209 161598 1003214
rect 161487 1003153 161492 1003209
rect 161548 1003153 161598 1003209
rect 209103 1003248 209169 1003251
rect 211791 1003248 211857 1003251
rect 316431 1003248 316497 1003251
rect 357423 1003248 357489 1003251
rect 362511 1003248 362577 1003251
rect 209103 1003246 209376 1003248
rect 209103 1003190 209108 1003246
rect 209164 1003190 209376 1003246
rect 209103 1003188 209376 1003190
rect 211488 1003246 211857 1003248
rect 211488 1003190 211796 1003246
rect 211852 1003190 211857 1003246
rect 211488 1003188 211857 1003190
rect 316128 1003246 316497 1003248
rect 316128 1003190 316436 1003246
rect 316492 1003190 316497 1003246
rect 316128 1003188 316497 1003190
rect 357216 1003246 357489 1003248
rect 357216 1003190 357428 1003246
rect 357484 1003190 357489 1003246
rect 357216 1003188 357489 1003190
rect 362208 1003246 362577 1003248
rect 362208 1003190 362516 1003246
rect 362572 1003190 362577 1003246
rect 362208 1003188 362577 1003190
rect 209103 1003185 209169 1003188
rect 211791 1003185 211857 1003188
rect 316431 1003185 316497 1003188
rect 357423 1003185 357489 1003188
rect 362511 1003185 362577 1003188
rect 161487 1003151 161598 1003153
rect 161487 1003148 161553 1003151
rect 308847 1002952 308913 1002955
rect 312111 1002952 312177 1002955
rect 308847 1002950 309024 1002952
rect 308847 1002894 308852 1002950
rect 308908 1002894 309024 1002950
rect 308847 1002892 309024 1002894
rect 312111 1002950 312288 1002952
rect 312111 1002894 312116 1002950
rect 312172 1002894 312288 1002950
rect 312111 1002892 312288 1002894
rect 308847 1002889 308913 1002892
rect 312111 1002889 312177 1002892
rect 308271 1002804 308337 1002807
rect 309327 1002804 309393 1002807
rect 358575 1002804 358641 1002807
rect 308271 1002802 308448 1002804
rect 308271 1002746 308276 1002802
rect 308332 1002746 308448 1002802
rect 308271 1002744 308448 1002746
rect 309327 1002802 309600 1002804
rect 309327 1002746 309332 1002802
rect 309388 1002746 309600 1002802
rect 309327 1002744 309600 1002746
rect 358368 1002802 358641 1002804
rect 358368 1002746 358580 1002802
rect 358636 1002746 358641 1002802
rect 358368 1002744 358641 1002746
rect 308271 1002741 308337 1002744
rect 309327 1002741 309393 1002744
rect 358575 1002741 358641 1002744
rect 153327 1002656 153393 1002659
rect 357999 1002656 358065 1002659
rect 153327 1002654 153504 1002656
rect 153327 1002598 153332 1002654
rect 153388 1002598 153504 1002654
rect 153327 1002596 153504 1002598
rect 357792 1002654 358065 1002656
rect 357792 1002598 358004 1002654
rect 358060 1002598 358065 1002654
rect 357792 1002596 358065 1002598
rect 153327 1002593 153393 1002596
rect 357999 1002593 358065 1002596
rect 151599 1002508 151665 1002511
rect 152655 1002508 152721 1002511
rect 361839 1002508 361905 1002511
rect 151599 1002506 151968 1002508
rect 151599 1002450 151604 1002506
rect 151660 1002450 151968 1002506
rect 151599 1002448 151968 1002450
rect 152655 1002506 153024 1002508
rect 152655 1002450 152660 1002506
rect 152716 1002450 153024 1002506
rect 152655 1002448 153024 1002450
rect 361632 1002506 361905 1002508
rect 361632 1002450 361844 1002506
rect 361900 1002450 361905 1002506
rect 361632 1002448 361905 1002450
rect 151599 1002445 151665 1002448
rect 152655 1002445 152721 1002448
rect 361839 1002445 361905 1002448
rect 151023 1002360 151089 1002363
rect 359055 1002360 359121 1002363
rect 362895 1002360 362961 1002363
rect 151023 1002358 151392 1002360
rect 151023 1002302 151028 1002358
rect 151084 1002302 151392 1002358
rect 151023 1002300 151392 1002302
rect 358944 1002358 359121 1002360
rect 358944 1002302 359060 1002358
rect 359116 1002302 359121 1002358
rect 358944 1002300 359121 1002302
rect 362688 1002358 362961 1002360
rect 362688 1002302 362900 1002358
rect 362956 1002302 362961 1002358
rect 362688 1002300 362961 1002302
rect 151023 1002297 151089 1002300
rect 359055 1002297 359121 1002300
rect 362895 1002297 362961 1002300
rect 361359 1002212 361425 1002215
rect 361056 1002210 361425 1002212
rect 361056 1002154 361364 1002210
rect 361420 1002154 361425 1002210
rect 361056 1002152 361425 1002154
rect 361359 1002149 361425 1002152
rect 356367 1001324 356433 1001327
rect 356160 1001322 356433 1001324
rect 356160 1001266 356372 1001322
rect 356428 1001266 356433 1001322
rect 356160 1001264 356433 1001266
rect 356367 1001261 356433 1001264
rect 357039 1001176 357105 1001179
rect 356736 1001174 357105 1001176
rect 356736 1001118 357044 1001174
rect 357100 1001118 357105 1001174
rect 356736 1001116 357105 1001118
rect 357039 1001113 357105 1001116
rect 359631 1000880 359697 1000883
rect 360207 1000880 360273 1000883
rect 359424 1000878 359697 1000880
rect 359424 1000822 359636 1000878
rect 359692 1000822 359697 1000878
rect 359424 1000820 359697 1000822
rect 360000 1000878 360273 1000880
rect 360000 1000822 360212 1000878
rect 360268 1000822 360273 1000878
rect 360000 1000820 360273 1000822
rect 359631 1000817 359697 1000820
rect 360207 1000817 360273 1000820
rect 155535 999400 155601 999403
rect 206895 999400 206961 999403
rect 258351 999400 258417 999403
rect 309903 999400 309969 999403
rect 364527 999400 364593 999403
rect 155535 999398 155712 999400
rect 155535 999342 155540 999398
rect 155596 999342 155712 999398
rect 155535 999340 155712 999342
rect 206895 999398 207168 999400
rect 206895 999342 206900 999398
rect 206956 999342 207168 999398
rect 206895 999340 207168 999342
rect 258351 999398 258528 999400
rect 258351 999342 258356 999398
rect 258412 999342 258528 999398
rect 258351 999340 258528 999342
rect 309903 999398 310176 999400
rect 309903 999342 309908 999398
rect 309964 999342 310176 999398
rect 309903 999340 310176 999342
rect 364320 999398 364593 999400
rect 364320 999342 364532 999398
rect 364588 999342 364593 999398
rect 364320 999340 364593 999342
rect 155535 999337 155601 999340
rect 206895 999337 206961 999340
rect 258351 999337 258417 999340
rect 309903 999337 309969 999340
rect 364527 999337 364593 999340
rect 314799 997920 314865 997923
rect 314496 997918 314865 997920
rect 314496 997862 314804 997918
rect 314860 997862 314865 997918
rect 314496 997860 314865 997862
rect 314799 997857 314865 997860
rect 365199 997920 365265 997923
rect 365199 997918 365472 997920
rect 365199 997862 365204 997918
rect 365260 997862 365472 997918
rect 365199 997860 365472 997862
rect 365199 997857 365265 997860
rect 270639 997180 270705 997183
rect 298095 997180 298161 997183
rect 270639 997178 298161 997180
rect 270639 997122 270644 997178
rect 270700 997122 298100 997178
rect 298156 997122 298161 997178
rect 270639 997120 298161 997122
rect 270639 997117 270705 997120
rect 298095 997117 298161 997120
rect 313743 997180 313809 997183
rect 313743 997178 313920 997180
rect 313743 997122 313748 997178
rect 313804 997122 313920 997178
rect 313743 997120 313920 997122
rect 313743 997117 313809 997120
rect 104655 996588 104721 996591
rect 205167 996588 205233 996591
rect 207951 996588 208017 996591
rect 311535 996588 311601 996591
rect 104655 996586 104928 996588
rect 104655 996530 104660 996586
rect 104716 996530 104928 996586
rect 104655 996528 104928 996530
rect 205167 996586 205536 996588
rect 205167 996530 205172 996586
rect 205228 996530 205536 996586
rect 205167 996528 205536 996530
rect 207951 996586 208224 996588
rect 207951 996530 207956 996586
rect 208012 996530 208224 996586
rect 207951 996528 208224 996530
rect 311535 996586 311712 996588
rect 311535 996530 311540 996586
rect 311596 996530 311712 996586
rect 311535 996528 311712 996530
rect 104655 996525 104721 996528
rect 205167 996525 205233 996528
rect 207951 996525 208017 996528
rect 311535 996525 311601 996528
rect 262479 996440 262545 996443
rect 262368 996438 262545 996440
rect 262368 996382 262484 996438
rect 262540 996382 262545 996438
rect 262368 996380 262545 996382
rect 262479 996377 262545 996380
rect 159183 996292 159249 996295
rect 158976 996290 159249 996292
rect 158976 996234 159188 996290
rect 159244 996234 159249 996290
rect 158976 996232 159249 996234
rect 159183 996229 159249 996232
rect 159759 996144 159825 996147
rect 159552 996142 159825 996144
rect 159552 996086 159764 996142
rect 159820 996086 159825 996142
rect 159552 996084 159825 996086
rect 159759 996081 159825 996084
rect 210159 996144 210225 996147
rect 257775 996144 257841 996147
rect 261999 996144 262065 996147
rect 263055 996144 263121 996147
rect 299535 996144 299601 996147
rect 210159 996142 210432 996144
rect 210159 996086 210164 996142
rect 210220 996086 210432 996142
rect 210159 996084 210432 996086
rect 257775 996142 257952 996144
rect 257775 996086 257780 996142
rect 257836 996086 257952 996142
rect 257775 996084 257952 996086
rect 261792 996142 262065 996144
rect 261792 996086 262004 996142
rect 262060 996086 262065 996142
rect 261792 996084 262065 996086
rect 262944 996142 263121 996144
rect 262944 996086 263060 996142
rect 263116 996086 263121 996142
rect 262944 996084 263121 996086
rect 210159 996081 210225 996084
rect 257775 996081 257841 996084
rect 261999 996081 262065 996084
rect 263055 996081 263121 996084
rect 297474 996142 299601 996144
rect 297474 996086 299540 996142
rect 299596 996086 299601 996142
rect 297474 996084 299601 996086
rect 99759 995996 99825 995999
rect 102831 995996 102897 995999
rect 108975 995996 109041 995999
rect 99759 995994 99936 995996
rect 99759 995938 99764 995994
rect 99820 995938 99936 995994
rect 99759 995936 99936 995938
rect 102831 995994 103200 995996
rect 102831 995938 102836 995994
rect 102892 995938 103200 995994
rect 102831 995936 103200 995938
rect 108672 995994 109041 995996
rect 108672 995938 108980 995994
rect 109036 995938 109041 995994
rect 108672 995936 109041 995938
rect 99759 995933 99825 995936
rect 102831 995933 102897 995936
rect 108975 995933 109041 995936
rect 109551 995996 109617 995999
rect 156591 995996 156657 995999
rect 160431 995996 160497 995999
rect 204015 995996 204081 995999
rect 210639 995996 210705 995999
rect 211791 995996 211857 995999
rect 219087 995996 219153 995999
rect 109551 995994 109728 995996
rect 109551 995938 109556 995994
rect 109612 995938 109728 995994
rect 109551 995936 109728 995938
rect 150018 995936 150240 995996
rect 156591 995994 156768 995996
rect 156591 995938 156596 995994
rect 156652 995938 156768 995994
rect 156591 995936 156768 995938
rect 160431 995994 160608 995996
rect 160431 995938 160436 995994
rect 160492 995938 160608 995994
rect 160431 995936 160608 995938
rect 204015 995994 204384 995996
rect 204015 995938 204020 995994
rect 204076 995938 204384 995994
rect 204015 995936 204384 995938
rect 210639 995994 210912 995996
rect 210639 995938 210644 995994
rect 210700 995938 210912 995994
rect 210639 995936 210912 995938
rect 211791 995994 212064 995996
rect 211791 995938 211796 995994
rect 211852 995938 212064 995994
rect 211791 995936 212064 995938
rect 212640 995936 212862 995996
rect 213696 995994 219153 995996
rect 213696 995938 219092 995994
rect 219148 995938 219153 995994
rect 213696 995936 219153 995938
rect 109551 995933 109617 995936
rect 98031 995846 98430 995848
rect 81039 995788 95025 995790
rect 81039 995785 81105 995788
rect 94959 995785 95025 995788
rect 81615 995700 81681 995703
rect 94959 995700 95025 995703
rect 81615 995698 95025 995700
rect 81615 995642 81620 995698
rect 81676 995642 94964 995698
rect 95020 995642 95025 995698
rect 81615 995640 95025 995642
rect 97794 995700 97854 995818
rect 98031 995790 98036 995846
rect 98092 995818 98430 995846
rect 100719 995848 100785 995851
rect 101199 995848 101265 995851
rect 102447 995848 102513 995851
rect 103983 995848 104049 995851
rect 107919 995848 107985 995851
rect 100719 995846 101088 995848
rect 98092 995790 98400 995818
rect 98031 995788 98400 995790
rect 98031 995785 98097 995788
rect 98850 995700 98910 995818
rect 100482 995700 100542 995818
rect 100719 995790 100724 995846
rect 100780 995790 101088 995846
rect 100719 995788 101088 995790
rect 101199 995846 101664 995848
rect 101199 995790 101204 995846
rect 101260 995790 101664 995846
rect 102447 995846 102720 995848
rect 101199 995788 101664 995790
rect 100719 995785 100785 995788
rect 101199 995785 101265 995788
rect 97794 995640 98910 995700
rect 99138 995640 100542 995700
rect 81615 995637 81681 995640
rect 94959 995637 95025 995640
rect 85359 995552 85425 995555
rect 85359 995550 88062 995552
rect 85359 995494 85364 995550
rect 85420 995494 88062 995550
rect 85359 995492 88062 995494
rect 85359 995489 85425 995492
rect 84783 995404 84849 995407
rect 88002 995404 88062 995492
rect 99138 995404 99198 995640
rect 84783 995402 86718 995404
rect 84783 995346 84788 995402
rect 84844 995346 86718 995402
rect 84783 995344 86718 995346
rect 88002 995344 99198 995404
rect 84783 995341 84849 995344
rect 86658 995108 86718 995344
rect 87759 995256 87825 995259
rect 102114 995256 102174 995818
rect 102447 995790 102452 995846
rect 102508 995790 102720 995846
rect 103983 995846 104352 995848
rect 102447 995788 102720 995790
rect 102447 995785 102513 995788
rect 102351 995700 102417 995703
rect 103746 995700 103806 995818
rect 103983 995790 103988 995846
rect 104044 995790 104352 995846
rect 103983 995788 104352 995790
rect 103983 995785 104049 995788
rect 105378 995703 105438 995818
rect 105954 995703 106014 995818
rect 106464 995788 106686 995848
rect 107919 995846 108192 995848
rect 102351 995698 103806 995700
rect 102351 995642 102356 995698
rect 102412 995642 103806 995698
rect 102351 995640 103806 995642
rect 105327 995698 105438 995703
rect 105327 995642 105332 995698
rect 105388 995642 105438 995698
rect 105327 995640 105438 995642
rect 105903 995698 106014 995703
rect 106626 995700 106686 995788
rect 105903 995642 105908 995698
rect 105964 995642 106014 995698
rect 105903 995640 106014 995642
rect 106242 995640 106686 995700
rect 102351 995637 102417 995640
rect 105327 995637 105393 995640
rect 105903 995637 105969 995640
rect 87759 995254 102174 995256
rect 87759 995198 87764 995254
rect 87820 995198 102174 995254
rect 87759 995196 102174 995198
rect 87759 995193 87825 995196
rect 97935 995108 98001 995111
rect 86658 995106 98001 995108
rect 86658 995050 97940 995106
rect 97996 995050 98001 995106
rect 86658 995048 98001 995050
rect 97935 995045 98001 995048
rect 89391 994960 89457 994963
rect 106242 994960 106302 995640
rect 106767 995256 106833 995259
rect 107010 995256 107070 995818
rect 107586 995703 107646 995818
rect 107919 995790 107924 995846
rect 107980 995790 108192 995846
rect 107919 995788 108192 995790
rect 107919 995785 107985 995788
rect 109218 995703 109278 995818
rect 107535 995698 107646 995703
rect 107535 995642 107540 995698
rect 107596 995642 107646 995698
rect 107535 995640 107646 995642
rect 109167 995698 109278 995703
rect 109167 995642 109172 995698
rect 109228 995642 109278 995698
rect 109167 995640 109278 995642
rect 110127 995700 110193 995703
rect 110274 995700 110334 995818
rect 110127 995698 110334 995700
rect 110127 995642 110132 995698
rect 110188 995642 110334 995698
rect 110127 995640 110334 995642
rect 107535 995637 107601 995640
rect 109167 995637 109233 995640
rect 110127 995637 110193 995640
rect 109359 995552 109425 995555
rect 110850 995552 110910 995818
rect 149154 995700 149214 995818
rect 150018 995700 150078 995936
rect 156591 995933 156657 995936
rect 160431 995933 160497 995936
rect 204015 995933 204081 995936
rect 210639 995933 210705 995936
rect 211791 995933 211857 995936
rect 154863 995848 154929 995851
rect 161487 995848 161553 995851
rect 183759 995848 183825 995851
rect 192495 995848 192561 995851
rect 195279 995848 195345 995851
rect 203055 995848 203121 995851
rect 203631 995848 203697 995851
rect 204687 995848 204753 995851
rect 154863 995846 155232 995848
rect 149154 995640 150078 995700
rect 109359 995550 110910 995552
rect 109359 995494 109364 995550
rect 109420 995494 110910 995550
rect 109359 995492 110910 995494
rect 133647 995552 133713 995555
rect 152418 995552 152478 995818
rect 133647 995550 152478 995552
rect 133647 995494 133652 995550
rect 133708 995494 152478 995550
rect 133647 995492 152478 995494
rect 109359 995489 109425 995492
rect 133647 995489 133713 995492
rect 149679 995404 149745 995407
rect 154050 995404 154110 995818
rect 149679 995402 154110 995404
rect 149679 995346 149684 995402
rect 149740 995346 154110 995402
rect 149679 995344 154110 995346
rect 149679 995341 149745 995344
rect 106767 995254 107070 995256
rect 106767 995198 106772 995254
rect 106828 995198 107070 995254
rect 106767 995196 107070 995198
rect 146799 995256 146865 995259
rect 154626 995256 154686 995818
rect 154863 995790 154868 995846
rect 154924 995790 155232 995846
rect 154863 995788 155232 995790
rect 154863 995785 154929 995788
rect 146799 995254 154686 995256
rect 146799 995198 146804 995254
rect 146860 995198 154686 995254
rect 146799 995196 154686 995198
rect 106767 995193 106833 995196
rect 146799 995193 146865 995196
rect 89391 994958 106302 994960
rect 89391 994902 89396 994958
rect 89452 994902 106302 994958
rect 89391 994900 106302 994902
rect 89391 994897 89457 994900
rect 132783 994516 132849 994519
rect 149679 994516 149745 994519
rect 132783 994514 149745 994516
rect 132783 994458 132788 994514
rect 132844 994458 149684 994514
rect 149740 994458 149745 994514
rect 132783 994456 149745 994458
rect 132783 994453 132849 994456
rect 149679 994453 149745 994456
rect 140751 994368 140817 994371
rect 156111 994368 156177 994371
rect 140751 994366 156177 994368
rect 140751 994310 140756 994366
rect 140812 994310 156116 994366
rect 156172 994310 156177 994366
rect 140751 994308 156177 994310
rect 140751 994305 140817 994308
rect 156111 994305 156177 994308
rect 136143 994220 136209 994223
rect 156258 994220 156318 995818
rect 157314 995407 157374 995818
rect 157263 995402 157374 995407
rect 157263 995346 157268 995402
rect 157324 995346 157374 995402
rect 157263 995344 157374 995346
rect 157263 995341 157329 995344
rect 156399 995256 156465 995259
rect 157890 995256 157950 995818
rect 158274 995788 158496 995848
rect 161487 995846 161760 995848
rect 161487 995790 161492 995846
rect 161548 995790 161760 995846
rect 183759 995846 189246 995848
rect 161487 995788 161760 995790
rect 158274 995700 158334 995788
rect 161487 995785 161553 995788
rect 158274 995640 158526 995700
rect 156399 995254 157950 995256
rect 156399 995198 156404 995254
rect 156460 995198 157950 995254
rect 156399 995196 157950 995198
rect 156399 995193 156465 995196
rect 136143 994218 156318 994220
rect 136143 994162 136148 994218
rect 136204 994162 156318 994218
rect 136143 994160 156318 994162
rect 136143 994157 136209 994160
rect 129711 994072 129777 994075
rect 158466 994072 158526 995640
rect 161679 995256 161745 995259
rect 162210 995256 162270 995818
rect 183759 995790 183764 995846
rect 183820 995790 189246 995846
rect 183759 995788 189246 995790
rect 183759 995785 183825 995788
rect 189186 995404 189246 995788
rect 192495 995846 195345 995848
rect 192495 995790 192500 995846
rect 192556 995790 195284 995846
rect 195340 995790 195345 995846
rect 192495 995788 195345 995790
rect 201120 995788 201534 995848
rect 192495 995785 192561 995788
rect 195279 995785 195345 995788
rect 197199 995700 197265 995703
rect 201474 995700 201534 995788
rect 202242 995700 202302 995818
rect 197199 995698 202302 995700
rect 197199 995642 197204 995698
rect 197260 995642 202302 995698
rect 197199 995640 202302 995642
rect 202434 995788 202848 995848
rect 203055 995846 203328 995848
rect 203055 995790 203060 995846
rect 203116 995790 203328 995846
rect 203055 995788 203328 995790
rect 203631 995846 203904 995848
rect 203631 995790 203636 995846
rect 203692 995790 203904 995846
rect 203631 995788 203904 995790
rect 204687 995846 204960 995848
rect 204687 995790 204692 995846
rect 204748 995790 204960 995846
rect 204687 995788 204960 995790
rect 205890 995788 206112 995848
rect 197199 995637 197265 995640
rect 189423 995552 189489 995555
rect 202434 995552 202494 995788
rect 203055 995785 203121 995788
rect 203631 995785 203697 995788
rect 204687 995785 204753 995788
rect 189423 995550 202494 995552
rect 189423 995494 189428 995550
rect 189484 995494 202494 995550
rect 189423 995492 202494 995494
rect 189423 995489 189489 995492
rect 205890 995404 205950 995788
rect 189186 995344 205950 995404
rect 161679 995254 162270 995256
rect 161679 995198 161684 995254
rect 161740 995198 162270 995254
rect 161679 995196 162270 995198
rect 198639 995256 198705 995259
rect 206562 995256 206622 995818
rect 207648 995788 207870 995848
rect 207810 995700 207870 995788
rect 198639 995254 206622 995256
rect 198639 995198 198644 995254
rect 198700 995198 206622 995254
rect 198639 995196 206622 995198
rect 207618 995640 207870 995700
rect 161679 995193 161745 995196
rect 198639 995193 198705 995196
rect 129711 994070 158526 994072
rect 129711 994014 129716 994070
rect 129772 994014 158526 994070
rect 129711 994012 158526 994014
rect 187311 994072 187377 994075
rect 207618 994072 207678 995640
rect 208770 995407 208830 995818
rect 208719 995402 208830 995407
rect 208719 995346 208724 995402
rect 208780 995346 208830 995402
rect 208719 995344 208830 995346
rect 208719 995341 208785 995344
rect 209826 995259 209886 995818
rect 212802 995700 212862 995936
rect 219087 995933 219153 995936
rect 254511 995996 254577 995999
rect 254895 995996 254961 995999
rect 261039 995996 261105 995999
rect 263247 995996 263313 995999
rect 254511 995994 254688 995996
rect 254511 995938 254516 995994
rect 254572 995938 254688 995994
rect 254511 995936 254688 995938
rect 254895 995994 255264 995996
rect 254895 995938 254900 995994
rect 254956 995938 255264 995994
rect 254895 995936 255264 995938
rect 261039 995994 261216 995996
rect 261039 995938 261044 995994
rect 261100 995938 261216 995994
rect 261039 995936 261216 995938
rect 263247 995994 263424 995996
rect 263247 995938 263252 995994
rect 263308 995938 263424 995994
rect 263247 995936 263424 995938
rect 254511 995933 254577 995936
rect 254895 995933 254961 995936
rect 261039 995933 261105 995936
rect 263247 995933 263313 995936
rect 213327 995848 213393 995851
rect 213120 995846 213393 995848
rect 213120 995790 213332 995846
rect 213388 995790 213393 995846
rect 213120 995788 213393 995790
rect 213327 995785 213393 995788
rect 239535 995848 239601 995851
rect 250479 995848 250545 995851
rect 256143 995848 256209 995851
rect 257103 995848 257169 995851
rect 259215 995848 259281 995851
rect 270735 995848 270801 995851
rect 239535 995846 250545 995848
rect 239535 995790 239540 995846
rect 239596 995790 250484 995846
rect 250540 995790 250545 995846
rect 239535 995788 250545 995790
rect 239535 995785 239601 995788
rect 250479 995785 250545 995788
rect 216015 995700 216081 995703
rect 212802 995698 216081 995700
rect 212802 995642 216020 995698
rect 216076 995642 216081 995698
rect 212802 995640 216081 995642
rect 216015 995637 216081 995640
rect 240783 995700 240849 995703
rect 251970 995700 252030 995818
rect 252738 995788 253152 995848
rect 256143 995846 256416 995848
rect 252738 995700 252798 995788
rect 240783 995698 250302 995700
rect 240783 995642 240788 995698
rect 240844 995642 250302 995698
rect 240783 995640 250302 995642
rect 251970 995640 252798 995700
rect 240783 995637 240849 995640
rect 243855 995552 243921 995555
rect 250095 995552 250161 995555
rect 243855 995550 250161 995552
rect 243855 995494 243860 995550
rect 243916 995494 250100 995550
rect 250156 995494 250161 995550
rect 243855 995492 250161 995494
rect 250242 995552 250302 995640
rect 254178 995552 254238 995818
rect 250242 995492 254238 995552
rect 243855 995489 243921 995492
rect 250095 995489 250161 995492
rect 240207 995404 240273 995407
rect 255810 995404 255870 995818
rect 256143 995790 256148 995846
rect 256204 995790 256416 995846
rect 257103 995846 257472 995848
rect 256143 995788 256416 995790
rect 256143 995785 256209 995788
rect 255951 995700 256017 995703
rect 256866 995700 256926 995818
rect 257103 995790 257108 995846
rect 257164 995790 257472 995846
rect 259215 995846 259680 995848
rect 257103 995788 257472 995790
rect 257103 995785 257169 995788
rect 255951 995698 256926 995700
rect 255951 995642 255956 995698
rect 256012 995642 256926 995698
rect 255951 995640 256926 995642
rect 255951 995637 256017 995640
rect 259074 995555 259134 995818
rect 259215 995790 259220 995846
rect 259276 995790 259680 995846
rect 259215 995788 259680 995790
rect 259215 995785 259281 995788
rect 259023 995550 259134 995555
rect 259023 995494 259028 995550
rect 259084 995494 259134 995550
rect 259023 995492 259134 995494
rect 259023 995489 259089 995492
rect 240207 995402 255870 995404
rect 240207 995346 240212 995402
rect 240268 995346 255870 995402
rect 240207 995344 255870 995346
rect 240207 995341 240273 995344
rect 260130 995259 260190 995818
rect 209775 995254 209886 995259
rect 209775 995198 209780 995254
rect 209836 995198 209886 995254
rect 209775 995196 209886 995198
rect 241743 995256 241809 995259
rect 256143 995256 256209 995259
rect 241743 995254 256209 995256
rect 241743 995198 241748 995254
rect 241804 995198 256148 995254
rect 256204 995198 256209 995254
rect 241743 995196 256209 995198
rect 209775 995193 209841 995196
rect 241743 995193 241809 995196
rect 256143 995193 256209 995196
rect 260079 995254 260190 995259
rect 260079 995198 260084 995254
rect 260140 995198 260190 995254
rect 260079 995196 260190 995198
rect 260079 995193 260145 995196
rect 250095 995108 250161 995111
rect 260706 995108 260766 995818
rect 263970 995552 264030 995818
rect 264480 995788 264894 995848
rect 265056 995846 270801 995848
rect 265056 995790 270740 995846
rect 270796 995790 270801 995846
rect 265056 995788 270801 995790
rect 264834 995700 264894 995788
rect 270735 995785 270801 995788
rect 287919 995848 287985 995851
rect 297474 995848 297534 996084
rect 299535 996081 299601 996084
rect 313167 996144 313233 996147
rect 314799 996144 314865 996147
rect 313167 996142 313440 996144
rect 313167 996086 313172 996142
rect 313228 996086 313440 996142
rect 313167 996084 313440 996086
rect 314799 996142 314976 996144
rect 314799 996086 314804 996142
rect 314860 996086 314976 996142
rect 314799 996084 314976 996086
rect 313167 996081 313233 996084
rect 314799 996081 314865 996084
rect 303951 995996 304017 995999
rect 303648 995994 304017 995996
rect 303648 995938 303956 995994
rect 304012 995938 304017 995994
rect 303648 995936 304017 995938
rect 303951 995933 304017 995936
rect 304335 995996 304401 995999
rect 305487 995996 305553 995999
rect 310287 995996 310353 995999
rect 319599 995996 319665 995999
rect 363951 995996 364017 995999
rect 304335 995994 304704 995996
rect 304335 995938 304340 995994
rect 304396 995938 304704 995994
rect 304335 995936 304704 995938
rect 305487 995994 305760 995996
rect 305487 995938 305492 995994
rect 305548 995938 305760 995994
rect 305487 995936 305760 995938
rect 310287 995994 310656 995996
rect 310287 995938 310292 995994
rect 310348 995938 310656 995994
rect 310287 995936 310656 995938
rect 316704 995994 319665 995996
rect 316704 995938 319604 995994
rect 319660 995938 319665 995994
rect 316704 995936 319665 995938
rect 363744 995994 364017 995996
rect 363744 995938 363956 995994
rect 364012 995938 364017 995994
rect 363744 995936 364017 995938
rect 304335 995933 304401 995936
rect 305487 995933 305553 995936
rect 310287 995933 310353 995936
rect 319599 995933 319665 995936
rect 363951 995933 364017 995936
rect 421551 995996 421617 995999
rect 421890 995996 421950 1015768
rect 435279 1006356 435345 1006359
rect 465615 1006356 465681 1006359
rect 435279 1006354 465681 1006356
rect 435279 1006298 435284 1006354
rect 435340 1006298 465620 1006354
rect 465676 1006298 465681 1006354
rect 435279 1006296 465681 1006298
rect 435279 1006293 435345 1006296
rect 465615 1006293 465681 1006296
rect 435183 1006060 435249 1006063
rect 466095 1006060 466161 1006063
rect 435183 1006058 466161 1006060
rect 435183 1006002 435188 1006058
rect 435244 1006002 466100 1006058
rect 466156 1006002 466161 1006058
rect 435183 1006000 466161 1006002
rect 435183 1005997 435249 1006000
rect 466095 1005997 466161 1006000
rect 435087 1005912 435153 1005915
rect 465231 1005912 465297 1005915
rect 435087 1005910 465297 1005912
rect 435087 1005854 435092 1005910
rect 435148 1005854 465236 1005910
rect 465292 1005854 465297 1005910
rect 435087 1005852 465297 1005854
rect 435087 1005849 435153 1005852
rect 465231 1005849 465297 1005852
rect 428655 1003248 428721 1003251
rect 502383 1003248 502449 1003251
rect 428448 1003246 428721 1003248
rect 428448 1003190 428660 1003246
rect 428716 1003190 428721 1003246
rect 428448 1003188 428721 1003190
rect 502176 1003246 502449 1003248
rect 502176 1003190 502388 1003246
rect 502444 1003190 502449 1003246
rect 502176 1003188 502449 1003190
rect 428655 1003185 428721 1003188
rect 502383 1003185 502449 1003188
rect 425391 1003100 425457 1003103
rect 428271 1003100 428337 1003103
rect 430287 1003100 430353 1003103
rect 501327 1003100 501393 1003103
rect 502959 1003100 503025 1003103
rect 555375 1003100 555441 1003103
rect 425184 1003098 425457 1003100
rect 425184 1003042 425396 1003098
rect 425452 1003042 425457 1003098
rect 425184 1003040 425457 1003042
rect 427968 1003098 428337 1003100
rect 427968 1003042 428276 1003098
rect 428332 1003042 428337 1003098
rect 427968 1003040 428337 1003042
rect 430176 1003098 430353 1003100
rect 430176 1003042 430292 1003098
rect 430348 1003042 430353 1003098
rect 430176 1003040 430353 1003042
rect 501120 1003098 501393 1003100
rect 501120 1003042 501332 1003098
rect 501388 1003042 501393 1003098
rect 501120 1003040 501393 1003042
rect 502752 1003098 503025 1003100
rect 502752 1003042 502964 1003098
rect 503020 1003042 503025 1003098
rect 502752 1003040 503025 1003042
rect 555264 1003098 555441 1003100
rect 555264 1003042 555380 1003098
rect 555436 1003042 555441 1003098
rect 555264 1003040 555441 1003042
rect 425391 1003037 425457 1003040
rect 428271 1003037 428337 1003040
rect 430287 1003037 430353 1003040
rect 501327 1003037 501393 1003040
rect 502959 1003037 503025 1003040
rect 555375 1003037 555441 1003040
rect 423855 1002952 423921 1002955
rect 426063 1002952 426129 1002955
rect 553743 1002952 553809 1002955
rect 554319 1002952 554385 1002955
rect 423648 1002950 423921 1002952
rect 423648 1002894 423860 1002950
rect 423916 1002894 423921 1002950
rect 423648 1002892 423921 1002894
rect 425760 1002950 426129 1002952
rect 425760 1002894 426068 1002950
rect 426124 1002894 426129 1002950
rect 425760 1002892 426129 1002894
rect 553632 1002950 553809 1002952
rect 553632 1002894 553748 1002950
rect 553804 1002894 553809 1002950
rect 553632 1002892 553809 1002894
rect 554208 1002950 554385 1002952
rect 554208 1002894 554324 1002950
rect 554380 1002894 554385 1002950
rect 554208 1002892 554385 1002894
rect 423855 1002889 423921 1002892
rect 426063 1002889 426129 1002892
rect 553743 1002889 553809 1002892
rect 554319 1002889 554385 1002892
rect 424335 1002804 424401 1002807
rect 424815 1002804 424881 1002807
rect 432015 1002804 432081 1002807
rect 554895 1002804 554961 1002807
rect 424128 1002802 424401 1002804
rect 424128 1002746 424340 1002802
rect 424396 1002746 424401 1002802
rect 424128 1002744 424401 1002746
rect 424704 1002802 424881 1002804
rect 424704 1002746 424820 1002802
rect 424876 1002746 424881 1002802
rect 424704 1002744 424881 1002746
rect 431712 1002802 432081 1002804
rect 431712 1002746 432020 1002802
rect 432076 1002746 432081 1002802
rect 431712 1002744 432081 1002746
rect 554688 1002802 554961 1002804
rect 554688 1002746 554900 1002802
rect 554956 1002746 554961 1002802
rect 554688 1002744 554961 1002746
rect 424335 1002741 424401 1002744
rect 424815 1002741 424881 1002744
rect 432015 1002741 432081 1002744
rect 554895 1002741 554961 1002744
rect 427599 1002656 427665 1002659
rect 429231 1002656 429297 1002659
rect 553263 1002656 553329 1002659
rect 427392 1002654 427665 1002656
rect 427392 1002598 427604 1002654
rect 427660 1002598 427665 1002654
rect 427392 1002596 427665 1002598
rect 429024 1002654 429297 1002656
rect 429024 1002598 429236 1002654
rect 429292 1002598 429297 1002654
rect 429024 1002596 429297 1002598
rect 553056 1002654 553329 1002656
rect 553056 1002598 553268 1002654
rect 553324 1002598 553329 1002654
rect 553056 1002596 553329 1002598
rect 427599 1002593 427665 1002596
rect 429231 1002593 429297 1002596
rect 553263 1002593 553329 1002596
rect 426639 1002508 426705 1002511
rect 427119 1002508 427185 1002511
rect 426336 1002506 426705 1002508
rect 426336 1002450 426644 1002506
rect 426700 1002450 426705 1002506
rect 426336 1002448 426705 1002450
rect 426912 1002506 427185 1002508
rect 426912 1002450 427124 1002506
rect 427180 1002450 427185 1002506
rect 426912 1002448 427185 1002450
rect 426639 1002445 426705 1002448
rect 427119 1002445 427185 1002448
rect 506319 1001028 506385 1001031
rect 506016 1001026 506385 1001028
rect 506016 1000970 506324 1001026
rect 506380 1000970 506385 1001026
rect 506016 1000968 506385 1000970
rect 506319 1000965 506385 1000968
rect 429903 1000880 429969 1000883
rect 430959 1000880 431025 1000883
rect 507855 1000880 507921 1000883
rect 552303 1000880 552369 1000883
rect 429600 1000878 429969 1000880
rect 429600 1000822 429908 1000878
rect 429964 1000822 429969 1000878
rect 429600 1000820 429969 1000822
rect 430656 1000878 431025 1000880
rect 430656 1000822 430964 1000878
rect 431020 1000822 431025 1000878
rect 430656 1000820 431025 1000822
rect 507648 1000878 507921 1000880
rect 507648 1000822 507860 1000878
rect 507916 1000822 507921 1000878
rect 507648 1000820 507921 1000822
rect 552000 1000878 552369 1000880
rect 552000 1000822 552308 1000878
rect 552364 1000822 552369 1000878
rect 552000 1000820 552369 1000822
rect 429903 1000817 429969 1000820
rect 430959 1000817 431025 1000820
rect 507855 1000817 507921 1000820
rect 552303 1000817 552369 1000820
rect 506895 1000732 506961 1000735
rect 506592 1000730 506961 1000732
rect 506592 1000674 506900 1000730
rect 506956 1000674 506961 1000730
rect 506592 1000672 506961 1000674
rect 506895 1000669 506961 1000672
rect 515535 1000288 515601 1000291
rect 523503 1000288 523569 1000291
rect 515535 1000286 523569 1000288
rect 515535 1000230 515540 1000286
rect 515596 1000230 523508 1000286
rect 523564 1000230 523569 1000286
rect 515535 1000228 523569 1000230
rect 515535 1000225 515601 1000228
rect 523503 1000225 523569 1000228
rect 512655 1000140 512721 1000143
rect 523599 1000140 523665 1000143
rect 512655 1000138 523665 1000140
rect 512655 1000082 512660 1000138
rect 512716 1000082 523604 1000138
rect 523660 1000082 523665 1000138
rect 512655 1000080 523665 1000082
rect 512655 1000077 512721 1000080
rect 523599 1000077 523665 1000080
rect 512271 999992 512337 999995
rect 523695 999992 523761 999995
rect 512271 999990 523761 999992
rect 512271 999934 512276 999990
rect 512332 999934 523700 999990
rect 523756 999934 523761 999990
rect 512271 999932 523761 999934
rect 512271 999929 512337 999932
rect 523695 999929 523761 999932
rect 504687 999844 504753 999847
rect 504384 999842 504753 999844
rect 504384 999786 504692 999842
rect 504748 999786 504753 999842
rect 504384 999784 504753 999786
rect 504687 999781 504753 999784
rect 512079 999844 512145 999847
rect 523983 999844 524049 999847
rect 512079 999842 524049 999844
rect 512079 999786 512084 999842
rect 512140 999786 523988 999842
rect 524044 999786 524049 999842
rect 512079 999784 524049 999786
rect 512079 999781 512145 999784
rect 523983 999781 524049 999784
rect 500751 999696 500817 999699
rect 500640 999694 500817 999696
rect 500640 999638 500756 999694
rect 500812 999638 500817 999694
rect 500640 999636 500817 999638
rect 500751 999633 500817 999636
rect 503631 999696 503697 999699
rect 512079 999696 512145 999699
rect 523791 999696 523857 999699
rect 503631 999694 503904 999696
rect 503631 999638 503636 999694
rect 503692 999638 503904 999694
rect 503631 999636 503904 999638
rect 512079 999694 523857 999696
rect 512079 999638 512084 999694
rect 512140 999638 523796 999694
rect 523852 999638 523857 999694
rect 512079 999636 523857 999638
rect 503631 999633 503697 999636
rect 512079 999633 512145 999636
rect 523791 999633 523857 999636
rect 501999 999548 502065 999551
rect 503631 999548 503697 999551
rect 501696 999546 502065 999548
rect 501696 999490 502004 999546
rect 502060 999490 502065 999546
rect 501696 999488 502065 999490
rect 503328 999546 503697 999548
rect 503328 999490 503636 999546
rect 503692 999490 503697 999546
rect 503328 999488 503697 999490
rect 501999 999485 502065 999488
rect 503631 999485 503697 999488
rect 512175 999548 512241 999551
rect 523887 999548 523953 999551
rect 512175 999546 523953 999548
rect 512175 999490 512180 999546
rect 512236 999490 523892 999546
rect 523948 999490 523953 999546
rect 512175 999488 523953 999490
rect 512175 999485 512241 999488
rect 523887 999485 523953 999488
rect 512079 999400 512145 999403
rect 524079 999400 524145 999403
rect 552879 999400 552945 999403
rect 512079 999398 524145 999400
rect 512079 999342 512084 999398
rect 512140 999342 524084 999398
rect 524140 999342 524145 999398
rect 512079 999340 524145 999342
rect 552480 999398 552945 999400
rect 552480 999342 552884 999398
rect 552940 999342 552945 999398
rect 552480 999340 552945 999342
rect 512079 999337 512145 999340
rect 524079 999337 524145 999340
rect 552879 999337 552945 999340
rect 558831 999252 558897 999255
rect 558528 999250 558897 999252
rect 558528 999194 558836 999250
rect 558892 999194 558897 999250
rect 558528 999192 558897 999194
rect 558831 999189 558897 999192
rect 557199 998808 557265 998811
rect 556896 998806 557265 998808
rect 556896 998750 557204 998806
rect 557260 998750 557265 998806
rect 556896 998748 557265 998750
rect 557199 998745 557265 998748
rect 555951 997920 556017 997923
rect 555744 997918 556017 997920
rect 555744 997862 555956 997918
rect 556012 997862 556017 997918
rect 555744 997860 556017 997862
rect 555951 997857 556017 997860
rect 558159 997772 558225 997775
rect 557952 997770 558225 997772
rect 557952 997714 558164 997770
rect 558220 997714 558225 997770
rect 557952 997712 558225 997714
rect 558159 997709 558225 997712
rect 557775 997624 557841 997627
rect 559407 997624 559473 997627
rect 557472 997622 557841 997624
rect 557472 997566 557780 997622
rect 557836 997566 557841 997622
rect 557472 997564 557841 997566
rect 559008 997622 559473 997624
rect 559008 997566 559412 997622
rect 559468 997566 559473 997622
rect 559008 997564 559473 997566
rect 557775 997561 557841 997564
rect 559407 997561 559473 997564
rect 505743 996588 505809 996591
rect 507471 996588 507537 996591
rect 505440 996586 505809 996588
rect 505440 996530 505748 996586
rect 505804 996530 505809 996586
rect 505440 996528 505809 996530
rect 507168 996586 507537 996588
rect 507168 996530 507476 996586
rect 507532 996530 507537 996586
rect 507168 996528 507537 996530
rect 505743 996525 505809 996528
rect 507471 996525 507537 996528
rect 432495 996292 432561 996295
rect 432495 996290 432864 996292
rect 432495 996234 432500 996290
rect 432556 996234 432864 996290
rect 432495 996232 432864 996234
rect 432495 996229 432561 996232
rect 432495 996144 432561 996147
rect 508911 996144 508977 996147
rect 432288 996142 432561 996144
rect 432288 996086 432500 996142
rect 432556 996086 432561 996142
rect 432288 996084 432561 996086
rect 508704 996142 508977 996144
rect 508704 996086 508916 996142
rect 508972 996086 508977 996142
rect 508704 996084 508977 996086
rect 432495 996081 432561 996084
rect 508911 996081 508977 996084
rect 509583 996144 509649 996147
rect 519855 996144 519921 996147
rect 528250 996144 528256 996146
rect 509583 996142 509856 996144
rect 509583 996086 509588 996142
rect 509644 996086 509856 996142
rect 509583 996084 509856 996086
rect 519855 996142 528256 996144
rect 519855 996086 519860 996142
rect 519916 996086 528256 996142
rect 519855 996084 528256 996086
rect 509583 996081 509649 996084
rect 519855 996081 519921 996084
rect 528250 996082 528256 996084
rect 528320 996082 528326 996146
rect 561039 996144 561105 996147
rect 561039 996142 561216 996144
rect 561039 996086 561044 996142
rect 561100 996086 561216 996142
rect 561039 996084 561216 996086
rect 561039 996081 561105 996084
rect 421551 995994 421950 995996
rect 421551 995938 421556 995994
rect 421612 995966 421950 995994
rect 430959 995996 431025 995999
rect 437871 995996 437937 995999
rect 508335 995996 508401 995999
rect 515535 995996 515601 995999
rect 430959 995994 431232 995996
rect 421612 995938 421920 995966
rect 421551 995936 421920 995938
rect 430959 995938 430964 995994
rect 431020 995938 431232 995994
rect 430959 995936 431232 995938
rect 434496 995994 437937 995996
rect 434496 995938 437876 995994
rect 437932 995938 437937 995994
rect 434496 995936 437937 995938
rect 508224 995994 508401 995996
rect 508224 995938 508340 995994
rect 508396 995938 508401 995994
rect 508224 995936 508401 995938
rect 511488 995994 515601 995996
rect 511488 995938 515540 995994
rect 515596 995938 515601 995994
rect 511488 995936 515601 995938
rect 421551 995933 421617 995936
rect 430959 995933 431025 995936
rect 437871 995933 437937 995936
rect 508335 995933 508401 995936
rect 515535 995933 515601 995936
rect 519759 995996 519825 995999
rect 519759 995994 528702 995996
rect 519759 995938 519764 995994
rect 519820 995938 528702 995994
rect 519759 995936 528702 995938
rect 519759 995933 519825 995936
rect 299343 995848 299409 995851
rect 305967 995848 306033 995851
rect 307599 995848 307665 995851
rect 360879 995848 360945 995851
rect 366159 995848 366225 995851
rect 366735 995848 366801 995851
rect 371535 995848 371601 995851
rect 287919 995846 297534 995848
rect 287919 995790 287924 995846
rect 287980 995790 297534 995846
rect 287919 995788 297534 995790
rect 298050 995846 299409 995848
rect 298050 995790 299348 995846
rect 299404 995790 299409 995846
rect 298050 995788 299409 995790
rect 287919 995785 287985 995788
rect 267855 995700 267921 995703
rect 264834 995698 267921 995700
rect 264834 995642 267860 995698
rect 267916 995642 267921 995698
rect 264834 995640 267921 995642
rect 267855 995637 267921 995640
rect 286767 995700 286833 995703
rect 298050 995700 298110 995788
rect 299343 995785 299409 995788
rect 286767 995698 298110 995700
rect 286767 995642 286772 995698
rect 286828 995642 298110 995698
rect 286767 995640 298110 995642
rect 298959 995700 299025 995703
rect 304098 995700 304158 995818
rect 305184 995788 305406 995848
rect 305346 995700 305406 995788
rect 305967 995846 306336 995848
rect 305967 995790 305972 995846
rect 306028 995790 306336 995846
rect 305967 995788 306336 995790
rect 306690 995788 306912 995848
rect 307599 995846 307968 995848
rect 305967 995785 306033 995788
rect 298959 995698 305406 995700
rect 298959 995642 298964 995698
rect 299020 995642 305406 995698
rect 298959 995640 305406 995642
rect 286767 995637 286833 995640
rect 298959 995637 299025 995640
rect 267951 995552 268017 995555
rect 263970 995550 268017 995552
rect 263970 995494 267956 995550
rect 268012 995494 268017 995550
rect 263970 995492 268017 995494
rect 267951 995489 268017 995492
rect 287439 995552 287505 995555
rect 299247 995552 299313 995555
rect 287439 995550 299313 995552
rect 287439 995494 287444 995550
rect 287500 995494 299252 995550
rect 299308 995494 299313 995550
rect 287439 995492 299313 995494
rect 287439 995489 287505 995492
rect 299247 995489 299313 995492
rect 299535 995552 299601 995555
rect 306690 995552 306750 995788
rect 299535 995550 306750 995552
rect 299535 995494 299540 995550
rect 299596 995494 306750 995550
rect 299535 995492 306750 995494
rect 299535 995489 299601 995492
rect 291471 995256 291537 995259
rect 307362 995256 307422 995818
rect 307599 995790 307604 995846
rect 307660 995790 307968 995846
rect 307599 995788 307968 995790
rect 307599 995785 307665 995788
rect 291471 995254 307422 995256
rect 291471 995198 291476 995254
rect 291532 995198 307422 995254
rect 291471 995196 307422 995198
rect 291471 995193 291537 995196
rect 250095 995106 260766 995108
rect 250095 995050 250100 995106
rect 250156 995050 260766 995106
rect 250095 995048 260766 995050
rect 250095 995045 250161 995048
rect 235791 994664 235857 994667
rect 247599 994664 247665 994667
rect 235791 994662 247665 994664
rect 235791 994606 235796 994662
rect 235852 994606 247604 994662
rect 247660 994606 247665 994662
rect 235791 994604 247665 994606
rect 235791 994601 235857 994604
rect 247599 994601 247665 994604
rect 232143 994516 232209 994519
rect 247503 994516 247569 994519
rect 232143 994514 247569 994516
rect 232143 994458 232148 994514
rect 232204 994458 247508 994514
rect 247564 994458 247569 994514
rect 232143 994456 247569 994458
rect 232143 994453 232209 994456
rect 247503 994453 247569 994456
rect 285999 994516 286065 994519
rect 311202 994516 311262 995818
rect 312834 995407 312894 995818
rect 315522 995700 315582 995818
rect 353952 995788 354366 995848
rect 360480 995846 360945 995848
rect 319695 995700 319761 995703
rect 315522 995698 319761 995700
rect 315522 995642 319700 995698
rect 319756 995642 319761 995698
rect 315522 995640 319761 995642
rect 354306 995700 354366 995788
rect 355074 995700 355134 995818
rect 360480 995790 360884 995846
rect 360940 995790 360945 995846
rect 365952 995846 366225 995848
rect 360480 995788 360945 995790
rect 360879 995785 360945 995788
rect 354306 995640 355134 995700
rect 319695 995637 319761 995640
rect 312783 995402 312894 995407
rect 312783 995346 312788 995402
rect 312844 995346 312894 995402
rect 312783 995344 312894 995346
rect 312783 995341 312849 995344
rect 363234 995256 363294 995818
rect 364866 995700 364926 995818
rect 365952 995790 366164 995846
rect 366220 995790 366225 995846
rect 365952 995788 366225 995790
rect 366528 995846 366801 995848
rect 366528 995790 366740 995846
rect 366796 995790 366801 995846
rect 366528 995788 366801 995790
rect 367008 995846 371601 995848
rect 367008 995790 371540 995846
rect 371596 995790 371601 995846
rect 367008 995788 371601 995790
rect 366159 995785 366225 995788
rect 366735 995785 366801 995788
rect 371535 995785 371601 995788
rect 383535 995848 383601 995851
rect 387471 995848 387537 995851
rect 472239 995848 472305 995851
rect 478383 995848 478449 995851
rect 499311 995848 499377 995851
rect 523695 995848 523761 995851
rect 528399 995848 528465 995851
rect 383535 995846 387537 995848
rect 383535 995790 383540 995846
rect 383596 995790 387476 995846
rect 387532 995790 387537 995846
rect 383535 995788 387537 995790
rect 383535 995785 383601 995788
rect 387471 995785 387537 995788
rect 368655 995700 368721 995703
rect 364866 995698 368721 995700
rect 364866 995642 368660 995698
rect 368716 995642 368721 995698
rect 364866 995640 368721 995642
rect 368655 995637 368721 995640
rect 383055 995700 383121 995703
rect 391791 995700 391857 995703
rect 383055 995698 391857 995700
rect 383055 995642 383060 995698
rect 383116 995642 391796 995698
rect 391852 995642 391857 995698
rect 383055 995640 391857 995642
rect 421410 995700 421470 995818
rect 422466 995700 422526 995818
rect 421410 995640 422526 995700
rect 433218 995788 433440 995848
rect 472239 995846 478449 995848
rect 433218 995700 433278 995788
rect 433890 995700 433950 995818
rect 472239 995790 472244 995846
rect 472300 995790 478388 995846
rect 478444 995790 478449 995846
rect 498912 995846 499377 995848
rect 472239 995788 478449 995790
rect 472239 995785 472305 995788
rect 478383 995785 478449 995788
rect 437775 995700 437841 995703
rect 433218 995640 433470 995700
rect 433890 995698 437841 995700
rect 433890 995642 437780 995698
rect 437836 995642 437841 995698
rect 433890 995640 437841 995642
rect 383055 995637 383121 995640
rect 391791 995637 391857 995640
rect 433410 995552 433470 995640
rect 437775 995637 437841 995640
rect 472047 995700 472113 995703
rect 482031 995700 482097 995703
rect 472047 995698 482097 995700
rect 472047 995642 472052 995698
rect 472108 995642 482036 995698
rect 482092 995642 482097 995698
rect 472047 995640 482097 995642
rect 498402 995700 498462 995818
rect 498912 995790 499316 995846
rect 499372 995790 499377 995846
rect 498912 995788 499377 995790
rect 499311 995785 499377 995788
rect 499458 995700 499518 995818
rect 498402 995640 499518 995700
rect 472047 995637 472113 995640
rect 482031 995637 482097 995640
rect 437967 995552 438033 995555
rect 433410 995550 438033 995552
rect 433410 995494 437972 995550
rect 438028 995494 438033 995550
rect 433410 995492 438033 995494
rect 437967 995489 438033 995492
rect 465615 995552 465681 995555
rect 477039 995552 477105 995555
rect 465615 995550 477105 995552
rect 465615 995494 465620 995550
rect 465676 995494 477044 995550
rect 477100 995494 477105 995550
rect 465615 995492 477105 995494
rect 465615 995489 465681 995492
rect 477039 995489 477105 995492
rect 499311 995552 499377 995555
rect 500034 995552 500094 995818
rect 501807 995552 501873 995555
rect 499311 995550 501873 995552
rect 499311 995494 499316 995550
rect 499372 995494 501812 995550
rect 501868 995494 501873 995550
rect 499311 995492 501873 995494
rect 504930 995552 504990 995818
rect 509250 995700 509310 995818
rect 510210 995788 510432 995848
rect 523695 995846 528465 995848
rect 509967 995700 510033 995703
rect 509250 995698 510033 995700
rect 509250 995642 509972 995698
rect 510028 995642 510033 995698
rect 509250 995640 510033 995642
rect 510210 995700 510270 995788
rect 510882 995700 510942 995818
rect 523695 995790 523700 995846
rect 523756 995790 528404 995846
rect 528460 995790 528465 995846
rect 523695 995788 528465 995790
rect 528642 995848 528702 995936
rect 532815 995848 532881 995851
rect 528642 995846 532881 995848
rect 528642 995790 532820 995846
rect 532876 995790 532881 995846
rect 550479 995848 550545 995851
rect 556527 995848 556593 995851
rect 569967 995848 570033 995851
rect 550479 995846 550944 995848
rect 528642 995788 532881 995790
rect 523695 995785 523761 995788
rect 528399 995785 528465 995788
rect 532815 995785 532881 995788
rect 515631 995700 515697 995703
rect 510210 995640 510462 995700
rect 510882 995698 515697 995700
rect 510882 995642 515636 995698
rect 515692 995642 515697 995698
rect 510882 995640 515697 995642
rect 509967 995637 510033 995640
rect 510255 995552 510321 995555
rect 504930 995550 510321 995552
rect 504930 995494 510260 995550
rect 510316 995494 510321 995550
rect 504930 995492 510321 995494
rect 510402 995552 510462 995640
rect 515631 995637 515697 995640
rect 523503 995700 523569 995703
rect 527823 995700 527889 995703
rect 533391 995700 533457 995703
rect 523503 995698 527889 995700
rect 523503 995642 523508 995698
rect 523564 995642 527828 995698
rect 527884 995642 527889 995698
rect 523503 995640 527889 995642
rect 523503 995637 523569 995640
rect 527823 995637 527889 995640
rect 528066 995698 533457 995700
rect 528066 995642 533396 995698
rect 533452 995642 533457 995698
rect 528066 995640 533457 995642
rect 515727 995552 515793 995555
rect 510402 995550 515793 995552
rect 510402 995494 515732 995550
rect 515788 995494 515793 995550
rect 510402 995492 515793 995494
rect 499311 995489 499377 995492
rect 501807 995489 501873 995492
rect 510255 995489 510321 995492
rect 515727 995489 515793 995492
rect 519663 995552 519729 995555
rect 528066 995552 528126 995640
rect 533391 995637 533457 995640
rect 519663 995550 528126 995552
rect 519663 995494 519668 995550
rect 519724 995494 528126 995550
rect 519663 995492 528126 995494
rect 519663 995489 519729 995492
rect 528250 995490 528256 995554
rect 528320 995552 528326 995554
rect 535311 995552 535377 995555
rect 528320 995550 535377 995552
rect 528320 995494 535316 995550
rect 535372 995494 535377 995550
rect 528320 995492 535377 995494
rect 549762 995552 549822 995818
rect 550338 995700 550398 995818
rect 550479 995790 550484 995846
rect 550540 995790 550944 995846
rect 556320 995846 556593 995848
rect 550479 995788 550944 995790
rect 550479 995785 550545 995788
rect 551394 995700 551454 995818
rect 556320 995790 556532 995846
rect 556588 995790 556593 995846
rect 556320 995788 556593 995790
rect 556527 995785 556593 995788
rect 559554 995703 559614 995818
rect 560130 995703 560190 995818
rect 560514 995788 560736 995848
rect 558927 995700 558993 995703
rect 550338 995698 558993 995700
rect 550338 995642 558932 995698
rect 558988 995642 558993 995698
rect 550338 995640 558993 995642
rect 559554 995698 559665 995703
rect 559554 995642 559604 995698
rect 559660 995642 559665 995698
rect 559554 995640 559665 995642
rect 560130 995698 560241 995703
rect 560130 995642 560180 995698
rect 560236 995642 560241 995698
rect 560130 995640 560241 995642
rect 560514 995700 560574 995788
rect 560514 995640 560766 995700
rect 558927 995637 558993 995640
rect 559599 995637 559665 995640
rect 560175 995637 560241 995640
rect 550479 995552 550545 995555
rect 549762 995550 550545 995552
rect 549762 995494 550484 995550
rect 550540 995494 550545 995550
rect 549762 995492 550545 995494
rect 528320 995490 528326 995492
rect 535311 995489 535377 995492
rect 550479 995489 550545 995492
rect 466095 995404 466161 995407
rect 477711 995404 477777 995407
rect 466095 995402 477777 995404
rect 466095 995346 466100 995402
rect 466156 995346 477716 995402
rect 477772 995346 477777 995402
rect 466095 995344 477777 995346
rect 560706 995404 560766 995640
rect 561762 995552 561822 995818
rect 562272 995788 562686 995848
rect 562848 995846 570033 995848
rect 562848 995790 569972 995846
rect 570028 995790 570033 995846
rect 562848 995788 570033 995790
rect 562626 995700 562686 995788
rect 569967 995785 570033 995788
rect 625935 995848 626001 995851
rect 629583 995848 629649 995851
rect 625935 995846 629649 995848
rect 625935 995790 625940 995846
rect 625996 995790 629588 995846
rect 629644 995790 629649 995846
rect 625935 995788 629649 995790
rect 625935 995785 626001 995788
rect 629583 995785 629649 995788
rect 569871 995700 569937 995703
rect 562626 995698 569937 995700
rect 562626 995642 569876 995698
rect 569932 995642 569937 995698
rect 562626 995640 569937 995642
rect 569871 995637 569937 995640
rect 569775 995552 569841 995555
rect 561762 995550 569841 995552
rect 561762 995494 569780 995550
rect 569836 995494 569841 995550
rect 561762 995492 569841 995494
rect 569775 995489 569841 995492
rect 567279 995404 567345 995407
rect 560706 995402 567345 995404
rect 560706 995346 567284 995402
rect 567340 995346 567345 995402
rect 560706 995344 567345 995346
rect 466095 995341 466161 995344
rect 477711 995341 477777 995344
rect 567279 995341 567345 995344
rect 385935 995256 386001 995259
rect 363234 995254 386001 995256
rect 363234 995198 385940 995254
rect 385996 995198 386001 995254
rect 363234 995196 386001 995198
rect 385935 995193 386001 995196
rect 396303 995256 396369 995259
rect 627663 995256 627729 995259
rect 396303 995254 627729 995256
rect 396303 995198 396308 995254
rect 396364 995198 627668 995254
rect 627724 995198 627729 995254
rect 396303 995196 627729 995198
rect 396303 995193 396369 995196
rect 627663 995193 627729 995196
rect 377295 994812 377361 994815
rect 390831 994812 390897 994815
rect 573903 994812 573969 994815
rect 634287 994812 634353 994815
rect 377295 994810 395454 994812
rect 377295 994754 377300 994810
rect 377356 994754 390836 994810
rect 390892 994754 395454 994810
rect 377295 994752 395454 994754
rect 377295 994749 377361 994752
rect 390831 994749 390897 994752
rect 285999 994514 311262 994516
rect 285999 994458 286004 994514
rect 286060 994458 311262 994514
rect 285999 994456 311262 994458
rect 373359 994516 373425 994519
rect 395151 994516 395217 994519
rect 373359 994514 395217 994516
rect 373359 994458 373364 994514
rect 373420 994458 395156 994514
rect 395212 994458 395217 994514
rect 373359 994456 395217 994458
rect 395394 994516 395454 994752
rect 573903 994810 634353 994812
rect 573903 994754 573908 994810
rect 573964 994754 634292 994810
rect 634348 994754 634353 994810
rect 573903 994752 634353 994754
rect 573903 994749 573969 994752
rect 634287 994749 634353 994752
rect 518319 994664 518385 994667
rect 534351 994664 534417 994667
rect 518319 994662 534417 994664
rect 518319 994606 518324 994662
rect 518380 994606 534356 994662
rect 534412 994606 534417 994662
rect 518319 994604 534417 994606
rect 518319 994601 518385 994604
rect 534351 994601 534417 994604
rect 573711 994664 573777 994667
rect 639183 994664 639249 994667
rect 573711 994662 639249 994664
rect 573711 994606 573716 994662
rect 573772 994606 639188 994662
rect 639244 994606 639249 994662
rect 573711 994604 639249 994606
rect 573711 994601 573777 994604
rect 639183 994601 639249 994604
rect 479823 994516 479889 994519
rect 531183 994516 531249 994519
rect 633039 994516 633105 994519
rect 395394 994514 633105 994516
rect 395394 994458 479828 994514
rect 479884 994458 531188 994514
rect 531244 994458 633044 994514
rect 633100 994458 633105 994514
rect 395394 994456 633105 994458
rect 285999 994453 286065 994456
rect 373359 994453 373425 994456
rect 395151 994453 395217 994456
rect 479823 994453 479889 994456
rect 531183 994453 531249 994456
rect 633039 994453 633105 994456
rect 296655 994368 296721 994371
rect 377295 994368 377361 994371
rect 296655 994366 377361 994368
rect 296655 994310 296660 994366
rect 296716 994310 377300 994366
rect 377356 994310 377361 994366
rect 296655 994308 377361 994310
rect 296655 994305 296721 994308
rect 377295 994305 377361 994308
rect 234351 994220 234417 994223
rect 259215 994220 259281 994223
rect 234351 994218 259281 994220
rect 234351 994162 234356 994218
rect 234412 994162 259220 994218
rect 259276 994162 259281 994218
rect 234351 994160 259281 994162
rect 234351 994157 234417 994160
rect 259215 994157 259281 994160
rect 294543 994220 294609 994223
rect 643311 994220 643377 994223
rect 294543 994218 643377 994220
rect 294543 994162 294548 994218
rect 294604 994162 643316 994218
rect 643372 994162 643377 994218
rect 294543 994160 643377 994162
rect 294543 994157 294609 994160
rect 643311 994157 643377 994160
rect 187311 994070 207678 994072
rect 187311 994014 187316 994070
rect 187372 994014 207678 994070
rect 187311 994012 207678 994014
rect 243183 994072 243249 994075
rect 650223 994072 650289 994075
rect 243183 994070 650289 994072
rect 243183 994014 243188 994070
rect 243244 994014 650228 994070
rect 650284 994014 650289 994070
rect 243183 994012 650289 994014
rect 129711 994009 129777 994012
rect 187311 994009 187377 994012
rect 243183 994009 243249 994012
rect 650223 994009 650289 994012
rect 88719 993924 88785 993927
rect 533679 993924 533745 993927
rect 88719 993922 533745 993924
rect 88719 993866 88724 993922
rect 88780 993866 533684 993922
rect 533740 993866 533745 993922
rect 88719 993864 533745 993866
rect 88719 993861 88785 993864
rect 533679 993861 533745 993864
rect 536751 993924 536817 993927
rect 640527 993924 640593 993927
rect 536751 993922 640593 993924
rect 536751 993866 536756 993922
rect 536812 993866 640532 993922
rect 640588 993866 640593 993922
rect 536751 993864 640593 993866
rect 536751 993861 536817 993864
rect 640527 993861 640593 993864
rect 78351 993776 78417 993779
rect 106767 993776 106833 993779
rect 134319 993776 134385 993779
rect 78351 993774 106833 993776
rect 78351 993718 78356 993774
rect 78412 993718 106772 993774
rect 106828 993718 106833 993774
rect 78351 993716 106833 993718
rect 78351 993713 78417 993716
rect 106767 993713 106833 993716
rect 134274 993774 134385 993776
rect 134274 993718 134324 993774
rect 134380 993718 134385 993774
rect 134274 993713 134385 993718
rect 140367 993776 140433 993779
rect 641103 993776 641169 993779
rect 140367 993774 641169 993776
rect 140367 993718 140372 993774
rect 140428 993718 641108 993774
rect 641164 993718 641169 993774
rect 140367 993716 641169 993718
rect 140367 993713 140433 993716
rect 641103 993713 641169 993716
rect 83439 993628 83505 993631
rect 92655 993628 92721 993631
rect 83439 993626 92721 993628
rect 83439 993570 83444 993626
rect 83500 993570 92660 993626
rect 92716 993570 92721 993626
rect 83439 993568 92721 993570
rect 83439 993565 83505 993568
rect 92655 993565 92721 993568
rect 126639 993628 126705 993631
rect 134274 993628 134334 993713
rect 186159 993628 186225 993631
rect 195471 993628 195537 993631
rect 126639 993626 195537 993628
rect 126639 993570 126644 993626
rect 126700 993570 186164 993626
rect 186220 993570 195476 993626
rect 195532 993570 195537 993626
rect 126639 993568 195537 993570
rect 126639 993565 126705 993568
rect 186159 993565 186225 993568
rect 195471 993565 195537 993568
rect 403119 993628 403185 993631
rect 479151 993628 479217 993631
rect 489135 993628 489201 993631
rect 403119 993626 489201 993628
rect 403119 993570 403124 993626
rect 403180 993570 479156 993626
rect 479212 993570 489140 993626
rect 489196 993570 489201 993626
rect 403119 993568 489201 993570
rect 403119 993565 403185 993568
rect 479151 993565 479217 993568
rect 489135 993565 489201 993568
rect 62031 992148 62097 992151
rect 83439 992148 83505 992151
rect 62031 992146 83505 992148
rect 62031 992090 62036 992146
rect 62092 992090 83444 992146
rect 83500 992090 83505 992146
rect 62031 992088 83505 992090
rect 62031 992085 62097 992088
rect 83439 992085 83505 992088
rect 655119 976756 655185 976759
rect 650208 976754 655185 976756
rect 650208 976698 655124 976754
rect 655180 976698 655185 976754
rect 650208 976696 655185 976698
rect 655119 976693 655185 976696
rect 59439 975424 59505 975427
rect 59439 975422 64416 975424
rect 59439 975366 59444 975422
rect 59500 975366 64416 975422
rect 59439 975364 64416 975366
rect 59439 975361 59505 975364
rect 42159 968764 42225 968767
rect 42298 968764 42304 968766
rect 42159 968762 42304 968764
rect 42159 968706 42164 968762
rect 42220 968706 42304 968762
rect 42159 968704 42304 968706
rect 42159 968701 42225 968704
rect 42298 968702 42304 968704
rect 42368 968702 42374 968766
rect 41775 967138 41841 967139
rect 41722 967136 41728 967138
rect 41684 967076 41728 967136
rect 41792 967134 41841 967138
rect 41836 967078 41841 967134
rect 41722 967074 41728 967076
rect 41792 967074 41841 967078
rect 41775 967073 41841 967074
rect 674511 966544 674577 966547
rect 675279 966544 675345 966547
rect 674511 966542 675345 966544
rect 674511 966486 674516 966542
rect 674572 966486 675284 966542
rect 675340 966486 675345 966542
rect 674511 966484 675345 966486
rect 674511 966481 674577 966484
rect 675279 966481 675345 966484
rect 675759 965804 675825 965807
rect 676666 965804 676672 965806
rect 675759 965802 676672 965804
rect 675759 965746 675764 965802
rect 675820 965746 676672 965802
rect 675759 965744 676672 965746
rect 675759 965741 675825 965744
rect 676666 965742 676672 965744
rect 676736 965742 676742 965806
rect 40762 965002 40768 965066
rect 40832 965064 40838 965066
rect 41775 965064 41841 965067
rect 655215 965064 655281 965067
rect 40832 965062 41841 965064
rect 40832 965006 41780 965062
rect 41836 965006 41841 965062
rect 40832 965004 41841 965006
rect 650208 965062 655281 965064
rect 650208 965006 655220 965062
rect 655276 965006 655281 965062
rect 650208 965004 655281 965006
rect 40832 965002 40838 965004
rect 41775 965001 41841 965004
rect 655215 965001 655281 965004
rect 674554 965002 674560 965066
rect 674624 965064 674630 965066
rect 675375 965064 675441 965067
rect 674624 965062 675441 965064
rect 674624 965006 675380 965062
rect 675436 965006 675441 965062
rect 674624 965004 675441 965006
rect 674624 965002 674630 965004
rect 675375 965001 675441 965004
rect 42159 964028 42225 964031
rect 42490 964028 42496 964030
rect 42159 964026 42496 964028
rect 42159 963970 42164 964026
rect 42220 963970 42496 964026
rect 42159 963968 42496 963970
rect 42159 963965 42225 963968
rect 42490 963966 42496 963968
rect 42560 963966 42566 964030
rect 40954 963374 40960 963438
rect 41024 963436 41030 963438
rect 41775 963436 41841 963439
rect 41024 963434 41841 963436
rect 41024 963378 41780 963434
rect 41836 963378 41841 963434
rect 41024 963376 41841 963378
rect 41024 963374 41030 963376
rect 41775 963373 41841 963376
rect 675759 963436 675825 963439
rect 675898 963436 675904 963438
rect 675759 963434 675904 963436
rect 675759 963378 675764 963434
rect 675820 963378 675904 963434
rect 675759 963376 675904 963378
rect 675759 963373 675825 963376
rect 675898 963374 675904 963376
rect 675968 963374 675974 963438
rect 41146 962634 41152 962698
rect 41216 962696 41222 962698
rect 41775 962696 41841 962699
rect 41216 962694 41841 962696
rect 41216 962638 41780 962694
rect 41836 962638 41841 962694
rect 41216 962636 41841 962638
rect 41216 962634 41222 962636
rect 41775 962633 41841 962636
rect 675663 962550 675729 962551
rect 675663 962546 675712 962550
rect 675776 962548 675782 962550
rect 675663 962490 675668 962546
rect 675663 962486 675712 962490
rect 675776 962488 675820 962548
rect 675776 962486 675782 962488
rect 675663 962485 675729 962486
rect 42159 962400 42225 962403
rect 43066 962400 43072 962402
rect 42159 962398 43072 962400
rect 42159 962342 42164 962398
rect 42220 962342 43072 962398
rect 42159 962340 43072 962342
rect 42159 962337 42225 962340
rect 43066 962338 43072 962340
rect 43136 962400 43142 962402
rect 62031 962400 62097 962403
rect 43136 962398 62097 962400
rect 43136 962342 62036 962398
rect 62092 962342 62097 962398
rect 43136 962340 62097 962342
rect 43136 962338 43142 962340
rect 62031 962337 62097 962340
rect 40378 962190 40384 962254
rect 40448 962252 40454 962254
rect 41871 962252 41937 962255
rect 40448 962250 41937 962252
rect 40448 962194 41876 962250
rect 41932 962194 41937 962250
rect 40448 962192 41937 962194
rect 40448 962190 40454 962192
rect 41871 962189 41937 962192
rect 673978 962190 673984 962254
rect 674048 962252 674054 962254
rect 675375 962252 675441 962255
rect 674048 962250 675441 962252
rect 674048 962194 675380 962250
rect 675436 962194 675441 962250
rect 674048 962192 675441 962194
rect 674048 962190 674054 962192
rect 675375 962189 675441 962192
rect 42447 962104 42513 962107
rect 42874 962104 42880 962106
rect 42447 962102 42880 962104
rect 42447 962046 42452 962102
rect 42508 962046 42880 962102
rect 42447 962044 42880 962046
rect 42447 962041 42513 962044
rect 42874 962042 42880 962044
rect 42944 962104 42950 962106
rect 61839 962104 61905 962107
rect 42944 962102 61905 962104
rect 42944 962046 61844 962102
rect 61900 962046 61905 962102
rect 42944 962044 61905 962046
rect 42944 962042 42950 962044
rect 61839 962041 61905 962044
rect 675759 961512 675825 961515
rect 676090 961512 676096 961514
rect 675759 961510 676096 961512
rect 675759 961454 675764 961510
rect 675820 961454 676096 961510
rect 675759 961452 676096 961454
rect 675759 961449 675825 961452
rect 676090 961450 676096 961452
rect 676160 961450 676166 961514
rect 59535 960920 59601 960923
rect 59535 960918 64416 960920
rect 59535 960862 59540 960918
rect 59596 960862 64416 960918
rect 59535 960860 64416 960862
rect 59535 960857 59601 960860
rect 675322 960710 675328 960774
rect 675392 960772 675398 960774
rect 675471 960772 675537 960775
rect 675392 960770 675537 960772
rect 675392 960714 675476 960770
rect 675532 960714 675537 960770
rect 675392 960712 675537 960714
rect 675392 960710 675398 960712
rect 675471 960709 675537 960712
rect 41530 959674 41536 959738
rect 41600 959736 41606 959738
rect 41775 959736 41841 959739
rect 41600 959734 41841 959736
rect 41600 959678 41780 959734
rect 41836 959678 41841 959734
rect 41600 959676 41841 959678
rect 41600 959674 41606 959676
rect 41775 959673 41841 959676
rect 674127 959292 674193 959295
rect 674362 959292 674368 959294
rect 674127 959290 674368 959292
rect 674127 959234 674132 959290
rect 674188 959234 674368 959290
rect 674127 959232 674368 959234
rect 674127 959229 674193 959232
rect 674362 959230 674368 959232
rect 674432 959292 674438 959294
rect 675087 959292 675153 959295
rect 674432 959290 675153 959292
rect 674432 959234 675092 959290
rect 675148 959234 675153 959290
rect 674432 959232 675153 959234
rect 674432 959230 674438 959232
rect 675087 959229 675153 959232
rect 41871 959146 41937 959147
rect 41871 959142 41920 959146
rect 41984 959144 41990 959146
rect 41871 959086 41876 959142
rect 41871 959082 41920 959086
rect 41984 959084 42028 959144
rect 41984 959082 41990 959084
rect 674746 959082 674752 959146
rect 674816 959144 674822 959146
rect 675471 959144 675537 959147
rect 674816 959142 675537 959144
rect 674816 959086 675476 959142
rect 675532 959086 675537 959142
rect 674816 959084 675537 959086
rect 674816 959082 674822 959084
rect 41871 959081 41937 959082
rect 675471 959081 675537 959084
rect 40570 958490 40576 958554
rect 40640 958552 40646 958554
rect 41775 958552 41841 958555
rect 40640 958550 41841 958552
rect 40640 958494 41780 958550
rect 41836 958494 41841 958550
rect 40640 958492 41841 958494
rect 40640 958490 40646 958492
rect 41775 958489 41841 958492
rect 675759 958404 675825 958407
rect 676474 958404 676480 958406
rect 675759 958402 676480 958404
rect 675759 958346 675764 958402
rect 675820 958346 676480 958402
rect 675759 958344 676480 958346
rect 675759 958341 675825 958344
rect 676474 958342 676480 958344
rect 676544 958342 676550 958406
rect 42159 957812 42225 957815
rect 42682 957812 42688 957814
rect 42159 957810 42688 957812
rect 42159 957754 42164 957810
rect 42220 957754 42688 957810
rect 42159 957752 42688 957754
rect 42159 957749 42225 957752
rect 42682 957750 42688 957752
rect 42752 957750 42758 957814
rect 675130 957602 675136 957666
rect 675200 957664 675206 957666
rect 675375 957664 675441 957667
rect 675200 957662 675441 957664
rect 675200 957606 675380 957662
rect 675436 957606 675441 957662
rect 675200 957604 675441 957606
rect 675200 957602 675206 957604
rect 675375 957601 675441 957604
rect 42063 956186 42129 956187
rect 42063 956182 42112 956186
rect 42176 956184 42182 956186
rect 42063 956126 42068 956182
rect 42063 956122 42112 956126
rect 42176 956124 42220 956184
rect 42176 956122 42182 956124
rect 42063 956121 42129 956122
rect 674938 955974 674944 956038
rect 675008 956036 675014 956038
rect 675471 956036 675537 956039
rect 675008 956034 675537 956036
rect 675008 955978 675476 956034
rect 675532 955978 675537 956034
rect 675008 955976 675537 955978
rect 675008 955974 675014 955976
rect 675471 955973 675537 955976
rect 674895 953520 674961 953523
rect 677050 953520 677056 953522
rect 674895 953518 677056 953520
rect 674895 953462 674900 953518
rect 674956 953462 677056 953518
rect 674895 953460 677056 953462
rect 674895 953457 674961 953460
rect 677050 953458 677056 953460
rect 677120 953458 677126 953522
rect 655311 953372 655377 953375
rect 650208 953370 655377 953372
rect 650208 953314 655316 953370
rect 655372 953314 655377 953370
rect 650208 953312 655377 953314
rect 655311 953309 655377 953312
rect 675183 953372 675249 953375
rect 676858 953372 676864 953374
rect 675183 953370 676864 953372
rect 675183 953314 675188 953370
rect 675244 953314 676864 953370
rect 675183 953312 676864 953314
rect 675183 953309 675249 953312
rect 676858 953310 676864 953312
rect 676928 953310 676934 953374
rect 59535 946712 59601 946715
rect 59535 946710 64416 946712
rect 59535 946654 59540 946710
rect 59596 946654 64416 946710
rect 59535 946652 64416 946654
rect 59535 946649 59601 946652
rect 42498 944643 42558 944906
rect 42498 944638 42609 944643
rect 42498 944582 42548 944638
rect 42604 944582 42609 944638
rect 42498 944580 42609 944582
rect 42543 944577 42609 944580
rect 42498 944199 42558 944314
rect 42498 944194 42609 944199
rect 42498 944138 42548 944194
rect 42604 944138 42609 944194
rect 42498 944136 42609 944138
rect 42543 944133 42609 944136
rect 42543 944048 42609 944051
rect 42498 944046 42609 944048
rect 42498 943990 42548 944046
rect 42604 943990 42609 944046
rect 42498 943985 42609 943990
rect 42498 943796 42558 943985
rect 40386 943015 40446 943278
rect 40386 943010 40497 943015
rect 42543 943012 42609 943015
rect 40386 942954 40436 943010
rect 40492 942954 40497 943010
rect 40386 942952 40497 942954
rect 40431 942949 40497 942952
rect 42498 943010 42609 943012
rect 42498 942954 42548 943010
rect 42604 942954 42609 943010
rect 42498 942949 42609 942954
rect 42498 942686 42558 942949
rect 42543 942420 42609 942423
rect 42498 942418 42609 942420
rect 42498 942362 42548 942418
rect 42604 942362 42609 942418
rect 42498 942357 42609 942362
rect 42498 942168 42558 942357
rect 40047 941976 40113 941979
rect 41775 941976 41841 941979
rect 40047 941974 41841 941976
rect 40047 941918 40052 941974
rect 40108 941918 41780 941974
rect 41836 941918 41841 941974
rect 40047 941916 41841 941918
rect 40047 941913 40113 941916
rect 41775 941913 41841 941916
rect 39951 941828 40017 941831
rect 40378 941828 40384 941830
rect 39951 941826 40384 941828
rect 39951 941770 39956 941826
rect 40012 941770 40384 941826
rect 39951 941768 40384 941770
rect 39951 941765 40017 941768
rect 40378 941766 40384 941768
rect 40448 941766 40454 941830
rect 47439 941680 47505 941683
rect 40416 941678 47505 941680
rect 40416 941650 47444 941678
rect 40386 941622 47444 941650
rect 47500 941622 47505 941678
rect 40386 941620 47505 941622
rect 40386 941386 40446 941620
rect 47439 941617 47505 941620
rect 653775 941532 653841 941535
rect 650208 941530 653841 941532
rect 650208 941474 653780 941530
rect 653836 941474 653841 941530
rect 650208 941472 653841 941474
rect 653775 941469 653841 941472
rect 40378 941322 40384 941386
rect 40448 941322 40454 941386
rect 42106 941322 42112 941386
rect 42176 941322 42182 941386
rect 42114 941058 42174 941322
rect 676866 940943 676926 941280
rect 41722 940878 41728 940942
rect 41792 940878 41798 940942
rect 676815 940938 676926 940943
rect 676815 940882 676820 940938
rect 676876 940882 676926 940938
rect 676815 940880 676926 940882
rect 41730 940540 41790 940878
rect 676815 940877 676881 940880
rect 676866 940499 676926 940762
rect 676866 940494 676977 940499
rect 676866 940438 676916 940494
rect 676972 940438 676977 940494
rect 676866 940436 676977 940438
rect 676911 940433 676977 940436
rect 40047 940348 40113 940351
rect 40002 940346 40113 940348
rect 40002 940290 40052 940346
rect 40108 940290 40113 940346
rect 40002 940285 40113 940290
rect 40002 940022 40062 940285
rect 674511 939904 674577 939907
rect 674754 939904 674814 940170
rect 674511 939902 674814 939904
rect 674511 939846 674516 939902
rect 674572 939846 674814 939902
rect 674511 939844 674814 939846
rect 674511 939841 674577 939844
rect 674415 939608 674481 939611
rect 674415 939606 674784 939608
rect 674415 939550 674420 939606
rect 674476 939550 674784 939606
rect 674415 939548 674784 939550
rect 674415 939545 674481 939548
rect 42682 939460 42688 939462
rect 42528 939400 42688 939460
rect 42682 939398 42688 939400
rect 42752 939398 42758 939462
rect 39951 939164 40017 939167
rect 673839 939164 673905 939167
rect 39951 939162 40062 939164
rect 39951 939106 39956 939162
rect 40012 939106 40062 939162
rect 39951 939101 40062 939106
rect 673839 939162 674784 939164
rect 673839 939106 673844 939162
rect 673900 939106 674784 939162
rect 673839 939104 674784 939106
rect 673839 939101 673905 939104
rect 40002 938912 40062 939101
rect 42298 938658 42304 938722
rect 42368 938658 42374 938722
rect 42306 938394 42366 938658
rect 676866 938279 676926 938542
rect 676815 938274 676926 938279
rect 676815 938218 676820 938274
rect 676876 938218 676926 938274
rect 676815 938216 676926 938218
rect 676815 938213 676881 938216
rect 674415 937980 674481 937983
rect 674415 937978 674784 937980
rect 674415 937922 674420 937978
rect 674476 937922 674784 937978
rect 674415 937920 674784 937922
rect 674415 937917 674481 937920
rect 42831 937832 42897 937835
rect 42528 937830 42897 937832
rect 42528 937774 42836 937830
rect 42892 937774 42897 937830
rect 42528 937772 42897 937774
rect 42831 937769 42897 937772
rect 40570 937622 40576 937686
rect 40640 937622 40646 937686
rect 674554 937622 674560 937686
rect 674624 937684 674630 937686
rect 674624 937624 674814 937684
rect 674624 937622 674630 937624
rect 40578 937284 40638 937622
rect 674754 937506 674814 937624
rect 676911 937240 676977 937243
rect 676866 937238 676977 937240
rect 676866 937182 676916 937238
rect 676972 937182 676977 937238
rect 676866 937177 676977 937182
rect 41914 937030 41920 937094
rect 41984 937030 41990 937094
rect 41922 936766 41982 937030
rect 676866 936914 676926 937177
rect 677050 936586 677056 936650
rect 677120 936586 677126 936650
rect 40762 936438 40768 936502
rect 40832 936438 40838 936502
rect 40770 936174 40830 936438
rect 677058 936322 677118 936586
rect 675898 936142 675904 936206
rect 675968 936142 675974 936206
rect 40954 935846 40960 935910
rect 41024 935846 41030 935910
rect 675906 935878 675966 936142
rect 40962 935656 41022 935846
rect 674746 935550 674752 935614
rect 674816 935550 674822 935614
rect 41530 935402 41536 935466
rect 41600 935402 41606 935466
rect 41538 935138 41598 935402
rect 674754 935286 674814 935550
rect 41146 934810 41152 934874
rect 41216 934810 41222 934874
rect 41154 934546 41214 934810
rect 674031 934724 674097 934727
rect 674031 934722 674784 934724
rect 674031 934666 674036 934722
rect 674092 934666 674784 934722
rect 674031 934664 674784 934666
rect 674031 934661 674097 934664
rect 42490 934366 42496 934430
rect 42560 934366 42566 934430
rect 676666 934366 676672 934430
rect 676736 934366 676742 934430
rect 42498 933954 42558 934366
rect 676674 934250 676734 934366
rect 675706 933774 675712 933838
rect 675776 933774 675782 933838
rect 675714 933658 675774 933774
rect 42498 933247 42558 933510
rect 673978 933330 673984 933394
rect 674048 933392 674054 933394
rect 674048 933332 674814 933392
rect 674048 933330 674054 933332
rect 42498 933242 42609 933247
rect 42498 933186 42548 933242
rect 42604 933186 42609 933242
rect 42498 933184 42609 933186
rect 42543 933181 42609 933184
rect 674754 933066 674814 933332
rect 35202 932655 35262 932918
rect 674938 932738 674944 932802
rect 675008 932738 675014 932802
rect 35202 932650 35313 932655
rect 35202 932594 35252 932650
rect 35308 932594 35313 932650
rect 674946 932622 675006 932738
rect 35202 932592 35313 932594
rect 35247 932589 35313 932592
rect 42498 932211 42558 932326
rect 35247 932208 35313 932211
rect 35202 932206 35313 932208
rect 35202 932150 35252 932206
rect 35308 932150 35313 932206
rect 35202 932145 35313 932150
rect 42498 932206 42609 932211
rect 42498 932150 42548 932206
rect 42604 932150 42609 932206
rect 42498 932148 42609 932150
rect 42543 932145 42609 932148
rect 59535 932208 59601 932211
rect 59535 932206 64416 932208
rect 59535 932150 59540 932206
rect 59596 932150 64416 932206
rect 59535 932148 64416 932150
rect 59535 932145 59601 932148
rect 675130 932146 675136 932210
rect 675200 932146 675206 932210
rect 35202 931882 35262 932145
rect 675138 932030 675198 932146
rect 676090 931702 676096 931766
rect 676160 931702 676166 931766
rect 676098 931438 676158 931702
rect 676474 931110 676480 931174
rect 676544 931110 676550 931174
rect 676482 930920 676542 931110
rect 676858 930666 676864 930730
rect 676928 930666 676934 930730
rect 676866 930402 676926 930666
rect 654447 929840 654513 929843
rect 650208 929838 654513 929840
rect 650208 929782 654452 929838
rect 654508 929782 654513 929838
rect 650208 929780 654513 929782
rect 654447 929777 654513 929780
rect 677058 929547 677118 929810
rect 677007 929542 677118 929547
rect 677007 929486 677012 929542
rect 677068 929486 677118 929542
rect 677007 929484 677118 929486
rect 677007 929481 677073 929484
rect 676866 928955 676926 929292
rect 676815 928950 676926 928955
rect 676815 928894 676820 928950
rect 676876 928894 676926 928950
rect 676815 928892 676926 928894
rect 676815 928889 676881 928892
rect 677058 928511 677118 928774
rect 676815 928508 676881 928511
rect 676815 928506 676926 928508
rect 676815 928450 676820 928506
rect 676876 928450 676926 928506
rect 676815 928445 676926 928450
rect 677007 928506 677118 928511
rect 677007 928450 677012 928506
rect 677068 928450 677118 928506
rect 677007 928448 677118 928450
rect 677007 928445 677073 928448
rect 676866 928182 676926 928445
rect 653967 918148 654033 918151
rect 650208 918146 654033 918148
rect 650208 918090 653972 918146
rect 654028 918090 654033 918146
rect 650208 918088 654033 918090
rect 653967 918085 654033 918088
rect 59535 917852 59601 917855
rect 59535 917850 64416 917852
rect 59535 917794 59540 917850
rect 59596 917794 64416 917850
rect 59535 917792 64416 917794
rect 59535 917789 59601 917792
rect 654447 906456 654513 906459
rect 650208 906454 654513 906456
rect 650208 906398 654452 906454
rect 654508 906398 654513 906454
rect 650208 906396 654513 906398
rect 654447 906393 654513 906396
rect 59535 903496 59601 903499
rect 59535 903494 64416 903496
rect 59535 903438 59540 903494
rect 59596 903438 64416 903494
rect 59535 903436 64416 903438
rect 59535 903433 59601 903436
rect 653775 894616 653841 894619
rect 650208 894614 653841 894616
rect 650208 894558 653780 894614
rect 653836 894558 653841 894614
rect 650208 894556 653841 894558
rect 653775 894553 653841 894556
rect 59535 889140 59601 889143
rect 59535 889138 64416 889140
rect 59535 889082 59540 889138
rect 59596 889082 64416 889138
rect 59535 889080 64416 889082
rect 59535 889077 59601 889080
rect 653967 882924 654033 882927
rect 650208 882922 654033 882924
rect 650208 882866 653972 882922
rect 654028 882866 654033 882922
rect 650208 882864 654033 882866
rect 653967 882861 654033 882864
rect 674170 876942 674176 877006
rect 674240 877004 674246 877006
rect 675375 877004 675441 877007
rect 674240 877002 675441 877004
rect 674240 876946 675380 877002
rect 675436 876946 675441 877002
rect 674240 876944 675441 876946
rect 674240 876942 674246 876944
rect 675375 876941 675441 876944
rect 675759 876560 675825 876563
rect 676090 876560 676096 876562
rect 675759 876558 676096 876560
rect 675759 876502 675764 876558
rect 675820 876502 676096 876558
rect 675759 876500 676096 876502
rect 675759 876497 675825 876500
rect 676090 876498 676096 876500
rect 676160 876498 676166 876562
rect 675087 875820 675153 875823
rect 675471 875822 675537 875823
rect 675322 875820 675328 875822
rect 675087 875818 675328 875820
rect 675087 875762 675092 875818
rect 675148 875762 675328 875818
rect 675087 875760 675328 875762
rect 675087 875757 675153 875760
rect 675322 875758 675328 875760
rect 675392 875758 675398 875822
rect 675471 875818 675520 875822
rect 675584 875820 675590 875822
rect 675471 875762 675476 875818
rect 675471 875758 675520 875762
rect 675584 875760 675628 875820
rect 675584 875758 675590 875760
rect 675471 875757 675537 875758
rect 674362 875610 674368 875674
rect 674432 875672 674438 875674
rect 675183 875672 675249 875675
rect 674432 875670 675249 875672
rect 674432 875614 675188 875670
rect 675244 875614 675249 875670
rect 674432 875612 675249 875614
rect 674432 875610 674438 875612
rect 675183 875609 675249 875612
rect 59535 874784 59601 874787
rect 59535 874782 64416 874784
rect 59535 874726 59540 874782
rect 59596 874726 64416 874782
rect 59535 874724 64416 874726
rect 59535 874721 59601 874724
rect 674554 873982 674560 874046
rect 674624 874044 674630 874046
rect 675471 874044 675537 874047
rect 674624 874042 675537 874044
rect 674624 873986 675476 874042
rect 675532 873986 675537 874042
rect 674624 873984 675537 873986
rect 674624 873982 674630 873984
rect 675471 873981 675537 873984
rect 674362 873538 674368 873602
rect 674432 873600 674438 873602
rect 675375 873600 675441 873603
rect 674432 873598 675441 873600
rect 674432 873542 675380 873598
rect 675436 873542 675441 873598
rect 674432 873540 675441 873542
rect 674432 873538 674438 873540
rect 675375 873537 675441 873540
rect 654447 871232 654513 871235
rect 650208 871230 654513 871232
rect 650208 871174 654452 871230
rect 654508 871174 654513 871230
rect 650208 871172 654513 871174
rect 654447 871169 654513 871172
rect 674938 869838 674944 869902
rect 675008 869900 675014 869902
rect 675375 869900 675441 869903
rect 675008 869898 675441 869900
rect 675008 869842 675380 869898
rect 675436 869842 675441 869898
rect 675008 869840 675441 869842
rect 675008 869838 675014 869840
rect 675375 869837 675441 869840
rect 675130 864658 675136 864722
rect 675200 864720 675206 864722
rect 675471 864720 675537 864723
rect 675200 864718 675537 864720
rect 675200 864662 675476 864718
rect 675532 864662 675537 864718
rect 675200 864660 675537 864662
rect 675200 864658 675206 864660
rect 675471 864657 675537 864660
rect 58575 860428 58641 860431
rect 58575 860426 64416 860428
rect 58575 860370 58580 860426
rect 58636 860370 64416 860426
rect 58575 860368 64416 860370
rect 58575 860365 58641 860368
rect 654159 859540 654225 859543
rect 650208 859538 654225 859540
rect 650208 859482 654164 859538
rect 654220 859482 654225 859538
rect 650208 859480 654225 859482
rect 654159 859477 654225 859480
rect 650127 848292 650193 848295
rect 650127 848290 650238 848292
rect 650127 848234 650132 848290
rect 650188 848234 650238 848290
rect 650127 848229 650238 848234
rect 650178 847670 650238 848229
rect 59535 846072 59601 846075
rect 59535 846070 64416 846072
rect 59535 846014 59540 846070
rect 59596 846014 64416 846070
rect 59535 846012 64416 846014
rect 59535 846009 59601 846012
rect 653967 836008 654033 836011
rect 650208 836006 654033 836008
rect 650208 835950 653972 836006
rect 654028 835950 654033 836006
rect 650208 835948 654033 835950
rect 653967 835945 654033 835948
rect 59535 831716 59601 831719
rect 59535 831714 64416 831716
rect 59535 831658 59540 831714
rect 59596 831658 64416 831714
rect 59535 831656 64416 831658
rect 59535 831653 59601 831656
rect 653967 824316 654033 824319
rect 650208 824314 654033 824316
rect 650208 824258 653972 824314
rect 654028 824258 654033 824314
rect 650208 824256 654033 824258
rect 653967 824253 654033 824256
rect 42543 819284 42609 819287
rect 42498 819282 42609 819284
rect 42498 819226 42548 819282
rect 42604 819226 42609 819282
rect 42498 819221 42609 819226
rect 42498 819106 42558 819221
rect 42831 818544 42897 818547
rect 42528 818542 42897 818544
rect 42528 818486 42836 818542
rect 42892 818486 42897 818542
rect 42528 818484 42897 818486
rect 42831 818481 42897 818484
rect 42543 818248 42609 818251
rect 42498 818246 42609 818248
rect 42498 818190 42548 818246
rect 42604 818190 42609 818246
rect 42498 818185 42609 818190
rect 42498 817922 42558 818185
rect 43215 817508 43281 817511
rect 42528 817506 43281 817508
rect 42528 817450 43220 817506
rect 43276 817450 43281 817506
rect 42528 817448 43281 817450
rect 43215 817445 43281 817448
rect 59535 817360 59601 817363
rect 59535 817358 64416 817360
rect 59535 817302 59540 817358
rect 59596 817302 64416 817358
rect 59535 817300 64416 817302
rect 59535 817297 59601 817300
rect 40431 817212 40497 817215
rect 40386 817210 40497 817212
rect 40386 817154 40436 817210
rect 40492 817154 40497 817210
rect 40386 817149 40497 817154
rect 40386 816886 40446 817149
rect 40335 816768 40401 816771
rect 40335 816766 41214 816768
rect 40335 816710 40340 816766
rect 40396 816710 41214 816766
rect 40335 816708 41214 816710
rect 40335 816705 40401 816708
rect 41154 816030 41214 816708
rect 40378 815966 40384 816030
rect 40448 815966 40454 816030
rect 41146 815966 41152 816030
rect 41216 815966 41222 816030
rect 40386 815880 40446 815966
rect 40386 815850 41376 815880
rect 40416 815820 41406 815850
rect 41346 815586 41406 815820
rect 41338 815522 41344 815586
rect 41408 815522 41414 815586
rect 41730 814995 41790 815258
rect 41679 814990 41790 814995
rect 41679 814934 41684 814990
rect 41740 814934 41790 814990
rect 41679 814932 41790 814934
rect 41679 814929 41745 814932
rect 42498 814403 42558 814666
rect 42498 814398 42609 814403
rect 42498 814342 42548 814398
rect 42604 814342 42609 814398
rect 42498 814340 42609 814342
rect 42543 814337 42609 814340
rect 40194 813959 40254 814222
rect 40194 813954 40305 813959
rect 40194 813898 40244 813954
rect 40300 813898 40305 813954
rect 40194 813896 40305 813898
rect 40239 813893 40305 813896
rect 41922 813367 41982 813630
rect 41922 813362 42033 813367
rect 41922 813306 41972 813362
rect 42028 813306 42033 813362
rect 41922 813304 42033 813306
rect 41967 813301 42033 813304
rect 42114 812775 42174 813038
rect 42063 812770 42174 812775
rect 42063 812714 42068 812770
rect 42124 812714 42174 812770
rect 42063 812712 42174 812714
rect 42063 812709 42129 812712
rect 654447 812624 654513 812627
rect 650208 812622 654513 812624
rect 41922 812331 41982 812594
rect 650208 812566 654452 812622
rect 654508 812566 654513 812622
rect 650208 812564 654513 812566
rect 654447 812561 654513 812564
rect 41871 812326 41982 812331
rect 41871 812270 41876 812326
rect 41932 812270 41982 812326
rect 41871 812268 41982 812270
rect 41871 812265 41937 812268
rect 40194 811739 40254 812002
rect 40143 811734 40254 811739
rect 40143 811678 40148 811734
rect 40204 811678 40254 811734
rect 40143 811676 40254 811678
rect 40143 811673 40209 811676
rect 43119 811440 43185 811443
rect 42528 811438 43185 811440
rect 42528 811382 43124 811438
rect 43180 811382 43185 811438
rect 42528 811380 43185 811382
rect 43119 811377 43185 811380
rect 41538 810555 41598 810966
rect 41487 810550 41598 810555
rect 41487 810494 41492 810550
rect 41548 810494 41598 810550
rect 41487 810492 41598 810494
rect 41487 810489 41553 810492
rect 42927 810404 42993 810407
rect 42528 810402 42993 810404
rect 42528 810346 42932 810402
rect 42988 810346 42993 810402
rect 42528 810344 42993 810346
rect 42927 810341 42993 810344
rect 42114 809519 42174 809782
rect 42114 809514 42225 809519
rect 42114 809458 42164 809514
rect 42220 809458 42225 809514
rect 42114 809456 42225 809458
rect 42159 809453 42225 809456
rect 41538 808927 41598 809264
rect 41538 808922 41649 808927
rect 41538 808866 41588 808922
rect 41644 808866 41649 808922
rect 41538 808864 41649 808866
rect 41583 808861 41649 808864
rect 41730 808483 41790 808746
rect 41730 808478 41841 808483
rect 41730 808422 41780 808478
rect 41836 808422 41841 808478
rect 41730 808420 41841 808422
rect 41775 808417 41841 808420
rect 43023 808184 43089 808187
rect 42528 808182 43089 808184
rect 42528 808126 43028 808182
rect 43084 808126 43089 808182
rect 42528 808124 43089 808126
rect 43023 808121 43089 808124
rect 42498 807296 42558 807636
rect 42498 807236 42750 807296
rect 35202 806855 35262 807118
rect 35151 806850 35262 806855
rect 42690 806852 42750 807236
rect 35151 806794 35156 806850
rect 35212 806794 35262 806850
rect 35151 806792 35262 806794
rect 42498 806792 42750 806852
rect 35151 806789 35217 806792
rect 42498 806556 42558 806792
rect 44655 806556 44721 806559
rect 42498 806554 44721 806556
rect 42498 806526 44660 806554
rect 42528 806498 44660 806526
rect 44716 806498 44721 806554
rect 42528 806496 44721 806498
rect 44655 806493 44721 806496
rect 35151 806408 35217 806411
rect 35151 806406 35262 806408
rect 35151 806350 35156 806406
rect 35212 806350 35262 806406
rect 35151 806345 35262 806350
rect 35202 806008 35262 806345
rect 59535 802856 59601 802859
rect 59535 802854 64416 802856
rect 59535 802798 59540 802854
rect 59596 802798 64416 802854
rect 59535 802796 64416 802798
rect 59535 802793 59601 802796
rect 40239 802116 40305 802119
rect 41530 802116 41536 802118
rect 40239 802114 41536 802116
rect 40239 802058 40244 802114
rect 40300 802058 41536 802114
rect 40239 802056 41536 802058
rect 40239 802053 40305 802056
rect 41530 802054 41536 802056
rect 41600 802054 41606 802118
rect 40143 801968 40209 801971
rect 40954 801968 40960 801970
rect 40143 801966 40960 801968
rect 40143 801910 40148 801966
rect 40204 801910 40960 801966
rect 40143 801908 40960 801910
rect 40143 801905 40209 801908
rect 40954 801906 40960 801908
rect 41024 801906 41030 801970
rect 650031 801376 650097 801379
rect 649986 801374 650097 801376
rect 649986 801318 650036 801374
rect 650092 801318 650097 801374
rect 649986 801313 650097 801318
rect 41487 800784 41553 800787
rect 42874 800784 42880 800786
rect 41487 800782 42880 800784
rect 41487 800726 41492 800782
rect 41548 800726 42880 800782
rect 41487 800724 42880 800726
rect 41487 800721 41553 800724
rect 42874 800722 42880 800724
rect 42944 800722 42950 800786
rect 649986 800754 650046 801313
rect 41583 800636 41649 800639
rect 41914 800636 41920 800638
rect 41583 800634 41920 800636
rect 41583 800578 41588 800634
rect 41644 800578 41920 800634
rect 41583 800576 41920 800578
rect 41583 800573 41649 800576
rect 41914 800574 41920 800576
rect 41984 800574 41990 800638
rect 41679 800488 41745 800491
rect 42490 800488 42496 800490
rect 41679 800486 42496 800488
rect 41679 800430 41684 800486
rect 41740 800430 42496 800486
rect 41679 800428 42496 800430
rect 41679 800425 41745 800428
rect 42490 800426 42496 800428
rect 42560 800426 42566 800490
rect 41775 800342 41841 800343
rect 42159 800342 42225 800343
rect 41722 800340 41728 800342
rect 41684 800280 41728 800340
rect 41792 800338 41841 800342
rect 42106 800340 42112 800342
rect 41836 800282 41841 800338
rect 41722 800278 41728 800280
rect 41792 800278 41841 800282
rect 42068 800280 42112 800340
rect 42176 800338 42225 800342
rect 42220 800282 42225 800338
rect 42106 800278 42112 800280
rect 42176 800278 42225 800282
rect 41775 800277 41841 800278
rect 42159 800277 42225 800278
rect 41914 796134 41920 796198
rect 41984 796196 41990 796198
rect 42735 796196 42801 796199
rect 41984 796194 42801 796196
rect 41984 796138 42740 796194
rect 42796 796138 42801 796194
rect 41984 796136 42801 796138
rect 41984 796134 41990 796136
rect 42735 796133 42801 796136
rect 40954 795986 40960 796050
rect 41024 796048 41030 796050
rect 41914 796048 41920 796050
rect 41024 795988 41920 796048
rect 41024 795986 41030 795988
rect 41914 795986 41920 795988
rect 41984 795986 41990 796050
rect 42063 794274 42129 794275
rect 42063 794272 42112 794274
rect 42020 794270 42112 794272
rect 42020 794214 42068 794270
rect 42020 794212 42112 794214
rect 42063 794210 42112 794212
rect 42176 794210 42182 794274
rect 42063 794209 42129 794210
rect 41775 793830 41841 793831
rect 41722 793766 41728 793830
rect 41792 793828 41841 793830
rect 41792 793826 41884 793828
rect 41836 793770 41884 793826
rect 41792 793768 41884 793770
rect 41792 793766 41841 793768
rect 41775 793765 41841 793766
rect 42106 792138 42112 792202
rect 42176 792200 42182 792202
rect 42447 792200 42513 792203
rect 42176 792198 42513 792200
rect 42176 792142 42452 792198
rect 42508 792142 42513 792198
rect 42176 792140 42513 792142
rect 42176 792138 42182 792140
rect 42447 792137 42513 792140
rect 42106 791842 42112 791906
rect 42176 791904 42182 791906
rect 42447 791904 42513 791907
rect 42831 791906 42897 791907
rect 42831 791904 42880 791906
rect 42176 791902 42513 791904
rect 42176 791846 42452 791902
rect 42508 791846 42513 791902
rect 42176 791844 42513 791846
rect 42788 791902 42880 791904
rect 42788 791846 42836 791902
rect 42788 791844 42880 791846
rect 42176 791842 42182 791844
rect 42447 791841 42513 791844
rect 42831 791842 42880 791844
rect 42944 791842 42950 791906
rect 42831 791841 42897 791842
rect 42490 791694 42496 791758
rect 42560 791756 42566 791758
rect 42927 791756 42993 791759
rect 42560 791754 42993 791756
rect 42560 791698 42932 791754
rect 42988 791698 42993 791754
rect 42560 791696 42993 791698
rect 42560 791694 42566 791696
rect 42927 791693 42993 791696
rect 42063 791166 42129 791167
rect 42063 791164 42112 791166
rect 42020 791162 42112 791164
rect 42176 791164 42182 791166
rect 43066 791164 43072 791166
rect 42020 791106 42068 791162
rect 42020 791104 42112 791106
rect 42063 791102 42112 791104
rect 42176 791104 43072 791164
rect 42176 791102 42182 791104
rect 43066 791102 43072 791104
rect 43136 791102 43142 791166
rect 42063 791101 42129 791102
rect 41775 790574 41841 790575
rect 41722 790510 41728 790574
rect 41792 790572 41841 790574
rect 42682 790572 42688 790574
rect 41792 790570 42688 790572
rect 41836 790514 42688 790570
rect 41792 790512 42688 790514
rect 41792 790510 41841 790512
rect 42682 790510 42688 790512
rect 42752 790510 42758 790574
rect 41775 790509 41841 790510
rect 41530 789326 41536 789390
rect 41600 789388 41606 789390
rect 42831 789388 42897 789391
rect 41600 789386 42897 789388
rect 41600 789330 42836 789386
rect 42892 789330 42897 789386
rect 41600 789328 42897 789330
rect 41600 789326 41606 789328
rect 42831 789325 42897 789328
rect 41914 789178 41920 789242
rect 41984 789240 41990 789242
rect 42735 789240 42801 789243
rect 41984 789238 42801 789240
rect 41984 789182 42740 789238
rect 42796 789182 42801 789238
rect 41984 789180 42801 789182
rect 41984 789178 41990 789180
rect 42735 789177 42801 789180
rect 654063 789092 654129 789095
rect 650208 789090 654129 789092
rect 650208 789034 654068 789090
rect 654124 789034 654129 789090
rect 650208 789032 654129 789034
rect 654063 789029 654129 789032
rect 59535 788648 59601 788651
rect 59535 788646 64416 788648
rect 59535 788590 59540 788646
rect 59596 788590 64416 788646
rect 59535 788588 64416 788590
rect 59535 788585 59601 788588
rect 673978 787994 673984 788058
rect 674048 788056 674054 788058
rect 675375 788056 675441 788059
rect 674048 788054 675441 788056
rect 674048 787998 675380 788054
rect 675436 787998 675441 788054
rect 674048 787996 675441 787998
rect 674048 787994 674054 787996
rect 675375 787993 675441 787996
rect 675322 787106 675328 787170
rect 675392 787168 675398 787170
rect 675471 787168 675537 787171
rect 675392 787166 675537 787168
rect 675392 787110 675476 787166
rect 675532 787110 675537 787166
rect 675392 787108 675537 787110
rect 675392 787106 675398 787108
rect 675471 787105 675537 787108
rect 675759 786724 675825 786727
rect 675898 786724 675904 786726
rect 675759 786722 675904 786724
rect 675759 786666 675764 786722
rect 675820 786666 675904 786722
rect 675759 786664 675904 786666
rect 675759 786661 675825 786664
rect 675898 786662 675904 786664
rect 675968 786662 675974 786726
rect 675759 784948 675825 784951
rect 676282 784948 676288 784950
rect 675759 784946 676288 784948
rect 675759 784890 675764 784946
rect 675820 784890 676288 784946
rect 675759 784888 676288 784890
rect 675759 784885 675825 784888
rect 676282 784886 676288 784888
rect 676352 784886 676358 784950
rect 675663 784210 675729 784211
rect 675663 784206 675712 784210
rect 675776 784208 675782 784210
rect 675663 784150 675668 784206
rect 675663 784146 675712 784150
rect 675776 784148 675820 784208
rect 675776 784146 675782 784148
rect 675663 784145 675729 784146
rect 675759 780656 675825 780659
rect 676666 780656 676672 780658
rect 675759 780654 676672 780656
rect 675759 780598 675764 780654
rect 675820 780598 676672 780654
rect 675759 780596 676672 780598
rect 675759 780593 675825 780596
rect 676666 780594 676672 780596
rect 676736 780594 676742 780658
rect 654063 777400 654129 777403
rect 650208 777398 654129 777400
rect 650208 777342 654068 777398
rect 654124 777342 654129 777398
rect 650208 777340 654129 777342
rect 654063 777337 654129 777340
rect 42735 775920 42801 775923
rect 42528 775918 42801 775920
rect 42528 775862 42740 775918
rect 42796 775862 42801 775918
rect 42528 775860 42801 775862
rect 42735 775857 42801 775860
rect 674511 775624 674577 775627
rect 677050 775624 677056 775626
rect 674511 775622 677056 775624
rect 674511 775566 674516 775622
rect 674572 775566 677056 775622
rect 674511 775564 677056 775566
rect 674511 775561 674577 775564
rect 677050 775562 677056 775564
rect 677120 775562 677126 775626
rect 674746 775414 674752 775478
rect 674816 775476 674822 775478
rect 675375 775476 675441 775479
rect 674816 775474 675441 775476
rect 674816 775418 675380 775474
rect 675436 775418 675441 775474
rect 674816 775416 675441 775418
rect 674816 775414 674822 775416
rect 675375 775413 675441 775416
rect 42735 775328 42801 775331
rect 42528 775326 42801 775328
rect 42528 775270 42740 775326
rect 42796 775270 42801 775326
rect 42528 775268 42801 775270
rect 42735 775265 42801 775268
rect 674703 775032 674769 775035
rect 676858 775032 676864 775034
rect 674703 775030 676864 775032
rect 674703 774974 674708 775030
rect 674764 774974 676864 775030
rect 674703 774972 676864 774974
rect 674703 774969 674769 774972
rect 676858 774970 676864 774972
rect 676928 774970 676934 775034
rect 42735 774810 42801 774813
rect 42528 774808 42801 774810
rect 42528 774752 42740 774808
rect 42796 774752 42801 774808
rect 42528 774750 42801 774752
rect 42735 774747 42801 774750
rect 43215 774292 43281 774295
rect 42528 774290 43281 774292
rect 42528 774234 43220 774290
rect 43276 774234 43281 774290
rect 42528 774232 43281 774234
rect 43215 774229 43281 774232
rect 59535 774144 59601 774147
rect 59535 774142 64416 774144
rect 59535 774086 59540 774142
rect 59596 774086 64416 774142
rect 59535 774084 64416 774086
rect 59535 774081 59601 774084
rect 676666 773786 676672 773850
rect 676736 773848 676742 773850
rect 676736 773788 676926 773848
rect 676736 773786 676742 773788
rect 43407 773700 43473 773703
rect 42528 773698 43473 773700
rect 42528 773642 43412 773698
rect 43468 773642 43473 773698
rect 42528 773640 43473 773642
rect 43407 773637 43473 773640
rect 675759 773700 675825 773703
rect 676666 773700 676672 773702
rect 675759 773698 676672 773700
rect 675759 773642 675764 773698
rect 675820 773642 676672 773698
rect 675759 773640 676672 773642
rect 675759 773637 675825 773640
rect 676666 773638 676672 773640
rect 676736 773638 676742 773702
rect 41146 773490 41152 773554
rect 41216 773490 41222 773554
rect 41154 773182 41214 773490
rect 676866 773256 676926 773788
rect 676674 773196 676926 773256
rect 41154 773152 41568 773182
rect 41184 773122 41598 773152
rect 41538 772962 41598 773122
rect 676674 773111 676734 773196
rect 676623 773106 676734 773111
rect 676623 773050 676628 773106
rect 676684 773050 676734 773106
rect 676623 773048 676734 773050
rect 676623 773045 676689 773048
rect 676858 773046 676864 773110
rect 676928 773108 676934 773110
rect 677818 773108 677824 773110
rect 676928 773048 677824 773108
rect 676928 773046 676934 773048
rect 677818 773046 677824 773048
rect 677888 773046 677894 773110
rect 41530 772898 41536 772962
rect 41600 772898 41606 772962
rect 674319 772960 674385 772963
rect 679162 772960 679168 772962
rect 674319 772958 679168 772960
rect 674319 772902 674324 772958
rect 674380 772902 679168 772958
rect 674319 772900 679168 772902
rect 674319 772897 674385 772900
rect 679162 772898 679168 772900
rect 679232 772898 679238 772962
rect 41338 772750 41344 772814
rect 41408 772750 41414 772814
rect 41346 772634 41406 772750
rect 674607 772664 674673 772667
rect 677242 772664 677248 772666
rect 674607 772662 677248 772664
rect 674607 772606 674612 772662
rect 674668 772606 677248 772662
rect 674607 772604 677248 772606
rect 674607 772601 674673 772604
rect 677242 772602 677248 772604
rect 677312 772602 677318 772666
rect 42927 772072 42993 772075
rect 42528 772070 42993 772072
rect 42528 772014 42932 772070
rect 42988 772014 42993 772070
rect 42528 772012 42993 772014
rect 42927 772009 42993 772012
rect 674746 771714 674752 771778
rect 674816 771776 674822 771778
rect 676474 771776 676480 771778
rect 674816 771716 676480 771776
rect 674816 771714 674822 771716
rect 676474 771714 676480 771716
rect 676544 771714 676550 771778
rect 41922 771187 41982 771524
rect 41922 771182 42033 771187
rect 41922 771126 41972 771182
rect 42028 771126 42033 771182
rect 41922 771124 42033 771126
rect 41967 771121 42033 771124
rect 40194 770743 40254 771006
rect 40194 770738 40305 770743
rect 40194 770682 40244 770738
rect 40300 770682 40305 770738
rect 40194 770680 40305 770682
rect 40239 770677 40305 770680
rect 41538 770151 41598 770414
rect 41487 770146 41598 770151
rect 41487 770090 41492 770146
rect 41548 770090 41598 770146
rect 41487 770088 41598 770090
rect 41487 770085 41553 770088
rect 41730 769559 41790 769896
rect 41730 769554 41841 769559
rect 41730 769498 41780 769554
rect 41836 769498 41841 769554
rect 41730 769496 41841 769498
rect 41775 769493 41841 769496
rect 41922 769115 41982 769378
rect 41871 769110 41982 769115
rect 41871 769054 41876 769110
rect 41932 769054 41982 769110
rect 41871 769052 41982 769054
rect 41871 769049 41937 769052
rect 40962 768670 41022 768786
rect 40954 768606 40960 768670
rect 41024 768606 41030 768670
rect 42498 767930 42558 768194
rect 42490 767866 42496 767930
rect 42560 767866 42566 767930
rect 41538 767487 41598 767750
rect 41538 767482 41649 767487
rect 41538 767426 41588 767482
rect 41644 767426 41649 767482
rect 41538 767424 41649 767426
rect 41583 767421 41649 767424
rect 43119 767188 43185 767191
rect 42528 767186 43185 767188
rect 42528 767130 43124 767186
rect 43180 767130 43185 767186
rect 42528 767128 43185 767130
rect 43119 767125 43185 767128
rect 42114 766303 42174 766566
rect 41679 766300 41745 766303
rect 41679 766298 41790 766300
rect 41679 766242 41684 766298
rect 41740 766242 41790 766298
rect 41679 766237 41790 766242
rect 42063 766298 42174 766303
rect 42063 766242 42068 766298
rect 42124 766242 42174 766298
rect 42063 766240 42174 766242
rect 42063 766237 42129 766240
rect 41730 766122 41790 766237
rect 43023 765560 43089 765563
rect 653967 765560 654033 765563
rect 42528 765558 43089 765560
rect 42528 765502 43028 765558
rect 43084 765502 43089 765558
rect 42528 765500 43089 765502
rect 650208 765558 654033 765560
rect 650208 765502 653972 765558
rect 654028 765502 654033 765558
rect 650208 765500 654033 765502
rect 43023 765497 43089 765500
rect 653967 765497 654033 765500
rect 42498 764672 42558 764938
rect 677775 764674 677841 764675
rect 42682 764672 42688 764674
rect 42498 764612 42688 764672
rect 42682 764610 42688 764612
rect 42752 764610 42758 764674
rect 677775 764670 677824 764674
rect 677888 764672 677894 764674
rect 677775 764614 677780 764670
rect 677775 764610 677824 764614
rect 677888 764612 677932 764672
rect 677888 764610 677894 764612
rect 677775 764609 677841 764610
rect 42498 764080 42558 764494
rect 677242 764462 677248 764526
rect 677312 764524 677318 764526
rect 677818 764524 677824 764526
rect 677312 764464 677824 764524
rect 677312 764462 677318 764464
rect 677818 764462 677824 764464
rect 677888 764462 677894 764526
rect 42498 764020 42750 764080
rect 35202 763639 35262 763902
rect 35151 763634 35262 763639
rect 42690 763636 42750 764020
rect 35151 763578 35156 763634
rect 35212 763578 35262 763634
rect 35151 763576 35262 763578
rect 42306 763576 42750 763636
rect 35151 763573 35217 763576
rect 42306 763340 42366 763576
rect 53295 763340 53361 763343
rect 42306 763310 42528 763340
rect 42690 763338 53361 763340
rect 42336 763280 42558 763310
rect 35151 763192 35217 763195
rect 42498 763192 42558 763280
rect 42690 763282 53300 763338
rect 53356 763282 53361 763338
rect 42690 763280 53361 763282
rect 42690 763192 42750 763280
rect 53295 763277 53361 763280
rect 35151 763190 35262 763192
rect 35151 763134 35156 763190
rect 35212 763134 35262 763190
rect 35151 763129 35262 763134
rect 42498 763132 42750 763192
rect 35202 762866 35262 763129
rect 674415 762896 674481 762899
rect 674415 762894 674784 762896
rect 674415 762838 674420 762894
rect 674476 762838 674784 762894
rect 674415 762836 674784 762838
rect 674415 762833 674481 762836
rect 674415 762304 674481 762307
rect 674415 762302 674784 762304
rect 674415 762246 674420 762302
rect 674476 762246 674784 762302
rect 674415 762244 674784 762246
rect 674415 762241 674481 762244
rect 674607 762008 674673 762011
rect 674607 762006 674814 762008
rect 674607 761950 674612 762006
rect 674668 761950 674814 762006
rect 674607 761948 674814 761950
rect 674607 761945 674673 761948
rect 674754 761830 674814 761948
rect 673839 761268 673905 761271
rect 673839 761266 674784 761268
rect 673839 761210 673844 761266
rect 673900 761210 674784 761266
rect 673839 761208 674784 761210
rect 673839 761205 673905 761208
rect 673839 760676 673905 760679
rect 673839 760674 674784 760676
rect 673839 760618 673844 760674
rect 673900 760618 674784 760674
rect 673839 760616 674784 760618
rect 673839 760613 673905 760616
rect 59535 759788 59601 759791
rect 677058 759790 677118 760202
rect 59535 759786 64416 759788
rect 59535 759730 59540 759786
rect 59596 759730 64416 759786
rect 59535 759728 64416 759730
rect 59535 759725 59601 759728
rect 677050 759726 677056 759790
rect 677120 759726 677126 759790
rect 676866 759346 676926 759610
rect 675514 759282 675520 759346
rect 675584 759282 675590 759346
rect 676858 759282 676864 759346
rect 676928 759282 676934 759346
rect 675522 759018 675582 759282
rect 675130 758838 675136 758902
rect 675200 758838 675206 758902
rect 675138 758574 675198 758838
rect 675130 758246 675136 758310
rect 675200 758308 675206 758310
rect 676623 758308 676689 758311
rect 675200 758306 676689 758308
rect 675200 758250 676628 758306
rect 676684 758250 676689 758306
rect 675200 758248 676689 758250
rect 675200 758246 675206 758248
rect 676623 758245 676689 758248
rect 674170 757950 674176 758014
rect 674240 758012 674246 758014
rect 674240 757952 674784 758012
rect 674240 757950 674246 757952
rect 40239 757716 40305 757719
rect 41146 757716 41152 757718
rect 40239 757714 41152 757716
rect 40239 757658 40244 757714
rect 40300 757658 41152 757714
rect 40239 757656 41152 757658
rect 40239 757653 40305 757656
rect 41146 757654 41152 757656
rect 41216 757654 41222 757718
rect 41487 757420 41553 757423
rect 42874 757420 42880 757422
rect 41487 757418 42880 757420
rect 41487 757362 41492 757418
rect 41548 757362 42880 757418
rect 41487 757360 42880 757362
rect 41487 757357 41553 757360
rect 42874 757358 42880 757360
rect 42944 757358 42950 757422
rect 41775 757272 41841 757275
rect 42106 757272 42112 757274
rect 41775 757270 42112 757272
rect 41775 757214 41780 757270
rect 41836 757214 42112 757270
rect 41775 757212 42112 757214
rect 41775 757209 41841 757212
rect 42106 757210 42112 757212
rect 42176 757210 42182 757274
rect 674554 757210 674560 757274
rect 674624 757272 674630 757274
rect 674754 757272 674814 757390
rect 674624 757212 674814 757272
rect 674624 757210 674630 757212
rect 41967 757126 42033 757127
rect 41914 757124 41920 757126
rect 41876 757064 41920 757124
rect 41984 757122 42033 757126
rect 42028 757066 42033 757122
rect 41914 757062 41920 757064
rect 41984 757062 42033 757066
rect 674746 757062 674752 757126
rect 674816 757062 674822 757126
rect 41967 757061 42033 757062
rect 674754 756872 674814 757062
rect 677242 756618 677248 756682
rect 677312 756618 677318 756682
rect 677250 756354 677310 756618
rect 676090 756026 676096 756090
rect 676160 756026 676166 756090
rect 676098 755762 676158 756026
rect 674362 755212 674368 755276
rect 674432 755274 674438 755276
rect 674432 755214 674784 755274
rect 674432 755212 674438 755214
rect 677818 754990 677824 755054
rect 677888 754990 677894 755054
rect 41871 754906 41937 754907
rect 41871 754904 41920 754906
rect 41828 754902 41920 754904
rect 41828 754846 41876 754902
rect 41828 754844 41920 754846
rect 41871 754842 41920 754844
rect 41984 754842 41990 754906
rect 41871 754841 41937 754842
rect 677826 754726 677886 754990
rect 649743 754460 649809 754463
rect 649743 754458 649854 754460
rect 649743 754402 649748 754458
rect 649804 754402 649854 754458
rect 649743 754397 649854 754402
rect 674746 754398 674752 754462
rect 674816 754460 674822 754462
rect 676474 754460 676480 754462
rect 674816 754400 676480 754460
rect 674816 754398 674822 754400
rect 676474 754398 676480 754400
rect 676544 754398 676550 754462
rect 677775 754460 677841 754463
rect 677775 754458 677886 754460
rect 677775 754402 677780 754458
rect 677836 754402 677886 754458
rect 677775 754397 677886 754402
rect 649794 753838 649854 754397
rect 677826 754134 677886 754397
rect 679162 753954 679168 754018
rect 679232 753954 679238 754018
rect 679170 753616 679230 753954
rect 673359 753128 673425 753131
rect 673359 753126 674784 753128
rect 673359 753070 673364 753126
rect 673420 753070 674784 753126
rect 673359 753068 674784 753070
rect 673359 753065 673425 753068
rect 673263 752536 673329 752539
rect 673263 752534 674784 752536
rect 673263 752478 673268 752534
rect 673324 752478 674784 752534
rect 673263 752476 674784 752478
rect 673263 752473 673329 752476
rect 673167 752092 673233 752095
rect 673167 752090 674814 752092
rect 673167 752034 673172 752090
rect 673228 752034 674814 752090
rect 673167 752032 674814 752034
rect 673167 752029 673233 752032
rect 674754 751988 674814 752032
rect 42927 751944 42993 751947
rect 43066 751944 43072 751946
rect 42927 751942 43072 751944
rect 42927 751886 42932 751942
rect 42988 751886 43072 751942
rect 42927 751884 43072 751886
rect 42927 751881 42993 751884
rect 43066 751882 43072 751884
rect 43136 751882 43142 751946
rect 42063 751796 42129 751799
rect 42682 751796 42688 751798
rect 42063 751794 42688 751796
rect 42063 751738 42068 751794
rect 42124 751738 42688 751794
rect 42063 751736 42688 751738
rect 42063 751733 42129 751736
rect 42682 751734 42688 751736
rect 42752 751734 42758 751798
rect 677058 751207 677118 751470
rect 677007 751202 677118 751207
rect 677007 751146 677012 751202
rect 677068 751146 677118 751202
rect 677007 751144 677118 751146
rect 677007 751141 677073 751144
rect 42927 751058 42993 751059
rect 42874 750994 42880 751058
rect 42944 751056 42993 751058
rect 42944 751054 43036 751056
rect 42988 750998 43036 751054
rect 42944 750996 43036 750998
rect 42944 750994 42993 750996
rect 42927 750993 42993 750994
rect 676866 750615 676926 750878
rect 676815 750610 676926 750615
rect 676815 750554 676820 750610
rect 676876 750554 676926 750610
rect 676815 750552 676926 750554
rect 677007 750612 677073 750615
rect 677007 750610 677118 750612
rect 677007 750554 677012 750610
rect 677068 750554 677118 750610
rect 676815 750549 676881 750552
rect 677007 750549 677118 750554
rect 677058 750360 677118 750549
rect 676815 750168 676881 750171
rect 676815 750166 676926 750168
rect 676815 750110 676820 750166
rect 676876 750110 676926 750166
rect 676815 750105 676926 750110
rect 42063 749874 42129 749875
rect 42063 749870 42112 749874
rect 42176 749872 42182 749874
rect 42063 749814 42068 749870
rect 42063 749810 42112 749814
rect 42176 749812 42220 749872
rect 676866 749842 676926 750105
rect 42176 749810 42182 749812
rect 42063 749809 42129 749810
rect 42447 749280 42513 749283
rect 43066 749280 43072 749282
rect 42447 749278 43072 749280
rect 42447 749222 42452 749278
rect 42508 749222 43072 749278
rect 42447 749220 43072 749222
rect 42447 749217 42513 749220
rect 43066 749218 43072 749220
rect 43136 749218 43142 749282
rect 41967 747802 42033 747803
rect 41914 747738 41920 747802
rect 41984 747800 42033 747802
rect 42298 747800 42304 747802
rect 41984 747798 42304 747800
rect 42028 747742 42304 747798
rect 41984 747740 42304 747742
rect 41984 747738 42033 747740
rect 42298 747738 42304 747740
rect 42368 747738 42374 747802
rect 41967 747737 42033 747738
rect 41775 747210 41841 747211
rect 41722 747146 41728 747210
rect 41792 747208 41841 747210
rect 41792 747206 41884 747208
rect 41836 747150 41884 747206
rect 41792 747148 41884 747150
rect 41792 747146 41841 747148
rect 41775 747145 41841 747146
rect 40954 746998 40960 747062
rect 41024 747060 41030 747062
rect 43119 747060 43185 747063
rect 41024 747058 43185 747060
rect 41024 747002 43124 747058
rect 43180 747002 43185 747058
rect 41024 747000 43185 747002
rect 41024 746998 41030 747000
rect 43119 746997 43185 747000
rect 41146 746850 41152 746914
rect 41216 746912 41222 746914
rect 43023 746912 43089 746915
rect 41216 746910 43089 746912
rect 41216 746854 43028 746910
rect 43084 746854 43089 746910
rect 41216 746852 43089 746854
rect 41216 746850 41222 746852
rect 43023 746849 43089 746852
rect 42063 746320 42129 746323
rect 42490 746320 42496 746322
rect 42063 746318 42496 746320
rect 42063 746262 42068 746318
rect 42124 746262 42496 746318
rect 42063 746260 42496 746262
rect 42063 746257 42129 746260
rect 42490 746258 42496 746260
rect 42560 746258 42566 746322
rect 59535 745580 59601 745583
rect 59535 745578 64416 745580
rect 59535 745522 59540 745578
rect 59596 745522 64416 745578
rect 59535 745520 64416 745522
rect 59535 745517 59601 745520
rect 674170 743150 674176 743214
rect 674240 743212 674246 743214
rect 675375 743212 675441 743215
rect 674240 743210 675441 743212
rect 674240 743154 675380 743210
rect 675436 743154 675441 743210
rect 674240 743152 675441 743154
rect 674240 743150 674246 743152
rect 675375 743149 675441 743152
rect 653967 742176 654033 742179
rect 650208 742174 654033 742176
rect 650208 742118 653972 742174
rect 654028 742118 654033 742174
rect 650208 742116 654033 742118
rect 653967 742113 654033 742116
rect 675471 742178 675537 742179
rect 675471 742174 675520 742178
rect 675584 742176 675590 742178
rect 675471 742118 675476 742174
rect 675471 742114 675520 742118
rect 675584 742116 675628 742176
rect 675584 742114 675590 742116
rect 675471 742113 675537 742114
rect 675759 741732 675825 741735
rect 676090 741732 676096 741734
rect 675759 741730 676096 741732
rect 675759 741674 675764 741730
rect 675820 741674 676096 741730
rect 675759 741672 676096 741674
rect 675759 741669 675825 741672
rect 676090 741670 676096 741672
rect 676160 741670 676166 741734
rect 676666 741670 676672 741734
rect 676736 741670 676742 741734
rect 676858 741670 676864 741734
rect 676928 741670 676934 741734
rect 675130 741522 675136 741586
rect 675200 741584 675206 741586
rect 676474 741584 676480 741586
rect 675200 741524 676480 741584
rect 675200 741522 675206 741524
rect 676474 741522 676480 741524
rect 676544 741522 676550 741586
rect 676674 741438 676734 741670
rect 676866 741438 676926 741670
rect 676666 741374 676672 741438
rect 676736 741374 676742 741438
rect 676858 741374 676864 741438
rect 676928 741374 676934 741438
rect 675130 740042 675136 740106
rect 675200 740104 675206 740106
rect 675375 740104 675441 740107
rect 675200 740102 675441 740104
rect 675200 740046 675380 740102
rect 675436 740046 675441 740102
rect 675200 740044 675441 740046
rect 675200 740042 675206 740044
rect 675375 740041 675441 740044
rect 674938 739154 674944 739218
rect 675008 739216 675014 739218
rect 675471 739216 675537 739219
rect 675008 739214 675537 739216
rect 675008 739158 675476 739214
rect 675532 739158 675537 739214
rect 675008 739156 675537 739158
rect 675008 739154 675014 739156
rect 675471 739153 675537 739156
rect 674362 738562 674368 738626
rect 674432 738624 674438 738626
rect 675375 738624 675441 738627
rect 674432 738622 675441 738624
rect 674432 738566 675380 738622
rect 675436 738566 675441 738622
rect 674432 738564 675441 738566
rect 674432 738562 674438 738564
rect 675375 738561 675441 738564
rect 41338 734270 41344 734334
rect 41408 734332 41414 734334
rect 42106 734332 42112 734334
rect 41408 734272 42112 734332
rect 41408 734270 41414 734272
rect 42106 734270 42112 734272
rect 42176 734270 42182 734334
rect 42831 732704 42897 732707
rect 42528 732702 42897 732704
rect 42528 732646 42836 732702
rect 42892 732646 42897 732702
rect 42528 732644 42897 732646
rect 42831 732641 42897 732644
rect 42831 732112 42897 732115
rect 42528 732110 42897 732112
rect 42528 732054 42836 732110
rect 42892 732054 42897 732110
rect 42528 732052 42897 732054
rect 42831 732049 42897 732052
rect 42831 731816 42897 731819
rect 42498 731814 42897 731816
rect 42498 731758 42836 731814
rect 42892 731758 42897 731814
rect 42498 731756 42897 731758
rect 42498 731638 42558 731756
rect 42831 731753 42897 731756
rect 43695 731076 43761 731079
rect 42528 731074 43761 731076
rect 42528 731018 43700 731074
rect 43756 731018 43761 731074
rect 42528 731016 43761 731018
rect 43695 731013 43761 731016
rect 59535 731076 59601 731079
rect 59535 731074 64416 731076
rect 59535 731018 59540 731074
rect 59596 731018 64416 731074
rect 59535 731016 64416 731018
rect 59535 731013 59601 731016
rect 43407 730484 43473 730487
rect 655215 730484 655281 730487
rect 42528 730482 43473 730484
rect 42528 730426 43412 730482
rect 43468 730426 43473 730482
rect 42528 730424 43473 730426
rect 650208 730482 655281 730484
rect 650208 730426 655220 730482
rect 655276 730426 655281 730482
rect 650208 730424 655281 730426
rect 43407 730421 43473 730424
rect 655215 730421 655281 730424
rect 41346 729598 41406 729936
rect 41338 729534 41344 729598
rect 41408 729534 41414 729598
rect 42114 729154 42174 729418
rect 42106 729090 42112 729154
rect 42176 729090 42182 729154
rect 41538 728711 41598 728826
rect 41487 728706 41598 728711
rect 41487 728650 41492 728706
rect 41548 728650 41598 728706
rect 41487 728648 41598 728650
rect 41487 728645 41553 728648
rect 42498 727971 42558 728308
rect 676666 728054 676672 728118
rect 676736 728116 676742 728118
rect 677818 728116 677824 728118
rect 676736 728056 677824 728116
rect 676736 728054 676742 728056
rect 677818 728054 677824 728056
rect 677888 728054 677894 728118
rect 42447 727966 42558 727971
rect 42447 727910 42452 727966
rect 42508 727910 42558 727966
rect 42447 727908 42558 727910
rect 42447 727905 42513 727908
rect 43066 727820 43072 727822
rect 42528 727760 43072 727820
rect 43066 727758 43072 727760
rect 43136 727758 43142 727822
rect 41538 726935 41598 727198
rect 41538 726930 41649 726935
rect 41538 726874 41588 726930
rect 41644 726874 41649 726930
rect 41538 726872 41649 726874
rect 41583 726869 41649 726872
rect 42498 726340 42558 726680
rect 43119 726340 43185 726343
rect 42498 726338 43185 726340
rect 42498 726282 43124 726338
rect 43180 726282 43185 726338
rect 42498 726280 43185 726282
rect 43119 726277 43185 726280
rect 41922 725899 41982 726162
rect 41871 725894 41982 725899
rect 41871 725838 41876 725894
rect 41932 725838 41982 725894
rect 41871 725836 41982 725838
rect 41871 725833 41937 725836
rect 41538 725306 41598 725570
rect 41530 725242 41536 725306
rect 41600 725242 41606 725306
rect 41730 724715 41790 725052
rect 41679 724710 41790 724715
rect 41679 724654 41684 724710
rect 41740 724654 41790 724710
rect 41679 724652 41790 724654
rect 41679 724649 41745 724652
rect 41730 724271 41790 724534
rect 41730 724266 41841 724271
rect 41730 724210 41780 724266
rect 41836 724210 41841 724266
rect 41730 724208 41841 724210
rect 41775 724205 41841 724208
rect 41922 723679 41982 723942
rect 41922 723674 42033 723679
rect 41922 723618 41972 723674
rect 42028 723618 42033 723674
rect 41922 723616 42033 723618
rect 41967 723613 42033 723616
rect 41154 723086 41214 723424
rect 41146 723022 41152 723086
rect 41216 723022 41222 723086
rect 41722 723022 41728 723086
rect 41792 723084 41798 723086
rect 42874 723084 42880 723086
rect 41792 723024 42880 723084
rect 41792 723022 41798 723024
rect 42874 723022 42880 723024
rect 42944 723022 42950 723086
rect 42114 722643 42174 722906
rect 42063 722638 42174 722643
rect 42063 722582 42068 722638
rect 42124 722582 42174 722638
rect 42063 722580 42174 722582
rect 42063 722577 42129 722580
rect 42114 722051 42174 722314
rect 42114 722046 42225 722051
rect 42114 721990 42164 722046
rect 42220 721990 42225 722046
rect 42114 721988 42225 721990
rect 42159 721985 42225 721988
rect 42447 722048 42513 722051
rect 43311 722048 43377 722051
rect 42447 722046 43377 722048
rect 42447 721990 42452 722046
rect 42508 721990 43316 722046
rect 43372 721990 43377 722046
rect 42447 721988 43377 721990
rect 42447 721985 42513 721988
rect 43311 721985 43377 721988
rect 42498 721607 42558 721796
rect 42447 721602 42558 721607
rect 42447 721546 42452 721602
rect 42508 721546 42558 721602
rect 42447 721544 42558 721546
rect 42447 721541 42513 721544
rect 42498 721012 42558 721278
rect 42498 720952 42750 721012
rect 35202 720423 35262 720686
rect 42690 720568 42750 720952
rect 35151 720418 35262 720423
rect 35151 720362 35156 720418
rect 35212 720362 35262 720418
rect 35151 720360 35262 720362
rect 42498 720508 42750 720568
rect 35151 720357 35217 720360
rect 42498 720124 42558 720508
rect 53487 720124 53553 720127
rect 42498 720122 53553 720124
rect 42498 720066 53492 720122
rect 53548 720066 53553 720122
rect 42498 720064 53553 720066
rect 53487 720061 53553 720064
rect 35151 719976 35217 719979
rect 35151 719974 35262 719976
rect 35151 719918 35156 719974
rect 35212 719918 35262 719974
rect 35151 719913 35262 719918
rect 35202 719650 35262 719913
rect 654255 718644 654321 718647
rect 650208 718642 654321 718644
rect 650208 718586 654260 718642
rect 654316 718586 654321 718642
rect 650208 718584 654321 718586
rect 654255 718581 654321 718584
rect 674607 718052 674673 718055
rect 674607 718050 674814 718052
rect 674607 717994 674612 718050
rect 674668 717994 674814 718050
rect 674607 717992 674814 717994
rect 674607 717989 674673 717992
rect 674754 717874 674814 717992
rect 674607 717608 674673 717611
rect 674607 717606 674814 717608
rect 674607 717550 674612 717606
rect 674668 717550 674814 717606
rect 674607 717548 674814 717550
rect 674607 717545 674673 717548
rect 674754 717282 674814 717548
rect 674607 717016 674673 717019
rect 674607 717014 674814 717016
rect 674607 716958 674612 717014
rect 674668 716958 674814 717014
rect 674607 716956 674814 716958
rect 674607 716953 674673 716956
rect 674754 716838 674814 716956
rect 59535 716720 59601 716723
rect 59535 716718 64416 716720
rect 59535 716662 59540 716718
rect 59596 716662 64416 716718
rect 59535 716660 64416 716662
rect 59535 716657 59601 716660
rect 673839 716276 673905 716279
rect 673839 716274 674784 716276
rect 673839 716218 673844 716274
rect 673900 716218 674784 716274
rect 673839 716216 674784 716218
rect 673839 716213 673905 716216
rect 673839 715684 673905 715687
rect 673839 715682 674784 715684
rect 673839 715626 673844 715682
rect 673900 715626 674784 715682
rect 673839 715624 674784 715626
rect 673839 715621 673905 715624
rect 677242 715474 677248 715538
rect 677312 715474 677318 715538
rect 676858 714882 676864 714946
rect 676928 714882 676934 714946
rect 676866 714618 676926 714882
rect 677103 714796 677169 714799
rect 677250 714796 677310 715474
rect 677103 714794 677310 714796
rect 677103 714738 677108 714794
rect 677164 714738 677310 714794
rect 677103 714736 677310 714738
rect 677103 714733 677169 714736
rect 675898 714290 675904 714354
rect 675968 714290 675974 714354
rect 42063 714056 42129 714059
rect 42682 714056 42688 714058
rect 42063 714054 42688 714056
rect 42063 713998 42068 714054
rect 42124 713998 42688 714054
rect 42063 713996 42688 713998
rect 42063 713993 42129 713996
rect 42682 713994 42688 713996
rect 42752 713994 42758 714058
rect 675906 714026 675966 714290
rect 41775 713910 41841 713911
rect 41722 713908 41728 713910
rect 41684 713848 41728 713908
rect 41792 713906 41841 713910
rect 41836 713850 41841 713906
rect 41722 713846 41728 713848
rect 41792 713846 41841 713850
rect 41775 713845 41841 713846
rect 42159 713908 42225 713911
rect 42298 713908 42304 713910
rect 42159 713906 42304 713908
rect 42159 713850 42164 713906
rect 42220 713850 42304 713906
rect 42159 713848 42304 713850
rect 42159 713845 42225 713848
rect 42298 713846 42304 713848
rect 42368 713846 42374 713910
rect 674746 713846 674752 713910
rect 674816 713846 674822 713910
rect 674754 713508 674814 713846
rect 42447 713318 42513 713319
rect 42447 713314 42496 713318
rect 42560 713316 42566 713318
rect 42447 713258 42452 713314
rect 42447 713254 42496 713258
rect 42560 713256 42604 713316
rect 42560 713254 42566 713256
rect 42447 713253 42513 713254
rect 673978 712958 673984 713022
rect 674048 713020 674054 713022
rect 674048 712960 674784 713020
rect 674048 712958 674054 712960
rect 676282 712662 676288 712726
rect 676352 712662 676358 712726
rect 676290 712398 676350 712662
rect 676474 712218 676480 712282
rect 676544 712218 676550 712282
rect 676482 711880 676542 712218
rect 677818 711626 677824 711690
rect 677888 711626 677894 711690
rect 43215 711392 43281 711395
rect 43695 711392 43761 711395
rect 43215 711390 43761 711392
rect 43215 711334 43220 711390
rect 43276 711334 43700 711390
rect 43756 711334 43761 711390
rect 677826 711362 677886 711626
rect 43215 711332 43761 711334
rect 43215 711329 43281 711332
rect 43695 711329 43761 711332
rect 41722 711034 41728 711098
rect 41792 711096 41798 711098
rect 43023 711096 43089 711099
rect 41792 711094 43089 711096
rect 41792 711038 43028 711094
rect 43084 711038 43089 711094
rect 41792 711036 43089 711038
rect 41792 711034 41798 711036
rect 43023 711033 43089 711036
rect 675322 711034 675328 711098
rect 675392 711034 675398 711098
rect 675330 710770 675390 711034
rect 675706 710590 675712 710654
rect 675776 710590 675782 710654
rect 675714 710252 675774 710590
rect 674607 709912 674673 709915
rect 674607 709910 674814 709912
rect 674607 709854 674612 709910
rect 674668 709854 674814 709910
rect 674607 709852 674814 709854
rect 674607 709849 674673 709852
rect 674754 709734 674814 709852
rect 674415 709172 674481 709175
rect 674415 709170 674784 709172
rect 674415 709114 674420 709170
rect 674476 709114 674784 709170
rect 674415 709112 674784 709114
rect 674415 709109 674481 709112
rect 41722 708666 41728 708730
rect 41792 708728 41798 708730
rect 42874 708728 42880 708730
rect 41792 708668 42880 708728
rect 41792 708666 41798 708668
rect 42874 708666 42880 708668
rect 42944 708666 42950 708730
rect 674415 708654 674481 708657
rect 674415 708652 674784 708654
rect 674415 708596 674420 708652
rect 674476 708596 674784 708652
rect 674415 708594 674784 708596
rect 674415 708591 674481 708594
rect 42063 708580 42129 708583
rect 42490 708580 42496 708582
rect 42063 708578 42496 708580
rect 42063 708522 42068 708578
rect 42124 708522 42496 708578
rect 42063 708520 42496 708522
rect 42063 708517 42129 708520
rect 42490 708518 42496 708520
rect 42560 708518 42566 708582
rect 673455 708136 673521 708139
rect 673455 708134 674784 708136
rect 673455 708078 673460 708134
rect 673516 708078 674784 708134
rect 673455 708076 674784 708078
rect 673455 708073 673521 708076
rect 41146 707926 41152 707990
rect 41216 707988 41222 707990
rect 41775 707988 41841 707991
rect 41216 707986 41841 707988
rect 41216 707930 41780 707986
rect 41836 707930 41841 707986
rect 41216 707928 41841 707930
rect 41216 707926 41222 707928
rect 41775 707925 41841 707928
rect 42735 707842 42801 707843
rect 42682 707778 42688 707842
rect 42752 707840 42801 707842
rect 42752 707838 42844 707840
rect 42796 707782 42844 707838
rect 42752 707780 42844 707782
rect 42752 707778 42801 707780
rect 42735 707777 42801 707778
rect 649839 707544 649905 707547
rect 649794 707542 649905 707544
rect 649794 707486 649844 707542
rect 649900 707486 649905 707542
rect 649794 707481 649905 707486
rect 673071 707544 673137 707547
rect 673071 707542 674784 707544
rect 673071 707486 673076 707542
rect 673132 707486 674784 707542
rect 673071 707484 674784 707486
rect 673071 707481 673137 707484
rect 42159 707396 42225 707399
rect 42298 707396 42304 707398
rect 42159 707394 42304 707396
rect 42159 707338 42164 707394
rect 42220 707338 42304 707394
rect 42159 707336 42304 707338
rect 42159 707333 42225 707336
rect 42298 707334 42304 707336
rect 42368 707334 42374 707398
rect 649794 706922 649854 707481
rect 674415 707026 674481 707029
rect 674415 707024 674784 707026
rect 674415 706968 674420 707024
rect 674476 706968 674784 707024
rect 674415 706966 674784 706968
rect 674415 706963 674481 706966
rect 677058 706215 677118 706478
rect 677007 706210 677118 706215
rect 677007 706154 677012 706210
rect 677068 706154 677118 706210
rect 677007 706152 677118 706154
rect 677007 706149 677073 706152
rect 676866 705623 676926 705886
rect 677103 705770 677169 705771
rect 677050 705768 677056 705770
rect 677012 705708 677056 705768
rect 677120 705766 677169 705770
rect 677164 705710 677169 705766
rect 677050 705706 677056 705708
rect 677120 705706 677169 705710
rect 677103 705705 677169 705706
rect 676815 705618 676926 705623
rect 676815 705562 676820 705618
rect 676876 705562 676926 705618
rect 676815 705560 676926 705562
rect 677007 705620 677073 705623
rect 677007 705618 677118 705620
rect 677007 705562 677012 705618
rect 677068 705562 677118 705618
rect 676815 705557 676881 705560
rect 677007 705557 677118 705562
rect 41530 705410 41536 705474
rect 41600 705472 41606 705474
rect 42447 705472 42513 705475
rect 41600 705470 42513 705472
rect 41600 705414 42452 705470
rect 42508 705414 42513 705470
rect 41600 705412 42513 705414
rect 41600 705410 41606 705412
rect 42447 705409 42513 705412
rect 677058 705368 677118 705557
rect 676815 705176 676881 705179
rect 676815 705174 676926 705176
rect 676815 705118 676820 705174
rect 676876 705118 676926 705174
rect 676815 705113 676926 705118
rect 676866 704850 676926 705113
rect 41871 704734 41937 704735
rect 41871 704732 41920 704734
rect 41828 704730 41920 704732
rect 41828 704674 41876 704730
rect 41828 704672 41920 704674
rect 41871 704670 41920 704672
rect 41984 704670 41990 704734
rect 41871 704669 41937 704670
rect 41775 704142 41841 704143
rect 41722 704078 41728 704142
rect 41792 704140 41841 704142
rect 41792 704138 41884 704140
rect 41836 704082 41884 704138
rect 41792 704080 41884 704082
rect 41792 704078 41841 704080
rect 41775 704077 41841 704078
rect 43023 703550 43089 703551
rect 43023 703548 43072 703550
rect 42980 703546 43072 703548
rect 42980 703490 43028 703546
rect 42980 703488 43072 703490
rect 43023 703486 43072 703488
rect 43136 703486 43142 703550
rect 43023 703485 43089 703486
rect 59535 702364 59601 702367
rect 59535 702362 64416 702364
rect 59535 702306 59540 702362
rect 59596 702306 64416 702362
rect 59535 702304 64416 702306
rect 59535 702301 59601 702304
rect 674746 697862 674752 697926
rect 674816 697924 674822 697926
rect 675375 697924 675441 697927
rect 674816 697922 675441 697924
rect 674816 697866 675380 697922
rect 675436 697866 675441 697922
rect 674816 697864 675441 697866
rect 674816 697862 674822 697864
rect 675375 697861 675441 697864
rect 675759 697332 675825 697335
rect 676666 697332 676672 697334
rect 675759 697330 676672 697332
rect 675759 697274 675764 697330
rect 675820 697274 676672 697330
rect 675759 697272 676672 697274
rect 675759 697269 675825 697272
rect 676666 697270 676672 697272
rect 676736 697270 676742 697334
rect 675375 696890 675441 696891
rect 675322 696888 675328 696890
rect 675284 696828 675328 696888
rect 675392 696886 675441 696890
rect 675436 696830 675441 696886
rect 675322 696826 675328 696828
rect 675392 696826 675441 696830
rect 675375 696825 675441 696826
rect 654447 695260 654513 695263
rect 650208 695258 654513 695260
rect 650208 695202 654452 695258
rect 654508 695202 654513 695258
rect 650208 695200 654513 695202
rect 654447 695197 654513 695200
rect 675759 694816 675825 694819
rect 675898 694816 675904 694818
rect 675759 694814 675904 694816
rect 675759 694758 675764 694814
rect 675820 694758 675904 694814
rect 675759 694756 675904 694758
rect 675759 694753 675825 694756
rect 675898 694754 675904 694756
rect 675968 694754 675974 694818
rect 674554 694310 674560 694374
rect 674624 694372 674630 694374
rect 675471 694372 675537 694375
rect 674624 694370 675537 694372
rect 674624 694314 675476 694370
rect 675532 694314 675537 694370
rect 674624 694312 675537 694314
rect 674624 694310 674630 694312
rect 675471 694309 675537 694312
rect 675759 693484 675825 693487
rect 676474 693484 676480 693486
rect 675759 693482 676480 693484
rect 675759 693426 675764 693482
rect 675820 693426 676480 693482
rect 675759 693424 676480 693426
rect 675759 693421 675825 693424
rect 676474 693422 676480 693424
rect 676544 693422 676550 693486
rect 675759 692004 675825 692007
rect 676282 692004 676288 692006
rect 675759 692002 676288 692004
rect 675759 691946 675764 692002
rect 675820 691946 676288 692002
rect 675759 691944 676288 691946
rect 675759 691941 675825 691944
rect 676282 691942 676288 691944
rect 676352 691942 676358 692006
rect 40762 690166 40768 690230
rect 40832 690228 40838 690230
rect 42106 690228 42112 690230
rect 40832 690168 42112 690228
rect 40832 690166 40838 690168
rect 42106 690166 42112 690168
rect 42176 690166 42182 690230
rect 42831 689488 42897 689491
rect 42528 689486 42897 689488
rect 42528 689430 42836 689486
rect 42892 689430 42897 689486
rect 42528 689428 42897 689430
rect 42831 689425 42897 689428
rect 42447 689192 42513 689195
rect 42447 689190 42558 689192
rect 42447 689134 42452 689190
rect 42508 689134 42558 689190
rect 42447 689129 42558 689134
rect 42498 688866 42558 689129
rect 42447 688600 42513 688603
rect 42447 688598 42558 688600
rect 42447 688542 42452 688598
rect 42508 688542 42558 688598
rect 42447 688537 42558 688542
rect 42498 688422 42558 688537
rect 59535 688008 59601 688011
rect 59535 688006 64416 688008
rect 59535 687950 59540 688006
rect 59596 687950 64416 688006
rect 59535 687948 64416 687950
rect 59535 687945 59601 687948
rect 42528 687800 43518 687860
rect 43215 687712 43281 687715
rect 42498 687710 43281 687712
rect 42498 687654 43220 687710
rect 43276 687654 43281 687710
rect 42498 687652 43281 687654
rect 42498 687238 42558 687652
rect 43215 687649 43281 687652
rect 43215 687564 43281 687567
rect 43458 687564 43518 687800
rect 43215 687562 43518 687564
rect 43215 687506 43220 687562
rect 43276 687506 43518 687562
rect 43215 687504 43518 687506
rect 43215 687501 43281 687504
rect 41338 686910 41344 686974
rect 41408 686910 41414 686974
rect 41346 686824 41406 686910
rect 41346 686794 42144 686824
rect 41376 686764 42174 686794
rect 42114 686530 42174 686764
rect 42106 686466 42112 686530
rect 42176 686466 42182 686530
rect 40770 685938 40830 686202
rect 40762 685874 40768 685938
rect 40832 685874 40838 685938
rect 41922 685495 41982 685610
rect 41871 685490 41982 685495
rect 41871 685434 41876 685490
rect 41932 685434 41982 685490
rect 41871 685432 41982 685434
rect 41871 685429 41937 685432
rect 42498 684903 42558 685166
rect 42447 684898 42558 684903
rect 42447 684842 42452 684898
rect 42508 684842 42558 684898
rect 42447 684840 42558 684842
rect 42447 684837 42513 684840
rect 40194 684311 40254 684574
rect 40194 684306 40305 684311
rect 40194 684250 40244 684306
rect 40300 684250 40305 684306
rect 40194 684248 40305 684250
rect 40239 684245 40305 684248
rect 41730 683719 41790 683982
rect 41679 683714 41790 683719
rect 41679 683658 41684 683714
rect 41740 683658 41790 683714
rect 41679 683656 41790 683658
rect 41679 683653 41745 683656
rect 655119 683568 655185 683571
rect 650208 683566 655185 683568
rect 41538 683127 41598 683538
rect 650208 683510 655124 683566
rect 655180 683510 655185 683566
rect 650208 683508 655185 683510
rect 655119 683505 655185 683508
rect 41538 683122 41649 683127
rect 41538 683066 41588 683122
rect 41644 683066 41649 683122
rect 41538 683064 41649 683066
rect 41583 683061 41649 683064
rect 41922 682683 41982 682946
rect 41922 682678 42033 682683
rect 41922 682622 41972 682678
rect 42028 682622 42033 682678
rect 41922 682620 42033 682622
rect 41967 682617 42033 682620
rect 42874 682384 42880 682386
rect 42528 682324 42880 682384
rect 42874 682322 42880 682324
rect 42944 682322 42950 682386
rect 42114 681499 42174 681910
rect 42114 681494 42225 681499
rect 42114 681438 42164 681494
rect 42220 681438 42225 681494
rect 42114 681436 42225 681438
rect 42159 681433 42225 681436
rect 40578 681055 40638 681318
rect 40527 681050 40638 681055
rect 40527 680994 40532 681050
rect 40588 680994 40638 681050
rect 40527 680992 40638 680994
rect 40527 680989 40593 680992
rect 43023 680756 43089 680759
rect 42528 680754 43089 680756
rect 42528 680698 43028 680754
rect 43084 680698 43089 680754
rect 42528 680696 43089 680698
rect 43023 680693 43089 680696
rect 40578 679871 40638 680208
rect 40578 679866 40689 679871
rect 40578 679810 40628 679866
rect 40684 679810 40689 679866
rect 40578 679808 40689 679810
rect 40623 679805 40689 679808
rect 41487 679868 41553 679871
rect 41487 679866 41598 679868
rect 41487 679810 41492 679866
rect 41548 679810 41598 679866
rect 41487 679805 41598 679810
rect 41538 679690 41598 679805
rect 43119 679128 43185 679131
rect 42528 679126 43185 679128
rect 42528 679070 43124 679126
rect 43180 679070 43185 679126
rect 42528 679068 43185 679070
rect 43119 679065 43185 679068
rect 42114 678391 42174 678580
rect 42063 678386 42174 678391
rect 42063 678330 42068 678386
rect 42124 678330 42174 678386
rect 42063 678328 42174 678330
rect 42063 678325 42129 678328
rect 42498 677796 42558 678062
rect 42498 677736 42750 677796
rect 35202 677207 35262 677470
rect 42690 677352 42750 677736
rect 42498 677292 42750 677352
rect 35202 677202 35313 677207
rect 35202 677146 35252 677202
rect 35308 677146 35313 677202
rect 35202 677144 35313 677146
rect 35247 677141 35313 677144
rect 42498 676908 42558 677292
rect 53679 676908 53745 676911
rect 42498 676906 53745 676908
rect 42498 676850 53684 676906
rect 53740 676850 53745 676906
rect 42498 676848 53745 676850
rect 53679 676845 53745 676848
rect 35247 676760 35313 676763
rect 35202 676758 35313 676760
rect 35202 676702 35252 676758
rect 35308 676702 35313 676758
rect 35202 676697 35313 676702
rect 35202 676434 35262 676697
rect 59535 673652 59601 673655
rect 59535 673650 64416 673652
rect 59535 673594 59540 673650
rect 59596 673594 64416 673650
rect 59535 673592 64416 673594
rect 59535 673589 59601 673592
rect 40239 673356 40305 673359
rect 43066 673356 43072 673358
rect 40239 673354 43072 673356
rect 40239 673298 40244 673354
rect 40300 673298 43072 673354
rect 40239 673296 43072 673298
rect 40239 673293 40305 673296
rect 43066 673294 43072 673296
rect 43136 673294 43142 673358
rect 674703 672912 674769 672915
rect 674703 672910 674814 672912
rect 674703 672854 674708 672910
rect 674764 672854 674814 672910
rect 674703 672849 674814 672854
rect 674754 672660 674814 672849
rect 674703 672320 674769 672323
rect 674703 672318 674814 672320
rect 674703 672262 674708 672318
rect 674764 672262 674814 672318
rect 674703 672257 674814 672262
rect 674754 672142 674814 672257
rect 674703 671876 674769 671879
rect 674703 671874 674814 671876
rect 674703 671818 674708 671874
rect 674764 671818 674814 671874
rect 674703 671813 674814 671818
rect 654447 671728 654513 671731
rect 650208 671726 654513 671728
rect 650208 671670 654452 671726
rect 654508 671670 654513 671726
rect 650208 671668 654513 671670
rect 654447 671665 654513 671668
rect 674754 671550 674814 671813
rect 40527 671138 40593 671139
rect 40527 671134 40576 671138
rect 40640 671136 40646 671138
rect 673839 671136 673905 671139
rect 40527 671078 40532 671134
rect 40527 671074 40576 671078
rect 40640 671076 40684 671136
rect 673839 671134 674814 671136
rect 673839 671078 673844 671134
rect 673900 671078 674814 671134
rect 673839 671076 674814 671078
rect 40640 671074 40646 671076
rect 40527 671073 40593 671074
rect 673839 671073 673905 671076
rect 674754 671032 674814 671076
rect 40623 670988 40689 670991
rect 40954 670988 40960 670990
rect 40623 670986 40960 670988
rect 40623 670930 40628 670986
rect 40684 670930 40960 670986
rect 40623 670928 40960 670930
rect 40623 670925 40689 670928
rect 40954 670926 40960 670928
rect 41024 670926 41030 670990
rect 41583 670988 41649 670991
rect 41722 670988 41728 670990
rect 41583 670986 41728 670988
rect 41583 670930 41588 670986
rect 41644 670930 41728 670986
rect 41583 670928 41728 670930
rect 41583 670925 41649 670928
rect 41722 670926 41728 670928
rect 41792 670926 41798 670990
rect 43119 670842 43185 670843
rect 43066 670840 43072 670842
rect 43028 670780 43072 670840
rect 43136 670838 43185 670842
rect 43180 670782 43185 670838
rect 43066 670778 43072 670780
rect 43136 670778 43185 670782
rect 43119 670777 43185 670778
rect 41775 670692 41841 670695
rect 42490 670692 42496 670694
rect 41775 670690 42496 670692
rect 41775 670634 41780 670690
rect 41836 670634 42496 670690
rect 41775 670632 42496 670634
rect 41775 670629 41841 670632
rect 42490 670630 42496 670632
rect 42560 670630 42566 670694
rect 677250 670250 677310 670514
rect 677050 670186 677056 670250
rect 677120 670186 677126 670250
rect 677242 670186 677248 670250
rect 677312 670186 677318 670250
rect 677058 669922 677118 670186
rect 676858 669594 676864 669658
rect 676928 669594 676934 669658
rect 676090 669150 676096 669214
rect 676160 669150 676166 669214
rect 676098 668886 676158 669150
rect 676866 669064 676926 669594
rect 677818 669064 677824 669066
rect 676866 669004 677824 669064
rect 677818 669002 677824 669004
rect 677888 669002 677894 669066
rect 41722 668558 41728 668622
rect 41792 668620 41798 668622
rect 42735 668620 42801 668623
rect 41792 668618 42801 668620
rect 41792 668562 42740 668618
rect 42796 668562 42801 668618
rect 41792 668560 42801 668562
rect 41792 668558 41798 668560
rect 42735 668557 42801 668560
rect 674703 668620 674769 668623
rect 674703 668618 674814 668620
rect 674703 668562 674708 668618
rect 674764 668562 674814 668618
rect 674703 668557 674814 668562
rect 42298 668410 42304 668474
rect 42368 668472 42374 668474
rect 43258 668472 43264 668474
rect 42368 668412 43264 668472
rect 42368 668410 42374 668412
rect 43258 668410 43264 668412
rect 43328 668410 43334 668474
rect 674754 668294 674814 668557
rect 674170 667744 674176 667808
rect 674240 667806 674246 667808
rect 674240 667746 674784 667806
rect 674240 667744 674246 667746
rect 675130 667522 675136 667586
rect 675200 667522 675206 667586
rect 675138 667258 675198 667522
rect 674415 666696 674481 666699
rect 674415 666694 674784 666696
rect 674415 666638 674420 666694
rect 674476 666638 674784 666694
rect 674415 666636 674784 666638
rect 674415 666633 674481 666636
rect 674223 666178 674289 666181
rect 674223 666176 674784 666178
rect 674223 666120 674228 666176
rect 674284 666120 674784 666176
rect 674223 666118 674784 666120
rect 674223 666115 674289 666118
rect 675514 665894 675520 665958
rect 675584 665894 675590 665958
rect 675522 665630 675582 665894
rect 674938 665302 674944 665366
rect 675008 665302 675014 665366
rect 674946 665038 675006 665302
rect 40954 664562 40960 664626
rect 41024 664624 41030 664626
rect 41775 664624 41841 664627
rect 41024 664622 41841 664624
rect 41024 664566 41780 664622
rect 41836 664566 41841 664622
rect 41024 664564 41841 664566
rect 41024 664562 41030 664564
rect 41775 664561 41841 664564
rect 674362 664488 674368 664552
rect 674432 664550 674438 664552
rect 674432 664490 674784 664550
rect 674432 664488 674438 664490
rect 42159 664180 42225 664183
rect 43066 664180 43072 664182
rect 42159 664178 43072 664180
rect 42159 664122 42164 664178
rect 42220 664122 43072 664178
rect 42159 664120 43072 664122
rect 42159 664117 42225 664120
rect 43066 664118 43072 664120
rect 43136 664118 43142 664182
rect 674703 664180 674769 664183
rect 674703 664178 674814 664180
rect 674703 664122 674708 664178
rect 674764 664122 674814 664178
rect 674703 664117 674814 664122
rect 674754 664002 674814 664117
rect 673839 663440 673905 663443
rect 673839 663438 674784 663440
rect 673839 663382 673844 663438
rect 673900 663382 674784 663438
rect 673839 663380 674784 663382
rect 673839 663377 673905 663380
rect 42447 662850 42513 662851
rect 42447 662846 42496 662850
rect 42560 662848 42566 662850
rect 673359 662848 673425 662851
rect 42447 662790 42452 662846
rect 42447 662786 42496 662790
rect 42560 662788 42604 662848
rect 673359 662846 674784 662848
rect 673359 662790 673364 662846
rect 673420 662790 674784 662846
rect 673359 662788 674784 662790
rect 42560 662786 42566 662788
rect 42447 662785 42513 662786
rect 673359 662785 673425 662788
rect 673263 662404 673329 662407
rect 673263 662402 674784 662404
rect 673263 662346 673268 662402
rect 673324 662346 674784 662402
rect 673263 662344 674784 662346
rect 673263 662341 673329 662344
rect 673839 661812 673905 661815
rect 673839 661810 674784 661812
rect 673839 661754 673844 661810
rect 673900 661754 674784 661810
rect 673839 661752 674784 661754
rect 673839 661749 673905 661752
rect 41775 661518 41841 661519
rect 41722 661454 41728 661518
rect 41792 661516 41841 661518
rect 41792 661514 41884 661516
rect 41836 661458 41884 661514
rect 41792 661456 41884 661458
rect 41792 661454 41841 661456
rect 41775 661453 41841 661454
rect 41871 661370 41937 661371
rect 41871 661368 41920 661370
rect 41828 661366 41920 661368
rect 41828 661310 41876 661366
rect 41828 661308 41920 661310
rect 41871 661306 41920 661308
rect 41984 661306 41990 661370
rect 41871 661305 41937 661306
rect 674754 660927 674814 661190
rect 674703 660922 674814 660927
rect 674703 660866 674708 660922
rect 674764 660866 674814 660922
rect 674703 660864 674814 660866
rect 674703 660861 674769 660864
rect 649935 660628 650001 660631
rect 649935 660626 650046 660628
rect 649935 660570 649940 660626
rect 649996 660570 650046 660626
rect 649935 660565 650046 660570
rect 40570 660270 40576 660334
rect 40640 660332 40646 660334
rect 41775 660332 41841 660335
rect 40640 660330 41841 660332
rect 40640 660274 41780 660330
rect 41836 660274 41841 660330
rect 40640 660272 41841 660274
rect 40640 660270 40646 660272
rect 41775 660269 41841 660272
rect 649986 660006 650046 660565
rect 675138 660483 675198 660746
rect 674703 660480 674769 660483
rect 674703 660478 674814 660480
rect 674703 660422 674708 660478
rect 674764 660422 674814 660478
rect 674703 660417 674814 660422
rect 675087 660478 675198 660483
rect 675087 660422 675092 660478
rect 675148 660422 675198 660478
rect 675087 660420 675198 660422
rect 675087 660417 675153 660420
rect 674754 660154 674814 660417
rect 675087 659888 675153 659891
rect 675087 659886 675198 659888
rect 675087 659830 675092 659886
rect 675148 659830 675198 659886
rect 675087 659825 675198 659830
rect 42874 659530 42880 659594
rect 42944 659592 42950 659594
rect 42944 659532 43134 659592
rect 675138 659562 675198 659825
rect 42944 659530 42950 659532
rect 43074 659151 43134 659532
rect 59535 659296 59601 659299
rect 59535 659294 64416 659296
rect 59535 659238 59540 659294
rect 59596 659238 64416 659294
rect 59535 659236 64416 659238
rect 59535 659233 59601 659236
rect 43074 659146 43185 659151
rect 43074 659090 43124 659146
rect 43180 659090 43185 659146
rect 43074 659088 43185 659090
rect 43119 659085 43185 659088
rect 677050 658790 677056 658854
rect 677120 658852 677126 658854
rect 677818 658852 677824 658854
rect 677120 658792 677824 658852
rect 677120 658790 677126 658792
rect 677818 658790 677824 658792
rect 677888 658790 677894 658854
rect 42159 656188 42225 656191
rect 42298 656188 42304 656190
rect 42159 656186 42304 656188
rect 42159 656130 42164 656186
rect 42220 656130 42304 656186
rect 42159 656128 42304 656130
rect 42159 656125 42225 656128
rect 42298 656126 42304 656128
rect 42368 656126 42374 656190
rect 674703 653672 674769 653675
rect 676282 653672 676288 653674
rect 674703 653670 676288 653672
rect 674703 653614 674708 653670
rect 674764 653614 676288 653670
rect 674703 653612 676288 653614
rect 674703 653609 674769 653612
rect 676282 653610 676288 653612
rect 676352 653610 676358 653674
rect 675130 652574 675136 652638
rect 675200 652636 675206 652638
rect 675375 652636 675441 652639
rect 675200 652634 675441 652636
rect 675200 652578 675380 652634
rect 675436 652578 675441 652634
rect 675200 652576 675441 652578
rect 675200 652574 675206 652576
rect 675375 652573 675441 652576
rect 674362 652130 674368 652194
rect 674432 652192 674438 652194
rect 675471 652192 675537 652195
rect 674432 652190 675537 652192
rect 674432 652134 675476 652190
rect 675532 652134 675537 652190
rect 674432 652132 675537 652134
rect 674432 652130 674438 652132
rect 675471 652129 675537 652132
rect 675471 651454 675537 651455
rect 675471 651450 675520 651454
rect 675584 651452 675590 651454
rect 675471 651394 675476 651450
rect 675471 651390 675520 651394
rect 675584 651392 675628 651452
rect 675584 651390 675590 651392
rect 675471 651389 675537 651390
rect 675663 649826 675729 649827
rect 675663 649822 675712 649826
rect 675776 649824 675782 649826
rect 675663 649766 675668 649822
rect 675663 649762 675712 649766
rect 675776 649764 675820 649824
rect 675776 649762 675782 649764
rect 675663 649761 675729 649762
rect 674938 648874 674944 648938
rect 675008 648936 675014 648938
rect 675471 648936 675537 648939
rect 675008 648934 675537 648936
rect 675008 648878 675476 648934
rect 675532 648878 675537 648934
rect 675008 648876 675537 648878
rect 675008 648874 675014 648876
rect 675471 648873 675537 648876
rect 654255 648344 654321 648347
rect 650208 648342 654321 648344
rect 650208 648286 654260 648342
rect 654316 648286 654321 648342
rect 650208 648284 654321 648286
rect 654255 648281 654321 648284
rect 42106 647098 42112 647162
rect 42176 647160 42182 647162
rect 43791 647160 43857 647163
rect 42176 647158 43857 647160
rect 42176 647102 43796 647158
rect 43852 647102 43857 647158
rect 42176 647100 43857 647102
rect 42176 647098 42182 647100
rect 43791 647097 43857 647100
rect 40762 646950 40768 647014
rect 40832 647012 40838 647014
rect 43599 647012 43665 647015
rect 40832 647010 43665 647012
rect 40832 646954 43604 647010
rect 43660 646954 43665 647010
rect 40832 646952 43665 646954
rect 40832 646950 40838 646952
rect 43599 646949 43665 646952
rect 42927 646272 42993 646275
rect 42528 646270 42993 646272
rect 42528 646214 42932 646270
rect 42988 646214 42993 646270
rect 42528 646212 42993 646214
rect 42927 646209 42993 646212
rect 42498 645535 42558 645724
rect 42447 645530 42558 645535
rect 42447 645474 42452 645530
rect 42508 645474 42558 645530
rect 42447 645472 42558 645474
rect 42447 645469 42513 645472
rect 673978 645322 673984 645386
rect 674048 645384 674054 645386
rect 675471 645384 675537 645387
rect 674048 645382 675537 645384
rect 674048 645326 675476 645382
rect 675532 645326 675537 645382
rect 674048 645324 675537 645326
rect 674048 645322 674054 645324
rect 675471 645321 675537 645324
rect 42927 645236 42993 645239
rect 42528 645234 42993 645236
rect 42528 645178 42932 645234
rect 42988 645178 42993 645234
rect 42528 645176 42993 645178
rect 42927 645173 42993 645176
rect 59535 644940 59601 644943
rect 59535 644938 64416 644940
rect 59535 644882 59540 644938
rect 59596 644882 64416 644938
rect 59535 644880 64416 644882
rect 59535 644877 59601 644880
rect 43407 644644 43473 644647
rect 42528 644642 43473 644644
rect 42528 644586 43412 644642
rect 43468 644586 43473 644642
rect 42528 644584 43473 644586
rect 43407 644581 43473 644584
rect 43215 644496 43281 644499
rect 42498 644494 43281 644496
rect 42498 644438 43220 644494
rect 43276 644438 43281 644494
rect 42498 644436 43281 644438
rect 42498 644096 42558 644436
rect 43215 644433 43281 644436
rect 43791 643608 43857 643611
rect 42528 643606 43857 643608
rect 42528 643550 43796 643606
rect 43852 643550 43857 643606
rect 42528 643548 43857 643550
rect 43791 643545 43857 643548
rect 43599 643016 43665 643019
rect 42528 643014 43665 643016
rect 42528 642958 43604 643014
rect 43660 642958 43665 643014
rect 42528 642956 43665 642958
rect 43599 642953 43665 642956
rect 41538 642279 41598 642468
rect 674127 642313 674193 642316
rect 673986 642311 674193 642313
rect 673986 642279 674132 642311
rect 41487 642274 41598 642279
rect 41487 642218 41492 642274
rect 41548 642218 41598 642274
rect 41487 642216 41598 642218
rect 673935 642274 674132 642279
rect 673935 642218 673940 642274
rect 673996 642255 674132 642274
rect 674188 642255 674193 642311
rect 673996 642253 674193 642255
rect 673996 642218 674046 642253
rect 674127 642250 674193 642253
rect 673935 642216 674046 642218
rect 41487 642213 41553 642216
rect 673935 642213 674001 642216
rect 42927 641980 42993 641983
rect 42528 641978 42993 641980
rect 42528 641922 42932 641978
rect 42988 641922 42993 641978
rect 42528 641920 42993 641922
rect 42927 641917 42993 641920
rect 39810 641095 39870 641358
rect 39810 641090 39921 641095
rect 39810 641034 39860 641090
rect 39916 641034 39921 641090
rect 39810 641032 39921 641034
rect 39855 641029 39921 641032
rect 41538 640503 41598 640840
rect 41538 640498 41649 640503
rect 41538 640442 41588 640498
rect 41644 640442 41649 640498
rect 41538 640440 41649 640442
rect 41583 640437 41649 640440
rect 675759 640352 675825 640355
rect 676282 640352 676288 640354
rect 675759 640350 676288 640352
rect 41730 640059 41790 640322
rect 675759 640294 675764 640350
rect 675820 640294 676288 640350
rect 675759 640292 676288 640294
rect 675759 640289 675825 640292
rect 676282 640290 676288 640292
rect 676352 640290 676358 640354
rect 41679 640054 41790 640059
rect 41679 639998 41684 640054
rect 41740 639998 41790 640054
rect 41679 639996 41790 639998
rect 41679 639993 41745 639996
rect 41922 639467 41982 639730
rect 41871 639462 41982 639467
rect 41871 639406 41876 639462
rect 41932 639406 41982 639462
rect 41871 639404 41982 639406
rect 41871 639401 41937 639404
rect 40194 638875 40254 639138
rect 40194 638870 40305 638875
rect 40194 638814 40244 638870
rect 40300 638814 40305 638870
rect 40194 638812 40305 638814
rect 40239 638809 40305 638812
rect 41346 638431 41406 638694
rect 675759 638576 675825 638579
rect 676090 638576 676096 638578
rect 675759 638574 676096 638576
rect 675759 638518 675764 638574
rect 675820 638518 676096 638574
rect 675759 638516 676096 638518
rect 675759 638513 675825 638516
rect 676090 638514 676096 638516
rect 676160 638514 676166 638578
rect 41295 638426 41406 638431
rect 41295 638370 41300 638426
rect 41356 638370 41406 638426
rect 41295 638368 41406 638370
rect 41295 638365 41361 638368
rect 43119 638132 43185 638135
rect 42528 638130 43185 638132
rect 42528 638074 43124 638130
rect 43180 638074 43185 638130
rect 42528 638072 43185 638074
rect 43119 638069 43185 638072
rect 42498 637244 42558 637510
rect 42874 637244 42880 637246
rect 42498 637184 42880 637244
rect 42874 637182 42880 637184
rect 42944 637182 42950 637246
rect 42114 636803 42174 637066
rect 42063 636798 42174 636803
rect 42063 636742 42068 636798
rect 42124 636742 42174 636798
rect 42063 636740 42174 636742
rect 42063 636737 42129 636740
rect 655311 636652 655377 636655
rect 650208 636650 655377 636652
rect 650208 636594 655316 636650
rect 655372 636594 655377 636650
rect 650208 636592 655377 636594
rect 655311 636589 655377 636592
rect 41922 636211 41982 636474
rect 41922 636206 42033 636211
rect 41922 636150 41972 636206
rect 42028 636150 42033 636206
rect 41922 636148 42033 636150
rect 41967 636145 42033 636148
rect 42114 635619 42174 635882
rect 42114 635614 42225 635619
rect 43023 635616 43089 635619
rect 42114 635558 42164 635614
rect 42220 635558 42225 635614
rect 42114 635556 42225 635558
rect 42159 635553 42225 635556
rect 42498 635614 43089 635616
rect 42498 635558 43028 635614
rect 43084 635558 43089 635614
rect 42498 635556 43089 635558
rect 42498 635438 42558 635556
rect 43023 635553 43089 635556
rect 42498 634580 42558 634846
rect 42498 634520 42750 634580
rect 35202 633991 35262 634254
rect 42690 634136 42750 634520
rect 35151 633986 35262 633991
rect 35151 633930 35156 633986
rect 35212 633930 35262 633986
rect 35151 633928 35262 633930
rect 42498 634076 42750 634136
rect 42498 633988 42558 634076
rect 56079 633988 56145 633991
rect 42498 633986 56145 633988
rect 42498 633930 56084 633986
rect 56140 633930 56145 633986
rect 42498 633928 56145 633930
rect 35151 633925 35217 633928
rect 42498 633810 42558 633928
rect 56079 633925 56145 633928
rect 35151 633544 35217 633547
rect 35151 633542 35262 633544
rect 35151 633486 35156 633542
rect 35212 633486 35262 633542
rect 35151 633481 35262 633486
rect 35202 633218 35262 633481
rect 59535 630584 59601 630587
rect 59535 630582 64416 630584
rect 59535 630526 59540 630582
rect 59596 630526 64416 630582
rect 59535 630524 64416 630526
rect 59535 630521 59601 630524
rect 40239 628068 40305 628071
rect 42298 628068 42304 628070
rect 40239 628066 42304 628068
rect 40239 628010 40244 628066
rect 40300 628010 42304 628066
rect 40239 628008 42304 628010
rect 40239 628005 40305 628008
rect 42298 628006 42304 628008
rect 42368 628006 42374 628070
rect 39855 627920 39921 627923
rect 40762 627920 40768 627922
rect 39855 627918 40768 627920
rect 39855 627862 39860 627918
rect 39916 627862 40768 627918
rect 39855 627860 40768 627862
rect 39855 627857 39921 627860
rect 40762 627858 40768 627860
rect 40832 627858 40838 627922
rect 41487 627920 41553 627923
rect 42490 627920 42496 627922
rect 41487 627918 42496 627920
rect 41487 627862 41492 627918
rect 41548 627862 42496 627918
rect 41487 627860 42496 627862
rect 41487 627857 41553 627860
rect 42490 627858 42496 627860
rect 42560 627858 42566 627922
rect 41295 627774 41361 627775
rect 41295 627772 41344 627774
rect 41252 627770 41344 627772
rect 41252 627714 41300 627770
rect 41252 627712 41344 627714
rect 41295 627710 41344 627712
rect 41408 627710 41414 627774
rect 41583 627772 41649 627775
rect 41722 627772 41728 627774
rect 41583 627770 41728 627772
rect 41583 627714 41588 627770
rect 41644 627714 41728 627770
rect 41583 627712 41728 627714
rect 41295 627709 41361 627710
rect 41583 627709 41649 627712
rect 41722 627710 41728 627712
rect 41792 627710 41798 627774
rect 674415 627698 674481 627701
rect 674415 627696 674784 627698
rect 674415 627640 674420 627696
rect 674476 627640 674784 627696
rect 674415 627638 674784 627640
rect 674415 627635 674481 627638
rect 41967 627478 42033 627479
rect 41914 627414 41920 627478
rect 41984 627476 42033 627478
rect 41984 627474 42076 627476
rect 42028 627418 42076 627474
rect 41984 627416 42076 627418
rect 41984 627414 42033 627416
rect 41967 627413 42033 627414
rect 674895 627328 674961 627331
rect 674895 627326 675006 627328
rect 674895 627270 674900 627326
rect 674956 627270 675006 627326
rect 674895 627265 675006 627270
rect 674946 627150 675006 627265
rect 674415 626588 674481 626591
rect 674415 626586 674784 626588
rect 674415 626530 674420 626586
rect 674476 626530 674784 626586
rect 674415 626528 674784 626530
rect 674415 626525 674481 626528
rect 677242 626378 677248 626442
rect 677312 626378 677318 626442
rect 677250 626040 677310 626378
rect 42106 625638 42112 625702
rect 42176 625700 42182 625702
rect 42682 625700 42688 625702
rect 42176 625640 42688 625700
rect 42176 625638 42182 625640
rect 42682 625638 42688 625640
rect 42752 625638 42758 625702
rect 674415 625552 674481 625555
rect 674415 625550 674784 625552
rect 674415 625494 674420 625550
rect 674476 625494 674784 625550
rect 674415 625492 674784 625494
rect 674415 625489 674481 625492
rect 42106 624898 42112 624962
rect 42176 624960 42182 624962
rect 42682 624960 42688 624962
rect 42176 624900 42688 624960
rect 42176 624898 42182 624900
rect 42682 624898 42688 624900
rect 42752 624898 42758 624962
rect 676866 624815 676926 624930
rect 654351 624812 654417 624815
rect 676815 624814 676926 624815
rect 676815 624812 676864 624814
rect 650208 624810 654417 624812
rect 650208 624754 654356 624810
rect 654412 624754 654417 624810
rect 650208 624752 654417 624754
rect 676736 624810 676864 624812
rect 676736 624754 676820 624810
rect 676736 624752 676864 624754
rect 654351 624749 654417 624752
rect 676815 624750 676864 624752
rect 676928 624750 676934 624814
rect 676815 624749 676881 624750
rect 677050 624602 677056 624666
rect 677120 624602 677126 624666
rect 675322 624158 675328 624222
rect 675392 624158 675398 624222
rect 675330 623894 675390 624158
rect 676911 624072 676977 624075
rect 677058 624072 677118 624602
rect 676911 624070 677118 624072
rect 676911 624014 676916 624070
rect 676972 624014 677118 624070
rect 676911 624012 677118 624014
rect 676911 624009 676977 624012
rect 42159 623480 42225 623483
rect 42874 623480 42880 623482
rect 42159 623478 42880 623480
rect 42159 623422 42164 623478
rect 42220 623422 42880 623478
rect 42159 623420 42880 623422
rect 42159 623417 42225 623420
rect 42874 623418 42880 623420
rect 42944 623418 42950 623482
rect 673935 623332 674001 623335
rect 673935 623330 674784 623332
rect 673935 623274 673940 623330
rect 673996 623274 674784 623330
rect 673935 623272 674784 623274
rect 673935 623269 674001 623272
rect 674746 623122 674752 623186
rect 674816 623122 674822 623186
rect 674754 622784 674814 623122
rect 675898 622530 675904 622594
rect 675968 622530 675974 622594
rect 675906 622266 675966 622530
rect 674511 622000 674577 622003
rect 674511 621998 674814 622000
rect 674511 621942 674516 621998
rect 674572 621942 674814 621998
rect 674511 621940 674814 621942
rect 674511 621937 674577 621940
rect 674754 621674 674814 621940
rect 42490 621494 42496 621558
rect 42560 621556 42566 621558
rect 43119 621556 43185 621559
rect 42560 621554 43185 621556
rect 42560 621498 43124 621554
rect 43180 621498 43185 621554
rect 42560 621496 43185 621498
rect 42560 621494 42566 621496
rect 43119 621493 43185 621496
rect 675087 621408 675153 621411
rect 675087 621406 675198 621408
rect 675087 621350 675092 621406
rect 675148 621350 675198 621406
rect 675087 621345 675198 621350
rect 675138 621082 675198 621345
rect 676666 620902 676672 620966
rect 676736 620902 676742 620966
rect 676674 620638 676734 620902
rect 674554 620310 674560 620374
rect 674624 620372 674630 620374
rect 674624 620312 674814 620372
rect 674624 620310 674630 620312
rect 674754 620046 674814 620312
rect 676474 619866 676480 619930
rect 676544 619866 676550 619930
rect 41722 619570 41728 619634
rect 41792 619632 41798 619634
rect 42447 619632 42513 619635
rect 41792 619630 42513 619632
rect 41792 619574 42452 619630
rect 42508 619574 42513 619630
rect 41792 619572 42513 619574
rect 41792 619570 41798 619572
rect 42447 619569 42513 619572
rect 676482 619454 676542 619866
rect 674607 619188 674673 619191
rect 674607 619186 674814 619188
rect 674607 619130 674612 619186
rect 674668 619130 674814 619186
rect 674607 619128 674814 619130
rect 674607 619125 674673 619128
rect 674754 619010 674814 619128
rect 41530 618386 41536 618450
rect 41600 618448 41606 618450
rect 41775 618448 41841 618451
rect 42682 618448 42688 618450
rect 41600 618446 42688 618448
rect 41600 618390 41780 618446
rect 41836 618390 42688 618446
rect 41600 618388 42688 618390
rect 41600 618386 41606 618388
rect 41775 618385 41841 618388
rect 42682 618386 42688 618388
rect 42752 618386 42758 618450
rect 674415 618448 674481 618451
rect 674415 618446 674784 618448
rect 674415 618390 674420 618446
rect 674476 618390 674784 618446
rect 674415 618388 674784 618390
rect 674415 618385 674481 618388
rect 41775 618302 41841 618303
rect 41722 618238 41728 618302
rect 41792 618300 41841 618302
rect 41792 618298 41884 618300
rect 41836 618242 41884 618298
rect 41792 618240 41884 618242
rect 41792 618238 41841 618240
rect 41775 618237 41841 618238
rect 41967 617858 42033 617859
rect 41914 617856 41920 617858
rect 41876 617796 41920 617856
rect 41984 617854 42033 617858
rect 42028 617798 42033 617854
rect 41914 617794 41920 617796
rect 41984 617794 42033 617798
rect 41967 617793 42033 617794
rect 674415 617856 674481 617859
rect 674415 617854 674784 617856
rect 674415 617798 674420 617854
rect 674476 617798 674784 617854
rect 674415 617796 674784 617798
rect 674415 617793 674481 617796
rect 674703 617560 674769 617563
rect 674703 617558 674814 617560
rect 674703 617502 674708 617558
rect 674764 617502 674814 617558
rect 674703 617497 674814 617502
rect 674754 617382 674814 617497
rect 673167 616820 673233 616823
rect 673167 616818 674784 616820
rect 673167 616762 673172 616818
rect 673228 616762 674784 616818
rect 673167 616760 674784 616762
rect 673167 616757 673233 616760
rect 41338 616610 41344 616674
rect 41408 616672 41414 616674
rect 41775 616672 41841 616675
rect 41408 616670 41841 616672
rect 41408 616614 41780 616670
rect 41836 616614 41841 616670
rect 41408 616612 41841 616614
rect 41408 616610 41414 616612
rect 41775 616609 41841 616612
rect 59535 616228 59601 616231
rect 59535 616226 64416 616228
rect 59535 616170 59540 616226
rect 59596 616170 64416 616226
rect 59535 616168 64416 616170
rect 59535 616165 59601 616168
rect 677058 615935 677118 616198
rect 677058 615930 677169 615935
rect 677058 615874 677108 615930
rect 677164 615874 677169 615930
rect 677058 615872 677169 615874
rect 677103 615869 677169 615872
rect 676866 615343 676926 615754
rect 676866 615338 676977 615343
rect 677103 615340 677169 615343
rect 676866 615282 676916 615338
rect 676972 615282 676977 615338
rect 676866 615280 676977 615282
rect 676911 615277 676977 615280
rect 677058 615338 677169 615340
rect 677058 615282 677108 615338
rect 677164 615282 677169 615338
rect 677058 615277 677169 615282
rect 677058 615162 677118 615277
rect 676911 614896 676977 614899
rect 676866 614894 676977 614896
rect 676866 614838 676916 614894
rect 676972 614838 676977 614894
rect 676866 614833 676977 614838
rect 676866 614570 676926 614833
rect 42159 613564 42225 613567
rect 42298 613564 42304 613566
rect 42159 613562 42304 613564
rect 42159 613506 42164 613562
rect 42220 613506 42304 613562
rect 42159 613504 42304 613506
rect 42159 613501 42225 613504
rect 42298 613502 42304 613504
rect 42368 613502 42374 613566
rect 654351 613120 654417 613123
rect 650208 613118 654417 613120
rect 650208 613062 654356 613118
rect 654412 613062 654417 613118
rect 650208 613060 654417 613062
rect 654351 613057 654417 613060
rect 40762 612762 40768 612826
rect 40832 612824 40838 612826
rect 41775 612824 41841 612827
rect 40832 612822 41841 612824
rect 40832 612766 41780 612822
rect 41836 612766 41841 612822
rect 40832 612764 41841 612766
rect 40832 612762 40838 612764
rect 41775 612761 41841 612764
rect 674170 607730 674176 607794
rect 674240 607792 674246 607794
rect 675375 607792 675441 607795
rect 674240 607790 675441 607792
rect 674240 607734 675380 607790
rect 675436 607734 675441 607790
rect 674240 607732 675441 607734
rect 674240 607730 674246 607732
rect 675375 607729 675441 607732
rect 674746 607138 674752 607202
rect 674816 607200 674822 607202
rect 675471 607200 675537 607203
rect 674816 607198 675537 607200
rect 674816 607142 675476 607198
rect 675532 607142 675537 607198
rect 674816 607140 675537 607142
rect 674816 607138 674822 607140
rect 675471 607137 675537 607140
rect 675322 606398 675328 606462
rect 675392 606460 675398 606462
rect 675471 606460 675537 606463
rect 675392 606458 675537 606460
rect 675392 606402 675476 606458
rect 675532 606402 675537 606458
rect 675392 606400 675537 606402
rect 675392 606398 675398 606400
rect 675471 606397 675537 606400
rect 41530 604770 41536 604834
rect 41600 604832 41606 604834
rect 42106 604832 42112 604834
rect 41600 604772 42112 604832
rect 41600 604770 41606 604772
rect 42106 604770 42112 604772
rect 42176 604770 42182 604834
rect 674554 604770 674560 604834
rect 674624 604832 674630 604834
rect 675375 604832 675441 604835
rect 674624 604830 675441 604832
rect 674624 604774 675380 604830
rect 675436 604774 675441 604830
rect 674624 604772 675441 604774
rect 674624 604770 674630 604772
rect 675375 604769 675441 604772
rect 42831 603056 42897 603059
rect 42528 603054 42897 603056
rect 42528 602998 42836 603054
rect 42892 602998 42897 603054
rect 42528 602996 42897 602998
rect 42831 602993 42897 602996
rect 42498 602316 42558 602582
rect 42735 602316 42801 602319
rect 42498 602314 42801 602316
rect 42498 602258 42740 602314
rect 42796 602258 42801 602314
rect 42498 602256 42801 602258
rect 42735 602253 42801 602256
rect 42159 602168 42225 602171
rect 42114 602166 42225 602168
rect 42114 602110 42164 602166
rect 42220 602110 42225 602166
rect 42114 602105 42225 602110
rect 42114 601990 42174 602105
rect 59535 601872 59601 601875
rect 59535 601870 64416 601872
rect 59535 601814 59540 601870
rect 59596 601814 64416 601870
rect 59535 601812 64416 601814
rect 59535 601809 59601 601812
rect 43983 601428 44049 601431
rect 654447 601428 654513 601431
rect 42528 601426 44049 601428
rect 42528 601370 43988 601426
rect 44044 601370 44049 601426
rect 42528 601368 44049 601370
rect 650208 601426 654513 601428
rect 650208 601370 654452 601426
rect 654508 601370 654513 601426
rect 650208 601368 654513 601370
rect 43983 601365 44049 601368
rect 654447 601365 654513 601368
rect 43311 601280 43377 601283
rect 42498 601278 43377 601280
rect 42498 601222 43316 601278
rect 43372 601222 43377 601278
rect 42498 601220 43377 601222
rect 42498 600880 42558 601220
rect 43311 601217 43377 601220
rect 43791 600392 43857 600395
rect 42528 600390 43857 600392
rect 42528 600334 43796 600390
rect 43852 600334 43857 600390
rect 42528 600332 43857 600334
rect 43791 600329 43857 600332
rect 675759 600244 675825 600247
rect 675898 600244 675904 600246
rect 675759 600242 675904 600244
rect 675759 600186 675764 600242
rect 675820 600186 675904 600242
rect 675759 600184 675904 600186
rect 675759 600181 675825 600184
rect 675898 600182 675904 600184
rect 675968 600182 675974 600246
rect 43599 599800 43665 599803
rect 42528 599798 43665 599800
rect 42528 599742 43604 599798
rect 43660 599742 43665 599798
rect 42528 599740 43665 599742
rect 43599 599737 43665 599740
rect 42498 599208 42558 599252
rect 43119 599208 43185 599211
rect 42498 599206 43185 599208
rect 42498 599150 43124 599206
rect 43180 599150 43185 599206
rect 42498 599148 43185 599150
rect 43119 599145 43185 599148
rect 42106 598998 42112 599062
rect 42176 599060 42182 599062
rect 43066 599060 43072 599062
rect 42176 599000 43072 599060
rect 42176 598998 42182 599000
rect 43066 598998 43072 599000
rect 43136 598998 43142 599062
rect 41922 598471 41982 598734
rect 41922 598466 42033 598471
rect 41922 598410 41972 598466
rect 42028 598410 42033 598466
rect 41922 598408 42033 598410
rect 41967 598405 42033 598408
rect 40578 597878 40638 598142
rect 40570 597814 40576 597878
rect 40640 597814 40646 597878
rect 41538 597287 41598 597624
rect 41538 597282 41649 597287
rect 41538 597226 41588 597282
rect 41644 597226 41649 597282
rect 41538 597224 41649 597226
rect 41583 597221 41649 597224
rect 41538 596843 41598 597106
rect 41487 596838 41598 596843
rect 41487 596782 41492 596838
rect 41548 596782 41598 596838
rect 41487 596780 41598 596782
rect 41487 596777 41553 596780
rect 41922 596251 41982 596514
rect 41871 596246 41982 596251
rect 41871 596190 41876 596246
rect 41932 596190 41982 596246
rect 41871 596188 41982 596190
rect 41871 596185 41937 596188
rect 40770 595658 40830 595996
rect 40762 595594 40768 595658
rect 40832 595594 40838 595658
rect 41730 595215 41790 595478
rect 675759 595360 675825 595363
rect 676666 595360 676672 595362
rect 675759 595358 676672 595360
rect 675759 595302 675764 595358
rect 675820 595302 676672 595358
rect 675759 595300 676672 595302
rect 675759 595297 675825 595300
rect 676666 595298 676672 595300
rect 676736 595298 676742 595362
rect 41730 595210 41841 595215
rect 41730 595154 41780 595210
rect 41836 595154 41841 595210
rect 41730 595152 41841 595154
rect 41775 595149 41841 595152
rect 41730 594623 41790 594886
rect 41679 594618 41790 594623
rect 41679 594562 41684 594618
rect 41740 594562 41790 594618
rect 41679 594560 41790 594562
rect 41679 594557 41745 594560
rect 41346 594030 41406 594368
rect 41338 593966 41344 594030
rect 41408 593966 41414 594030
rect 42114 593587 42174 593850
rect 42114 593582 42225 593587
rect 42114 593526 42164 593582
rect 42220 593526 42225 593582
rect 42114 593524 42225 593526
rect 42159 593521 42225 593524
rect 675759 593436 675825 593439
rect 676474 593436 676480 593438
rect 675759 593434 676480 593436
rect 675759 593378 675764 593434
rect 675820 593378 676480 593434
rect 675759 593376 676480 593378
rect 675759 593373 675825 593376
rect 676474 593374 676480 593376
rect 676544 593374 676550 593438
rect 42114 592995 42174 593258
rect 42063 592990 42174 592995
rect 42063 592934 42068 592990
rect 42124 592934 42174 592990
rect 42063 592932 42174 592934
rect 42063 592929 42129 592932
rect 42831 592770 42897 592773
rect 42528 592768 42897 592770
rect 42528 592712 42836 592768
rect 42892 592712 42897 592768
rect 42528 592710 42897 592712
rect 42831 592707 42897 592710
rect 42498 591958 42558 592222
rect 42490 591894 42496 591958
rect 42560 591894 42566 591958
rect 42498 591364 42558 591630
rect 42498 591304 42750 591364
rect 30594 590774 30654 591112
rect 42690 590920 42750 591304
rect 42498 590860 42750 590920
rect 30586 590710 30592 590774
rect 30656 590710 30662 590774
rect 42498 590624 42558 590860
rect 53775 590624 53841 590627
rect 42498 590622 53841 590624
rect 42498 590594 53780 590622
rect 42528 590566 53780 590594
rect 53836 590566 53841 590622
rect 42528 590564 53841 590566
rect 53775 590561 53841 590564
rect 30586 590266 30592 590330
rect 30656 590266 30662 590330
rect 30594 590002 30654 590266
rect 654447 589588 654513 589591
rect 650208 589586 654513 589588
rect 650208 589530 654452 589586
rect 654508 589530 654513 589586
rect 650208 589528 654513 589530
rect 654447 589525 654513 589528
rect 42490 588342 42496 588406
rect 42560 588404 42566 588406
rect 42735 588404 42801 588407
rect 42560 588402 42801 588404
rect 42560 588346 42740 588402
rect 42796 588346 42801 588402
rect 42560 588344 42801 588346
rect 42560 588342 42566 588344
rect 42735 588341 42801 588344
rect 59535 587516 59601 587519
rect 59535 587514 64416 587516
rect 59535 587458 59540 587514
rect 59596 587458 64416 587514
rect 59535 587456 64416 587458
rect 59535 587453 59601 587456
rect 41583 584704 41649 584707
rect 42298 584704 42304 584706
rect 41583 584702 42304 584704
rect 41583 584646 41588 584702
rect 41644 584646 42304 584702
rect 41583 584644 42304 584646
rect 41583 584641 41649 584644
rect 42298 584642 42304 584644
rect 42368 584642 42374 584706
rect 41679 584558 41745 584559
rect 41679 584556 41728 584558
rect 41636 584554 41728 584556
rect 41636 584498 41684 584554
rect 41636 584496 41728 584498
rect 41679 584494 41728 584496
rect 41792 584494 41798 584558
rect 42490 584494 42496 584558
rect 42560 584556 42566 584558
rect 42831 584556 42897 584559
rect 42560 584554 42897 584556
rect 42560 584498 42836 584554
rect 42892 584498 42897 584554
rect 42560 584496 42897 584498
rect 42560 584494 42566 584496
rect 41679 584493 41745 584494
rect 42831 584493 42897 584496
rect 42063 584410 42129 584411
rect 42063 584408 42112 584410
rect 42020 584406 42112 584408
rect 42020 584350 42068 584406
rect 42020 584348 42112 584350
rect 42063 584346 42112 584348
rect 42176 584346 42182 584410
rect 42063 584345 42129 584346
rect 41967 584262 42033 584263
rect 41914 584198 41920 584262
rect 41984 584260 42033 584262
rect 42159 584260 42225 584263
rect 42874 584260 42880 584262
rect 41984 584258 42076 584260
rect 42028 584202 42076 584258
rect 41984 584200 42076 584202
rect 42159 584258 42880 584260
rect 42159 584202 42164 584258
rect 42220 584202 42880 584258
rect 42159 584200 42880 584202
rect 41984 584198 42033 584200
rect 41967 584197 42033 584198
rect 42159 584197 42225 584200
rect 42874 584198 42880 584200
rect 42944 584198 42950 584262
rect 674607 582188 674673 582191
rect 674754 582188 674814 582454
rect 674607 582186 674814 582188
rect 674607 582130 674612 582186
rect 674668 582130 674814 582186
rect 674607 582128 674814 582130
rect 674607 582125 674673 582128
rect 41871 582042 41937 582043
rect 41871 582038 41920 582042
rect 41984 582040 41990 582042
rect 41871 581982 41876 582038
rect 41871 581978 41920 581982
rect 41984 581980 42028 582040
rect 41984 581978 41990 581980
rect 41871 581977 41937 581978
rect 674415 581966 674481 581969
rect 674415 581964 674784 581966
rect 674415 581908 674420 581964
rect 674476 581908 674784 581964
rect 674415 581906 674784 581908
rect 674415 581903 674481 581906
rect 674607 581596 674673 581599
rect 674607 581594 674814 581596
rect 674607 581538 674612 581594
rect 674668 581538 674814 581594
rect 674607 581536 674814 581538
rect 674607 581533 674673 581536
rect 674754 581418 674814 581536
rect 674415 580856 674481 580859
rect 674415 580854 674784 580856
rect 674415 580798 674420 580854
rect 674476 580798 674784 580854
rect 674415 580796 674784 580798
rect 674415 580793 674481 580796
rect 41338 580202 41344 580266
rect 41408 580264 41414 580266
rect 41775 580264 41841 580267
rect 41408 580262 41841 580264
rect 41408 580206 41780 580262
rect 41836 580206 41841 580262
rect 41408 580204 41841 580206
rect 41408 580202 41414 580204
rect 41775 580201 41841 580204
rect 673839 580264 673905 580267
rect 673839 580262 674784 580264
rect 673839 580206 673844 580262
rect 673900 580206 674784 580262
rect 673839 580204 674784 580206
rect 673839 580201 673905 580204
rect 672015 579820 672081 579823
rect 672015 579818 677280 579820
rect 672015 579762 672020 579818
rect 672076 579790 677280 579818
rect 672076 579762 677310 579790
rect 672015 579760 677310 579762
rect 672015 579757 672081 579760
rect 676815 579524 676881 579527
rect 677250 579526 677310 579760
rect 677050 579524 677056 579526
rect 676815 579522 677056 579524
rect 676815 579466 676820 579522
rect 676876 579466 677056 579522
rect 676815 579464 677056 579466
rect 676815 579461 676926 579464
rect 677050 579462 677056 579464
rect 677120 579462 677126 579526
rect 677242 579462 677248 579526
rect 677312 579462 677318 579526
rect 676866 579198 676926 579461
rect 42682 578870 42688 578934
rect 42752 578932 42758 578934
rect 43066 578932 43072 578934
rect 42752 578872 43072 578932
rect 42752 578870 42758 578872
rect 43066 578870 43072 578872
rect 43136 578870 43142 578934
rect 675514 578870 675520 578934
rect 675584 578870 675590 578934
rect 675522 578606 675582 578870
rect 42063 578488 42129 578491
rect 42874 578488 42880 578490
rect 42063 578486 42880 578488
rect 42063 578430 42068 578486
rect 42124 578430 42880 578486
rect 42063 578428 42880 578430
rect 42063 578425 42129 578428
rect 42874 578426 42880 578428
rect 42944 578426 42950 578490
rect 676282 578426 676288 578490
rect 676352 578426 676358 578490
rect 42298 578278 42304 578342
rect 42368 578340 42374 578342
rect 42927 578340 42993 578343
rect 42368 578338 42993 578340
rect 42368 578282 42932 578338
rect 42988 578282 42993 578338
rect 42368 578280 42993 578282
rect 42368 578278 42374 578280
rect 42927 578277 42993 578280
rect 676290 578162 676350 578426
rect 654447 577896 654513 577899
rect 650208 577894 654513 577896
rect 650208 577838 654452 577894
rect 654508 577838 654513 577894
rect 650208 577836 654513 577838
rect 654447 577833 654513 577836
rect 675130 577834 675136 577898
rect 675200 577834 675206 577898
rect 42159 577600 42225 577603
rect 42490 577600 42496 577602
rect 42159 577598 42496 577600
rect 42159 577542 42164 577598
rect 42220 577542 42496 577598
rect 42159 577540 42496 577542
rect 42159 577537 42225 577540
rect 42490 577538 42496 577540
rect 42560 577538 42566 577602
rect 675138 577570 675198 577834
rect 675706 577242 675712 577306
rect 675776 577242 675782 577306
rect 675714 576978 675774 577242
rect 673978 576502 673984 576566
rect 674048 576564 674054 576566
rect 674048 576504 674784 576564
rect 674048 576502 674054 576504
rect 676090 576206 676096 576270
rect 676160 576206 676166 576270
rect 676098 575942 676158 576206
rect 674362 575318 674368 575382
rect 674432 575380 674438 575382
rect 674432 575320 674784 575380
rect 674432 575318 674438 575320
rect 674938 575170 674944 575234
rect 675008 575170 675014 575234
rect 42063 574936 42129 574939
rect 42682 574936 42688 574938
rect 42063 574934 42688 574936
rect 42063 574878 42068 574934
rect 42124 574878 42688 574934
rect 42063 574876 42688 574878
rect 42063 574873 42129 574876
rect 42682 574874 42688 574876
rect 42752 574874 42758 574938
rect 674946 574906 675006 575170
rect 42063 574642 42129 574643
rect 41530 574578 41536 574642
rect 41600 574578 41606 574642
rect 42063 574638 42112 574642
rect 42176 574640 42182 574642
rect 42063 574582 42068 574638
rect 42063 574578 42112 574582
rect 42176 574580 42220 574640
rect 42176 574578 42182 574580
rect 41538 574494 41598 574578
rect 42063 574577 42129 574578
rect 41530 574430 41536 574494
rect 41600 574492 41606 574494
rect 41775 574492 41841 574495
rect 41600 574490 41841 574492
rect 41600 574434 41780 574490
rect 41836 574434 41841 574490
rect 41600 574432 41841 574434
rect 41600 574430 41606 574432
rect 41775 574429 41841 574432
rect 673263 574344 673329 574347
rect 673263 574342 674784 574344
rect 673263 574286 673268 574342
rect 673324 574286 674784 574342
rect 673263 574284 674784 574286
rect 673263 574281 673329 574284
rect 41775 574050 41841 574051
rect 41722 574048 41728 574050
rect 41684 573988 41728 574048
rect 41792 574046 41841 574050
rect 41836 573990 41841 574046
rect 41722 573986 41728 573988
rect 41792 573986 41841 573990
rect 41775 573985 41841 573986
rect 673839 573752 673905 573755
rect 673839 573750 674784 573752
rect 673839 573694 673844 573750
rect 673900 573694 674784 573750
rect 673839 573692 674784 573694
rect 673839 573689 673905 573692
rect 673839 573308 673905 573311
rect 673839 573306 674784 573308
rect 673839 573250 673844 573306
rect 673900 573250 674784 573306
rect 673839 573248 674784 573250
rect 673839 573245 673905 573248
rect 40570 573098 40576 573162
rect 40640 573160 40646 573162
rect 43215 573160 43281 573163
rect 40640 573158 43281 573160
rect 40640 573102 43220 573158
rect 43276 573102 43281 573158
rect 40640 573100 43281 573102
rect 40640 573098 40646 573100
rect 43215 573097 43281 573100
rect 59535 573012 59601 573015
rect 59535 573010 64416 573012
rect 59535 572954 59540 573010
rect 59596 572954 64416 573010
rect 59535 572952 64416 572954
rect 59535 572949 59601 572952
rect 673743 572716 673809 572719
rect 673743 572714 674784 572716
rect 673743 572658 673748 572714
rect 673804 572658 674784 572714
rect 673743 572656 674784 572658
rect 673743 572653 673809 572656
rect 673839 572124 673905 572127
rect 673839 572122 674784 572124
rect 673839 572066 673844 572122
rect 673900 572066 674784 572122
rect 673839 572064 674784 572066
rect 673839 572061 673905 572064
rect 674415 571606 674481 571609
rect 674415 571604 674784 571606
rect 674415 571548 674420 571604
rect 674476 571548 674784 571604
rect 674415 571546 674784 571548
rect 674415 571543 674481 571546
rect 677058 570795 677118 571058
rect 677007 570790 677118 570795
rect 677007 570734 677012 570790
rect 677068 570734 677118 570790
rect 677007 570732 677118 570734
rect 677007 570729 677073 570732
rect 40762 570434 40768 570498
rect 40832 570496 40838 570498
rect 41775 570496 41841 570499
rect 40832 570494 41841 570496
rect 40832 570438 41780 570494
rect 41836 570438 41841 570494
rect 40832 570436 41841 570438
rect 40832 570434 40838 570436
rect 41775 570433 41841 570436
rect 676866 570203 676926 570466
rect 676815 570198 676926 570203
rect 676815 570142 676820 570198
rect 676876 570142 676926 570198
rect 676815 570140 676926 570142
rect 676815 570137 676881 570140
rect 676815 569756 676881 569759
rect 676815 569754 676926 569756
rect 676815 569698 676820 569754
rect 676876 569698 676926 569754
rect 676815 569693 676926 569698
rect 676866 569430 676926 569693
rect 677058 569611 677118 569948
rect 677007 569606 677118 569611
rect 677007 569550 677012 569606
rect 677068 569550 677118 569606
rect 677007 569548 677118 569550
rect 677007 569545 677073 569548
rect 654447 566204 654513 566207
rect 650208 566202 654513 566204
rect 650208 566146 654452 566202
rect 654508 566146 654513 566202
rect 650208 566144 654513 566146
rect 654447 566141 654513 566144
rect 41530 564958 41536 565022
rect 41600 565020 41606 565022
rect 41722 565020 41728 565022
rect 41600 564960 41728 565020
rect 41600 564958 41606 564960
rect 41722 564958 41728 564960
rect 41792 564958 41798 565022
rect 674362 562590 674368 562654
rect 674432 562652 674438 562654
rect 675471 562652 675537 562655
rect 674432 562650 675537 562652
rect 674432 562594 675476 562650
rect 675532 562594 675537 562650
rect 674432 562592 675537 562594
rect 674432 562590 674438 562592
rect 675471 562589 675537 562592
rect 675471 561766 675537 561767
rect 675471 561762 675520 561766
rect 675584 561764 675590 561766
rect 675471 561706 675476 561762
rect 675471 561702 675520 561706
rect 675584 561704 675628 561764
rect 675584 561702 675590 561704
rect 675471 561701 675537 561702
rect 675130 561406 675136 561470
rect 675200 561468 675206 561470
rect 675375 561468 675441 561471
rect 675200 561466 675441 561468
rect 675200 561410 675380 561466
rect 675436 561410 675441 561466
rect 675200 561408 675441 561410
rect 675200 561406 675206 561408
rect 675375 561405 675441 561408
rect 42498 559692 42558 559810
rect 42831 559692 42897 559695
rect 42498 559690 42897 559692
rect 42498 559634 42836 559690
rect 42892 559634 42897 559690
rect 42498 559632 42897 559634
rect 42831 559629 42897 559632
rect 43023 559396 43089 559399
rect 42528 559394 43089 559396
rect 42528 559338 43028 559394
rect 43084 559338 43089 559394
rect 42528 559336 43089 559338
rect 43023 559333 43089 559336
rect 40186 559038 40192 559102
rect 40256 559100 40262 559102
rect 43503 559100 43569 559103
rect 40256 559098 43569 559100
rect 40256 559042 43508 559098
rect 43564 559042 43569 559098
rect 40256 559040 43569 559042
rect 40256 559038 40262 559040
rect 43503 559037 43569 559040
rect 59535 558952 59601 558955
rect 59535 558950 64416 558952
rect 59535 558894 59540 558950
rect 59596 558894 64416 558950
rect 59535 558892 64416 558894
rect 59535 558889 59601 558892
rect 674938 558890 674944 558954
rect 675008 558952 675014 558954
rect 675471 558952 675537 558955
rect 675008 558950 675537 558952
rect 675008 558894 675476 558950
rect 675532 558894 675537 558950
rect 675008 558892 675537 558894
rect 675008 558890 675014 558892
rect 675471 558889 675537 558892
rect 42927 558804 42993 558807
rect 42528 558802 42993 558804
rect 42528 558746 42932 558802
rect 42988 558746 42993 558802
rect 42528 558744 42993 558746
rect 42927 558741 42993 558744
rect 43695 558508 43761 558511
rect 42306 558506 43761 558508
rect 42306 558450 43700 558506
rect 43756 558450 43761 558506
rect 42306 558448 43761 558450
rect 42306 558182 42366 558448
rect 43695 558445 43761 558448
rect 43983 558064 44049 558067
rect 42498 558062 44049 558064
rect 42498 558006 43988 558062
rect 44044 558006 44049 558062
rect 42498 558004 44049 558006
rect 42498 557738 42558 558004
rect 43983 558001 44049 558004
rect 43407 557176 43473 557179
rect 43791 557176 43857 557179
rect 42528 557174 43857 557176
rect 42528 557118 43412 557174
rect 43468 557118 43796 557174
rect 43852 557118 43857 557174
rect 42528 557116 43857 557118
rect 43407 557113 43473 557116
rect 43791 557113 43857 557116
rect 40186 556818 40192 556882
rect 40256 556818 40262 556882
rect 40194 556554 40254 556818
rect 41538 555847 41598 556110
rect 41538 555842 41649 555847
rect 41538 555786 41588 555842
rect 41644 555786 41649 555842
rect 41538 555784 41649 555786
rect 41583 555781 41649 555784
rect 41922 555255 41982 555518
rect 41871 555250 41982 555255
rect 41871 555194 41876 555250
rect 41932 555194 41982 555250
rect 41871 555192 41982 555194
rect 41871 555189 41937 555192
rect 40770 554662 40830 554926
rect 40762 554598 40768 554662
rect 40832 554598 40838 554662
rect 654447 554512 654513 554515
rect 650208 554510 654513 554512
rect 41538 554071 41598 554482
rect 650208 554454 654452 554510
rect 654508 554454 654513 554510
rect 650208 554452 654513 554454
rect 654447 554449 654513 554452
rect 675759 554512 675825 554515
rect 676858 554512 676864 554514
rect 675759 554510 676864 554512
rect 675759 554454 675764 554510
rect 675820 554454 676864 554510
rect 675759 554452 676864 554454
rect 675759 554449 675825 554452
rect 676858 554450 676864 554452
rect 676928 554450 676934 554514
rect 41487 554066 41598 554071
rect 41487 554010 41492 554066
rect 41548 554010 41598 554066
rect 41487 554008 41598 554010
rect 41487 554005 41553 554008
rect 42114 553627 42174 553890
rect 42114 553622 42225 553627
rect 42114 553566 42164 553622
rect 42220 553566 42225 553622
rect 42114 553564 42225 553566
rect 42159 553561 42225 553564
rect 42498 553035 42558 553298
rect 42447 553030 42558 553035
rect 42447 552974 42452 553030
rect 42508 552974 42558 553030
rect 42447 552972 42558 552974
rect 42447 552969 42513 552972
rect 40962 552442 41022 552854
rect 40954 552378 40960 552442
rect 41024 552378 41030 552442
rect 41922 551999 41982 552262
rect 41922 551994 42033 551999
rect 41922 551938 41972 551994
rect 42028 551938 42033 551994
rect 41922 551936 42033 551938
rect 41967 551933 42033 551936
rect 41730 551407 41790 551670
rect 41730 551402 41841 551407
rect 41730 551346 41780 551402
rect 41836 551346 41841 551402
rect 41730 551344 41841 551346
rect 41775 551341 41841 551344
rect 42498 550812 42558 551152
rect 43119 550812 43185 550815
rect 42498 550810 43185 550812
rect 42498 550754 43124 550810
rect 43180 550754 43185 550810
rect 42498 550752 43185 550754
rect 43119 550749 43185 550752
rect 42114 550371 42174 550634
rect 42063 550366 42174 550371
rect 42063 550310 42068 550366
rect 42124 550310 42174 550366
rect 42063 550308 42174 550310
rect 42063 550305 42129 550308
rect 41346 549779 41406 550042
rect 41346 549774 41457 549779
rect 41346 549718 41396 549774
rect 41452 549718 41457 549774
rect 41346 549716 41457 549718
rect 41391 549713 41457 549716
rect 41730 549187 41790 549524
rect 41679 549182 41790 549187
rect 41679 549126 41684 549182
rect 41740 549126 41790 549182
rect 41679 549124 41790 549126
rect 41679 549121 41745 549124
rect 43119 549036 43185 549039
rect 42528 549034 43185 549036
rect 42528 548978 43124 549034
rect 43180 548978 43185 549034
rect 42528 548976 43185 548978
rect 43119 548973 43185 548976
rect 42498 548148 42558 548414
rect 42498 548088 42750 548148
rect 35202 547559 35262 547896
rect 42690 547704 42750 548088
rect 35151 547554 35262 547559
rect 35151 547498 35156 547554
rect 35212 547498 35262 547554
rect 35151 547496 35262 547498
rect 42498 547644 42750 547704
rect 35151 547493 35217 547496
rect 42498 547408 42558 547644
rect 44559 547408 44625 547411
rect 42498 547406 44625 547408
rect 42498 547378 44564 547406
rect 42528 547350 44564 547378
rect 44620 547350 44625 547406
rect 42528 547348 44625 547350
rect 44559 547345 44625 547348
rect 35151 547112 35217 547115
rect 35151 547110 35262 547112
rect 35151 547054 35156 547110
rect 35212 547054 35262 547110
rect 35151 547049 35262 547054
rect 35202 546786 35262 547049
rect 42682 544596 42688 544598
rect 42114 544536 42688 544596
rect 42114 544450 42174 544536
rect 42682 544534 42688 544536
rect 42752 544534 42758 544598
rect 42106 544386 42112 544450
rect 42176 544386 42182 544450
rect 59535 544448 59601 544451
rect 59535 544446 64416 544448
rect 59535 544390 59540 544446
rect 59596 544390 64416 544446
rect 59535 544388 64416 544390
rect 59535 544385 59601 544388
rect 654447 542672 654513 542675
rect 650208 542670 654513 542672
rect 650208 542614 654452 542670
rect 654508 542614 654513 542670
rect 650208 542612 654513 542614
rect 654447 542609 654513 542612
rect 42874 541574 42880 541638
rect 42944 541636 42950 541638
rect 43023 541636 43089 541639
rect 42944 541634 43089 541636
rect 42944 541578 43028 541634
rect 43084 541578 43089 541634
rect 42944 541576 43089 541578
rect 42944 541574 42950 541576
rect 43023 541573 43089 541576
rect 41487 541488 41553 541491
rect 43066 541488 43072 541490
rect 41487 541486 43072 541488
rect 41487 541430 41492 541486
rect 41548 541430 43072 541486
rect 41487 541428 43072 541430
rect 41487 541425 41553 541428
rect 43066 541426 43072 541428
rect 43136 541426 43142 541490
rect 41391 541342 41457 541343
rect 41338 541340 41344 541342
rect 41300 541280 41344 541340
rect 41408 541338 41457 541342
rect 41452 541282 41457 541338
rect 41338 541278 41344 541280
rect 41408 541278 41457 541282
rect 41391 541277 41457 541278
rect 41679 541342 41745 541343
rect 41679 541338 41728 541342
rect 41792 541340 41798 541342
rect 41679 541282 41684 541338
rect 41679 541278 41728 541282
rect 41792 541280 41836 541340
rect 41792 541278 41798 541280
rect 41679 541277 41745 541278
rect 41914 541130 41920 541194
rect 41984 541192 41990 541194
rect 42159 541192 42225 541195
rect 41984 541190 42225 541192
rect 41984 541134 42164 541190
rect 42220 541134 42225 541190
rect 41984 541132 42225 541134
rect 41984 541130 41990 541132
rect 42159 541129 42225 541132
rect 41775 541044 41841 541047
rect 42298 541044 42304 541046
rect 41775 541042 42304 541044
rect 41775 540986 41780 541042
rect 41836 540986 42304 541042
rect 41775 540984 42304 540986
rect 41775 540981 41841 540984
rect 42298 540982 42304 540984
rect 42368 540982 42374 541046
rect 42298 538022 42304 538086
rect 42368 538084 42374 538086
rect 43023 538084 43089 538087
rect 42368 538082 43089 538084
rect 42368 538026 43028 538082
rect 43084 538026 43089 538082
rect 42368 538024 43089 538026
rect 42368 538022 42374 538024
rect 43023 538021 43089 538024
rect 676866 537199 676926 537462
rect 674799 537196 674865 537199
rect 674754 537194 674865 537196
rect 674754 537138 674804 537194
rect 674860 537138 674865 537194
rect 674754 537133 674865 537138
rect 676815 537194 676926 537199
rect 676815 537138 676820 537194
rect 676876 537138 676926 537194
rect 676815 537136 676926 537138
rect 676815 537133 676881 537136
rect 42063 537048 42129 537051
rect 42874 537048 42880 537050
rect 42063 537046 42880 537048
rect 42063 536990 42068 537046
rect 42124 536990 42880 537046
rect 42063 536988 42880 536990
rect 42063 536985 42129 536988
rect 42874 536986 42880 536988
rect 42944 536986 42950 537050
rect 674754 536870 674814 537133
rect 674799 536604 674865 536607
rect 674754 536602 674865 536604
rect 674754 536546 674804 536602
rect 674860 536546 674865 536602
rect 674754 536541 674865 536546
rect 674754 536426 674814 536541
rect 674799 536160 674865 536163
rect 674754 536158 674865 536160
rect 674754 536102 674804 536158
rect 674860 536102 674865 536158
rect 674754 536097 674865 536102
rect 674754 535834 674814 536097
rect 677250 535127 677310 535242
rect 677250 535122 677361 535127
rect 677250 535066 677300 535122
rect 677356 535066 677361 535122
rect 677250 535064 677361 535066
rect 677295 535061 677361 535064
rect 677242 534914 677248 534978
rect 677312 534914 677318 534978
rect 677250 534828 677310 534914
rect 677250 534798 677472 534828
rect 677280 534768 677502 534798
rect 677442 534535 677502 534768
rect 677050 534470 677056 534534
rect 677120 534470 677126 534534
rect 677391 534530 677502 534535
rect 677391 534474 677396 534530
rect 677452 534474 677502 534530
rect 677391 534472 677502 534474
rect 41775 534386 41841 534387
rect 41722 534322 41728 534386
rect 41792 534384 41841 534386
rect 41792 534382 41884 534384
rect 41836 534326 41884 534382
rect 41792 534324 41884 534326
rect 41792 534322 41841 534324
rect 41775 534321 41841 534322
rect 677058 534236 677118 534470
rect 677391 534469 677457 534472
rect 676896 534206 677118 534236
rect 676866 534176 677088 534206
rect 676866 533943 676926 534176
rect 675322 533878 675328 533942
rect 675392 533878 675398 533942
rect 676866 533938 676977 533943
rect 676866 533882 676916 533938
rect 676972 533882 676977 533938
rect 676866 533880 676977 533882
rect 41967 533794 42033 533795
rect 41914 533730 41920 533794
rect 41984 533792 42033 533794
rect 41984 533790 42076 533792
rect 42028 533734 42076 533790
rect 41984 533732 42076 533734
rect 41984 533730 42033 533732
rect 41967 533729 42033 533730
rect 675330 533614 675390 533878
rect 676911 533877 676977 533880
rect 676666 533434 676672 533498
rect 676736 533434 676742 533498
rect 676674 533170 676734 533434
rect 42063 532758 42129 532759
rect 42063 532756 42112 532758
rect 42020 532754 42112 532756
rect 42020 532698 42068 532754
rect 42020 532696 42112 532698
rect 42063 532694 42112 532696
rect 42176 532694 42182 532758
rect 42063 532693 42129 532694
rect 40954 532546 40960 532610
rect 41024 532608 41030 532610
rect 42927 532608 42993 532611
rect 41024 532606 42993 532608
rect 41024 532550 42932 532606
rect 42988 532550 42993 532606
rect 41024 532548 42993 532550
rect 41024 532546 41030 532548
rect 42927 532545 42993 532548
rect 674170 532546 674176 532610
rect 674240 532608 674246 532610
rect 674240 532548 674784 532608
rect 674240 532546 674246 532548
rect 674554 532250 674560 532314
rect 674624 532312 674630 532314
rect 674624 532252 674814 532312
rect 674624 532250 674630 532252
rect 674754 531986 674814 532252
rect 41775 531870 41841 531871
rect 41722 531806 41728 531870
rect 41792 531868 41841 531870
rect 41792 531866 41884 531868
rect 41836 531810 41884 531866
rect 41792 531808 41884 531810
rect 41792 531806 41841 531808
rect 675898 531806 675904 531870
rect 675968 531806 675974 531870
rect 41775 531805 41841 531806
rect 675906 531542 675966 531806
rect 41338 531214 41344 531278
rect 41408 531276 41414 531278
rect 41775 531276 41841 531279
rect 41408 531274 41841 531276
rect 41408 531218 41780 531274
rect 41836 531218 41841 531274
rect 41408 531216 41841 531218
rect 41408 531214 41414 531216
rect 41775 531213 41841 531216
rect 676474 531214 676480 531278
rect 676544 531214 676550 531278
rect 654063 530980 654129 530983
rect 650208 530978 654129 530980
rect 650208 530922 654068 530978
rect 654124 530922 654129 530978
rect 676482 530950 676542 531214
rect 650208 530920 654129 530922
rect 654063 530917 654129 530920
rect 674746 530622 674752 530686
rect 674816 530622 674822 530686
rect 674754 530358 674814 530622
rect 40762 530030 40768 530094
rect 40832 530092 40838 530094
rect 43023 530092 43089 530095
rect 40832 530090 43089 530092
rect 40832 530034 43028 530090
rect 43084 530034 43089 530090
rect 40832 530032 43089 530034
rect 40832 530030 40838 530032
rect 43023 530029 43089 530032
rect 59535 530092 59601 530095
rect 59535 530090 64416 530092
rect 59535 530034 59540 530090
rect 59596 530034 64416 530090
rect 59535 530032 64416 530034
rect 59535 530029 59601 530032
rect 673647 529944 673713 529947
rect 673647 529942 674814 529944
rect 673647 529886 673652 529942
rect 673708 529886 674814 529942
rect 673647 529884 674814 529886
rect 673647 529881 673713 529884
rect 674754 529840 674814 529884
rect 42159 529500 42225 529503
rect 43066 529500 43072 529502
rect 42159 529498 43072 529500
rect 42159 529442 42164 529498
rect 42220 529442 43072 529498
rect 42159 529440 43072 529442
rect 42159 529437 42225 529440
rect 43066 529438 43072 529440
rect 43136 529438 43142 529502
rect 673551 529352 673617 529355
rect 673551 529350 674784 529352
rect 673551 529294 673556 529350
rect 673612 529294 674784 529350
rect 673551 529292 674784 529294
rect 673551 529289 673617 529292
rect 674799 529056 674865 529059
rect 674754 529054 674865 529056
rect 674754 528998 674804 529054
rect 674860 528998 674865 529054
rect 674754 528993 674865 528998
rect 674754 528730 674814 528993
rect 674799 528464 674865 528467
rect 674754 528462 674865 528464
rect 674754 528406 674804 528462
rect 674860 528406 674865 528462
rect 674754 528401 674865 528406
rect 674754 528212 674814 528401
rect 673359 527724 673425 527727
rect 673359 527722 674784 527724
rect 673359 527666 673364 527722
rect 673420 527666 674784 527722
rect 673359 527664 674784 527666
rect 673359 527661 673425 527664
rect 673071 527132 673137 527135
rect 673071 527130 674784 527132
rect 673071 527074 673076 527130
rect 673132 527074 674784 527130
rect 673071 527072 674784 527074
rect 673071 527069 673137 527072
rect 673167 526688 673233 526691
rect 673167 526686 674814 526688
rect 673167 526630 673172 526686
rect 673228 526630 674814 526686
rect 673167 526628 674814 526630
rect 673167 526625 673233 526628
rect 674754 526584 674814 526628
rect 677058 525803 677118 526066
rect 677007 525798 677118 525803
rect 677007 525742 677012 525798
rect 677068 525742 677118 525798
rect 677007 525740 677118 525742
rect 677007 525737 677073 525740
rect 676866 525211 676926 525474
rect 676815 525206 676926 525211
rect 676815 525150 676820 525206
rect 676876 525150 676926 525206
rect 676815 525148 676926 525150
rect 677007 525208 677073 525211
rect 677007 525206 677118 525208
rect 677007 525150 677012 525206
rect 677068 525150 677118 525206
rect 676815 525145 676881 525148
rect 677007 525145 677118 525150
rect 677058 524956 677118 525145
rect 676815 524764 676881 524767
rect 676815 524762 676926 524764
rect 676815 524706 676820 524762
rect 676876 524706 676926 524762
rect 676815 524701 676926 524706
rect 676866 524438 676926 524701
rect 43119 524172 43185 524175
rect 43311 524172 43377 524175
rect 43119 524170 43377 524172
rect 43119 524114 43124 524170
rect 43180 524114 43316 524170
rect 43372 524114 43377 524170
rect 43119 524112 43377 524114
rect 43119 524109 43185 524112
rect 43311 524109 43377 524112
rect 654447 519288 654513 519291
rect 650208 519286 654513 519288
rect 650208 519230 654452 519286
rect 654508 519230 654513 519286
rect 650208 519228 654513 519230
rect 654447 519225 654513 519228
rect 59535 515736 59601 515739
rect 59535 515734 64416 515736
rect 59535 515678 59540 515734
rect 59596 515678 64416 515734
rect 59535 515676 64416 515678
rect 59535 515673 59601 515676
rect 42159 509964 42225 509967
rect 42298 509964 42304 509966
rect 42159 509962 42304 509964
rect 42159 509906 42164 509962
rect 42220 509906 42304 509962
rect 42159 509904 42304 509906
rect 42159 509901 42225 509904
rect 42298 509902 42304 509904
rect 42368 509902 42374 509966
rect 654447 507448 654513 507451
rect 650208 507446 654513 507448
rect 650208 507390 654452 507446
rect 654508 507390 654513 507446
rect 650208 507388 654513 507390
rect 654447 507385 654513 507388
rect 42159 504046 42225 504047
rect 42106 504044 42112 504046
rect 42068 503984 42112 504044
rect 42176 504042 42225 504046
rect 42220 503986 42225 504042
rect 42106 503982 42112 503984
rect 42176 503982 42225 503986
rect 42159 503981 42225 503982
rect 59535 501232 59601 501235
rect 59535 501230 64416 501232
rect 59535 501174 59540 501230
rect 59596 501174 64416 501230
rect 59535 501172 64416 501174
rect 59535 501169 59601 501172
rect 654351 495756 654417 495759
rect 650208 495754 654417 495756
rect 650208 495698 654356 495754
rect 654412 495698 654417 495754
rect 650208 495696 654417 495698
rect 654351 495693 654417 495696
rect 674946 493243 675006 493506
rect 674895 493238 675006 493243
rect 674895 493182 674900 493238
rect 674956 493182 675006 493238
rect 674895 493180 675006 493182
rect 675087 493240 675153 493243
rect 675087 493238 675198 493240
rect 675087 493182 675092 493238
rect 675148 493182 675198 493238
rect 674895 493177 674961 493180
rect 675087 493177 675198 493182
rect 675138 492914 675198 493177
rect 673839 492352 673905 492355
rect 673839 492350 674784 492352
rect 673839 492294 673844 492350
rect 673900 492294 674784 492350
rect 673839 492292 674784 492294
rect 673839 492289 673905 492292
rect 677295 492204 677361 492207
rect 677250 492202 677361 492204
rect 677250 492146 677300 492202
rect 677356 492146 677361 492202
rect 677250 492141 677361 492146
rect 677250 491878 677310 492141
rect 677442 491023 677502 491286
rect 677391 491018 677502 491023
rect 677391 490962 677396 491018
rect 677452 490962 677502 491018
rect 677391 490960 677502 490962
rect 677391 490957 677457 490960
rect 677250 490579 677310 490694
rect 677199 490574 677310 490579
rect 677199 490518 677204 490574
rect 677260 490518 677310 490574
rect 677199 490516 677310 490518
rect 677199 490513 677265 490516
rect 676866 489987 676926 490250
rect 675130 489922 675136 489986
rect 675200 489922 675206 489986
rect 676866 489982 676977 489987
rect 676866 489926 676916 489982
rect 676972 489926 676977 489982
rect 676866 489924 676977 489926
rect 42106 489626 42112 489690
rect 42176 489626 42182 489690
rect 675138 489658 675198 489922
rect 676911 489921 676977 489924
rect 42114 489392 42174 489626
rect 42298 489392 42304 489394
rect 42114 489332 42304 489392
rect 42298 489330 42304 489332
rect 42368 489330 42374 489394
rect 674511 489392 674577 489395
rect 674511 489390 674814 489392
rect 674511 489334 674516 489390
rect 674572 489334 674814 489390
rect 674511 489332 674814 489334
rect 674511 489329 674577 489332
rect 674754 489066 674814 489332
rect 674362 488590 674368 488654
rect 674432 488652 674438 488654
rect 674432 488592 674784 488652
rect 674432 488590 674438 488592
rect 674223 488060 674289 488063
rect 674223 488058 674784 488060
rect 674223 488002 674228 488058
rect 674284 488002 674784 488058
rect 674223 488000 674784 488002
rect 674223 487997 674289 488000
rect 674415 487468 674481 487471
rect 674415 487466 674784 487468
rect 674415 487410 674420 487466
rect 674476 487410 674784 487466
rect 674415 487408 674784 487410
rect 674415 487405 674481 487408
rect 674607 487172 674673 487175
rect 674607 487170 674814 487172
rect 674607 487114 674612 487170
rect 674668 487114 674814 487170
rect 674607 487112 674814 487114
rect 674607 487109 674673 487112
rect 674754 486994 674814 487112
rect 58575 486876 58641 486879
rect 58575 486874 64416 486876
rect 58575 486818 58580 486874
rect 58636 486818 64416 486874
rect 58575 486816 64416 486818
rect 58575 486813 58641 486816
rect 675514 486666 675520 486730
rect 675584 486666 675590 486730
rect 675522 486402 675582 486666
rect 674938 486074 674944 486138
rect 675008 486074 675014 486138
rect 674946 485810 675006 486074
rect 674799 485544 674865 485547
rect 674754 485542 674865 485544
rect 674754 485486 674804 485542
rect 674860 485486 674865 485542
rect 674754 485481 674865 485486
rect 674754 485366 674814 485481
rect 674319 484804 674385 484807
rect 674319 484802 674784 484804
rect 674319 484746 674324 484802
rect 674380 484746 674784 484802
rect 674319 484744 674784 484746
rect 674319 484741 674385 484744
rect 673263 484212 673329 484215
rect 673263 484210 674784 484212
rect 673263 484154 673268 484210
rect 673324 484154 674784 484210
rect 673263 484152 674784 484154
rect 673263 484149 673329 484152
rect 654255 484064 654321 484067
rect 650208 484062 654321 484064
rect 650208 484006 654260 484062
rect 654316 484006 654321 484062
rect 650208 484004 654321 484006
rect 654255 484001 654321 484004
rect 42063 483768 42129 483771
rect 42298 483768 42304 483770
rect 42063 483766 42304 483768
rect 42063 483710 42068 483766
rect 42124 483710 42304 483766
rect 42063 483708 42304 483710
rect 42063 483705 42129 483708
rect 42298 483706 42304 483708
rect 42368 483706 42374 483770
rect 673743 483768 673809 483771
rect 673743 483766 674814 483768
rect 673743 483710 673748 483766
rect 673804 483710 674814 483766
rect 673743 483708 674814 483710
rect 673743 483705 673809 483708
rect 674754 483664 674814 483708
rect 676858 483410 676864 483474
rect 676928 483410 676934 483474
rect 676866 483146 676926 483410
rect 673839 482584 673905 482587
rect 673839 482582 674784 482584
rect 673839 482526 673844 482582
rect 673900 482526 674784 482582
rect 673839 482524 674784 482526
rect 673839 482521 673905 482524
rect 677058 481699 677118 482036
rect 677007 481694 677118 481699
rect 677007 481638 677012 481694
rect 677068 481638 677118 481694
rect 677007 481636 677118 481638
rect 677007 481633 677073 481636
rect 676866 481255 676926 481518
rect 676815 481250 676926 481255
rect 676815 481194 676820 481250
rect 676876 481194 676926 481250
rect 676815 481192 676926 481194
rect 676815 481189 676881 481192
rect 677058 480811 677118 480926
rect 676815 480808 676881 480811
rect 676815 480806 676926 480808
rect 676815 480750 676820 480806
rect 676876 480750 676926 480806
rect 676815 480745 676926 480750
rect 677007 480806 677118 480811
rect 677007 480750 677012 480806
rect 677068 480750 677118 480806
rect 677007 480748 677118 480750
rect 677007 480745 677073 480748
rect 676866 480408 676926 480745
rect 59535 472520 59601 472523
rect 59535 472518 64416 472520
rect 59535 472462 59540 472518
rect 59596 472462 64416 472518
rect 59535 472460 64416 472462
rect 59535 472457 59601 472460
rect 654447 472224 654513 472227
rect 650208 472222 654513 472224
rect 650208 472166 654452 472222
rect 654508 472166 654513 472222
rect 650208 472164 654513 472166
rect 654447 472161 654513 472164
rect 42063 463936 42129 463939
rect 42063 463934 42174 463936
rect 42063 463878 42068 463934
rect 42124 463878 42174 463934
rect 42063 463873 42174 463878
rect 42114 463790 42174 463873
rect 42106 463726 42112 463790
rect 42176 463726 42182 463790
rect 654447 460532 654513 460535
rect 650208 460530 654513 460532
rect 650208 460474 654452 460530
rect 654508 460474 654513 460530
rect 650208 460472 654513 460474
rect 654447 460469 654513 460472
rect 59535 458164 59601 458167
rect 59535 458162 64416 458164
rect 59535 458106 59540 458162
rect 59596 458106 64416 458162
rect 59535 458104 64416 458106
rect 59535 458101 59601 458104
rect 654351 448840 654417 448843
rect 650208 448838 654417 448840
rect 650208 448782 654356 448838
rect 654412 448782 654417 448838
rect 650208 448780 654417 448782
rect 654351 448777 654417 448780
rect 59535 443808 59601 443811
rect 59535 443806 64416 443808
rect 59535 443750 59540 443806
rect 59596 443750 64416 443806
rect 59535 443748 64416 443750
rect 59535 443745 59601 443748
rect 654447 437000 654513 437003
rect 650208 436998 654513 437000
rect 650208 436942 654452 436998
rect 654508 436942 654513 436998
rect 650208 436940 654513 436942
rect 654447 436937 654513 436940
rect 42831 432264 42897 432267
rect 42528 432262 42897 432264
rect 42528 432206 42836 432262
rect 42892 432206 42897 432262
rect 42528 432204 42897 432206
rect 42831 432201 42897 432204
rect 42543 431968 42609 431971
rect 42498 431966 42609 431968
rect 42498 431910 42548 431966
rect 42604 431910 42609 431966
rect 42498 431905 42609 431910
rect 42498 431716 42558 431905
rect 41871 431376 41937 431379
rect 41871 431374 41982 431376
rect 41871 431318 41876 431374
rect 41932 431318 41982 431374
rect 41871 431313 41982 431318
rect 41922 431198 41982 431313
rect 42927 430636 42993 430639
rect 42528 430634 42993 430636
rect 42528 430578 42932 430634
rect 42988 430578 42993 430634
rect 42528 430576 42993 430578
rect 42927 430573 42993 430576
rect 43215 430192 43281 430195
rect 42498 430190 43281 430192
rect 42498 430134 43220 430190
rect 43276 430134 43281 430190
rect 42498 430132 43281 430134
rect 42498 430088 42558 430132
rect 43215 430129 43281 430132
rect 43119 429748 43185 429751
rect 42498 429746 43185 429748
rect 42498 429690 43124 429746
rect 43180 429690 43185 429746
rect 42498 429688 43185 429690
rect 42498 429600 42558 429688
rect 43119 429685 43185 429688
rect 40416 429570 42558 429600
rect 40386 429540 42528 429570
rect 40386 429306 40446 429540
rect 59535 429452 59601 429455
rect 59535 429450 64416 429452
rect 59535 429394 59540 429450
rect 59596 429394 64416 429450
rect 59535 429392 64416 429394
rect 59535 429389 59601 429392
rect 40378 429242 40384 429306
rect 40448 429242 40454 429306
rect 43503 429008 43569 429011
rect 40608 429006 43569 429008
rect 40608 428978 43508 429006
rect 40578 428950 43508 428978
rect 43564 428950 43569 429006
rect 40578 428948 43569 428950
rect 40578 428714 40638 428948
rect 43503 428945 43569 428948
rect 40570 428650 40576 428714
rect 40640 428650 40646 428714
rect 40770 428122 40830 428460
rect 40762 428058 40768 428122
rect 40832 428058 40838 428122
rect 42498 427679 42558 427942
rect 42498 427674 42609 427679
rect 42498 427618 42548 427674
rect 42604 427618 42609 427674
rect 42498 427616 42609 427618
rect 42543 427613 42609 427616
rect 40962 427086 41022 427350
rect 40954 427022 40960 427086
rect 41024 427022 41030 427086
rect 41346 426494 41406 426832
rect 41338 426430 41344 426494
rect 41408 426430 41414 426494
rect 42114 426050 42174 426314
rect 42106 425986 42112 426050
rect 42176 425986 42182 426050
rect 40194 425459 40254 425722
rect 40194 425454 40305 425459
rect 654447 425456 654513 425459
rect 40194 425398 40244 425454
rect 40300 425398 40305 425454
rect 40194 425396 40305 425398
rect 650208 425454 654513 425456
rect 650208 425398 654452 425454
rect 654508 425398 654513 425454
rect 650208 425396 654513 425398
rect 40239 425393 40305 425396
rect 654447 425393 654513 425396
rect 41154 424866 41214 425204
rect 41146 424802 41152 424866
rect 41216 424802 41222 424866
rect 41538 424422 41598 424686
rect 41530 424358 41536 424422
rect 41600 424358 41606 424422
rect 43119 424124 43185 424127
rect 42528 424122 43185 424124
rect 42528 424066 43124 424122
rect 43180 424066 43185 424122
rect 42528 424064 43185 424066
rect 43119 424061 43185 424064
rect 42306 423387 42366 423576
rect 42306 423382 42417 423387
rect 42306 423326 42356 423382
rect 42412 423326 42417 423382
rect 42306 423324 42417 423326
rect 42351 423321 42417 423324
rect 40002 422795 40062 423058
rect 39951 422790 40062 422795
rect 39951 422734 39956 422790
rect 40012 422734 40062 422790
rect 39951 422732 40062 422734
rect 39951 422729 40017 422732
rect 40194 422203 40254 422466
rect 40143 422198 40254 422203
rect 40143 422142 40148 422198
rect 40204 422142 40254 422198
rect 40143 422140 40254 422142
rect 40143 422137 40209 422140
rect 40002 421611 40062 421874
rect 40002 421606 40113 421611
rect 40002 421550 40052 421606
rect 40108 421550 40113 421606
rect 40002 421548 40113 421550
rect 40047 421545 40113 421548
rect 42927 421460 42993 421463
rect 42528 421458 42993 421460
rect 42528 421402 42932 421458
rect 42988 421402 42993 421458
rect 42528 421400 42993 421402
rect 42927 421397 42993 421400
rect 42498 420572 42558 420838
rect 42498 420512 42750 420572
rect 35202 419983 35262 420246
rect 42690 420128 42750 420512
rect 35151 419978 35262 419983
rect 35151 419922 35156 419978
rect 35212 419922 35262 419978
rect 35151 419920 35262 419922
rect 42498 420068 42750 420128
rect 35151 419917 35217 419920
rect 42498 419539 42558 420068
rect 35151 419536 35217 419539
rect 35151 419534 35262 419536
rect 35151 419478 35156 419534
rect 35212 419478 35262 419534
rect 35151 419473 35262 419478
rect 42447 419534 42558 419539
rect 42447 419478 42452 419534
rect 42508 419478 42558 419534
rect 42447 419476 42558 419478
rect 42447 419473 42513 419476
rect 35202 419210 35262 419473
rect 58383 415096 58449 415099
rect 58383 415094 64416 415096
rect 58383 415038 58388 415094
rect 58444 415038 64416 415094
rect 58383 415036 64416 415038
rect 58383 415033 58449 415036
rect 653871 413616 653937 413619
rect 650208 413614 653937 413616
rect 650208 413558 653876 413614
rect 653932 413558 653937 413614
rect 650208 413556 653937 413558
rect 653871 413553 653937 413556
rect 42298 409262 42304 409326
rect 42368 409324 42374 409326
rect 43023 409324 43089 409327
rect 42368 409322 43089 409324
rect 42368 409266 43028 409322
rect 43084 409266 43089 409322
rect 42368 409264 43089 409266
rect 42368 409262 42374 409264
rect 43023 409261 43089 409264
rect 41914 408966 41920 409030
rect 41984 409028 41990 409030
rect 42490 409028 42496 409030
rect 41984 408968 42496 409028
rect 41984 408966 41990 408968
rect 42490 408966 42496 408968
rect 42560 408966 42566 409030
rect 41914 408818 41920 408882
rect 41984 408880 41990 408882
rect 42490 408880 42496 408882
rect 41984 408820 42496 408880
rect 41984 408818 41990 408820
rect 42490 408818 42496 408820
rect 42560 408818 42566 408882
rect 42351 408142 42417 408143
rect 42298 408078 42304 408142
rect 42368 408140 42417 408142
rect 42368 408138 42460 408140
rect 42412 408082 42460 408138
rect 42368 408080 42460 408082
rect 42368 408078 42417 408080
rect 42351 408077 42417 408078
rect 42063 406070 42129 406071
rect 42063 406066 42112 406070
rect 42176 406068 42182 406070
rect 42063 406010 42068 406066
rect 42063 406006 42112 406010
rect 42176 406008 42220 406068
rect 42176 406006 42182 406008
rect 42063 406005 42129 406006
rect 674703 405476 674769 405479
rect 674703 405474 674814 405476
rect 674703 405418 674708 405474
rect 674764 405418 674814 405474
rect 674703 405413 674814 405418
rect 674754 405298 674814 405413
rect 673839 404736 673905 404739
rect 673839 404734 674784 404736
rect 673839 404678 673844 404734
rect 673900 404678 674784 404734
rect 673839 404676 674784 404678
rect 673839 404673 673905 404676
rect 674703 404440 674769 404443
rect 674703 404438 674814 404440
rect 674703 404382 674708 404438
rect 674764 404382 674814 404438
rect 674703 404377 674814 404382
rect 42063 404294 42129 404295
rect 42063 404292 42112 404294
rect 42020 404290 42112 404292
rect 42020 404234 42068 404290
rect 42020 404232 42112 404234
rect 42063 404230 42112 404232
rect 42176 404230 42182 404294
rect 42063 404229 42129 404230
rect 674754 404188 674814 404377
rect 677391 403996 677457 403999
rect 677391 403994 677502 403996
rect 677391 403938 677396 403994
rect 677452 403938 677502 403994
rect 677391 403933 677502 403938
rect 41775 403850 41841 403851
rect 41722 403786 41728 403850
rect 41792 403848 41841 403850
rect 41792 403846 41884 403848
rect 41836 403790 41884 403846
rect 41792 403788 41884 403790
rect 41792 403786 41841 403788
rect 41775 403785 41841 403786
rect 677442 403670 677502 403933
rect 673839 403108 673905 403111
rect 673839 403106 674784 403108
rect 673839 403050 673844 403106
rect 673900 403050 674784 403106
rect 673839 403048 674784 403050
rect 673839 403045 673905 403048
rect 677199 402812 677265 402815
rect 677199 402810 677310 402812
rect 677199 402754 677204 402810
rect 677260 402754 677310 402810
rect 677199 402749 677310 402754
rect 41530 402602 41536 402666
rect 41600 402664 41606 402666
rect 41775 402664 41841 402667
rect 41600 402662 41841 402664
rect 41600 402606 41780 402662
rect 41836 402606 41841 402662
rect 41600 402604 41841 402606
rect 41600 402602 41606 402604
rect 41775 402601 41841 402604
rect 677250 402560 677310 402749
rect 676911 402220 676977 402223
rect 676866 402218 676977 402220
rect 676866 402162 676916 402218
rect 676972 402162 676977 402218
rect 676866 402157 676977 402162
rect 676866 402042 676926 402157
rect 41338 401862 41344 401926
rect 41408 401924 41414 401926
rect 41775 401924 41841 401927
rect 41408 401922 41841 401924
rect 41408 401866 41780 401922
rect 41836 401866 41841 401922
rect 41408 401864 41841 401866
rect 41408 401862 41414 401864
rect 41775 401861 41841 401864
rect 654447 401776 654513 401779
rect 650208 401774 654513 401776
rect 650208 401718 654452 401774
rect 654508 401718 654513 401774
rect 650208 401716 654513 401718
rect 654447 401713 654513 401716
rect 675138 401335 675198 401450
rect 675087 401330 675198 401335
rect 675087 401274 675092 401330
rect 675148 401274 675198 401330
rect 675087 401272 675198 401274
rect 675087 401269 675153 401272
rect 57615 400740 57681 400743
rect 57615 400738 64416 400740
rect 57615 400682 57620 400738
rect 57676 400682 64416 400738
rect 57615 400680 64416 400682
rect 57615 400677 57681 400680
rect 674554 400530 674560 400594
rect 674624 400592 674630 400594
rect 674754 400592 674814 400858
rect 674624 400532 674814 400592
rect 674624 400530 674630 400532
rect 675330 400151 675390 400414
rect 40762 400086 40768 400150
rect 40832 400148 40838 400150
rect 41775 400148 41841 400151
rect 40832 400146 41841 400148
rect 40832 400090 41780 400146
rect 41836 400090 41841 400146
rect 40832 400088 41841 400090
rect 675330 400146 675441 400151
rect 675330 400090 675380 400146
rect 675436 400090 675441 400146
rect 675330 400088 675441 400090
rect 40832 400086 40838 400088
rect 41775 400085 41841 400088
rect 675375 400085 675441 400088
rect 674127 399852 674193 399855
rect 674127 399850 674784 399852
rect 674127 399794 674132 399850
rect 674188 399794 674784 399850
rect 674127 399792 674784 399794
rect 674127 399789 674193 399792
rect 41146 399494 41152 399558
rect 41216 399556 41222 399558
rect 41775 399556 41841 399559
rect 41216 399554 41841 399556
rect 41216 399498 41780 399554
rect 41836 399498 41841 399554
rect 41216 399496 41841 399498
rect 41216 399494 41222 399496
rect 41775 399493 41841 399496
rect 674362 399198 674368 399262
rect 674432 399260 674438 399262
rect 674432 399200 674784 399260
rect 674432 399198 674438 399200
rect 40954 398754 40960 398818
rect 41024 398816 41030 398818
rect 41775 398816 41841 398819
rect 41024 398814 41841 398816
rect 41024 398758 41780 398814
rect 41836 398758 41841 398814
rect 41024 398756 41841 398758
rect 41024 398754 41030 398756
rect 41775 398753 41841 398756
rect 674170 398754 674176 398818
rect 674240 398816 674246 398818
rect 674240 398756 674784 398816
rect 674240 398754 674246 398756
rect 675138 397931 675198 398194
rect 675138 397926 675249 397931
rect 675138 397870 675188 397926
rect 675244 397870 675249 397926
rect 675138 397868 675249 397870
rect 675183 397865 675249 397868
rect 674223 397632 674289 397635
rect 674223 397630 674784 397632
rect 674223 397574 674228 397630
rect 674284 397574 674784 397630
rect 674223 397572 674784 397574
rect 674223 397569 674289 397572
rect 674946 396895 675006 397158
rect 674895 396890 675006 396895
rect 674895 396834 674900 396890
rect 674956 396834 675006 396890
rect 674895 396832 675006 396834
rect 674895 396829 674961 396832
rect 673935 396596 674001 396599
rect 673935 396594 674784 396596
rect 673935 396538 673940 396594
rect 673996 396538 674784 396594
rect 673935 396536 674784 396538
rect 673935 396533 674001 396536
rect 674511 395856 674577 395859
rect 674754 395856 674814 395974
rect 674511 395854 674814 395856
rect 674511 395798 674516 395854
rect 674572 395798 674814 395854
rect 674511 395796 674814 395798
rect 674511 395793 674577 395796
rect 674946 395267 675006 395530
rect 674946 395262 675057 395267
rect 674946 395206 674996 395262
rect 675052 395206 675057 395262
rect 674946 395204 675057 395206
rect 674991 395201 675057 395204
rect 674754 394675 674814 394938
rect 674754 394670 674865 394675
rect 674754 394614 674804 394670
rect 674860 394614 674865 394670
rect 674754 394612 674865 394614
rect 674799 394609 674865 394612
rect 674607 394228 674673 394231
rect 674754 394228 674814 394346
rect 674607 394226 674814 394228
rect 674607 394170 674612 394226
rect 674668 394170 674814 394226
rect 674607 394168 674814 394170
rect 674607 394165 674673 394168
rect 677058 393491 677118 393902
rect 677058 393486 677169 393491
rect 677058 393430 677108 393486
rect 677164 393430 677169 393486
rect 677058 393428 677169 393430
rect 677103 393425 677169 393428
rect 676866 393047 676926 393310
rect 676866 393042 676977 393047
rect 677103 393044 677169 393047
rect 676866 392986 676916 393042
rect 676972 392986 676977 393042
rect 676866 392984 676977 392986
rect 676911 392981 676977 392984
rect 677058 393042 677169 393044
rect 677058 392986 677108 393042
rect 677164 392986 677169 393042
rect 677058 392981 677169 392986
rect 677058 392718 677118 392981
rect 676911 392600 676977 392603
rect 676866 392598 676977 392600
rect 676866 392542 676916 392598
rect 676972 392542 676977 392598
rect 676866 392537 676977 392542
rect 676866 392200 676926 392537
rect 654447 390084 654513 390087
rect 650208 390082 654513 390084
rect 650208 390026 654452 390082
rect 654508 390026 654513 390082
rect 650208 390024 654513 390026
rect 654447 390021 654513 390024
rect 42351 389344 42417 389347
rect 42306 389342 42417 389344
rect 42306 389286 42356 389342
rect 42412 389286 42417 389342
rect 42306 389281 42417 389286
rect 42306 389018 42366 389281
rect 42639 388752 42705 388755
rect 42498 388750 42705 388752
rect 42498 388694 42644 388750
rect 42700 388694 42705 388750
rect 42498 388692 42705 388694
rect 42498 388574 42558 388692
rect 42639 388689 42705 388692
rect 42639 388012 42705 388015
rect 42528 388010 42705 388012
rect 42528 387954 42644 388010
rect 42700 387954 42705 388010
rect 42528 387952 42705 387954
rect 42639 387949 42705 387952
rect 42498 387272 42558 387390
rect 43407 387272 43473 387275
rect 42498 387270 43473 387272
rect 42498 387214 43412 387270
rect 43468 387214 43473 387270
rect 42498 387212 43473 387214
rect 43407 387209 43473 387212
rect 42927 387124 42993 387127
rect 42498 387122 42993 387124
rect 42498 387066 42932 387122
rect 42988 387066 42993 387122
rect 42498 387064 42993 387066
rect 42498 386946 42558 387064
rect 42927 387061 42993 387064
rect 59247 386384 59313 386387
rect 59247 386382 64416 386384
rect 40386 386090 40446 386354
rect 59247 386326 59252 386382
rect 59308 386326 64416 386382
rect 59247 386324 64416 386326
rect 59247 386321 59313 386324
rect 40378 386026 40384 386090
rect 40448 386026 40454 386090
rect 40570 386026 40576 386090
rect 40640 386026 40646 386090
rect 40578 385762 40638 386026
rect 40770 384906 40830 385318
rect 40762 384842 40768 384906
rect 40832 384842 40838 384906
rect 42735 384756 42801 384759
rect 42528 384754 42801 384756
rect 42528 384698 42740 384754
rect 42796 384698 42801 384754
rect 42528 384696 42801 384698
rect 42735 384693 42801 384696
rect 40962 383870 41022 384134
rect 40954 383806 40960 383870
rect 41024 383806 41030 383870
rect 41346 383278 41406 383616
rect 41338 383214 41344 383278
rect 41408 383214 41414 383278
rect 41538 382834 41598 383098
rect 41530 382770 41536 382834
rect 41600 382770 41606 382834
rect 42306 382243 42366 382506
rect 42306 382238 42417 382243
rect 42306 382182 42356 382238
rect 42412 382182 42417 382238
rect 42306 382180 42417 382182
rect 42351 382177 42417 382180
rect 41154 381650 41214 381988
rect 41146 381586 41152 381650
rect 41216 381586 41222 381650
rect 42114 381206 42174 381470
rect 42106 381142 42112 381206
rect 42176 381142 42182 381206
rect 40002 380615 40062 380878
rect 39951 380610 40062 380615
rect 39951 380554 39956 380610
rect 40012 380554 40062 380610
rect 39951 380552 40062 380554
rect 39951 380549 40017 380552
rect 40002 380171 40062 380360
rect 40002 380166 40113 380171
rect 40002 380110 40052 380166
rect 40108 380110 40113 380166
rect 40002 380108 40113 380110
rect 40047 380105 40113 380108
rect 42298 380106 42304 380170
rect 42368 380168 42374 380170
rect 42874 380168 42880 380170
rect 42368 380108 42880 380168
rect 42368 380106 42374 380108
rect 42874 380106 42880 380108
rect 42944 380106 42950 380170
rect 43023 379872 43089 379875
rect 42528 379870 43089 379872
rect 42528 379814 43028 379870
rect 43084 379814 43089 379870
rect 42528 379812 43089 379814
rect 43023 379809 43089 379812
rect 42498 378986 42558 379250
rect 42490 378922 42496 378986
rect 42560 378922 42566 378986
rect 674362 378774 674368 378838
rect 674432 378836 674438 378838
rect 675471 378836 675537 378839
rect 674432 378834 675537 378836
rect 674432 378778 675476 378834
rect 675532 378778 675537 378834
rect 674432 378776 675537 378778
rect 674432 378774 674438 378776
rect 675471 378773 675537 378776
rect 40194 378395 40254 378732
rect 654447 378540 654513 378543
rect 650208 378538 654513 378540
rect 650208 378482 654452 378538
rect 654508 378482 654513 378538
rect 650208 378480 654513 378482
rect 654447 378477 654513 378480
rect 40194 378390 40305 378395
rect 40194 378334 40244 378390
rect 40300 378334 40305 378390
rect 40194 378332 40305 378334
rect 40239 378329 40305 378332
rect 42927 378244 42993 378247
rect 42528 378242 42993 378244
rect 42528 378186 42932 378242
rect 42988 378186 42993 378242
rect 42528 378184 42993 378186
rect 42927 378181 42993 378184
rect 42639 377652 42705 377655
rect 42528 377650 42705 377652
rect 42528 377594 42644 377650
rect 42700 377594 42705 377650
rect 42528 377592 42705 377594
rect 42639 377589 42705 377592
rect 35202 376767 35262 377104
rect 35151 376762 35262 376767
rect 35151 376706 35156 376762
rect 35212 376706 35262 376762
rect 35151 376704 35262 376706
rect 35151 376701 35217 376704
rect 42639 376616 42705 376619
rect 42528 376614 42705 376616
rect 42528 376558 42644 376614
rect 42700 376558 42705 376614
rect 42528 376556 42705 376558
rect 42639 376553 42705 376556
rect 35151 376320 35217 376323
rect 35151 376318 35262 376320
rect 35151 376262 35156 376318
rect 35212 376262 35262 376318
rect 35151 376257 35262 376262
rect 35202 375994 35262 376257
rect 675087 374544 675153 374547
rect 675322 374544 675328 374546
rect 675087 374542 675328 374544
rect 675087 374486 675092 374542
rect 675148 374486 675328 374542
rect 675087 374484 675328 374486
rect 675087 374481 675153 374484
rect 675322 374482 675328 374484
rect 675392 374482 675398 374546
rect 673743 374396 673809 374399
rect 676858 374396 676864 374398
rect 673743 374394 676864 374396
rect 673743 374338 673748 374394
rect 673804 374338 676864 374394
rect 673743 374336 676864 374338
rect 673743 374333 673809 374336
rect 676858 374334 676864 374336
rect 676928 374334 676934 374398
rect 675183 374100 675249 374103
rect 675514 374100 675520 374102
rect 675183 374098 675520 374100
rect 675183 374042 675188 374098
rect 675244 374042 675520 374098
rect 675183 374040 675520 374042
rect 675183 374037 675249 374040
rect 675514 374038 675520 374040
rect 675584 374038 675590 374102
rect 674554 373890 674560 373954
rect 674624 373952 674630 373954
rect 675471 373952 675537 373955
rect 674624 373950 675537 373952
rect 674624 373894 675476 373950
rect 675532 373894 675537 373950
rect 674624 373892 675537 373894
rect 674624 373890 674630 373892
rect 675471 373889 675537 373892
rect 673359 373360 673425 373363
rect 677050 373360 677056 373362
rect 673359 373358 677056 373360
rect 673359 373302 673364 373358
rect 673420 373302 677056 373358
rect 673359 373300 677056 373302
rect 673359 373297 673425 373300
rect 677050 373298 677056 373300
rect 677120 373298 677126 373362
rect 674170 371966 674176 372030
rect 674240 372028 674246 372030
rect 675375 372028 675441 372031
rect 674240 372026 675441 372028
rect 674240 371970 675380 372026
rect 675436 371970 675441 372026
rect 674240 371968 675441 371970
rect 674240 371966 674246 371968
rect 675375 371965 675441 371968
rect 59535 371880 59601 371883
rect 59535 371878 64416 371880
rect 59535 371822 59540 371878
rect 59596 371822 64416 371878
rect 59535 371820 64416 371822
rect 59535 371817 59601 371820
rect 42106 368710 42112 368774
rect 42176 368710 42182 368774
rect 42114 368478 42174 368710
rect 42106 368414 42112 368478
rect 42176 368414 42182 368478
rect 654447 366552 654513 366555
rect 650208 366550 654513 366552
rect 650208 366494 654452 366550
rect 654508 366494 654513 366550
rect 650208 366492 654513 366494
rect 654447 366489 654513 366492
rect 41530 362790 41536 362854
rect 41600 362852 41606 362854
rect 41775 362852 41841 362855
rect 41600 362850 41841 362852
rect 41600 362794 41780 362850
rect 41836 362794 41841 362850
rect 41600 362792 41841 362794
rect 41600 362790 41606 362792
rect 41775 362789 41841 362792
rect 42159 361964 42225 361967
rect 42298 361964 42304 361966
rect 42159 361962 42304 361964
rect 42159 361906 42164 361962
rect 42220 361906 42304 361962
rect 42159 361904 42304 361906
rect 42159 361901 42225 361904
rect 42298 361902 42304 361904
rect 42368 361964 42374 361966
rect 42874 361964 42880 361966
rect 42368 361904 42880 361964
rect 42368 361902 42374 361904
rect 42874 361902 42880 361904
rect 42944 361902 42950 361966
rect 42255 361224 42321 361227
rect 42490 361224 42496 361226
rect 42255 361222 42496 361224
rect 42255 361166 42260 361222
rect 42316 361166 42496 361222
rect 42255 361164 42496 361166
rect 42255 361161 42321 361164
rect 42490 361162 42496 361164
rect 42560 361162 42566 361226
rect 41722 360570 41728 360634
rect 41792 360632 41798 360634
rect 42159 360632 42225 360635
rect 42874 360632 42880 360634
rect 41792 360630 42880 360632
rect 41792 360574 42164 360630
rect 42220 360574 42880 360630
rect 41792 360572 42880 360574
rect 41792 360570 41798 360572
rect 42159 360569 42225 360572
rect 42874 360570 42880 360572
rect 42944 360570 42950 360634
rect 674415 360040 674481 360043
rect 674415 360038 674784 360040
rect 674415 359982 674420 360038
rect 674476 359982 674784 360038
rect 674415 359980 674784 359982
rect 674415 359977 674481 359980
rect 674703 359744 674769 359747
rect 674703 359742 674814 359744
rect 674703 359686 674708 359742
rect 674764 359686 674814 359742
rect 674703 359681 674814 359686
rect 674754 359566 674814 359681
rect 42063 359450 42129 359451
rect 42063 359446 42112 359450
rect 42176 359448 42182 359450
rect 42063 359390 42068 359446
rect 42063 359386 42112 359390
rect 42176 359388 42220 359448
rect 42176 359386 42182 359388
rect 42063 359385 42129 359386
rect 674415 359004 674481 359007
rect 674415 359002 674784 359004
rect 674415 358946 674420 359002
rect 674476 358946 674784 359002
rect 674415 358944 674784 358946
rect 674415 358941 674481 358944
rect 41338 358646 41344 358710
rect 41408 358708 41414 358710
rect 41775 358708 41841 358711
rect 41408 358706 41841 358708
rect 41408 358650 41780 358706
rect 41836 358650 41841 358706
rect 41408 358648 41841 358650
rect 41408 358646 41414 358648
rect 41775 358645 41841 358648
rect 673839 358412 673905 358415
rect 673839 358410 674784 358412
rect 673839 358354 673844 358410
rect 673900 358354 674784 358410
rect 673839 358352 674784 358354
rect 673839 358349 673905 358352
rect 59535 357672 59601 357675
rect 677058 357674 677118 357938
rect 59535 357670 64416 357672
rect 59535 357614 59540 357670
rect 59596 357614 64416 357670
rect 59535 357612 64416 357614
rect 59535 357609 59601 357612
rect 677050 357610 677056 357674
rect 677120 357610 677126 357674
rect 677434 357672 677440 357674
rect 677250 357612 677440 357672
rect 677250 357376 677310 357612
rect 677434 357610 677440 357612
rect 677504 357610 677510 357674
rect 676896 357346 677310 357376
rect 676866 357316 677280 357346
rect 676866 357082 676926 357316
rect 676858 357018 676864 357082
rect 676928 357018 676934 357082
rect 40762 356870 40768 356934
rect 40832 356932 40838 356934
rect 41775 356932 41841 356935
rect 40832 356930 41841 356932
rect 40832 356874 41780 356930
rect 41836 356874 41841 356930
rect 40832 356872 41841 356874
rect 40832 356870 40838 356872
rect 41775 356869 41841 356872
rect 677250 356638 677310 356754
rect 677242 356574 677248 356638
rect 677312 356574 677318 356638
rect 41146 356426 41152 356490
rect 41216 356488 41222 356490
rect 41775 356488 41841 356491
rect 41216 356486 41841 356488
rect 41216 356430 41780 356486
rect 41836 356430 41841 356486
rect 41216 356428 41841 356430
rect 41216 356426 41222 356428
rect 41775 356425 41841 356428
rect 674946 356047 675006 356310
rect 674895 356042 675006 356047
rect 674895 355986 674900 356042
rect 674956 355986 675006 356042
rect 674895 355984 675006 355986
rect 674895 355981 674961 355984
rect 674170 355686 674176 355750
rect 674240 355748 674246 355750
rect 674240 355688 674784 355748
rect 674240 355686 674246 355688
rect 40954 355538 40960 355602
rect 41024 355600 41030 355602
rect 41775 355600 41841 355603
rect 41024 355598 41841 355600
rect 41024 355542 41780 355598
rect 41836 355542 41841 355598
rect 41024 355540 41841 355542
rect 41024 355538 41030 355540
rect 41775 355537 41841 355540
rect 675138 355011 675198 355126
rect 675138 355006 675249 355011
rect 675138 354950 675188 355006
rect 675244 354950 675249 355006
rect 675138 354948 675249 354950
rect 675183 354945 675249 354948
rect 655215 354860 655281 354863
rect 650208 354858 655281 354860
rect 650208 354802 655220 354858
rect 655276 354802 655281 354858
rect 650208 354800 655281 354802
rect 655215 354797 655281 354800
rect 674946 354419 675006 354682
rect 674946 354414 675057 354419
rect 674946 354358 674996 354414
rect 675052 354358 675057 354414
rect 674946 354356 675057 354358
rect 674991 354353 675057 354356
rect 673935 354120 674001 354123
rect 673935 354118 674784 354120
rect 673935 354062 673940 354118
rect 673996 354062 674784 354118
rect 673935 354060 674784 354062
rect 673935 354057 674001 354060
rect 677058 353235 677118 353498
rect 677058 353230 677169 353235
rect 677058 353174 677108 353230
rect 677164 353174 677169 353230
rect 677058 353172 677169 353174
rect 677103 353169 677169 353172
rect 675330 352791 675390 353054
rect 675279 352786 675390 352791
rect 675279 352730 675284 352786
rect 675340 352730 675390 352786
rect 675279 352728 675390 352730
rect 675279 352725 675345 352728
rect 675138 352199 675198 352462
rect 675087 352194 675198 352199
rect 675087 352138 675092 352194
rect 675148 352138 675198 352194
rect 675087 352136 675198 352138
rect 675087 352133 675153 352136
rect 674319 351900 674385 351903
rect 674319 351898 674784 351900
rect 674319 351842 674324 351898
rect 674380 351842 674784 351898
rect 674319 351840 674784 351842
rect 674319 351837 674385 351840
rect 676866 351163 676926 351352
rect 676866 351158 676977 351163
rect 676866 351102 676916 351158
rect 676972 351102 676977 351158
rect 676866 351100 676977 351102
rect 676911 351097 676977 351100
rect 674127 350864 674193 350867
rect 674127 350862 674784 350864
rect 674127 350806 674132 350862
rect 674188 350806 674784 350862
rect 674127 350804 674784 350806
rect 674127 350801 674193 350804
rect 674754 350127 674814 350242
rect 674703 350122 674814 350127
rect 674703 350066 674708 350122
rect 674764 350066 674814 350122
rect 674703 350064 674814 350066
rect 674703 350061 674769 350064
rect 674031 349680 674097 349683
rect 674754 349680 674814 349724
rect 674031 349678 674814 349680
rect 674031 349622 674036 349678
rect 674092 349622 674814 349678
rect 674031 349620 674814 349622
rect 674031 349617 674097 349620
rect 674511 348940 674577 348943
rect 674754 348940 674814 349206
rect 674511 348938 674814 348940
rect 674511 348882 674516 348938
rect 674572 348882 674814 348938
rect 674511 348880 674814 348882
rect 674511 348877 674577 348880
rect 677058 348351 677118 348614
rect 677007 348346 677118 348351
rect 677007 348290 677012 348346
rect 677068 348290 677118 348346
rect 677007 348288 677118 348290
rect 677007 348285 677073 348288
rect 676866 347759 676926 348096
rect 676815 347754 676926 347759
rect 676815 347698 676820 347754
rect 676876 347698 676926 347754
rect 676815 347696 676926 347698
rect 676815 347693 676881 347696
rect 677058 347315 677118 347578
rect 676815 347312 676881 347315
rect 676815 347310 676926 347312
rect 676815 347254 676820 347310
rect 676876 347254 676926 347310
rect 676815 347249 676926 347254
rect 677007 347310 677118 347315
rect 677007 347254 677012 347310
rect 677068 347254 677118 347310
rect 677007 347252 677118 347254
rect 677007 347249 677073 347252
rect 676866 346986 676926 347249
rect 42831 345906 42897 345909
rect 42528 345904 42897 345906
rect 42528 345848 42836 345904
rect 42892 345848 42897 345904
rect 42528 345846 42897 345848
rect 42831 345843 42897 345846
rect 42831 345388 42897 345391
rect 42528 345386 42897 345388
rect 42528 345330 42836 345386
rect 42892 345330 42897 345386
rect 42528 345328 42897 345330
rect 42831 345325 42897 345328
rect 676666 345178 676672 345242
rect 676736 345240 676742 345242
rect 677103 345240 677169 345243
rect 676736 345238 677169 345240
rect 676736 345182 677108 345238
rect 677164 345182 677169 345238
rect 676736 345180 677169 345182
rect 676736 345178 676742 345180
rect 677103 345177 677169 345180
rect 42831 344796 42897 344799
rect 42528 344794 42897 344796
rect 42528 344738 42836 344794
rect 42892 344738 42897 344794
rect 42528 344736 42897 344738
rect 42831 344733 42897 344736
rect 42498 344204 42558 344248
rect 43407 344204 43473 344207
rect 42498 344202 43473 344204
rect 42498 344146 43412 344202
rect 43468 344146 43473 344202
rect 42498 344144 43473 344146
rect 43407 344141 43473 344144
rect 676474 344142 676480 344206
rect 676544 344204 676550 344206
rect 676911 344204 676977 344207
rect 676544 344202 676977 344204
rect 676544 344146 676916 344202
rect 676972 344146 676977 344202
rect 676544 344144 676977 344146
rect 676544 344142 676550 344144
rect 676911 344141 676977 344144
rect 43215 343760 43281 343763
rect 42528 343758 43281 343760
rect 42528 343702 43220 343758
rect 43276 343702 43281 343758
rect 42528 343700 43281 343702
rect 43215 343697 43281 343700
rect 58383 343168 58449 343171
rect 654447 343168 654513 343171
rect 58383 343166 64416 343168
rect 40386 343022 40446 343138
rect 58383 343110 58388 343166
rect 58444 343110 64416 343166
rect 58383 343108 64416 343110
rect 650208 343166 654513 343168
rect 650208 343110 654452 343166
rect 654508 343110 654513 343166
rect 650208 343108 654513 343110
rect 58383 343105 58449 343108
rect 654447 343105 654513 343108
rect 40378 342958 40384 343022
rect 40448 342958 40454 343022
rect 40570 342810 40576 342874
rect 40640 342810 40646 342874
rect 40578 342546 40638 342810
rect 40770 341838 40830 342102
rect 40762 341774 40768 341838
rect 40832 341774 40838 341838
rect 42831 341540 42897 341543
rect 42528 341538 42897 341540
rect 42528 341482 42836 341538
rect 42892 341482 42897 341538
rect 42528 341480 42897 341482
rect 42831 341477 42897 341480
rect 40962 340654 41022 340918
rect 40954 340590 40960 340654
rect 41024 340590 41030 340654
rect 41346 340210 41406 340474
rect 41338 340146 41344 340210
rect 41408 340146 41414 340210
rect 42114 339618 42174 339882
rect 42106 339554 42112 339618
rect 42176 339554 42182 339618
rect 41730 339027 41790 339290
rect 41730 339022 41841 339027
rect 41730 338966 41780 339022
rect 41836 338966 41841 339022
rect 41730 338964 41841 338966
rect 41775 338961 41841 338964
rect 41154 338582 41214 338846
rect 41146 338518 41152 338582
rect 41216 338518 41222 338582
rect 41538 337990 41598 338254
rect 41530 337926 41536 337990
rect 41600 337926 41606 337990
rect 42306 337547 42366 337662
rect 42255 337542 42366 337547
rect 42255 337486 42260 337542
rect 42316 337486 42366 337542
rect 42255 337484 42366 337486
rect 42255 337481 42321 337484
rect 40002 336955 40062 337218
rect 40002 336950 40113 336955
rect 40002 336894 40052 336950
rect 40108 336894 40113 336950
rect 40002 336892 40113 336894
rect 40047 336889 40113 336892
rect 40194 336363 40254 336626
rect 40143 336358 40254 336363
rect 40143 336302 40148 336358
rect 40204 336302 40254 336358
rect 40143 336300 40254 336302
rect 40143 336297 40209 336300
rect 42682 336064 42688 336066
rect 42528 336004 42688 336064
rect 42682 336002 42688 336004
rect 42752 336002 42758 336066
rect 41730 335178 41790 335590
rect 41722 335114 41728 335178
rect 41792 335114 41798 335178
rect 675279 335030 675345 335031
rect 675279 335026 675328 335030
rect 675392 335028 675398 335030
rect 42498 334735 42558 334998
rect 675279 334970 675284 335026
rect 675279 334966 675328 334970
rect 675392 334968 675436 335028
rect 675392 334966 675398 334968
rect 675279 334965 675345 334966
rect 42498 334730 42609 334735
rect 42498 334674 42548 334730
rect 42604 334674 42609 334730
rect 42498 334672 42609 334674
rect 42543 334669 42609 334672
rect 675471 334586 675537 334587
rect 675471 334582 675520 334586
rect 675584 334584 675590 334586
rect 675471 334526 675476 334582
rect 675471 334522 675520 334526
rect 675584 334524 675628 334584
rect 675584 334522 675590 334524
rect 675471 334521 675537 334522
rect 42498 334140 42558 334406
rect 42498 334080 42750 334140
rect 35202 333551 35262 333888
rect 42690 333696 42750 334080
rect 35151 333546 35262 333551
rect 35151 333490 35156 333546
rect 35212 333490 35262 333546
rect 35151 333488 35262 333490
rect 42498 333636 42750 333696
rect 35151 333485 35217 333488
rect 42498 333400 42558 333636
rect 43215 333400 43281 333403
rect 42498 333398 43281 333400
rect 42498 333370 43220 333398
rect 42528 333342 43220 333370
rect 43276 333342 43281 333398
rect 42528 333340 43281 333342
rect 43215 333337 43281 333340
rect 35151 333104 35217 333107
rect 35151 333102 35262 333104
rect 35151 333046 35156 333102
rect 35212 333046 35262 333102
rect 35151 333041 35262 333046
rect 35202 332778 35262 333041
rect 654447 331624 654513 331627
rect 650208 331622 654513 331624
rect 650208 331566 654452 331622
rect 654508 331566 654513 331622
rect 650208 331564 654513 331566
rect 654447 331561 654513 331564
rect 673978 331118 673984 331182
rect 674048 331180 674054 331182
rect 675087 331180 675153 331183
rect 674048 331178 675153 331180
rect 674048 331122 675092 331178
rect 675148 331122 675153 331178
rect 674048 331120 675153 331122
rect 674048 331118 674054 331120
rect 675087 331117 675153 331120
rect 675759 330588 675825 330591
rect 676474 330588 676480 330590
rect 675759 330586 676480 330588
rect 675759 330530 675764 330586
rect 675820 330530 676480 330586
rect 675759 330528 676480 330530
rect 675759 330525 675825 330528
rect 676474 330526 676480 330528
rect 676544 330526 676550 330590
rect 674991 329552 675057 329555
rect 675322 329552 675328 329554
rect 674991 329550 675328 329552
rect 674991 329494 674996 329550
rect 675052 329494 675328 329550
rect 674991 329492 675328 329494
rect 674991 329489 675057 329492
rect 675322 329490 675328 329492
rect 675392 329490 675398 329554
rect 57807 328812 57873 328815
rect 57807 328810 64416 328812
rect 57807 328754 57812 328810
rect 57868 328754 64416 328810
rect 57807 328752 64416 328754
rect 57807 328749 57873 328752
rect 674170 328306 674176 328370
rect 674240 328368 674246 328370
rect 675375 328368 675441 328371
rect 674240 328366 675441 328368
rect 674240 328310 675380 328366
rect 675436 328310 675441 328366
rect 674240 328308 675441 328310
rect 674240 328306 674246 328308
rect 675375 328305 675441 328308
rect 675759 326888 675825 326891
rect 676666 326888 676672 326890
rect 675759 326886 676672 326888
rect 675759 326830 675764 326886
rect 675820 326830 676672 326886
rect 675759 326828 676672 326830
rect 675759 326825 675825 326828
rect 676666 326826 676672 326828
rect 676736 326826 676742 326890
rect 42682 324754 42688 324818
rect 42752 324816 42758 324818
rect 42831 324816 42897 324819
rect 42752 324814 42897 324816
rect 42752 324758 42836 324814
rect 42892 324758 42897 324814
rect 42752 324756 42897 324758
rect 42752 324754 42758 324756
rect 42831 324753 42897 324756
rect 41775 320526 41841 320527
rect 41722 320462 41728 320526
rect 41792 320524 41841 320526
rect 41792 320522 41884 320524
rect 41836 320466 41884 320522
rect 41792 320464 41884 320466
rect 41792 320462 41841 320464
rect 41775 320461 41841 320462
rect 42063 319786 42129 319787
rect 42063 319782 42112 319786
rect 42176 319784 42182 319786
rect 655119 319784 655185 319787
rect 42063 319726 42068 319782
rect 42063 319722 42112 319726
rect 42176 319724 42220 319784
rect 650208 319782 655185 319784
rect 650208 319726 655124 319782
rect 655180 319726 655185 319782
rect 650208 319724 655185 319726
rect 42176 319722 42182 319724
rect 42063 319721 42129 319722
rect 655119 319721 655185 319724
rect 41722 318390 41728 318454
rect 41792 318452 41798 318454
rect 42159 318452 42225 318455
rect 42490 318452 42496 318454
rect 41792 318450 42496 318452
rect 41792 318394 42164 318450
rect 42220 318394 42496 318450
rect 41792 318392 42496 318394
rect 41792 318390 41798 318392
rect 42159 318389 42225 318392
rect 42490 318390 42496 318392
rect 42560 318390 42566 318454
rect 41914 317946 41920 318010
rect 41984 318008 41990 318010
rect 42063 318008 42129 318011
rect 42874 318008 42880 318010
rect 41984 318006 42880 318008
rect 41984 317950 42068 318006
rect 42124 317950 42880 318006
rect 41984 317948 42880 317950
rect 41984 317946 41990 317948
rect 42063 317945 42129 317948
rect 42874 317946 42880 317948
rect 42944 317946 42950 318010
rect 41530 316170 41536 316234
rect 41600 316232 41606 316234
rect 41775 316232 41841 316235
rect 41600 316230 41841 316232
rect 41600 316174 41780 316230
rect 41836 316174 41841 316230
rect 41600 316172 41841 316174
rect 41600 316170 41606 316172
rect 41775 316169 41841 316172
rect 41338 315430 41344 315494
rect 41408 315492 41414 315494
rect 41775 315492 41841 315495
rect 41408 315490 41841 315492
rect 41408 315434 41780 315490
rect 41836 315434 41841 315490
rect 41408 315432 41841 315434
rect 41408 315430 41414 315432
rect 41775 315429 41841 315432
rect 674415 315048 674481 315051
rect 674415 315046 674784 315048
rect 674415 314990 674420 315046
rect 674476 314990 674784 315046
rect 674415 314988 674784 314990
rect 674415 314985 674481 314988
rect 674703 314752 674769 314755
rect 674703 314750 674814 314752
rect 674703 314694 674708 314750
rect 674764 314694 674814 314750
rect 674703 314689 674814 314694
rect 57999 314604 58065 314607
rect 57999 314602 64416 314604
rect 57999 314546 58004 314602
rect 58060 314546 64416 314602
rect 674754 314574 674814 314689
rect 57999 314544 64416 314546
rect 57999 314541 58065 314544
rect 674415 314012 674481 314015
rect 674415 314010 674784 314012
rect 674415 313954 674420 314010
rect 674476 313954 674784 314010
rect 674415 313952 674784 313954
rect 674415 313949 674481 313952
rect 40762 313654 40768 313718
rect 40832 313716 40838 313718
rect 41871 313716 41937 313719
rect 40832 313714 41937 313716
rect 40832 313658 41876 313714
rect 41932 313658 41937 313714
rect 40832 313656 41937 313658
rect 40832 313654 40838 313656
rect 41871 313653 41937 313656
rect 677050 313654 677056 313718
rect 677120 313654 677126 313718
rect 677058 313390 677118 313654
rect 41146 313210 41152 313274
rect 41216 313272 41222 313274
rect 41775 313272 41841 313275
rect 41216 313270 41841 313272
rect 41216 313214 41780 313270
rect 41836 313214 41841 313270
rect 41216 313212 41841 313214
rect 41216 313210 41222 313212
rect 41775 313209 41841 313212
rect 677250 312534 677310 312946
rect 677242 312470 677248 312534
rect 677312 312470 677318 312534
rect 40954 312322 40960 312386
rect 41024 312384 41030 312386
rect 41775 312384 41841 312387
rect 41024 312382 41841 312384
rect 41024 312326 41780 312382
rect 41836 312326 41841 312382
rect 41024 312324 41841 312326
rect 41024 312322 41030 312324
rect 41775 312321 41841 312324
rect 677442 312090 677502 312354
rect 677434 312026 677440 312090
rect 677504 312026 677510 312090
rect 677058 311498 677118 311762
rect 677050 311434 677056 311498
rect 677120 311434 677126 311498
rect 674031 311348 674097 311351
rect 674031 311346 674784 311348
rect 674031 311290 674036 311346
rect 674092 311290 674784 311346
rect 674031 311288 674784 311290
rect 674031 311285 674097 311288
rect 674170 310694 674176 310758
rect 674240 310756 674246 310758
rect 674240 310696 674784 310756
rect 674240 310694 674246 310696
rect 675138 310019 675198 310134
rect 675087 310014 675198 310019
rect 675087 309958 675092 310014
rect 675148 309958 675198 310014
rect 675087 309956 675198 309958
rect 675087 309953 675153 309956
rect 674319 309646 674385 309649
rect 674319 309644 674784 309646
rect 674319 309588 674324 309644
rect 674380 309588 674784 309644
rect 674319 309586 674784 309588
rect 674319 309583 674385 309586
rect 674946 308835 675006 309098
rect 674946 308830 675057 308835
rect 674946 308774 674996 308830
rect 675052 308774 675057 308830
rect 674946 308772 675057 308774
rect 674991 308769 675057 308772
rect 677058 308243 677118 308506
rect 677007 308238 677118 308243
rect 677007 308182 677012 308238
rect 677068 308182 677118 308238
rect 677007 308180 677118 308182
rect 677007 308177 677073 308180
rect 655311 307944 655377 307947
rect 650208 307942 655377 307944
rect 650208 307886 655316 307942
rect 655372 307886 655377 307942
rect 650208 307884 655377 307886
rect 655311 307881 655377 307884
rect 674946 307799 675006 307988
rect 674895 307794 675006 307799
rect 674895 307738 674900 307794
rect 674956 307738 675006 307794
rect 674895 307736 675006 307738
rect 674895 307733 674961 307736
rect 674754 307207 674814 307470
rect 674754 307202 674865 307207
rect 674754 307146 674804 307202
rect 674860 307146 674865 307202
rect 674754 307144 674865 307146
rect 674799 307141 674865 307144
rect 674607 306760 674673 306763
rect 674754 306760 674814 306878
rect 674607 306758 674814 306760
rect 674607 306702 674612 306758
rect 674668 306702 674814 306758
rect 674607 306700 674814 306702
rect 674607 306697 674673 306700
rect 676866 306023 676926 306360
rect 676866 306018 676977 306023
rect 676866 305962 676916 306018
rect 676972 305962 676977 306018
rect 676866 305960 676977 305962
rect 676911 305957 676977 305960
rect 674127 305872 674193 305875
rect 674127 305870 674784 305872
rect 674127 305814 674132 305870
rect 674188 305814 674784 305870
rect 674127 305812 674784 305814
rect 674127 305809 674193 305812
rect 674754 305135 674814 305250
rect 674703 305130 674814 305135
rect 674703 305074 674708 305130
rect 674764 305074 674814 305130
rect 674703 305072 674814 305074
rect 674703 305069 674769 305072
rect 674511 304540 674577 304543
rect 674754 304540 674814 304732
rect 674511 304538 674814 304540
rect 674511 304482 674516 304538
rect 674572 304482 674814 304538
rect 674511 304480 674814 304482
rect 674511 304477 674577 304480
rect 674223 304244 674289 304247
rect 674223 304242 674784 304244
rect 674223 304186 674228 304242
rect 674284 304186 674784 304242
rect 674223 304184 674784 304186
rect 674223 304181 674289 304184
rect 674415 303652 674481 303655
rect 674415 303650 674784 303652
rect 674415 303594 674420 303650
rect 674476 303594 674784 303650
rect 674415 303592 674784 303594
rect 674415 303589 674481 303592
rect 676866 302767 676926 303104
rect 676815 302762 676926 302767
rect 676815 302706 676820 302762
rect 676876 302706 676926 302762
rect 676815 302704 676926 302706
rect 676815 302701 676881 302704
rect 42831 302690 42897 302693
rect 42528 302688 42897 302690
rect 42528 302632 42836 302688
rect 42892 302632 42897 302688
rect 42528 302630 42897 302632
rect 42831 302627 42897 302630
rect 674415 302616 674481 302619
rect 674415 302614 674784 302616
rect 674415 302558 674420 302614
rect 674476 302558 674784 302614
rect 674415 302556 674784 302558
rect 674415 302553 674481 302556
rect 42447 302320 42513 302323
rect 676815 302320 676881 302323
rect 42447 302318 42558 302320
rect 42447 302262 42452 302318
rect 42508 302262 42558 302318
rect 42447 302257 42558 302262
rect 676815 302318 676926 302320
rect 676815 302262 676820 302318
rect 676876 302262 676926 302318
rect 676815 302257 676926 302262
rect 42498 302142 42558 302257
rect 676866 301994 676926 302257
rect 42831 301580 42897 301583
rect 42528 301578 42897 301580
rect 42528 301522 42836 301578
rect 42892 301522 42897 301578
rect 42528 301520 42897 301522
rect 42831 301517 42897 301520
rect 42498 300988 42558 301032
rect 43119 300988 43185 300991
rect 42498 300986 43185 300988
rect 42498 300930 43124 300986
rect 43180 300930 43185 300986
rect 42498 300928 43185 300930
rect 43119 300925 43185 300928
rect 43215 300544 43281 300547
rect 42528 300542 43281 300544
rect 42528 300486 43220 300542
rect 43276 300486 43281 300542
rect 42528 300484 43281 300486
rect 43215 300481 43281 300484
rect 59439 300100 59505 300103
rect 59439 300098 64416 300100
rect 59439 300042 59444 300098
rect 59500 300042 64416 300098
rect 59439 300040 64416 300042
rect 59439 300037 59505 300040
rect 40386 299806 40446 299922
rect 40378 299742 40384 299806
rect 40448 299742 40454 299806
rect 40570 299594 40576 299658
rect 40640 299656 40646 299658
rect 42298 299656 42304 299658
rect 40640 299596 42304 299656
rect 40640 299594 40646 299596
rect 42298 299594 42304 299596
rect 42368 299594 42374 299658
rect 42306 299404 42366 299594
rect 675898 299446 675904 299510
rect 675968 299508 675974 299510
rect 676911 299508 676977 299511
rect 675968 299506 676977 299508
rect 675968 299450 676916 299506
rect 676972 299450 676977 299506
rect 675968 299448 676977 299450
rect 675968 299446 675974 299448
rect 676911 299445 676977 299448
rect 676666 299298 676672 299362
rect 676736 299360 676742 299362
rect 677007 299360 677073 299363
rect 676736 299358 677073 299360
rect 676736 299302 677012 299358
rect 677068 299302 677073 299358
rect 676736 299300 677073 299302
rect 676736 299298 676742 299300
rect 677007 299297 677073 299300
rect 40962 298622 41022 298886
rect 40954 298558 40960 298622
rect 41024 298558 41030 298622
rect 41730 298031 41790 298294
rect 41730 298026 41841 298031
rect 41730 297970 41780 298026
rect 41836 297970 41841 298026
rect 41730 297968 41841 297970
rect 41775 297965 41841 297968
rect 40770 297438 40830 297776
rect 40762 297374 40768 297438
rect 40832 297374 40838 297438
rect 41346 296994 41406 297258
rect 41338 296930 41344 296994
rect 41408 296930 41414 296994
rect 42114 296550 42174 296666
rect 42106 296486 42112 296550
rect 42176 296486 42182 296550
rect 654543 296252 654609 296255
rect 650208 296250 654609 296252
rect 650208 296194 654548 296250
rect 654604 296194 654609 296250
rect 650208 296192 654609 296194
rect 654543 296189 654609 296192
rect 42306 295811 42366 296148
rect 42255 295806 42366 295811
rect 42255 295750 42260 295806
rect 42316 295750 42366 295806
rect 42255 295748 42366 295750
rect 42255 295745 42321 295748
rect 41154 295366 41214 295630
rect 41146 295302 41152 295366
rect 41216 295302 41222 295366
rect 41538 294774 41598 295038
rect 41530 294710 41536 294774
rect 41600 294710 41606 294774
rect 42306 294331 42366 294520
rect 42306 294326 42417 294331
rect 42306 294270 42356 294326
rect 42412 294270 42417 294326
rect 42306 294268 42417 294270
rect 42351 294265 42417 294268
rect 40194 293739 40254 294002
rect 40194 293734 40305 293739
rect 40194 293678 40244 293734
rect 40300 293678 40305 293734
rect 40194 293676 40305 293678
rect 40239 293673 40305 293676
rect 40002 293147 40062 293410
rect 40002 293142 40113 293147
rect 40002 293086 40052 293142
rect 40108 293086 40113 293142
rect 40002 293084 40113 293086
rect 40047 293081 40113 293084
rect 40002 292555 40062 292818
rect 39951 292550 40062 292555
rect 39951 292494 39956 292550
rect 40012 292494 40062 292550
rect 39951 292492 40062 292494
rect 39951 292489 40017 292492
rect 40194 292111 40254 292374
rect 40143 292106 40254 292111
rect 40143 292050 40148 292106
rect 40204 292050 40254 292106
rect 40143 292048 40254 292050
rect 40143 292045 40209 292048
rect 42682 291812 42688 291814
rect 42528 291752 42688 291812
rect 42682 291750 42688 291752
rect 42752 291750 42758 291814
rect 42498 290924 42558 291190
rect 42498 290864 42750 290924
rect 35202 290483 35262 290746
rect 35151 290478 35262 290483
rect 42690 290480 42750 290864
rect 35151 290422 35156 290478
rect 35212 290422 35262 290478
rect 35151 290420 35262 290422
rect 42498 290420 42750 290480
rect 35151 290417 35217 290420
rect 42498 290184 42558 290420
rect 42831 290184 42897 290187
rect 42498 290182 42897 290184
rect 42498 290154 42836 290182
rect 42528 290126 42836 290154
rect 42892 290126 42897 290182
rect 42528 290124 42897 290126
rect 42831 290121 42897 290124
rect 675279 290038 675345 290039
rect 675279 290034 675328 290038
rect 675392 290036 675398 290038
rect 675279 289978 675284 290034
rect 675279 289974 675328 289978
rect 675392 289976 675436 290036
rect 675392 289974 675398 289976
rect 675279 289973 675345 289974
rect 35151 289888 35217 289891
rect 35151 289886 35262 289888
rect 35151 289830 35156 289886
rect 35212 289830 35262 289886
rect 35151 289825 35262 289830
rect 35202 289562 35262 289825
rect 673935 289594 674001 289595
rect 673935 289590 673984 289594
rect 674048 289592 674054 289594
rect 673935 289534 673940 289590
rect 673935 289530 673984 289534
rect 674048 289532 674092 289592
rect 674048 289530 674054 289532
rect 673935 289529 674001 289530
rect 58095 285892 58161 285895
rect 58095 285890 64416 285892
rect 58095 285834 58100 285890
rect 58156 285834 64416 285890
rect 58095 285832 64416 285834
rect 58095 285829 58161 285832
rect 674362 284942 674368 285006
rect 674432 285004 674438 285006
rect 675087 285004 675153 285007
rect 674432 285002 675153 285004
rect 674432 284946 675092 285002
rect 675148 284946 675153 285002
rect 674432 284944 675153 284946
rect 674432 284942 674438 284944
rect 675087 284941 675153 284944
rect 42351 284856 42417 284859
rect 42490 284856 42496 284858
rect 42351 284854 42496 284856
rect 42351 284798 42356 284854
rect 42412 284798 42496 284854
rect 42351 284796 42496 284798
rect 42351 284793 42417 284796
rect 42490 284794 42496 284796
rect 42560 284794 42566 284858
rect 675759 284856 675825 284859
rect 675898 284856 675904 284858
rect 675759 284854 675904 284856
rect 675759 284798 675764 284854
rect 675820 284798 675904 284854
rect 675759 284796 675904 284798
rect 675759 284793 675825 284796
rect 675898 284794 675904 284796
rect 675968 284794 675974 284858
rect 654063 284708 654129 284711
rect 650208 284706 654129 284708
rect 650208 284650 654068 284706
rect 654124 284650 654129 284706
rect 650208 284648 654129 284650
rect 654063 284645 654129 284648
rect 673935 284710 674001 284711
rect 673935 284706 673984 284710
rect 674048 284708 674054 284710
rect 673935 284650 673940 284706
rect 673935 284646 673984 284650
rect 674048 284648 674092 284708
rect 674048 284646 674054 284648
rect 673935 284645 674001 284646
rect 674170 283610 674176 283674
rect 674240 283672 674246 283674
rect 675375 283672 675441 283675
rect 674240 283670 675441 283672
rect 674240 283614 675380 283670
rect 675436 283614 675441 283670
rect 674240 283612 675441 283614
rect 674240 283610 674246 283612
rect 675375 283609 675441 283612
rect 675759 281896 675825 281899
rect 676666 281896 676672 281898
rect 675759 281894 676672 281896
rect 675759 281838 675764 281894
rect 675820 281838 676672 281894
rect 675759 281836 676672 281838
rect 675759 281833 675825 281836
rect 676666 281834 676672 281836
rect 676736 281834 676742 281898
rect 42351 281600 42417 281603
rect 42490 281600 42496 281602
rect 42351 281598 42496 281600
rect 42351 281542 42356 281598
rect 42412 281542 42496 281598
rect 42351 281540 42496 281542
rect 42351 281537 42417 281540
rect 42490 281538 42496 281540
rect 42560 281538 42566 281602
rect 42159 278640 42225 278643
rect 42682 278640 42688 278642
rect 42159 278638 42688 278640
rect 42159 278582 42164 278638
rect 42220 278582 42688 278638
rect 42159 278580 42688 278582
rect 42159 278577 42225 278580
rect 42682 278578 42688 278580
rect 42752 278578 42758 278642
rect 368559 278640 368625 278643
rect 383823 278640 383889 278643
rect 257730 278638 368625 278640
rect 257730 278582 368564 278638
rect 368620 278582 368625 278638
rect 257730 278580 368625 278582
rect 257583 278492 257649 278495
rect 257730 278492 257790 278580
rect 368559 278577 368625 278580
rect 368706 278638 383889 278640
rect 368706 278582 383828 278638
rect 383884 278582 383889 278638
rect 368706 278580 383889 278582
rect 257583 278490 257790 278492
rect 257583 278434 257588 278490
rect 257644 278434 257790 278490
rect 257583 278432 257790 278434
rect 293967 278492 294033 278495
rect 299535 278492 299601 278495
rect 293967 278490 299601 278492
rect 293967 278434 293972 278490
rect 294028 278434 299540 278490
rect 299596 278434 299601 278490
rect 293967 278432 299601 278434
rect 257583 278429 257649 278432
rect 293967 278429 294033 278432
rect 299535 278429 299601 278432
rect 299727 278492 299793 278495
rect 300399 278492 300465 278495
rect 299727 278490 300465 278492
rect 299727 278434 299732 278490
rect 299788 278434 300404 278490
rect 300460 278434 300465 278490
rect 299727 278432 300465 278434
rect 299727 278429 299793 278432
rect 300399 278429 300465 278432
rect 315279 278492 315345 278495
rect 368706 278492 368766 278580
rect 383823 278577 383889 278580
rect 417474 278580 428910 278640
rect 417474 278495 417534 278580
rect 428850 278495 428910 278580
rect 515394 278580 515646 278640
rect 315279 278490 368766 278492
rect 315279 278434 315284 278490
rect 315340 278434 368766 278490
rect 315279 278432 368766 278434
rect 368847 278492 368913 278495
rect 397455 278492 397521 278495
rect 368847 278490 397521 278492
rect 368847 278434 368852 278490
rect 368908 278434 397460 278490
rect 397516 278434 397521 278490
rect 368847 278432 397521 278434
rect 315279 278429 315345 278432
rect 368847 278429 368913 278432
rect 397455 278429 397521 278432
rect 417423 278490 417534 278495
rect 417423 278434 417428 278490
rect 417484 278434 417534 278490
rect 417423 278432 417534 278434
rect 428847 278490 428913 278495
rect 428847 278434 428852 278490
rect 428908 278434 428913 278490
rect 417423 278429 417489 278432
rect 428847 278429 428913 278434
rect 429039 278492 429105 278495
rect 440655 278492 440721 278495
rect 429039 278490 440721 278492
rect 429039 278434 429044 278490
rect 429100 278434 440660 278490
rect 440716 278434 440721 278490
rect 429039 278432 440721 278434
rect 429039 278429 429105 278432
rect 440655 278429 440721 278432
rect 489615 278492 489681 278495
rect 495375 278492 495441 278495
rect 489615 278490 495441 278492
rect 489615 278434 489620 278490
rect 489676 278434 495380 278490
rect 495436 278434 495441 278490
rect 489615 278432 495441 278434
rect 489615 278429 489681 278432
rect 495375 278429 495441 278432
rect 501327 278492 501393 278495
rect 515394 278492 515454 278580
rect 501327 278490 515454 278492
rect 501327 278434 501332 278490
rect 501388 278434 515454 278490
rect 501327 278432 515454 278434
rect 515586 278492 515646 278580
rect 551298 278580 558846 278640
rect 551298 278495 551358 278580
rect 525519 278492 525585 278495
rect 515586 278490 525585 278492
rect 515586 278434 525524 278490
rect 525580 278434 525585 278490
rect 515586 278432 525585 278434
rect 501327 278429 501393 278432
rect 525519 278429 525585 278432
rect 551247 278490 551358 278495
rect 551247 278434 551252 278490
rect 551308 278434 551358 278490
rect 551247 278432 551358 278434
rect 551247 278429 551313 278432
rect 299535 278344 299601 278347
rect 300303 278344 300369 278347
rect 299535 278342 300369 278344
rect 299535 278286 299540 278342
rect 299596 278286 300308 278342
rect 300364 278286 300369 278342
rect 299535 278284 300369 278286
rect 299535 278281 299601 278284
rect 300303 278281 300369 278284
rect 303375 278344 303441 278347
rect 467535 278344 467601 278347
rect 303375 278342 467601 278344
rect 303375 278286 303380 278342
rect 303436 278286 467540 278342
rect 467596 278286 467601 278342
rect 303375 278284 467601 278286
rect 558786 278344 558846 278580
rect 578754 278580 590334 278640
rect 578754 278344 578814 278580
rect 590274 278494 590334 278580
rect 590266 278430 590272 278494
rect 590336 278430 590342 278494
rect 604858 278430 604864 278494
rect 604928 278492 604934 278494
rect 610479 278492 610545 278495
rect 604928 278490 610545 278492
rect 604928 278434 610484 278490
rect 610540 278434 610545 278490
rect 604928 278432 610545 278434
rect 604928 278430 604934 278432
rect 610479 278429 610545 278432
rect 610767 278492 610833 278495
rect 625071 278492 625137 278495
rect 610767 278490 625137 278492
rect 610767 278434 610772 278490
rect 610828 278434 625076 278490
rect 625132 278434 625137 278490
rect 610767 278432 625137 278434
rect 610767 278429 610833 278432
rect 625071 278429 625137 278432
rect 631023 278492 631089 278495
rect 631023 278490 645054 278492
rect 631023 278434 631028 278490
rect 631084 278434 645054 278490
rect 631023 278432 645054 278434
rect 631023 278429 631089 278432
rect 558786 278284 578814 278344
rect 303375 278281 303441 278284
rect 467535 278281 467601 278284
rect 590458 278282 590464 278346
rect 590528 278344 590534 278346
rect 604858 278344 604864 278346
rect 590528 278284 604864 278344
rect 590528 278282 590534 278284
rect 604858 278282 604864 278284
rect 604928 278282 604934 278346
rect 644994 278344 645054 278432
rect 645178 278344 645184 278346
rect 644994 278284 645184 278344
rect 645178 278282 645184 278284
rect 645248 278282 645254 278346
rect 304527 278196 304593 278199
rect 474735 278196 474801 278199
rect 304527 278194 474801 278196
rect 304527 278138 304532 278194
rect 304588 278138 474740 278194
rect 474796 278138 474801 278194
rect 304527 278136 474801 278138
rect 304527 278133 304593 278136
rect 474735 278133 474801 278136
rect 645178 278134 645184 278198
rect 645248 278134 645254 278198
rect 305199 278048 305265 278051
rect 481839 278048 481905 278051
rect 305199 278046 481905 278048
rect 305199 277990 305204 278046
rect 305260 277990 481844 278046
rect 481900 277990 481905 278046
rect 305199 277988 481905 277990
rect 645186 278048 645246 278134
rect 645999 278048 646065 278051
rect 645186 278046 646065 278048
rect 645186 277990 646004 278046
rect 646060 277990 646065 278046
rect 645186 277988 646065 277990
rect 305199 277985 305265 277988
rect 481839 277985 481905 277988
rect 645999 277985 646065 277988
rect 299631 277900 299697 277903
rect 300399 277900 300465 277903
rect 299631 277898 300465 277900
rect 299631 277842 299636 277898
rect 299692 277842 300404 277898
rect 300460 277842 300465 277898
rect 299631 277840 300465 277842
rect 299631 277837 299697 277840
rect 300399 277837 300465 277840
rect 306351 277900 306417 277903
rect 488943 277900 489009 277903
rect 306351 277898 489009 277900
rect 306351 277842 306356 277898
rect 306412 277842 488948 277898
rect 489004 277842 489009 277898
rect 306351 277840 489009 277842
rect 306351 277837 306417 277840
rect 488943 277837 489009 277840
rect 299535 277752 299601 277755
rect 300303 277752 300369 277755
rect 299535 277750 300369 277752
rect 299535 277694 299540 277750
rect 299596 277694 300308 277750
rect 300364 277694 300369 277750
rect 299535 277692 300369 277694
rect 299535 277689 299601 277692
rect 300303 277689 300369 277692
rect 307119 277752 307185 277755
rect 496143 277752 496209 277755
rect 307119 277750 496209 277752
rect 307119 277694 307124 277750
rect 307180 277694 496148 277750
rect 496204 277694 496209 277750
rect 307119 277692 496209 277694
rect 307119 277689 307185 277692
rect 496143 277689 496209 277692
rect 308367 277604 308433 277607
rect 507087 277604 507153 277607
rect 308367 277602 507153 277604
rect 308367 277546 308372 277602
rect 308428 277546 507092 277602
rect 507148 277546 507153 277602
rect 308367 277544 507153 277546
rect 308367 277541 308433 277544
rect 507087 277541 507153 277544
rect 309519 277456 309585 277459
rect 517743 277456 517809 277459
rect 309519 277454 517809 277456
rect 309519 277398 309524 277454
rect 309580 277398 517748 277454
rect 517804 277398 517809 277454
rect 309519 277396 517809 277398
rect 309519 277393 309585 277396
rect 517743 277393 517809 277396
rect 310959 277308 311025 277311
rect 528495 277308 528561 277311
rect 310959 277306 528561 277308
rect 310959 277250 310964 277306
rect 311020 277250 528500 277306
rect 528556 277250 528561 277306
rect 310959 277248 528561 277250
rect 310959 277245 311025 277248
rect 528495 277245 528561 277248
rect 312303 277160 312369 277163
rect 539247 277160 539313 277163
rect 312303 277158 539313 277160
rect 312303 277102 312308 277158
rect 312364 277102 539252 277158
rect 539308 277102 539313 277158
rect 312303 277100 539313 277102
rect 312303 277097 312369 277100
rect 539247 277097 539313 277100
rect 206031 277012 206097 277015
rect 378255 277012 378321 277015
rect 206031 277010 378321 277012
rect 206031 276954 206036 277010
rect 206092 276954 378260 277010
rect 378316 276954 378321 277010
rect 206031 276952 378321 276954
rect 206031 276949 206097 276952
rect 378255 276949 378321 276952
rect 378447 277012 378513 277015
rect 383055 277012 383121 277015
rect 378447 277010 383121 277012
rect 378447 276954 378452 277010
rect 378508 276954 383060 277010
rect 383116 276954 383121 277010
rect 378447 276952 383121 276954
rect 378447 276949 378513 276952
rect 383055 276949 383121 276952
rect 383247 277012 383313 277015
rect 396687 277012 396753 277015
rect 383247 277010 396753 277012
rect 383247 276954 383252 277010
rect 383308 276954 396692 277010
rect 396748 276954 396753 277010
rect 383247 276952 396753 276954
rect 383247 276949 383313 276952
rect 396687 276949 396753 276952
rect 321903 276864 321969 276867
rect 617679 276864 617745 276867
rect 321903 276862 617745 276864
rect 321903 276806 321908 276862
rect 321964 276806 617684 276862
rect 617740 276806 617745 276862
rect 321903 276804 617745 276806
rect 321903 276801 321969 276804
rect 617679 276801 617745 276804
rect 325551 276716 325617 276719
rect 635535 276716 635601 276719
rect 325551 276714 635601 276716
rect 325551 276658 325556 276714
rect 325612 276658 635540 276714
rect 635596 276658 635601 276714
rect 325551 276656 635601 276658
rect 325551 276653 325617 276656
rect 635535 276653 635601 276656
rect 42063 276570 42129 276571
rect 42063 276566 42112 276570
rect 42176 276568 42182 276570
rect 324687 276568 324753 276571
rect 642735 276568 642801 276571
rect 42063 276510 42068 276566
rect 42063 276506 42112 276510
rect 42176 276508 42220 276568
rect 324687 276566 642801 276568
rect 324687 276510 324692 276566
rect 324748 276510 642740 276566
rect 642796 276510 642801 276566
rect 324687 276508 642801 276510
rect 42176 276506 42182 276508
rect 42063 276505 42129 276506
rect 324687 276505 324753 276508
rect 642735 276505 642801 276508
rect 262863 276420 262929 276423
rect 374127 276420 374193 276423
rect 262863 276418 374193 276420
rect 262863 276362 262868 276418
rect 262924 276362 374132 276418
rect 374188 276362 374193 276418
rect 262863 276360 374193 276362
rect 262863 276357 262929 276360
rect 374127 276357 374193 276360
rect 374319 276420 374385 276423
rect 637935 276420 638001 276423
rect 374319 276418 638001 276420
rect 374319 276362 374324 276418
rect 374380 276362 637940 276418
rect 637996 276362 638001 276418
rect 374319 276360 638001 276362
rect 374319 276357 374385 276360
rect 637935 276357 638001 276360
rect 318639 276272 318705 276275
rect 592719 276272 592785 276275
rect 318639 276270 592785 276272
rect 318639 276214 318644 276270
rect 318700 276214 592724 276270
rect 592780 276214 592785 276270
rect 318639 276212 592785 276214
rect 318639 276209 318705 276212
rect 592719 276209 592785 276212
rect 269391 276124 269457 276127
rect 325455 276124 325521 276127
rect 269391 276122 325521 276124
rect 269391 276066 269396 276122
rect 269452 276066 325460 276122
rect 325516 276066 325521 276122
rect 269391 276064 325521 276066
rect 269391 276061 269457 276064
rect 325455 276061 325521 276064
rect 325647 276124 325713 276127
rect 607023 276124 607089 276127
rect 325647 276122 607089 276124
rect 325647 276066 325652 276122
rect 325708 276066 607028 276122
rect 607084 276066 607089 276122
rect 325647 276064 607089 276066
rect 325647 276061 325713 276064
rect 607023 276061 607089 276064
rect 319791 275976 319857 275979
rect 599823 275976 599889 275979
rect 319791 275974 599889 275976
rect 319791 275918 319796 275974
rect 319852 275918 599828 275974
rect 599884 275918 599889 275974
rect 319791 275916 599889 275918
rect 319791 275913 319857 275916
rect 599823 275913 599889 275916
rect 320847 275828 320913 275831
rect 610575 275828 610641 275831
rect 320847 275826 610641 275828
rect 320847 275770 320852 275826
rect 320908 275770 610580 275826
rect 610636 275770 610641 275826
rect 320847 275768 610641 275770
rect 320847 275765 320913 275768
rect 610575 275765 610641 275768
rect 322863 275680 322929 275683
rect 624879 275680 624945 275683
rect 322863 275678 624945 275680
rect 322863 275622 322868 275678
rect 322924 275622 624884 275678
rect 624940 275622 624945 275678
rect 322863 275620 624945 275622
rect 322863 275617 322929 275620
rect 624879 275617 624945 275620
rect 264399 275532 264465 275535
rect 602223 275532 602289 275535
rect 264399 275530 602289 275532
rect 264399 275474 264404 275530
rect 264460 275474 602228 275530
rect 602284 275474 602289 275530
rect 264399 275472 602289 275474
rect 264399 275469 264465 275472
rect 602223 275469 602289 275472
rect 265935 275384 266001 275387
rect 616527 275384 616593 275387
rect 265935 275382 616593 275384
rect 265935 275326 265940 275382
rect 265996 275326 616532 275382
rect 616588 275326 616593 275382
rect 265935 275324 616593 275326
rect 265935 275321 266001 275324
rect 616527 275321 616593 275324
rect 267087 275236 267153 275239
rect 623631 275236 623697 275239
rect 267087 275234 623697 275236
rect 267087 275178 267092 275234
rect 267148 275178 623636 275234
rect 623692 275178 623697 275234
rect 267087 275176 623697 275178
rect 267087 275173 267153 275176
rect 623631 275173 623697 275176
rect 267183 275088 267249 275091
rect 627279 275088 627345 275091
rect 267183 275086 627345 275088
rect 267183 275030 267188 275086
rect 267244 275030 627284 275086
rect 627340 275030 627345 275086
rect 267183 275028 627345 275030
rect 267183 275025 267249 275028
rect 627279 275025 627345 275028
rect 261615 274940 261681 274943
rect 373359 274940 373425 274943
rect 261615 274938 373425 274940
rect 261615 274882 261620 274938
rect 261676 274882 373364 274938
rect 373420 274882 373425 274938
rect 261615 274880 373425 274882
rect 261615 274877 261681 274880
rect 373359 274877 373425 274880
rect 378063 274940 378129 274943
rect 382671 274940 382737 274943
rect 378063 274938 382737 274940
rect 378063 274882 378068 274938
rect 378124 274882 382676 274938
rect 382732 274882 382737 274938
rect 378063 274880 382737 274882
rect 378063 274877 378129 274880
rect 382671 274877 382737 274880
rect 383247 274940 383313 274943
rect 645135 274940 645201 274943
rect 383247 274938 645201 274940
rect 383247 274882 383252 274938
rect 383308 274882 645140 274938
rect 645196 274882 645201 274938
rect 383247 274880 645201 274882
rect 383247 274877 383313 274880
rect 645135 274877 645201 274880
rect 41967 274794 42033 274795
rect 41914 274730 41920 274794
rect 41984 274792 42033 274794
rect 254127 274792 254193 274795
rect 520143 274792 520209 274795
rect 41984 274790 42076 274792
rect 42028 274734 42076 274790
rect 41984 274732 42076 274734
rect 254127 274790 520209 274792
rect 254127 274734 254132 274790
rect 254188 274734 520148 274790
rect 520204 274734 520209 274790
rect 254127 274732 520209 274734
rect 41984 274730 42033 274732
rect 41967 274729 42033 274730
rect 254127 274729 254193 274732
rect 520143 274729 520209 274732
rect 41722 274582 41728 274646
rect 41792 274644 41798 274646
rect 42159 274644 42225 274647
rect 42874 274644 42880 274646
rect 41792 274642 42880 274644
rect 41792 274586 42164 274642
rect 42220 274586 42880 274642
rect 41792 274584 42880 274586
rect 41792 274582 41798 274584
rect 42159 274581 42225 274584
rect 42874 274582 42880 274584
rect 42944 274582 42950 274646
rect 253935 274644 254001 274647
rect 516591 274644 516657 274647
rect 253935 274642 516657 274644
rect 253935 274586 253940 274642
rect 253996 274586 516596 274642
rect 516652 274586 516657 274642
rect 253935 274584 516657 274586
rect 253935 274581 254001 274584
rect 516591 274581 516657 274584
rect 252399 274496 252465 274499
rect 505935 274496 506001 274499
rect 252399 274494 506001 274496
rect 252399 274438 252404 274494
rect 252460 274438 505940 274494
rect 505996 274438 506001 274494
rect 252399 274436 506001 274438
rect 252399 274433 252465 274436
rect 505935 274433 506001 274436
rect 251823 274348 251889 274351
rect 498831 274348 498897 274351
rect 251823 274346 498897 274348
rect 251823 274290 251828 274346
rect 251884 274290 498836 274346
rect 498892 274290 498897 274346
rect 251823 274288 498897 274290
rect 251823 274285 251889 274288
rect 498831 274285 498897 274288
rect 250671 274200 250737 274203
rect 491631 274200 491697 274203
rect 250671 274198 491697 274200
rect 250671 274142 250676 274198
rect 250732 274142 491636 274198
rect 491692 274142 491697 274198
rect 250671 274140 491697 274142
rect 250671 274137 250737 274140
rect 491631 274137 491697 274140
rect 249807 274052 249873 274055
rect 484431 274052 484497 274055
rect 249807 274050 484497 274052
rect 249807 273994 249812 274050
rect 249868 273994 484436 274050
rect 484492 273994 484497 274050
rect 249807 273992 484497 273994
rect 249807 273989 249873 273992
rect 484431 273989 484497 273992
rect 263343 273904 263409 273907
rect 382959 273904 383025 273907
rect 403119 273904 403185 273907
rect 263343 273902 383025 273904
rect 263343 273846 263348 273902
rect 263404 273846 382964 273902
rect 383020 273846 383025 273902
rect 263343 273844 383025 273846
rect 263343 273841 263409 273844
rect 382959 273841 383025 273844
rect 390210 273902 403185 273904
rect 390210 273846 403124 273902
rect 403180 273846 403185 273902
rect 440751 273904 440817 273907
rect 457935 273904 458001 273907
rect 504015 273904 504081 273907
rect 440751 273902 458001 273904
rect 390210 273844 403185 273846
rect 256815 273756 256881 273759
rect 378063 273756 378129 273759
rect 256815 273754 378129 273756
rect 256815 273698 256820 273754
rect 256876 273698 378068 273754
rect 378124 273698 378129 273754
rect 256815 273696 378129 273698
rect 256815 273693 256881 273696
rect 378063 273693 378129 273696
rect 378255 273756 378321 273759
rect 390210 273756 390270 273844
rect 403119 273841 403185 273844
rect 437826 273807 438078 273867
rect 440751 273846 440756 273902
rect 440812 273846 457940 273902
rect 457996 273846 458001 273902
rect 440751 273844 458001 273846
rect 440751 273841 440817 273844
rect 457935 273841 458001 273844
rect 498114 273844 498366 273904
rect 437826 273756 437886 273807
rect 378255 273754 390270 273756
rect 378255 273698 378260 273754
rect 378316 273698 390270 273754
rect 378255 273696 390270 273698
rect 417474 273696 437886 273756
rect 438018 273756 438078 273807
rect 440559 273756 440625 273759
rect 438018 273754 440625 273756
rect 438018 273698 440564 273754
rect 440620 273698 440625 273754
rect 438018 273696 440625 273698
rect 378255 273693 378321 273696
rect 417327 273645 417393 273648
rect 417474 273645 417534 273696
rect 440559 273693 440625 273696
rect 477946 273694 477952 273758
rect 478016 273756 478022 273758
rect 489615 273756 489681 273759
rect 498114 273756 498174 273844
rect 478016 273696 478206 273756
rect 478016 273694 478022 273696
rect 417327 273643 417534 273645
rect 88431 273608 88497 273611
rect 372975 273608 373041 273611
rect 88431 273606 373041 273608
rect 88431 273550 88436 273606
rect 88492 273550 372980 273606
rect 373036 273550 373041 273606
rect 88431 273548 373041 273550
rect 88431 273545 88497 273548
rect 372975 273545 373041 273548
rect 373167 273608 373233 273611
rect 382191 273608 382257 273611
rect 373167 273606 382257 273608
rect 373167 273550 373172 273606
rect 373228 273550 382196 273606
rect 382252 273550 382257 273606
rect 373167 273548 382257 273550
rect 373167 273545 373233 273548
rect 382191 273545 382257 273548
rect 382959 273608 383025 273611
rect 397359 273608 397425 273611
rect 382959 273606 397425 273608
rect 382959 273550 382964 273606
rect 383020 273550 397364 273606
rect 397420 273550 397425 273606
rect 417327 273587 417332 273643
rect 417388 273587 417534 273643
rect 417327 273585 417534 273587
rect 417327 273582 417393 273585
rect 382959 273548 397425 273550
rect 382959 273545 383025 273548
rect 397359 273545 397425 273548
rect 83631 273460 83697 273463
rect 375663 273460 375729 273463
rect 83631 273458 375729 273460
rect 83631 273402 83636 273458
rect 83692 273402 375668 273458
rect 375724 273402 375729 273458
rect 83631 273400 375729 273402
rect 83631 273397 83697 273400
rect 375663 273397 375729 273400
rect 375855 273460 375921 273463
rect 384399 273460 384465 273463
rect 375855 273458 384465 273460
rect 375855 273402 375860 273458
rect 375916 273402 384404 273458
rect 384460 273402 384465 273458
rect 375855 273400 384465 273402
rect 375855 273397 375921 273400
rect 384399 273397 384465 273400
rect 385359 273460 385425 273463
rect 407482 273460 407488 273462
rect 385359 273458 407488 273460
rect 385359 273402 385364 273458
rect 385420 273402 407488 273458
rect 385359 273400 407488 273402
rect 385359 273397 385425 273400
rect 407482 273398 407488 273400
rect 407552 273398 407558 273462
rect 458031 273460 458097 273463
rect 477946 273460 477952 273462
rect 458031 273458 477952 273460
rect 458031 273402 458036 273458
rect 458092 273402 477952 273458
rect 458031 273400 477952 273402
rect 458031 273397 458097 273400
rect 477946 273398 477952 273400
rect 478016 273398 478022 273462
rect 478146 273460 478206 273696
rect 489615 273754 498174 273756
rect 489615 273698 489620 273754
rect 489676 273698 498174 273754
rect 489615 273696 498174 273698
rect 498306 273756 498366 273844
rect 504015 273902 518334 273904
rect 504015 273846 504020 273902
rect 504076 273846 518334 273902
rect 504015 273844 518334 273846
rect 504015 273841 504081 273844
rect 503919 273756 503985 273759
rect 498306 273754 503985 273756
rect 498306 273698 503924 273754
rect 503980 273698 503985 273754
rect 498306 273696 503985 273698
rect 518274 273756 518334 273844
rect 529839 273756 529905 273759
rect 548751 273756 548817 273759
rect 518274 273696 518526 273756
rect 489615 273693 489681 273696
rect 503919 273693 503985 273696
rect 489615 273460 489681 273463
rect 478146 273458 489681 273460
rect 478146 273402 489620 273458
rect 489676 273402 489681 273458
rect 478146 273400 489681 273402
rect 518466 273460 518526 273696
rect 529839 273754 548817 273756
rect 529839 273698 529844 273754
rect 529900 273698 548756 273754
rect 548812 273698 548817 273754
rect 529839 273696 548817 273698
rect 529839 273693 529905 273696
rect 548751 273693 548817 273696
rect 529839 273460 529905 273463
rect 518466 273458 529905 273460
rect 518466 273402 529844 273458
rect 529900 273402 529905 273458
rect 518466 273400 529905 273402
rect 489615 273397 489681 273400
rect 529839 273397 529905 273400
rect 259407 273312 259473 273315
rect 563055 273312 563121 273315
rect 259407 273310 563121 273312
rect 259407 273254 259412 273310
rect 259468 273254 563060 273310
rect 563116 273254 563121 273310
rect 259407 273252 563121 273254
rect 259407 273249 259473 273252
rect 563055 273249 563121 273252
rect 86031 273164 86097 273167
rect 377295 273164 377361 273167
rect 86031 273162 377361 273164
rect 86031 273106 86036 273162
rect 86092 273106 377300 273162
rect 377356 273106 377361 273162
rect 86031 273104 377361 273106
rect 86031 273101 86097 273104
rect 377295 273101 377361 273104
rect 378063 273164 378129 273167
rect 397359 273164 397425 273167
rect 378063 273162 397425 273164
rect 378063 273106 378068 273162
rect 378124 273106 397364 273162
rect 397420 273106 397425 273162
rect 378063 273104 397425 273106
rect 378063 273101 378129 273104
rect 397359 273101 397425 273104
rect 397551 273164 397617 273167
rect 409018 273164 409024 273166
rect 397551 273162 409024 273164
rect 397551 273106 397556 273162
rect 397612 273106 409024 273162
rect 397551 273104 409024 273106
rect 397551 273101 397617 273104
rect 409018 273102 409024 273104
rect 409088 273102 409094 273166
rect 41530 272954 41536 273018
rect 41600 273016 41606 273018
rect 41775 273016 41841 273019
rect 41600 273014 41841 273016
rect 41600 272958 41780 273014
rect 41836 272958 41841 273014
rect 41600 272956 41841 272958
rect 41600 272954 41606 272956
rect 41775 272953 41841 272956
rect 81327 273016 81393 273019
rect 373167 273016 373233 273019
rect 81327 273014 373233 273016
rect 81327 272958 81332 273014
rect 81388 272958 373172 273014
rect 373228 272958 373233 273014
rect 81327 272956 373233 272958
rect 81327 272953 81393 272956
rect 373167 272953 373233 272956
rect 373359 273016 373425 273019
rect 387663 273016 387729 273019
rect 373359 273014 387729 273016
rect 373359 272958 373364 273014
rect 373420 272958 387668 273014
rect 387724 272958 387729 273014
rect 373359 272956 387729 272958
rect 373359 272953 373425 272956
rect 387663 272953 387729 272956
rect 394095 273016 394161 273019
rect 410554 273016 410560 273018
rect 394095 273014 410560 273016
rect 394095 272958 394100 273014
rect 394156 272958 410560 273014
rect 394095 272956 410560 272958
rect 394095 272953 394161 272956
rect 410554 272954 410560 272956
rect 410624 272954 410630 273018
rect 78927 272868 78993 272871
rect 375855 272868 375921 272871
rect 383343 272868 383409 272871
rect 78927 272866 375921 272868
rect 78927 272810 78932 272866
rect 78988 272810 375860 272866
rect 375916 272810 375921 272866
rect 78927 272808 375921 272810
rect 78927 272805 78993 272808
rect 375855 272805 375921 272808
rect 376002 272866 383409 272868
rect 376002 272810 383348 272866
rect 383404 272810 383409 272866
rect 376002 272808 383409 272810
rect 76527 272720 76593 272723
rect 376002 272720 376062 272808
rect 383343 272805 383409 272808
rect 387567 272868 387633 272871
rect 393135 272868 393201 272871
rect 387567 272866 392958 272868
rect 387567 272810 387572 272866
rect 387628 272810 392958 272866
rect 387567 272808 392958 272810
rect 387567 272805 387633 272808
rect 76527 272718 376062 272720
rect 76527 272662 76532 272718
rect 76588 272662 376062 272718
rect 76527 272660 376062 272662
rect 376143 272720 376209 272723
rect 392898 272720 392958 272808
rect 393135 272866 408894 272868
rect 393135 272810 393140 272866
rect 393196 272810 408894 272866
rect 393135 272808 408894 272810
rect 393135 272805 393201 272808
rect 395823 272720 395889 272723
rect 408591 272720 408657 272723
rect 376143 272718 392766 272720
rect 376143 272662 376148 272718
rect 376204 272662 392766 272718
rect 376143 272660 392766 272662
rect 392898 272660 395694 272720
rect 76527 272657 76593 272660
rect 376143 272657 376209 272660
rect 70575 272572 70641 272575
rect 348687 272572 348753 272575
rect 381999 272572 382065 272575
rect 70575 272570 348753 272572
rect 70575 272514 70580 272570
rect 70636 272514 348692 272570
rect 348748 272514 348753 272570
rect 70575 272512 348753 272514
rect 70575 272509 70641 272512
rect 348687 272509 348753 272512
rect 358530 272570 382065 272572
rect 358530 272514 382004 272570
rect 382060 272514 382065 272570
rect 358530 272512 382065 272514
rect 71727 272424 71793 272427
rect 358530 272424 358590 272512
rect 381999 272509 382065 272512
rect 382191 272572 382257 272575
rect 384879 272572 384945 272575
rect 382191 272570 384945 272572
rect 382191 272514 382196 272570
rect 382252 272514 384884 272570
rect 384940 272514 384945 272570
rect 382191 272512 384945 272514
rect 392706 272572 392766 272660
rect 394287 272572 394353 272575
rect 392706 272570 394353 272572
rect 392706 272514 394292 272570
rect 394348 272514 394353 272570
rect 392706 272512 394353 272514
rect 395634 272572 395694 272660
rect 395823 272718 408657 272720
rect 395823 272662 395828 272718
rect 395884 272662 408596 272718
rect 408652 272662 408657 272718
rect 395823 272660 408657 272662
rect 408834 272720 408894 272808
rect 411130 272720 411136 272722
rect 408834 272660 411136 272720
rect 395823 272657 395889 272660
rect 408591 272657 408657 272660
rect 411130 272658 411136 272660
rect 411200 272658 411206 272722
rect 396975 272572 397041 272575
rect 395634 272570 397041 272572
rect 395634 272514 396980 272570
rect 397036 272514 397041 272570
rect 395634 272512 397041 272514
rect 382191 272509 382257 272512
rect 384879 272509 384945 272512
rect 394287 272509 394353 272512
rect 396975 272509 397041 272512
rect 398415 272572 398481 272575
rect 408495 272572 408561 272575
rect 398415 272570 408561 272572
rect 398415 272514 398420 272570
rect 398476 272514 408500 272570
rect 408556 272514 408561 272570
rect 398415 272512 408561 272514
rect 398415 272509 398481 272512
rect 408495 272509 408561 272512
rect 71727 272422 358590 272424
rect 71727 272366 71732 272422
rect 71788 272366 358590 272422
rect 71727 272364 358590 272366
rect 358671 272424 358737 272427
rect 381231 272424 381297 272427
rect 358671 272422 381297 272424
rect 358671 272366 358676 272422
rect 358732 272366 381236 272422
rect 381292 272366 381297 272422
rect 358671 272364 381297 272366
rect 71727 272361 71793 272364
rect 358671 272361 358737 272364
rect 381231 272361 381297 272364
rect 381423 272424 381489 272427
rect 385935 272424 386001 272427
rect 381423 272422 386001 272424
rect 381423 272366 381428 272422
rect 381484 272366 385940 272422
rect 385996 272366 386001 272422
rect 381423 272364 386001 272366
rect 381423 272361 381489 272364
rect 385935 272361 386001 272364
rect 389679 272424 389745 272427
rect 397551 272424 397617 272427
rect 389679 272422 397617 272424
rect 389679 272366 389684 272422
rect 389740 272366 397556 272422
rect 397612 272366 397617 272422
rect 389679 272364 397617 272366
rect 389679 272361 389745 272364
rect 397551 272361 397617 272364
rect 400143 272424 400209 272427
rect 408399 272424 408465 272427
rect 400143 272422 408465 272424
rect 400143 272366 400148 272422
rect 400204 272366 408404 272422
rect 408460 272366 408465 272422
rect 400143 272364 408465 272366
rect 400143 272361 400209 272364
rect 408399 272361 408465 272364
rect 41338 272214 41344 272278
rect 41408 272276 41414 272278
rect 41775 272276 41841 272279
rect 41408 272274 41841 272276
rect 41408 272218 41780 272274
rect 41836 272218 41841 272274
rect 41408 272216 41841 272218
rect 41408 272214 41414 272216
rect 41775 272213 41841 272216
rect 74127 272276 74193 272279
rect 383247 272276 383313 272279
rect 74127 272274 383313 272276
rect 74127 272218 74132 272274
rect 74188 272218 383252 272274
rect 383308 272218 383313 272274
rect 74127 272216 383313 272218
rect 74127 272213 74193 272216
rect 383247 272213 383313 272216
rect 386607 272276 386673 272279
rect 409786 272276 409792 272278
rect 386607 272274 409792 272276
rect 386607 272218 386612 272274
rect 386668 272218 409792 272274
rect 386607 272216 409792 272218
rect 386607 272213 386673 272216
rect 409786 272214 409792 272216
rect 409856 272214 409862 272278
rect 69423 272128 69489 272131
rect 358671 272128 358737 272131
rect 69423 272126 358737 272128
rect 69423 272070 69428 272126
rect 69484 272070 358676 272126
rect 358732 272070 358737 272126
rect 69423 272068 358737 272070
rect 69423 272065 69489 272068
rect 358671 272065 358737 272068
rect 372783 272128 372849 272131
rect 376335 272128 376401 272131
rect 372783 272126 376401 272128
rect 372783 272070 372788 272126
rect 372844 272070 376340 272126
rect 376396 272070 376401 272126
rect 372783 272068 376401 272070
rect 372783 272065 372849 272068
rect 376335 272065 376401 272068
rect 377295 272128 377361 272131
rect 379983 272128 380049 272131
rect 377295 272126 380049 272128
rect 377295 272070 377300 272126
rect 377356 272070 379988 272126
rect 380044 272070 380049 272126
rect 377295 272068 380049 272070
rect 377295 272065 377361 272068
rect 379983 272065 380049 272068
rect 380175 272128 380241 272131
rect 392463 272128 392529 272131
rect 380175 272126 392529 272128
rect 380175 272070 380180 272126
rect 380236 272070 392468 272126
rect 392524 272070 392529 272126
rect 380175 272068 392529 272070
rect 380175 272065 380241 272068
rect 392463 272065 392529 272068
rect 402735 272128 402801 272131
rect 408591 272128 408657 272131
rect 409978 272128 409984 272130
rect 402735 272126 408318 272128
rect 402735 272070 402740 272126
rect 402796 272070 408318 272126
rect 402735 272068 408318 272070
rect 402735 272065 402801 272068
rect 90831 271980 90897 271983
rect 369039 271980 369105 271983
rect 388143 271980 388209 271983
rect 90831 271978 369105 271980
rect 90831 271922 90836 271978
rect 90892 271922 369044 271978
rect 369100 271922 369105 271978
rect 90831 271920 369105 271922
rect 90831 271917 90897 271920
rect 369039 271917 369105 271920
rect 369282 271978 388209 271980
rect 369282 271922 388148 271978
rect 388204 271922 388209 271978
rect 369282 271920 388209 271922
rect 93231 271832 93297 271835
rect 369282 271832 369342 271920
rect 388143 271917 388209 271920
rect 389583 271980 389649 271983
rect 408058 271980 408064 271982
rect 389583 271978 408064 271980
rect 389583 271922 389588 271978
rect 389644 271922 408064 271978
rect 389583 271920 408064 271922
rect 389583 271917 389649 271920
rect 408058 271918 408064 271920
rect 408128 271918 408134 271982
rect 389391 271832 389457 271835
rect 93231 271830 369342 271832
rect 93231 271774 93236 271830
rect 93292 271774 369342 271830
rect 93231 271772 369342 271774
rect 369474 271830 389457 271832
rect 369474 271774 389396 271830
rect 389452 271774 389457 271830
rect 369474 271772 389457 271774
rect 93231 271769 93297 271772
rect 96783 271684 96849 271687
rect 369474 271684 369534 271772
rect 389391 271769 389457 271772
rect 390831 271832 390897 271835
rect 406138 271832 406144 271834
rect 390831 271830 406144 271832
rect 390831 271774 390836 271830
rect 390892 271774 406144 271830
rect 390831 271772 406144 271774
rect 390831 271769 390897 271772
rect 406138 271770 406144 271772
rect 406208 271770 406214 271834
rect 96783 271682 369534 271684
rect 96783 271626 96788 271682
rect 96844 271626 369534 271682
rect 96783 271624 369534 271626
rect 370383 271684 370449 271687
rect 380559 271684 380625 271687
rect 370383 271682 380625 271684
rect 370383 271626 370388 271682
rect 370444 271626 380564 271682
rect 380620 271626 380625 271682
rect 370383 271624 380625 271626
rect 96783 271621 96849 271624
rect 370383 271621 370449 271624
rect 380559 271621 380625 271624
rect 381327 271684 381393 271687
rect 382863 271684 382929 271687
rect 381327 271682 382929 271684
rect 381327 271626 381332 271682
rect 381388 271626 382868 271682
rect 382924 271626 382929 271682
rect 381327 271624 382929 271626
rect 381327 271621 381393 271624
rect 382863 271621 382929 271624
rect 383055 271684 383121 271687
rect 397263 271684 397329 271687
rect 383055 271682 397329 271684
rect 383055 271626 383060 271682
rect 383116 271626 397268 271682
rect 397324 271626 397329 271682
rect 383055 271624 397329 271626
rect 383055 271621 383121 271624
rect 397263 271621 397329 271624
rect 401871 271684 401937 271687
rect 407055 271684 407121 271687
rect 401871 271682 407121 271684
rect 401871 271626 401876 271682
rect 401932 271626 407060 271682
rect 407116 271626 407121 271682
rect 401871 271624 407121 271626
rect 401871 271621 401937 271624
rect 407055 271621 407121 271624
rect 100335 271536 100401 271539
rect 389871 271536 389937 271539
rect 100335 271534 389937 271536
rect 100335 271478 100340 271534
rect 100396 271478 389876 271534
rect 389932 271478 389937 271534
rect 100335 271476 389937 271478
rect 100335 271473 100401 271476
rect 389871 271473 389937 271476
rect 395151 271536 395217 271539
rect 406714 271536 406720 271538
rect 395151 271534 406720 271536
rect 395151 271478 395156 271534
rect 395212 271478 406720 271534
rect 395151 271476 406720 271478
rect 395151 271473 395217 271476
rect 406714 271474 406720 271476
rect 406784 271474 406790 271538
rect 408258 271536 408318 272068
rect 408591 272126 409984 272128
rect 408591 272070 408596 272126
rect 408652 272070 409984 272126
rect 408591 272068 409984 272070
rect 408591 272065 408657 272068
rect 409978 272066 409984 272068
rect 410048 272066 410054 272130
rect 408495 271832 408561 271835
rect 410362 271832 410368 271834
rect 408495 271830 410368 271832
rect 408495 271774 408500 271830
rect 408556 271774 410368 271830
rect 408495 271772 410368 271774
rect 408495 271769 408561 271772
rect 410362 271770 410368 271772
rect 410432 271770 410438 271834
rect 408399 271684 408465 271687
rect 410170 271684 410176 271686
rect 408399 271682 410176 271684
rect 408399 271626 408404 271682
rect 408460 271626 410176 271682
rect 408399 271624 410176 271626
rect 408399 271621 408465 271624
rect 410170 271622 410176 271624
rect 410240 271622 410246 271686
rect 410746 271536 410752 271538
rect 408258 271476 410752 271536
rect 410746 271474 410752 271476
rect 410816 271474 410822 271538
rect 72975 271388 73041 271391
rect 328186 271388 328192 271390
rect 72975 271386 328192 271388
rect 72975 271330 72980 271386
rect 73036 271330 328192 271386
rect 72975 271328 328192 271330
rect 72975 271325 73041 271328
rect 328186 271326 328192 271328
rect 328256 271326 328262 271390
rect 373839 271388 373905 271391
rect 566511 271388 566577 271391
rect 373839 271386 566577 271388
rect 373839 271330 373844 271386
rect 373900 271330 566516 271386
rect 566572 271330 566577 271386
rect 373839 271328 566577 271330
rect 373839 271325 373905 271328
rect 566511 271325 566577 271328
rect 82575 271240 82641 271243
rect 211983 271240 212049 271243
rect 82575 271238 212049 271240
rect 82575 271182 82580 271238
rect 82636 271182 211988 271238
rect 212044 271182 212049 271238
rect 82575 271180 212049 271182
rect 82575 271177 82641 271180
rect 211983 271177 212049 271180
rect 324495 271240 324561 271243
rect 328623 271240 328689 271243
rect 324495 271238 328689 271240
rect 324495 271182 324500 271238
rect 324556 271182 328628 271238
rect 328684 271182 328689 271238
rect 324495 271180 328689 271182
rect 324495 271177 324561 271180
rect 328623 271177 328689 271180
rect 348687 271240 348753 271243
rect 381615 271240 381681 271243
rect 348687 271238 381681 271240
rect 348687 271182 348692 271238
rect 348748 271182 381620 271238
rect 381676 271182 381681 271238
rect 348687 271180 381681 271182
rect 348687 271177 348753 271180
rect 381615 271177 381681 271180
rect 381754 271178 381760 271242
rect 381824 271240 381830 271242
rect 381903 271240 381969 271243
rect 381824 271238 381969 271240
rect 381824 271182 381908 271238
rect 381964 271182 381969 271238
rect 381824 271180 381969 271182
rect 381824 271178 381830 271180
rect 381903 271177 381969 271180
rect 383439 271240 383505 271243
rect 385551 271240 385617 271243
rect 383439 271238 385617 271240
rect 383439 271182 383444 271238
rect 383500 271182 385556 271238
rect 385612 271182 385617 271238
rect 383439 271180 385617 271182
rect 383439 271177 383505 271180
rect 385551 271177 385617 271180
rect 386415 271240 386481 271243
rect 388719 271240 388785 271243
rect 386415 271238 388785 271240
rect 386415 271182 386420 271238
rect 386476 271182 388724 271238
rect 388780 271182 388785 271238
rect 386415 271180 388785 271182
rect 386415 271177 386481 271180
rect 388719 271177 388785 271180
rect 396879 271240 396945 271243
rect 406906 271240 406912 271242
rect 396879 271238 406912 271240
rect 396879 271182 396884 271238
rect 396940 271182 406912 271238
rect 396879 271180 406912 271182
rect 396879 271177 396945 271180
rect 406906 271178 406912 271180
rect 406976 271178 406982 271242
rect 407055 271240 407121 271243
rect 409402 271240 409408 271242
rect 407055 271238 409408 271240
rect 407055 271182 407060 271238
rect 407116 271182 409408 271238
rect 407055 271180 409408 271182
rect 407055 271177 407121 271180
rect 409402 271178 409408 271180
rect 409472 271178 409478 271242
rect 87183 271092 87249 271095
rect 211695 271092 211761 271095
rect 87183 271090 211761 271092
rect 87183 271034 87188 271090
rect 87244 271034 211700 271090
rect 211756 271034 211761 271090
rect 87183 271032 211761 271034
rect 87183 271029 87249 271032
rect 211695 271029 211761 271032
rect 265455 271092 265521 271095
rect 336879 271092 336945 271095
rect 265455 271090 336945 271092
rect 265455 271034 265460 271090
rect 265516 271034 336884 271090
rect 336940 271034 336945 271090
rect 265455 271032 336945 271034
rect 265455 271029 265521 271032
rect 336879 271029 336945 271032
rect 369039 271092 369105 271095
rect 387471 271092 387537 271095
rect 369039 271090 387537 271092
rect 369039 271034 369044 271090
rect 369100 271034 387476 271090
rect 387532 271034 387537 271090
rect 369039 271032 387537 271034
rect 369039 271029 369105 271032
rect 387471 271029 387537 271032
rect 387663 271092 387729 271095
rect 394479 271092 394545 271095
rect 387663 271090 394545 271092
rect 387663 271034 387668 271090
rect 387724 271034 394484 271090
rect 394540 271034 394545 271090
rect 387663 271032 394545 271034
rect 387663 271029 387729 271032
rect 394479 271029 394545 271032
rect 399471 271092 399537 271095
rect 407866 271092 407872 271094
rect 399471 271090 407872 271092
rect 399471 271034 399476 271090
rect 399532 271034 407872 271090
rect 399471 271032 407872 271034
rect 399471 271029 399537 271032
rect 407866 271030 407872 271032
rect 407936 271030 407942 271094
rect 77775 270944 77841 270947
rect 315279 270944 315345 270947
rect 77775 270942 315345 270944
rect 77775 270886 77780 270942
rect 77836 270886 315284 270942
rect 315340 270886 315345 270942
rect 77775 270884 315345 270886
rect 77775 270881 77841 270884
rect 315279 270881 315345 270884
rect 325263 270944 325329 270947
rect 328431 270944 328497 270947
rect 325263 270942 328497 270944
rect 325263 270886 325268 270942
rect 325324 270886 328436 270942
rect 328492 270886 328497 270942
rect 325263 270884 328497 270886
rect 325263 270881 325329 270884
rect 328431 270881 328497 270884
rect 328570 270882 328576 270946
rect 328640 270944 328646 270946
rect 329007 270944 329073 270947
rect 328640 270942 329073 270944
rect 328640 270886 329012 270942
rect 329068 270886 329073 270942
rect 328640 270884 329073 270886
rect 328640 270882 328646 270884
rect 329007 270881 329073 270884
rect 332559 270944 332625 270947
rect 339183 270944 339249 270947
rect 332559 270942 339249 270944
rect 332559 270886 332564 270942
rect 332620 270886 339188 270942
rect 339244 270886 339249 270942
rect 332559 270884 339249 270886
rect 332559 270881 332625 270884
rect 339183 270881 339249 270884
rect 372975 270944 373041 270947
rect 378351 270944 378417 270947
rect 372975 270942 378417 270944
rect 372975 270886 372980 270942
rect 373036 270886 378356 270942
rect 378412 270886 378417 270942
rect 372975 270884 378417 270886
rect 372975 270881 373041 270884
rect 378351 270881 378417 270884
rect 378543 270944 378609 270947
rect 394479 270944 394545 270947
rect 378543 270942 394545 270944
rect 378543 270886 378548 270942
rect 378604 270886 394484 270942
rect 394540 270886 394545 270942
rect 378543 270884 394545 270886
rect 378543 270881 378609 270884
rect 394479 270881 394545 270884
rect 397839 270944 397905 270947
rect 406330 270944 406336 270946
rect 397839 270942 406336 270944
rect 397839 270886 397844 270942
rect 397900 270886 406336 270942
rect 397839 270884 406336 270886
rect 397839 270881 397905 270884
rect 406330 270882 406336 270884
rect 406400 270882 406406 270946
rect 260655 270796 260721 270799
rect 393807 270796 393873 270799
rect 260655 270794 393873 270796
rect 260655 270738 260660 270794
rect 260716 270738 393812 270794
rect 393868 270738 393873 270794
rect 260655 270736 393873 270738
rect 260655 270733 260721 270736
rect 393807 270733 393873 270736
rect 394042 270734 394048 270798
rect 394112 270796 394118 270798
rect 395631 270796 395697 270799
rect 394112 270794 395697 270796
rect 394112 270738 395636 270794
rect 395692 270738 395697 270794
rect 394112 270736 395697 270738
rect 394112 270734 394118 270736
rect 395631 270733 395697 270736
rect 395770 270734 395776 270798
rect 395840 270796 395846 270798
rect 395919 270796 395985 270799
rect 395840 270794 395985 270796
rect 395840 270738 395924 270794
rect 395980 270738 395985 270794
rect 395840 270736 395985 270738
rect 395840 270734 395846 270736
rect 395919 270733 395985 270736
rect 401199 270796 401265 270799
rect 406522 270796 406528 270798
rect 401199 270794 406528 270796
rect 401199 270738 401204 270794
rect 401260 270738 406528 270794
rect 401199 270736 406528 270738
rect 401199 270733 401265 270736
rect 406522 270734 406528 270736
rect 406592 270734 406598 270798
rect 429135 270796 429201 270799
rect 449199 270796 449265 270799
rect 429135 270794 449265 270796
rect 429135 270738 429140 270794
rect 429196 270738 449204 270794
rect 449260 270738 449265 270794
rect 429135 270736 449265 270738
rect 429135 270733 429201 270736
rect 449199 270733 449265 270736
rect 40954 270586 40960 270650
rect 41024 270648 41030 270650
rect 41775 270648 41841 270651
rect 41024 270646 41841 270648
rect 41024 270590 41780 270646
rect 41836 270590 41841 270646
rect 41024 270588 41841 270590
rect 41024 270586 41030 270588
rect 41775 270585 41841 270588
rect 41914 270586 41920 270650
rect 41984 270648 41990 270650
rect 43119 270648 43185 270651
rect 41984 270646 43185 270648
rect 41984 270590 43124 270646
rect 43180 270590 43185 270646
rect 41984 270588 43185 270590
rect 41984 270586 41990 270588
rect 43119 270585 43185 270588
rect 201519 270648 201585 270651
rect 317487 270648 317553 270651
rect 201519 270646 317553 270648
rect 201519 270590 201524 270646
rect 201580 270590 317492 270646
rect 317548 270590 317553 270646
rect 201519 270588 317553 270590
rect 201519 270585 201585 270588
rect 317487 270585 317553 270588
rect 317679 270648 317745 270651
rect 325263 270648 325329 270651
rect 317679 270646 325329 270648
rect 317679 270590 317684 270646
rect 317740 270590 325268 270646
rect 325324 270590 325329 270646
rect 317679 270588 325329 270590
rect 317679 270585 317745 270588
rect 325263 270585 325329 270588
rect 325455 270648 325521 270651
rect 634287 270648 634353 270651
rect 325455 270646 634353 270648
rect 325455 270590 325460 270646
rect 325516 270590 634292 270646
rect 634348 270590 634353 270646
rect 325455 270588 634353 270590
rect 325455 270585 325521 270588
rect 634287 270585 634353 270588
rect 258927 270500 258993 270503
rect 370479 270500 370545 270503
rect 370671 270502 370737 270503
rect 258927 270498 370545 270500
rect 258927 270442 258932 270498
rect 258988 270442 370484 270498
rect 370540 270442 370545 270498
rect 258927 270440 370545 270442
rect 258927 270437 258993 270440
rect 370479 270437 370545 270440
rect 370618 270438 370624 270502
rect 370688 270500 370737 270502
rect 370863 270500 370929 270503
rect 371194 270500 371200 270502
rect 370688 270498 370780 270500
rect 370732 270442 370780 270498
rect 370688 270440 370780 270442
rect 370863 270498 371200 270500
rect 370863 270442 370868 270498
rect 370924 270442 371200 270498
rect 370863 270440 371200 270442
rect 370688 270438 370737 270440
rect 370671 270437 370737 270438
rect 370863 270437 370929 270440
rect 371194 270438 371200 270440
rect 371264 270438 371270 270502
rect 371439 270500 371505 270503
rect 371578 270500 371584 270502
rect 371439 270498 371584 270500
rect 371439 270442 371444 270498
rect 371500 270442 371584 270498
rect 371439 270440 371584 270442
rect 371439 270437 371505 270440
rect 371578 270438 371584 270440
rect 371648 270438 371654 270502
rect 371727 270500 371793 270503
rect 378543 270500 378609 270503
rect 371727 270498 378609 270500
rect 371727 270442 371732 270498
rect 371788 270442 378548 270498
rect 378604 270442 378609 270498
rect 371727 270440 378609 270442
rect 371727 270437 371793 270440
rect 378543 270437 378609 270440
rect 378831 270500 378897 270503
rect 379215 270500 379281 270503
rect 378831 270498 379281 270500
rect 378831 270442 378836 270498
rect 378892 270442 379220 270498
rect 379276 270442 379281 270498
rect 378831 270440 379281 270442
rect 378831 270437 378897 270440
rect 379215 270437 379281 270440
rect 379407 270500 379473 270503
rect 388623 270500 388689 270503
rect 379407 270498 388689 270500
rect 379407 270442 379412 270498
rect 379468 270442 388628 270498
rect 388684 270442 388689 270498
rect 379407 270440 388689 270442
rect 379407 270437 379473 270440
rect 388623 270437 388689 270440
rect 388815 270500 388881 270503
rect 440655 270500 440721 270503
rect 388815 270498 440721 270500
rect 388815 270442 388820 270498
rect 388876 270442 440660 270498
rect 440716 270442 440721 270498
rect 388815 270440 440721 270442
rect 388815 270437 388881 270440
rect 440655 270437 440721 270440
rect 460719 270500 460785 270503
rect 544431 270500 544497 270503
rect 460719 270498 544497 270500
rect 460719 270442 460724 270498
rect 460780 270442 544436 270498
rect 544492 270442 544497 270498
rect 460719 270440 544497 270442
rect 460719 270437 460785 270440
rect 544431 270437 544497 270440
rect 564399 270500 564465 270503
rect 623055 270500 623121 270503
rect 564399 270498 623121 270500
rect 564399 270442 564404 270498
rect 564460 270442 623060 270498
rect 623116 270442 623121 270498
rect 564399 270440 623121 270442
rect 564399 270437 564465 270440
rect 623055 270437 623121 270440
rect 318159 270352 318225 270355
rect 338703 270352 338769 270355
rect 469071 270352 469137 270355
rect 318159 270350 338622 270352
rect 318159 270294 318164 270350
rect 318220 270294 338622 270350
rect 318159 270292 338622 270294
rect 318159 270289 318225 270292
rect 318927 270204 318993 270207
rect 338562 270204 338622 270292
rect 338703 270350 469137 270352
rect 338703 270294 338708 270350
rect 338764 270294 469076 270350
rect 469132 270294 469137 270350
rect 338703 270292 469137 270294
rect 338703 270289 338769 270292
rect 469071 270289 469137 270292
rect 469551 270352 469617 270355
rect 499503 270352 499569 270355
rect 469551 270350 499569 270352
rect 469551 270294 469556 270350
rect 469612 270294 499508 270350
rect 499564 270294 499569 270350
rect 469551 270292 499569 270294
rect 469551 270289 469617 270292
rect 499503 270289 499569 270292
rect 499642 270290 499648 270354
rect 499712 270352 499718 270354
rect 509487 270352 509553 270355
rect 519471 270352 519537 270355
rect 499712 270350 509553 270352
rect 499712 270294 509492 270350
rect 509548 270294 509553 270350
rect 499712 270292 509553 270294
rect 499712 270290 499718 270292
rect 509487 270289 509553 270292
rect 509634 270350 519537 270352
rect 509634 270294 519476 270350
rect 519532 270294 519537 270350
rect 509634 270292 519537 270294
rect 469359 270204 469425 270207
rect 318927 270202 338430 270204
rect 318927 270146 318932 270202
rect 318988 270146 338430 270202
rect 318927 270144 338430 270146
rect 338562 270202 469425 270204
rect 338562 270146 469364 270202
rect 469420 270146 469425 270202
rect 338562 270144 469425 270146
rect 318927 270141 318993 270144
rect 41146 269994 41152 270058
rect 41216 270056 41222 270058
rect 41775 270056 41841 270059
rect 41216 270054 41841 270056
rect 41216 269998 41780 270054
rect 41836 269998 41841 270054
rect 41216 269996 41841 269998
rect 41216 269994 41222 269996
rect 41775 269993 41841 269996
rect 268143 270056 268209 270059
rect 314415 270056 314481 270059
rect 268143 270054 314481 270056
rect 268143 269998 268148 270054
rect 268204 269998 314420 270054
rect 314476 269998 314481 270054
rect 268143 269996 314481 269998
rect 268143 269993 268209 269996
rect 314415 269993 314481 269996
rect 320175 270056 320241 270059
rect 338370 270056 338430 270144
rect 469359 270141 469425 270144
rect 469551 270204 469617 270207
rect 499695 270204 499761 270207
rect 469551 270202 499761 270204
rect 469551 270146 469556 270202
rect 469612 270146 499700 270202
rect 499756 270146 499761 270202
rect 469551 270144 499761 270146
rect 469551 270141 469617 270144
rect 499695 270141 499761 270144
rect 428943 270056 429009 270059
rect 320175 270054 338238 270056
rect 320175 269998 320180 270054
rect 320236 269998 338238 270054
rect 320175 269996 338238 269998
rect 338370 270054 429009 270056
rect 338370 269998 428948 270054
rect 429004 269998 429009 270054
rect 338370 269996 429009 269998
rect 320175 269993 320241 269996
rect 261999 269908 262065 269911
rect 318063 269908 318129 269911
rect 261999 269906 318129 269908
rect 261999 269850 262004 269906
rect 262060 269850 318068 269906
rect 318124 269850 318129 269906
rect 261999 269848 318129 269850
rect 261999 269845 262065 269848
rect 318063 269845 318129 269848
rect 319695 269908 319761 269911
rect 327183 269908 327249 269911
rect 319695 269906 327249 269908
rect 319695 269850 319700 269906
rect 319756 269850 327188 269906
rect 327244 269850 327249 269906
rect 319695 269848 327249 269850
rect 319695 269845 319761 269848
rect 327183 269845 327249 269848
rect 328431 269908 328497 269911
rect 338031 269908 338097 269911
rect 328431 269906 338097 269908
rect 328431 269850 328436 269906
rect 328492 269850 338036 269906
rect 338092 269850 338097 269906
rect 328431 269848 338097 269850
rect 338178 269908 338238 269996
rect 428943 269993 429009 269996
rect 429231 270056 429297 270059
rect 469167 270056 469233 270059
rect 429231 270054 469233 270056
rect 429231 269998 429236 270054
rect 429292 269998 469172 270054
rect 469228 269998 469233 270054
rect 429231 269996 469233 269998
rect 429231 269993 429297 269996
rect 469167 269993 469233 269996
rect 469647 270056 469713 270059
rect 499599 270056 499665 270059
rect 469647 270054 499665 270056
rect 469647 269998 469652 270054
rect 469708 269998 499604 270054
rect 499660 269998 499665 270054
rect 469647 269996 499665 269998
rect 469647 269993 469713 269996
rect 499599 269993 499665 269996
rect 499791 270056 499857 270059
rect 509634 270056 509694 270292
rect 519471 270289 519537 270292
rect 519663 270352 519729 270355
rect 582063 270352 582129 270355
rect 519663 270350 582129 270352
rect 519663 270294 519668 270350
rect 519724 270294 582068 270350
rect 582124 270294 582129 270350
rect 519663 270292 582129 270294
rect 519663 270289 519729 270292
rect 582063 270289 582129 270292
rect 519855 270204 519921 270207
rect 589167 270204 589233 270207
rect 519855 270202 589233 270204
rect 519855 270146 519860 270202
rect 519916 270146 589172 270202
rect 589228 270146 589233 270202
rect 519855 270144 589233 270146
rect 519855 270141 519921 270144
rect 589167 270141 589233 270144
rect 499791 270054 509694 270056
rect 499791 269998 499796 270054
rect 499852 269998 509694 270054
rect 499791 269996 509694 269998
rect 519759 270056 519825 270059
rect 596367 270056 596433 270059
rect 519759 270054 596433 270056
rect 519759 269998 519764 270054
rect 519820 269998 596372 270054
rect 596428 269998 596433 270054
rect 519759 269996 596433 269998
rect 499791 269993 499857 269996
rect 519759 269993 519825 269996
rect 596367 269993 596433 269996
rect 674415 270056 674481 270059
rect 674415 270054 674784 270056
rect 674415 269998 674420 270054
rect 674476 269998 674784 270054
rect 674415 269996 674784 269998
rect 674415 269993 674481 269996
rect 429039 269908 429105 269911
rect 338178 269906 429105 269908
rect 338178 269850 429044 269906
rect 429100 269850 429105 269906
rect 338178 269848 429105 269850
rect 328431 269845 328497 269848
rect 338031 269845 338097 269848
rect 429039 269845 429105 269848
rect 449199 269908 449265 269911
rect 469263 269908 469329 269911
rect 449199 269906 469329 269908
rect 449199 269850 449204 269906
rect 449260 269850 469268 269906
rect 469324 269850 469329 269906
rect 449199 269848 469329 269850
rect 449199 269845 449265 269848
rect 469263 269845 469329 269848
rect 529839 269908 529905 269911
rect 603375 269908 603441 269911
rect 529839 269906 603441 269908
rect 529839 269850 529844 269906
rect 529900 269850 603380 269906
rect 603436 269850 603441 269906
rect 529839 269848 603441 269850
rect 529839 269845 529905 269848
rect 603375 269845 603441 269848
rect 261135 269760 261201 269763
rect 577263 269760 577329 269763
rect 261135 269758 577329 269760
rect 261135 269702 261140 269758
rect 261196 269702 577268 269758
rect 577324 269702 577329 269758
rect 261135 269700 577329 269702
rect 261135 269697 261201 269700
rect 577263 269697 577329 269700
rect 674703 269760 674769 269763
rect 674703 269758 674814 269760
rect 674703 269702 674708 269758
rect 674764 269702 674814 269758
rect 674703 269697 674814 269702
rect 264879 269612 264945 269615
rect 605775 269612 605841 269615
rect 264879 269610 605841 269612
rect 264879 269554 264884 269610
rect 264940 269554 605780 269610
rect 605836 269554 605841 269610
rect 674754 269582 674814 269697
rect 264879 269552 605841 269554
rect 264879 269549 264945 269552
rect 605775 269549 605841 269552
rect 266607 269464 266673 269467
rect 620079 269464 620145 269467
rect 266607 269462 620145 269464
rect 266607 269406 266612 269462
rect 266668 269406 620084 269462
rect 620140 269406 620145 269462
rect 266607 269404 620145 269406
rect 266607 269401 266673 269404
rect 620079 269401 620145 269404
rect 267663 269316 267729 269319
rect 630831 269316 630897 269319
rect 267663 269314 630897 269316
rect 267663 269258 267668 269314
rect 267724 269258 630836 269314
rect 630892 269258 630897 269314
rect 267663 269256 630897 269258
rect 267663 269253 267729 269256
rect 630831 269253 630897 269256
rect 40762 269106 40768 269170
rect 40832 269168 40838 269170
rect 41775 269168 41841 269171
rect 40832 269166 41841 269168
rect 40832 269110 41780 269166
rect 41836 269110 41841 269166
rect 40832 269108 41841 269110
rect 40832 269106 40838 269108
rect 41775 269105 41841 269108
rect 253359 269168 253425 269171
rect 513039 269168 513105 269171
rect 253359 269166 513105 269168
rect 253359 269110 253364 269166
rect 253420 269110 513044 269166
rect 513100 269110 513105 269166
rect 253359 269108 513105 269110
rect 253359 269105 253425 269108
rect 513039 269105 513105 269108
rect 519471 269168 519537 269171
rect 529839 269168 529905 269171
rect 519471 269166 529905 269168
rect 519471 269110 519476 269166
rect 519532 269110 529844 269166
rect 529900 269110 529905 269166
rect 519471 269108 529905 269110
rect 519471 269105 519537 269108
rect 529839 269105 529905 269108
rect 674703 269168 674769 269171
rect 674703 269166 674814 269168
rect 674703 269110 674708 269166
rect 674764 269110 674814 269166
rect 674703 269105 674814 269110
rect 260559 269020 260625 269023
rect 371247 269020 371313 269023
rect 260559 269018 371313 269020
rect 260559 268962 260564 269018
rect 260620 268962 371252 269018
rect 371308 268962 371313 269018
rect 260559 268960 371313 268962
rect 260559 268957 260625 268960
rect 371247 268957 371313 268960
rect 371439 269020 371505 269023
rect 379791 269020 379857 269023
rect 379983 269022 380049 269023
rect 379983 269020 380032 269022
rect 371439 269018 379857 269020
rect 371439 268962 371444 269018
rect 371500 268962 379796 269018
rect 379852 268962 379857 269018
rect 371439 268960 379857 268962
rect 379940 269018 380032 269020
rect 379940 268962 379988 269018
rect 379940 268960 380032 268962
rect 371439 268957 371505 268960
rect 379791 268957 379857 268960
rect 379983 268958 380032 268960
rect 380096 268958 380102 269022
rect 380271 269020 380337 269023
rect 640335 269020 640401 269023
rect 380271 269018 640401 269020
rect 380271 268962 380276 269018
rect 380332 268962 640340 269018
rect 640396 268962 640401 269018
rect 674754 268990 674814 269105
rect 380271 268960 640401 268962
rect 379983 268957 380049 268958
rect 380271 268957 380337 268960
rect 640335 268957 640401 268960
rect 316719 268872 316785 268875
rect 574863 268872 574929 268875
rect 316719 268870 574929 268872
rect 316719 268814 316724 268870
rect 316780 268814 574868 268870
rect 574924 268814 574929 268870
rect 316719 268812 574929 268814
rect 316719 268809 316785 268812
rect 574863 268809 574929 268812
rect 252879 268724 252945 268727
rect 499450 268724 499456 268726
rect 252879 268722 499456 268724
rect 252879 268666 252884 268722
rect 252940 268666 499456 268722
rect 252879 268664 499456 268666
rect 252879 268661 252945 268664
rect 499450 268662 499456 268664
rect 499520 268662 499526 268726
rect 499599 268724 499665 268727
rect 519759 268724 519825 268727
rect 499599 268722 519825 268724
rect 499599 268666 499604 268722
rect 499660 268666 519764 268722
rect 519820 268666 519825 268722
rect 499599 268664 519825 268666
rect 499599 268661 499665 268664
rect 519759 268661 519825 268664
rect 677242 268662 677248 268726
rect 677312 268662 677318 268726
rect 255855 268576 255921 268579
rect 276346 268576 276352 268578
rect 255855 268574 276352 268576
rect 255855 268518 255860 268574
rect 255916 268518 276352 268574
rect 255855 268516 276352 268518
rect 255855 268513 255921 268516
rect 276346 268514 276352 268516
rect 276416 268514 276422 268578
rect 297999 268576 298065 268579
rect 317679 268576 317745 268579
rect 297999 268574 317745 268576
rect 297999 268518 298004 268574
rect 298060 268518 317684 268574
rect 317740 268518 317745 268574
rect 297999 268516 317745 268518
rect 297999 268513 298065 268516
rect 317679 268513 317745 268516
rect 317871 268576 317937 268579
rect 567759 268576 567825 268579
rect 317871 268574 567825 268576
rect 317871 268518 317876 268574
rect 317932 268518 567764 268574
rect 567820 268518 567825 268574
rect 317871 268516 567825 268518
rect 317871 268513 317937 268516
rect 567759 268513 567825 268516
rect 252015 268428 252081 268431
rect 499407 268428 499473 268431
rect 252015 268426 499473 268428
rect 252015 268370 252020 268426
rect 252076 268370 499412 268426
rect 499468 268370 499473 268426
rect 252015 268368 499473 268370
rect 252015 268365 252081 268368
rect 499407 268365 499473 268368
rect 499695 268428 499761 268431
rect 519855 268428 519921 268431
rect 499695 268426 519921 268428
rect 499695 268370 499700 268426
rect 499756 268370 519860 268426
rect 519916 268370 519921 268426
rect 677250 268398 677310 268662
rect 499695 268368 519921 268370
rect 499695 268365 499761 268368
rect 519855 268365 519921 268368
rect 211503 268280 211569 268283
rect 254607 268280 254673 268283
rect 211503 268278 254673 268280
rect 211503 268222 211508 268278
rect 211564 268222 254612 268278
rect 254668 268222 254673 268278
rect 211503 268220 254673 268222
rect 211503 268217 211569 268220
rect 254607 268217 254673 268220
rect 265071 268280 265137 268283
rect 377103 268280 377169 268283
rect 265071 268278 377169 268280
rect 265071 268222 265076 268278
rect 265132 268222 377108 268278
rect 377164 268222 377169 268278
rect 265071 268220 377169 268222
rect 265071 268217 265137 268220
rect 377103 268217 377169 268220
rect 377338 268218 377344 268282
rect 377408 268280 377414 268282
rect 388719 268280 388785 268283
rect 377408 268278 388785 268280
rect 377408 268222 388724 268278
rect 388780 268222 388785 268278
rect 377408 268220 388785 268222
rect 377408 268218 377414 268220
rect 388719 268217 388785 268220
rect 388911 268280 388977 268283
rect 403695 268280 403761 268283
rect 388911 268278 403761 268280
rect 388911 268222 388916 268278
rect 388972 268222 403700 268278
rect 403756 268222 403761 268278
rect 388911 268220 403761 268222
rect 388911 268217 388977 268220
rect 403695 268217 403761 268220
rect 403887 268280 403953 268283
rect 404602 268280 404608 268282
rect 403887 268278 404608 268280
rect 403887 268222 403892 268278
rect 403948 268222 404608 268278
rect 403887 268220 404608 268222
rect 403887 268217 403953 268220
rect 404602 268218 404608 268220
rect 404672 268218 404678 268282
rect 404847 268280 404913 268283
rect 405562 268280 405568 268282
rect 404847 268278 405568 268280
rect 404847 268222 404852 268278
rect 404908 268222 405568 268278
rect 404847 268220 405568 268222
rect 404847 268217 404913 268220
rect 405562 268218 405568 268220
rect 405632 268218 405638 268282
rect 405711 268280 405777 268283
rect 405946 268280 405952 268282
rect 405711 268278 405952 268280
rect 405711 268222 405716 268278
rect 405772 268222 405952 268278
rect 405711 268220 405952 268222
rect 405711 268217 405777 268220
rect 405946 268218 405952 268220
rect 406016 268218 406022 268282
rect 406095 268280 406161 268283
rect 626031 268280 626097 268283
rect 406095 268278 626097 268280
rect 406095 268222 406100 268278
rect 406156 268222 626036 268278
rect 626092 268222 626097 268278
rect 406095 268220 626097 268222
rect 406095 268217 406161 268220
rect 626031 268217 626097 268220
rect 250287 268132 250353 268135
rect 488079 268132 488145 268135
rect 250287 268130 488145 268132
rect 250287 268074 250292 268130
rect 250348 268074 488084 268130
rect 488140 268074 488145 268130
rect 250287 268072 488145 268074
rect 250287 268069 250353 268072
rect 488079 268069 488145 268072
rect 488271 268132 488337 268135
rect 499311 268132 499377 268135
rect 488271 268130 499377 268132
rect 488271 268074 488276 268130
rect 488332 268074 499316 268130
rect 499372 268074 499377 268130
rect 488271 268072 499377 268074
rect 488271 268069 488337 268072
rect 499311 268069 499377 268072
rect 499503 268132 499569 268135
rect 519663 268132 519729 268135
rect 499503 268130 519729 268132
rect 499503 268074 499508 268130
rect 499564 268074 519668 268130
rect 519724 268074 519729 268130
rect 499503 268072 519729 268074
rect 499503 268069 499569 268072
rect 519663 268069 519729 268072
rect 212271 267984 212337 267987
rect 263727 267984 263793 267987
rect 212271 267982 263793 267984
rect 212271 267926 212276 267982
rect 212332 267926 263732 267982
rect 263788 267926 263793 267982
rect 212271 267924 263793 267926
rect 212271 267921 212337 267924
rect 263727 267921 263793 267924
rect 269199 267984 269265 267987
rect 297999 267984 298065 267987
rect 269199 267982 298065 267984
rect 269199 267926 269204 267982
rect 269260 267926 298004 267982
rect 298060 267926 298065 267982
rect 269199 267924 298065 267926
rect 269199 267921 269265 267924
rect 297999 267921 298065 267924
rect 298191 267984 298257 267987
rect 315855 267984 315921 267987
rect 317871 267984 317937 267987
rect 298191 267982 300606 267984
rect 298191 267926 298196 267982
rect 298252 267926 300606 267982
rect 298191 267924 300606 267926
rect 298191 267921 298257 267924
rect 255087 267836 255153 267839
rect 256623 267836 256689 267839
rect 267759 267836 267825 267839
rect 276207 267836 276273 267839
rect 255087 267834 255294 267836
rect 255087 267778 255092 267834
rect 255148 267778 255294 267834
rect 255087 267776 255294 267778
rect 255087 267773 255153 267776
rect 255234 267688 255294 267776
rect 256623 267834 267825 267836
rect 256623 267778 256628 267834
rect 256684 267778 267764 267834
rect 267820 267778 267825 267834
rect 256623 267776 267825 267778
rect 256623 267773 256689 267776
rect 267759 267773 267825 267776
rect 276162 267834 276273 267836
rect 276162 267778 276212 267834
rect 276268 267778 276273 267834
rect 276162 267773 276273 267778
rect 297807 267836 297873 267839
rect 298383 267836 298449 267839
rect 297807 267834 298449 267836
rect 297807 267778 297812 267834
rect 297868 267778 298388 267834
rect 298444 267778 298449 267834
rect 297807 267776 298449 267778
rect 300546 267836 300606 267924
rect 315855 267982 317937 267984
rect 315855 267926 315860 267982
rect 315916 267926 317876 267982
rect 317932 267926 317937 267982
rect 315855 267924 317937 267926
rect 315855 267921 315921 267924
rect 317871 267921 317937 267924
rect 318063 267984 318129 267987
rect 325743 267984 325809 267987
rect 318063 267982 325809 267984
rect 318063 267926 318068 267982
rect 318124 267926 325748 267982
rect 325804 267926 325809 267982
rect 318063 267924 325809 267926
rect 318063 267921 318129 267924
rect 325743 267921 325809 267924
rect 327087 267984 327153 267987
rect 327226 267984 327232 267986
rect 327087 267982 327232 267984
rect 327087 267926 327092 267982
rect 327148 267926 327232 267982
rect 327087 267924 327232 267926
rect 327087 267921 327153 267924
rect 327226 267922 327232 267924
rect 327296 267922 327302 267986
rect 329146 267922 329152 267986
rect 329216 267984 329222 267986
rect 336207 267984 336273 267987
rect 329216 267982 336273 267984
rect 329216 267926 336212 267982
rect 336268 267926 336273 267982
rect 329216 267924 336273 267926
rect 329216 267922 329222 267924
rect 336207 267921 336273 267924
rect 336399 267984 336465 267987
rect 560655 267984 560721 267987
rect 336399 267982 560721 267984
rect 336399 267926 336404 267982
rect 336460 267926 560660 267982
rect 560716 267926 560721 267982
rect 336399 267924 560721 267926
rect 336399 267921 336465 267924
rect 560655 267921 560721 267924
rect 300546 267776 371070 267836
rect 297807 267773 297873 267776
rect 298383 267773 298449 267776
rect 276162 267688 276222 267773
rect 255234 267628 276222 267688
rect 276346 267626 276352 267690
rect 276416 267688 276422 267690
rect 328762 267688 328768 267690
rect 276416 267628 328768 267688
rect 276416 267626 276422 267628
rect 328762 267626 328768 267628
rect 328832 267626 328838 267690
rect 352762 267626 352768 267690
rect 352832 267688 352838 267690
rect 370810 267688 370816 267690
rect 352832 267628 370816 267688
rect 352832 267626 352838 267628
rect 370810 267626 370816 267628
rect 370880 267626 370886 267690
rect 371010 267688 371070 267776
rect 371194 267774 371200 267838
rect 371264 267836 371270 267838
rect 377146 267836 377152 267838
rect 371264 267776 377152 267836
rect 371264 267774 371270 267776
rect 377146 267774 377152 267776
rect 377216 267774 377222 267838
rect 377391 267836 377457 267839
rect 388815 267836 388881 267839
rect 377391 267834 388881 267836
rect 377391 267778 377396 267834
rect 377452 267778 388820 267834
rect 388876 267778 388881 267834
rect 377391 267776 388881 267778
rect 377391 267773 377457 267776
rect 388815 267773 388881 267776
rect 389007 267838 389073 267839
rect 389007 267834 389056 267838
rect 389120 267836 389126 267838
rect 389007 267778 389012 267834
rect 389007 267774 389056 267778
rect 389120 267776 389164 267836
rect 389295 267834 389361 267839
rect 389295 267778 389300 267834
rect 389356 267778 389361 267834
rect 389120 267774 389126 267776
rect 389007 267773 389073 267774
rect 389295 267773 389361 267778
rect 397551 267836 397617 267839
rect 413103 267836 413169 267839
rect 397551 267834 413169 267836
rect 397551 267778 397556 267834
rect 397612 267778 413108 267834
rect 413164 267778 413169 267834
rect 397551 267776 413169 267778
rect 397551 267773 397617 267776
rect 413103 267773 413169 267776
rect 413295 267836 413361 267839
rect 614223 267836 614289 267839
rect 413295 267834 614289 267836
rect 413295 267778 413300 267834
rect 413356 267778 614228 267834
rect 614284 267778 614289 267834
rect 413295 267776 614289 267778
rect 413295 267773 413361 267776
rect 614223 267773 614289 267776
rect 389298 267688 389358 267773
rect 371010 267628 389358 267688
rect 389434 267626 389440 267690
rect 389504 267688 389510 267690
rect 639087 267688 639153 267691
rect 677250 267690 677310 267880
rect 389504 267686 639153 267688
rect 389504 267630 639092 267686
rect 639148 267630 639153 267686
rect 389504 267628 639153 267630
rect 389504 267626 389510 267628
rect 639087 267625 639153 267628
rect 677242 267626 677248 267690
rect 677312 267626 677318 267690
rect 677434 267478 677440 267542
rect 677504 267478 677510 267542
rect 677442 267392 677502 267478
rect 676896 267362 677502 267392
rect 676866 267332 677472 267362
rect 676866 267098 676926 267332
rect 676858 267034 676864 267098
rect 676928 267034 676934 267098
rect 677050 267034 677056 267098
rect 677120 267034 677126 267098
rect 677058 266770 677118 267034
rect 674511 266060 674577 266063
rect 674754 266060 674814 266252
rect 674511 266058 674814 266060
rect 674511 266002 674516 266058
rect 674572 266002 674814 266058
rect 674511 266000 674814 266002
rect 674511 265997 674577 266000
rect 413391 265912 413457 265915
rect 609423 265912 609489 265915
rect 413391 265910 609489 265912
rect 413391 265854 413396 265910
rect 413452 265854 609428 265910
rect 609484 265854 609489 265910
rect 413391 265852 609489 265854
rect 413391 265849 413457 265852
rect 609423 265849 609489 265852
rect 413103 265616 413169 265619
rect 628431 265616 628497 265619
rect 413103 265614 628497 265616
rect 413103 265558 413108 265614
rect 413164 265558 628436 265614
rect 628492 265558 628497 265614
rect 413103 265556 628497 265558
rect 413103 265553 413169 265556
rect 628431 265553 628497 265556
rect 677058 265471 677118 265734
rect 412815 265468 412881 265471
rect 632079 265468 632145 265471
rect 412815 265466 632145 265468
rect 412815 265410 412820 265466
rect 412876 265410 632084 265466
rect 632140 265410 632145 265466
rect 412815 265408 632145 265410
rect 677058 265466 677169 265471
rect 677058 265410 677108 265466
rect 677164 265410 677169 265466
rect 677058 265408 677169 265410
rect 412815 265405 412881 265408
rect 632079 265405 632145 265408
rect 677103 265405 677169 265408
rect 412911 265320 412977 265323
rect 527343 265320 527409 265323
rect 412911 265318 527409 265320
rect 412911 265262 412916 265318
rect 412972 265262 527348 265318
rect 527404 265262 527409 265318
rect 412911 265260 527409 265262
rect 412911 265257 412977 265260
rect 527343 265257 527409 265260
rect 412719 265172 412785 265175
rect 530895 265172 530961 265175
rect 412719 265170 530961 265172
rect 412719 265114 412724 265170
rect 412780 265114 530900 265170
rect 530956 265114 530961 265170
rect 412719 265112 530961 265114
rect 412719 265109 412785 265112
rect 530895 265109 530961 265112
rect 675138 265027 675198 265142
rect 412623 265024 412689 265027
rect 537999 265024 538065 265027
rect 412623 265022 538065 265024
rect 412623 264966 412628 265022
rect 412684 264966 538004 265022
rect 538060 264966 538065 265022
rect 412623 264964 538065 264966
rect 675138 265022 675249 265027
rect 675138 264966 675188 265022
rect 675244 264966 675249 265022
rect 675138 264964 675249 264966
rect 412623 264961 412689 264964
rect 537999 264961 538065 264964
rect 675183 264961 675249 264964
rect 378927 264913 378993 264916
rect 378882 264911 378993 264913
rect 267855 264876 267921 264879
rect 276495 264876 276561 264879
rect 267855 264874 276561 264876
rect 267855 264818 267860 264874
rect 267916 264818 276500 264874
rect 276556 264818 276561 264874
rect 267855 264816 276561 264818
rect 267855 264813 267921 264816
rect 276495 264813 276561 264816
rect 308079 264876 308145 264879
rect 378882 264876 378932 264911
rect 308079 264874 378932 264876
rect 308079 264818 308084 264874
rect 308140 264855 378932 264874
rect 378988 264855 378993 264911
rect 385071 264911 385137 264916
rect 308140 264850 378993 264855
rect 379119 264876 379185 264879
rect 385071 264876 385076 264911
rect 379119 264874 385076 264876
rect 308140 264818 378942 264850
rect 308079 264816 378942 264818
rect 379119 264818 379124 264874
rect 379180 264855 385076 264874
rect 385132 264855 385137 264911
rect 379180 264850 385137 264855
rect 406479 264913 406545 264916
rect 407247 264913 407313 264916
rect 406479 264911 406590 264913
rect 406479 264855 406484 264911
rect 406540 264876 406590 264911
rect 407247 264911 407358 264913
rect 407098 264876 407104 264878
rect 406540 264855 407104 264876
rect 406479 264850 407104 264855
rect 379180 264818 385134 264850
rect 379119 264816 385134 264818
rect 406530 264816 407104 264850
rect 308079 264813 308145 264816
rect 379119 264813 379185 264816
rect 407098 264814 407104 264816
rect 407168 264814 407174 264878
rect 407247 264855 407252 264911
rect 407308 264855 407358 264911
rect 407727 264911 407793 264916
rect 407727 264878 407732 264911
rect 407247 264850 407358 264855
rect 407098 264518 407104 264582
rect 407168 264580 407174 264582
rect 407298 264580 407358 264850
rect 407674 264814 407680 264878
rect 407788 264855 407793 264911
rect 407744 264850 407793 264855
rect 408111 264911 408177 264916
rect 408111 264855 408116 264911
rect 408172 264855 408177 264911
rect 408783 264913 408849 264916
rect 409551 264913 409617 264916
rect 410799 264913 410865 264916
rect 411183 264913 411249 264916
rect 408783 264911 408894 264913
rect 408111 264850 408177 264855
rect 407744 264816 407790 264850
rect 407744 264814 407750 264816
rect 408114 264728 408174 264850
rect 408250 264814 408256 264878
rect 408320 264876 408326 264878
rect 408783 264876 408788 264911
rect 408320 264855 408788 264876
rect 408844 264855 408894 264911
rect 408320 264816 408894 264855
rect 409551 264911 409662 264913
rect 409551 264855 409556 264911
rect 409612 264878 409662 264911
rect 410754 264911 410865 264913
rect 409551 264850 409600 264855
rect 408320 264814 408326 264816
rect 409594 264814 409600 264850
rect 409664 264814 409670 264878
rect 410754 264855 410804 264911
rect 410860 264855 410865 264911
rect 411138 264911 411249 264913
rect 410754 264850 410865 264855
rect 408442 264728 408448 264730
rect 408114 264668 408448 264728
rect 408442 264666 408448 264668
rect 408512 264666 408518 264730
rect 410754 264728 410814 264850
rect 410938 264814 410944 264878
rect 411008 264876 411014 264878
rect 411138 264876 411188 264911
rect 411008 264855 411188 264876
rect 411244 264855 411249 264911
rect 411008 264850 411249 264855
rect 413295 264876 413361 264879
rect 555855 264876 555921 264879
rect 413295 264874 555921 264876
rect 411008 264816 411198 264850
rect 413295 264818 413300 264874
rect 413356 264818 555860 264874
rect 555916 264818 555921 264874
rect 413295 264816 555921 264818
rect 411008 264814 411014 264816
rect 413295 264813 413361 264816
rect 555855 264813 555921 264816
rect 411322 264728 411328 264730
rect 410754 264668 411328 264728
rect 411322 264666 411328 264668
rect 411392 264666 411398 264730
rect 407168 264520 407358 264580
rect 407168 264518 407174 264520
rect 675138 264435 675198 264624
rect 675087 264430 675198 264435
rect 675087 264374 675092 264430
rect 675148 264374 675198 264430
rect 675087 264372 675198 264374
rect 675087 264369 675153 264372
rect 674170 264074 674176 264138
rect 674240 264136 674246 264138
rect 674240 264076 674784 264136
rect 674240 264074 674246 264076
rect 676866 263251 676926 263514
rect 676866 263246 676977 263251
rect 676866 263190 676916 263246
rect 676972 263190 676977 263246
rect 676866 263188 676977 263190
rect 676911 263185 676977 263188
rect 675330 262807 675390 262996
rect 675279 262802 675390 262807
rect 675279 262746 675284 262802
rect 675340 262746 675390 262802
rect 675279 262744 675390 262746
rect 675279 262741 675345 262744
rect 674319 262508 674385 262511
rect 674319 262506 674784 262508
rect 674319 262450 674324 262506
rect 674380 262450 674784 262506
rect 674319 262448 674784 262450
rect 674319 262445 674385 262448
rect 207183 261324 207249 261327
rect 211842 261324 211902 261812
rect 674754 261771 674814 261886
rect 674754 261766 674865 261771
rect 674754 261710 674804 261766
rect 674860 261710 674865 261766
rect 674754 261708 674865 261710
rect 674799 261705 674865 261708
rect 207183 261322 211902 261324
rect 207183 261266 207188 261322
rect 207244 261266 211902 261322
rect 207183 261264 211902 261266
rect 207183 261261 207249 261264
rect 674754 261179 674814 261368
rect 674703 261174 674814 261179
rect 674703 261118 674708 261174
rect 674764 261118 674814 261174
rect 674703 261116 674814 261118
rect 674703 261113 674769 261116
rect 674127 260880 674193 260883
rect 674127 260878 674784 260880
rect 674127 260822 674132 260878
rect 674188 260822 674784 260878
rect 674127 260820 674784 260822
rect 674127 260817 674193 260820
rect 674946 260143 675006 260258
rect 674895 260138 675006 260143
rect 674895 260082 674900 260138
rect 674956 260082 675006 260138
rect 674895 260080 675006 260082
rect 674895 260077 674961 260080
rect 42543 259696 42609 259699
rect 42498 259694 42609 259696
rect 42498 259638 42548 259694
rect 42604 259638 42609 259694
rect 42498 259633 42609 259638
rect 42498 259518 42558 259633
rect 674607 259548 674673 259551
rect 674754 259548 674814 259740
rect 674607 259546 674814 259548
rect 674607 259490 674612 259546
rect 674668 259490 674814 259546
rect 674607 259488 674814 259490
rect 674607 259485 674673 259488
rect 674946 258959 675006 259222
rect 42639 258956 42705 258959
rect 42528 258954 42705 258956
rect 42528 258898 42644 258954
rect 42700 258898 42705 258954
rect 42528 258896 42705 258898
rect 674946 258954 675057 258959
rect 674946 258898 674996 258954
rect 675052 258898 675057 258954
rect 674946 258896 675057 258898
rect 42639 258893 42705 258896
rect 674991 258893 675057 258896
rect 677058 258367 677118 258630
rect 677007 258362 677118 258367
rect 42498 258219 42558 258334
rect 677007 258306 677012 258362
rect 677068 258306 677118 258362
rect 677007 258304 677118 258306
rect 677007 258301 677073 258304
rect 42498 258214 42609 258219
rect 42498 258158 42548 258214
rect 42604 258158 42609 258214
rect 42498 258156 42609 258158
rect 42543 258153 42609 258156
rect 42306 257624 42366 257890
rect 676866 257775 676926 258112
rect 676815 257770 676926 257775
rect 676815 257714 676820 257770
rect 676876 257714 676926 257770
rect 676815 257712 676926 257714
rect 677007 257772 677073 257775
rect 677007 257770 677118 257772
rect 677007 257714 677012 257770
rect 677068 257714 677118 257770
rect 676815 257709 676881 257712
rect 677007 257709 677118 257714
rect 42543 257624 42609 257627
rect 42306 257622 42609 257624
rect 42306 257566 42548 257622
rect 42604 257566 42609 257622
rect 677058 257594 677118 257709
rect 42306 257564 42609 257566
rect 42543 257561 42609 257564
rect 43215 257328 43281 257331
rect 42528 257326 43281 257328
rect 42528 257270 43220 257326
rect 43276 257270 43281 257326
rect 42528 257268 43281 257270
rect 43215 257265 43281 257268
rect 676815 257328 676881 257331
rect 676815 257326 676926 257328
rect 676815 257270 676820 257326
rect 676876 257270 676926 257326
rect 676815 257265 676926 257270
rect 40378 256970 40384 257034
rect 40448 256970 40454 257034
rect 676866 257002 676926 257265
rect 40386 256736 40446 256970
rect 43407 256736 43473 256739
rect 40386 256734 43473 256736
rect 40386 256706 43412 256734
rect 40416 256678 43412 256706
rect 43468 256678 43473 256734
rect 40416 256676 43473 256678
rect 43407 256673 43473 256676
rect 42298 256378 42304 256442
rect 42368 256378 42374 256442
rect 42306 256292 42366 256378
rect 42306 256262 42528 256292
rect 42336 256232 42558 256262
rect 42498 255848 42558 256232
rect 43311 255848 43377 255851
rect 42498 255846 43377 255848
rect 42498 255790 43316 255846
rect 43372 255790 43377 255846
rect 42498 255788 43377 255790
rect 43311 255785 43377 255788
rect 40578 255406 40638 255670
rect 40570 255342 40576 255406
rect 40640 255342 40646 255406
rect 207279 255404 207345 255407
rect 211842 255404 211902 255880
rect 207279 255402 211902 255404
rect 207279 255346 207284 255402
rect 207340 255346 211902 255402
rect 207279 255344 211902 255346
rect 207279 255341 207345 255344
rect 43023 255108 43089 255111
rect 42528 255106 43089 255108
rect 42528 255050 43028 255106
rect 43084 255050 43089 255106
rect 42528 255048 43089 255050
rect 43023 255045 43089 255048
rect 40386 254222 40446 254560
rect 40378 254158 40384 254222
rect 40448 254158 40454 254222
rect 40770 253778 40830 254042
rect 40762 253714 40768 253778
rect 40832 253714 40838 253778
rect 41346 253334 41406 253450
rect 41338 253270 41344 253334
rect 41408 253270 41414 253334
rect 675706 253270 675712 253334
rect 675776 253332 675782 253334
rect 676911 253332 676977 253335
rect 675776 253330 676977 253332
rect 675776 253274 676916 253330
rect 676972 253274 676977 253330
rect 675776 253272 676977 253274
rect 675776 253270 675782 253272
rect 676911 253269 676977 253272
rect 675898 253122 675904 253186
rect 675968 253184 675974 253186
rect 677103 253184 677169 253187
rect 675968 253182 677169 253184
rect 675968 253126 677108 253182
rect 677164 253126 677169 253182
rect 675968 253124 677169 253126
rect 675968 253122 675974 253124
rect 677103 253121 677169 253124
rect 41730 252595 41790 252932
rect 41730 252590 41841 252595
rect 41730 252534 41780 252590
rect 41836 252534 41841 252590
rect 41730 252532 41841 252534
rect 41775 252529 41841 252532
rect 40962 252150 41022 252414
rect 40954 252086 40960 252150
rect 41024 252086 41030 252150
rect 41154 251558 41214 251822
rect 41146 251494 41152 251558
rect 41216 251494 41222 251558
rect 41538 251114 41598 251304
rect 41530 251050 41536 251114
rect 41600 251050 41606 251114
rect 40194 250523 40254 250786
rect 40194 250518 40305 250523
rect 40194 250462 40244 250518
rect 40300 250462 40305 250518
rect 40194 250460 40305 250462
rect 40239 250457 40305 250460
rect 40002 249931 40062 250194
rect 39951 249926 40062 249931
rect 39951 249870 39956 249926
rect 40012 249870 40062 249926
rect 39951 249868 40062 249870
rect 39951 249865 40017 249868
rect 40002 249339 40062 249676
rect 40002 249334 40113 249339
rect 40002 249278 40052 249334
rect 40108 249278 40113 249334
rect 40002 249276 40113 249278
rect 40047 249273 40113 249276
rect 207087 249336 207153 249339
rect 211842 249336 211902 249896
rect 207087 249334 211902 249336
rect 207087 249278 207092 249334
rect 207148 249278 211902 249334
rect 207087 249276 211902 249278
rect 207087 249273 207153 249276
rect 40194 248895 40254 249158
rect 40143 248890 40254 248895
rect 40143 248834 40148 248890
rect 40204 248834 40254 248890
rect 40143 248832 40254 248834
rect 40143 248829 40209 248832
rect 43119 248596 43185 248599
rect 42528 248594 43185 248596
rect 42528 248538 43124 248594
rect 43180 248538 43185 248594
rect 42528 248536 43185 248538
rect 43119 248533 43185 248536
rect 42498 247859 42558 248048
rect 42498 247854 42609 247859
rect 407674 247856 407680 247858
rect 42498 247798 42548 247854
rect 42604 247798 42609 247854
rect 42498 247796 42609 247798
rect 42543 247793 42609 247796
rect 406914 247796 407680 247856
rect 163983 247708 164049 247711
rect 187215 247708 187281 247711
rect 163983 247706 187281 247708
rect 163983 247650 163988 247706
rect 164044 247650 187220 247706
rect 187276 247650 187281 247706
rect 163983 247648 187281 247650
rect 163983 247645 164049 247648
rect 187215 247645 187281 247648
rect 196911 247708 196977 247711
rect 208719 247708 208785 247711
rect 196911 247706 208785 247708
rect 196911 247650 196916 247706
rect 196972 247650 208724 247706
rect 208780 247650 208785 247706
rect 196911 247648 208785 247650
rect 196911 247645 196977 247648
rect 208719 247645 208785 247648
rect 175503 247560 175569 247563
rect 197391 247560 197457 247563
rect 405946 247560 405952 247562
rect 175503 247558 197310 247560
rect 35202 247267 35262 247530
rect 175503 247502 175508 247558
rect 175564 247502 197310 247558
rect 175503 247500 197310 247502
rect 175503 247497 175569 247500
rect 181263 247412 181329 247415
rect 196911 247412 196977 247415
rect 181263 247410 196977 247412
rect 181263 247354 181268 247410
rect 181324 247354 196916 247410
rect 196972 247354 196977 247410
rect 181263 247352 196977 247354
rect 197250 247412 197310 247500
rect 197391 247558 405952 247560
rect 197391 247502 197396 247558
rect 197452 247502 405952 247558
rect 197391 247500 405952 247502
rect 197391 247497 197457 247500
rect 405946 247498 405952 247500
rect 406016 247498 406022 247562
rect 406914 247560 406974 247796
rect 407674 247794 407680 247796
rect 407744 247794 407750 247858
rect 408442 247646 408448 247710
rect 408512 247708 408518 247710
rect 410938 247708 410944 247710
rect 408512 247648 410944 247708
rect 408512 247646 408518 247648
rect 410938 247646 410944 247648
rect 411008 247646 411014 247710
rect 406098 247500 406974 247560
rect 406098 247412 406158 247500
rect 409594 247412 409600 247414
rect 197250 247352 225918 247412
rect 181263 247349 181329 247352
rect 196911 247349 196977 247352
rect 35202 247262 35313 247267
rect 42543 247264 42609 247267
rect 35202 247206 35252 247262
rect 35308 247206 35313 247262
rect 35202 247204 35313 247206
rect 35247 247201 35313 247204
rect 42498 247262 42609 247264
rect 42498 247206 42548 247262
rect 42604 247206 42609 247262
rect 42498 247201 42609 247206
rect 187023 247264 187089 247267
rect 196911 247264 196977 247267
rect 187023 247262 196977 247264
rect 187023 247206 187028 247262
rect 187084 247206 196916 247262
rect 196972 247206 196977 247262
rect 187023 247204 196977 247206
rect 187023 247201 187089 247204
rect 196911 247201 196977 247204
rect 210114 247204 225534 247264
rect 42498 246938 42558 247201
rect 181359 247118 181425 247119
rect 181306 247116 181312 247118
rect 146562 247079 146814 247116
rect 146946 247079 166782 247116
rect 146562 247056 166782 247079
rect 181268 247056 181312 247116
rect 181376 247114 181425 247118
rect 181420 247058 181425 247114
rect 35247 246820 35313 246823
rect 146562 246820 146622 247056
rect 146754 247019 147006 247056
rect 35202 246818 35313 246820
rect 35202 246762 35252 246818
rect 35308 246762 35313 246818
rect 35202 246757 35313 246762
rect 106626 246760 146622 246820
rect 166722 246820 166782 247056
rect 181306 247054 181312 247056
rect 181376 247054 181425 247058
rect 181359 247053 181425 247054
rect 187215 247116 187281 247119
rect 197007 247116 197073 247119
rect 187215 247114 197073 247116
rect 187215 247058 187220 247114
rect 187276 247058 197012 247114
rect 197068 247058 197073 247114
rect 187215 247056 197073 247058
rect 187215 247053 187281 247056
rect 197007 247053 197073 247056
rect 207226 247054 207232 247118
rect 207296 247116 207302 247118
rect 210114 247116 210174 247204
rect 207296 247056 210174 247116
rect 210351 247116 210417 247119
rect 210351 247114 225342 247116
rect 210351 247058 210356 247114
rect 210412 247058 225342 247114
rect 210351 247056 225342 247058
rect 207296 247054 207302 247056
rect 210351 247053 210417 247056
rect 166863 246968 166929 246971
rect 166863 246966 224766 246968
rect 166863 246910 166868 246966
rect 166924 246910 224766 246966
rect 166863 246908 224766 246910
rect 166863 246905 166929 246908
rect 210159 246820 210225 246823
rect 223119 246820 223185 246823
rect 166722 246818 210225 246820
rect 166722 246762 210164 246818
rect 210220 246762 210225 246818
rect 166722 246760 210225 246762
rect 35202 246420 35262 246757
rect 80463 246672 80529 246675
rect 48450 246670 80529 246672
rect 48450 246614 80468 246670
rect 80524 246614 80529 246670
rect 48450 246612 80529 246614
rect 42874 246462 42880 246526
rect 42944 246524 42950 246526
rect 48450 246524 48510 246612
rect 80463 246609 80529 246612
rect 86511 246672 86577 246675
rect 106626 246672 106686 246760
rect 210159 246757 210225 246760
rect 210498 246818 223185 246820
rect 210498 246762 223124 246818
rect 223180 246762 223185 246818
rect 210498 246760 223185 246762
rect 224706 246820 224766 246908
rect 225282 246823 225342 247056
rect 225474 246968 225534 247204
rect 225858 247116 225918 247352
rect 227442 247352 406158 247412
rect 406386 247352 409600 247412
rect 227442 247116 227502 247352
rect 406386 247264 406446 247352
rect 409594 247350 409600 247352
rect 409664 247350 409670 247414
rect 225858 247056 227502 247116
rect 227586 247204 367806 247264
rect 225474 246908 226110 246968
rect 224847 246820 224913 246823
rect 224706 246818 224913 246820
rect 224706 246762 224852 246818
rect 224908 246762 224913 246818
rect 224706 246760 224913 246762
rect 225282 246818 225393 246823
rect 225282 246762 225332 246818
rect 225388 246762 225393 246818
rect 225282 246760 225393 246762
rect 226050 246820 226110 246908
rect 227586 246820 227646 247204
rect 228210 247056 367230 247116
rect 228210 246968 228270 247056
rect 228162 246908 228270 246968
rect 228354 246908 246462 246968
rect 228162 246823 228222 246908
rect 228354 246823 228414 246908
rect 246402 246823 246462 246908
rect 248178 246908 285006 246968
rect 248178 246823 248238 246908
rect 284946 246823 285006 246908
rect 285378 246908 307950 246968
rect 226050 246760 227646 246820
rect 228111 246818 228222 246823
rect 228111 246762 228116 246818
rect 228172 246762 228222 246818
rect 228111 246760 228222 246762
rect 228303 246818 228414 246823
rect 228303 246762 228308 246818
rect 228364 246762 228414 246818
rect 228303 246760 228414 246762
rect 228591 246820 228657 246823
rect 246159 246820 246225 246823
rect 228591 246818 246225 246820
rect 228591 246762 228596 246818
rect 228652 246762 246164 246818
rect 246220 246762 246225 246818
rect 228591 246760 246225 246762
rect 246402 246818 246513 246823
rect 246402 246762 246452 246818
rect 246508 246762 246513 246818
rect 246402 246760 246513 246762
rect 86511 246670 106686 246672
rect 86511 246614 86516 246670
rect 86572 246614 106686 246670
rect 86511 246612 106686 246614
rect 172719 246672 172785 246675
rect 207226 246672 207232 246674
rect 172719 246670 207232 246672
rect 172719 246614 172724 246670
rect 172780 246614 207232 246670
rect 172719 246612 207232 246614
rect 86511 246609 86577 246612
rect 172719 246609 172785 246612
rect 207226 246610 207232 246612
rect 207296 246610 207302 246674
rect 42944 246464 48510 246524
rect 53679 246524 53745 246527
rect 197295 246524 197361 246527
rect 210255 246524 210321 246527
rect 53679 246522 197361 246524
rect 53679 246466 53684 246522
rect 53740 246466 197300 246522
rect 197356 246466 197361 246522
rect 53679 246464 197361 246466
rect 42944 246462 42950 246464
rect 53679 246461 53745 246464
rect 197295 246461 197361 246464
rect 197442 246522 210321 246524
rect 197442 246466 210260 246522
rect 210316 246466 210321 246522
rect 197442 246464 210321 246466
rect 53295 246376 53361 246379
rect 196719 246376 196785 246379
rect 53295 246374 196785 246376
rect 53295 246318 53300 246374
rect 53356 246318 196724 246374
rect 196780 246318 196785 246374
rect 53295 246316 196785 246318
rect 53295 246313 53361 246316
rect 196719 246313 196785 246316
rect 196911 246376 196977 246379
rect 197442 246376 197502 246464
rect 210255 246461 210321 246464
rect 196911 246374 197502 246376
rect 196911 246318 196916 246374
rect 196972 246318 197502 246374
rect 196911 246316 197502 246318
rect 197583 246376 197649 246379
rect 210351 246376 210417 246379
rect 197583 246374 210417 246376
rect 197583 246318 197588 246374
rect 197644 246318 210356 246374
rect 210412 246318 210417 246374
rect 197583 246316 210417 246318
rect 196911 246313 196977 246316
rect 197583 246313 197649 246316
rect 210351 246313 210417 246316
rect 44655 246228 44721 246231
rect 197199 246228 197265 246231
rect 44655 246226 197265 246228
rect 44655 246170 44660 246226
rect 44716 246170 197204 246226
rect 197260 246170 197265 246226
rect 44655 246168 197265 246170
rect 44655 246165 44721 246168
rect 197199 246165 197265 246168
rect 65103 246080 65169 246083
rect 210351 246080 210417 246083
rect 65103 246078 210417 246080
rect 65103 246022 65108 246078
rect 65164 246022 210356 246078
rect 210412 246022 210417 246078
rect 65103 246020 210417 246022
rect 65103 246017 65169 246020
rect 210351 246017 210417 246020
rect 181359 245934 181425 245935
rect 181306 245932 181312 245934
rect 181268 245872 181312 245932
rect 181376 245930 181425 245934
rect 181420 245874 181425 245930
rect 181306 245870 181312 245872
rect 181376 245870 181425 245874
rect 181359 245869 181425 245870
rect 189999 245932 190065 245935
rect 197583 245932 197649 245935
rect 189999 245930 197649 245932
rect 189999 245874 190004 245930
rect 190060 245874 197588 245930
rect 197644 245874 197649 245930
rect 189999 245872 197649 245874
rect 189999 245869 190065 245872
rect 197583 245869 197649 245872
rect 149583 245784 149649 245787
rect 210351 245784 210417 245787
rect 149583 245782 210417 245784
rect 149583 245726 149588 245782
rect 149644 245726 210356 245782
rect 210412 245726 210417 245782
rect 149583 245724 210417 245726
rect 149583 245721 149649 245724
rect 210351 245721 210417 245724
rect 197199 245636 197265 245639
rect 210351 245636 210417 245639
rect 197199 245634 210417 245636
rect 197199 245578 197204 245634
rect 197260 245578 210356 245634
rect 210412 245578 210417 245634
rect 197199 245576 210417 245578
rect 197199 245573 197265 245576
rect 210351 245573 210417 245576
rect 155343 245488 155409 245491
rect 210498 245488 210558 246760
rect 223119 246757 223185 246760
rect 224847 246757 224913 246760
rect 225327 246757 225393 246760
rect 228111 246757 228177 246760
rect 228303 246757 228369 246760
rect 228591 246757 228657 246760
rect 246159 246757 246225 246760
rect 246447 246757 246513 246760
rect 247311 246820 247377 246823
rect 247791 246820 247857 246823
rect 247311 246818 247857 246820
rect 247311 246762 247316 246818
rect 247372 246762 247796 246818
rect 247852 246762 247857 246818
rect 247311 246760 247857 246762
rect 247311 246757 247377 246760
rect 247791 246757 247857 246760
rect 248175 246818 248241 246823
rect 248175 246762 248180 246818
rect 248236 246762 248241 246818
rect 248175 246757 248241 246762
rect 248367 246820 248433 246823
rect 260943 246820 261009 246823
rect 248367 246818 261009 246820
rect 248367 246762 248372 246818
rect 248428 246762 260948 246818
rect 261004 246762 261009 246818
rect 248367 246760 261009 246762
rect 248367 246757 248433 246760
rect 260943 246757 261009 246760
rect 269199 246820 269265 246823
rect 281295 246820 281361 246823
rect 269199 246818 281361 246820
rect 269199 246762 269204 246818
rect 269260 246762 281300 246818
rect 281356 246762 281361 246818
rect 269199 246760 281361 246762
rect 269199 246757 269265 246760
rect 281295 246757 281361 246760
rect 284943 246818 285009 246823
rect 284943 246762 284948 246818
rect 285004 246762 285009 246818
rect 284943 246757 285009 246762
rect 285231 246820 285297 246823
rect 285378 246820 285438 246908
rect 307890 246823 307950 246908
rect 308082 246908 328590 246968
rect 308082 246823 308142 246908
rect 328530 246823 328590 246908
rect 328962 246908 348606 246968
rect 328962 246823 329022 246908
rect 348546 246823 348606 246908
rect 349074 246908 366846 246968
rect 349074 246823 349134 246908
rect 366786 246823 366846 246908
rect 285231 246818 285438 246820
rect 285231 246762 285236 246818
rect 285292 246762 285438 246818
rect 285231 246760 285438 246762
rect 287535 246820 287601 246823
rect 307407 246820 307473 246823
rect 287535 246818 307473 246820
rect 287535 246762 287540 246818
rect 287596 246762 307412 246818
rect 307468 246762 307473 246818
rect 287535 246760 307473 246762
rect 285231 246757 285297 246760
rect 287535 246757 287601 246760
rect 307407 246757 307473 246760
rect 307887 246818 307953 246823
rect 307887 246762 307892 246818
rect 307948 246762 307953 246818
rect 307887 246757 307953 246762
rect 308079 246818 308145 246823
rect 308079 246762 308084 246818
rect 308140 246762 308145 246818
rect 308079 246757 308145 246762
rect 311151 246820 311217 246823
rect 328335 246820 328401 246823
rect 311151 246818 328401 246820
rect 311151 246762 311156 246818
rect 311212 246762 328340 246818
rect 328396 246762 328401 246818
rect 311151 246760 328401 246762
rect 311151 246757 311217 246760
rect 328335 246757 328401 246760
rect 328527 246818 328593 246823
rect 328527 246762 328532 246818
rect 328588 246762 328593 246818
rect 328527 246757 328593 246762
rect 328911 246818 329022 246823
rect 328911 246762 328916 246818
rect 328972 246762 329022 246818
rect 328911 246760 329022 246762
rect 329295 246820 329361 246823
rect 342543 246820 342609 246823
rect 329295 246818 342609 246820
rect 329295 246762 329300 246818
rect 329356 246762 342548 246818
rect 342604 246762 342609 246818
rect 329295 246760 342609 246762
rect 348546 246818 348657 246823
rect 348546 246762 348596 246818
rect 348652 246762 348657 246818
rect 348546 246760 348657 246762
rect 328911 246757 328977 246760
rect 329295 246757 329361 246760
rect 342543 246757 342609 246760
rect 348591 246757 348657 246760
rect 349071 246818 349137 246823
rect 349071 246762 349076 246818
rect 349132 246762 349137 246818
rect 349071 246757 349137 246762
rect 349647 246820 349713 246823
rect 366447 246820 366513 246823
rect 349647 246818 366513 246820
rect 349647 246762 349652 246818
rect 349708 246762 366452 246818
rect 366508 246762 366513 246818
rect 349647 246760 366513 246762
rect 366786 246818 366897 246823
rect 366786 246762 366836 246818
rect 366892 246762 366897 246818
rect 366786 246760 366897 246762
rect 367170 246820 367230 247056
rect 367311 246820 367377 246823
rect 367170 246818 367377 246820
rect 367170 246762 367316 246818
rect 367372 246762 367377 246818
rect 367170 246760 367377 246762
rect 367746 246820 367806 247204
rect 370434 247204 406446 247264
rect 369519 246820 369585 246823
rect 367746 246818 369585 246820
rect 367746 246762 369524 246818
rect 369580 246762 369585 246818
rect 367746 246760 369585 246762
rect 349647 246757 349713 246760
rect 366447 246757 366513 246760
rect 366831 246757 366897 246760
rect 367311 246757 367377 246760
rect 369519 246757 369585 246760
rect 370287 246820 370353 246823
rect 370434 246820 370494 247204
rect 407866 247202 407872 247266
rect 407936 247264 407942 247266
rect 408634 247264 408640 247266
rect 407936 247204 408640 247264
rect 407936 247202 407942 247204
rect 408634 247202 408640 247204
rect 408704 247202 408710 247266
rect 410746 247202 410752 247266
rect 410816 247264 410822 247266
rect 412143 247264 412209 247267
rect 410816 247262 412209 247264
rect 410816 247206 412148 247262
rect 412204 247206 412209 247262
rect 410816 247204 412209 247206
rect 410816 247202 410822 247204
rect 412143 247201 412209 247204
rect 407098 247116 407104 247118
rect 370818 247056 407104 247116
rect 370287 246818 370494 246820
rect 370287 246762 370292 246818
rect 370348 246762 370494 246818
rect 370287 246760 370494 246762
rect 370671 246820 370737 246823
rect 370818 246820 370878 247056
rect 407098 247054 407104 247056
rect 407168 247054 407174 247118
rect 408442 247116 408448 247118
rect 407874 247056 408448 247116
rect 405562 246968 405568 246970
rect 373458 246908 389070 246968
rect 373458 246823 373518 246908
rect 389010 246823 389070 246908
rect 389298 246908 405568 246968
rect 389298 246823 389358 246908
rect 405562 246906 405568 246908
rect 405632 246906 405638 246970
rect 406714 246968 406720 246970
rect 406338 246908 406720 246968
rect 406338 246823 406398 246908
rect 406714 246906 406720 246908
rect 406784 246906 406790 246970
rect 406906 246906 406912 246970
rect 406976 246968 406982 246970
rect 406976 246908 407166 246968
rect 406976 246906 406982 246908
rect 370671 246818 370878 246820
rect 370671 246762 370676 246818
rect 370732 246762 370878 246818
rect 370671 246760 370878 246762
rect 373455 246818 373521 246823
rect 373455 246762 373460 246818
rect 373516 246762 373521 246818
rect 370287 246757 370353 246760
rect 370671 246757 370737 246760
rect 373455 246757 373521 246762
rect 389007 246818 389073 246823
rect 389007 246762 389012 246818
rect 389068 246762 389073 246818
rect 389007 246757 389073 246762
rect 389295 246818 389361 246823
rect 389295 246762 389300 246818
rect 389356 246762 389361 246818
rect 389295 246757 389361 246762
rect 390255 246820 390321 246823
rect 405903 246820 405969 246823
rect 406095 246822 406161 246823
rect 406095 246820 406144 246822
rect 390255 246818 405969 246820
rect 390255 246762 390260 246818
rect 390316 246762 405908 246818
rect 405964 246762 405969 246818
rect 390255 246760 405969 246762
rect 406052 246818 406144 246820
rect 406052 246762 406100 246818
rect 406052 246760 406144 246762
rect 390255 246757 390321 246760
rect 405903 246757 405969 246760
rect 406095 246758 406144 246760
rect 406208 246758 406214 246822
rect 406338 246818 406449 246823
rect 406767 246822 406833 246823
rect 406338 246762 406388 246818
rect 406444 246762 406449 246818
rect 406338 246760 406449 246762
rect 406095 246757 406161 246758
rect 406383 246757 406449 246760
rect 406522 246758 406528 246822
rect 406592 246820 406598 246822
rect 406592 246786 406638 246820
rect 406592 246781 406641 246786
rect 406575 246725 406580 246758
rect 406636 246725 406641 246781
rect 406714 246758 406720 246822
rect 406784 246820 406833 246822
rect 406959 246820 407025 246823
rect 407106 246820 407166 246908
rect 406784 246818 406876 246820
rect 406828 246762 406876 246818
rect 406784 246760 406876 246762
rect 406959 246818 407166 246820
rect 406959 246762 406964 246818
rect 407020 246762 407166 246818
rect 406959 246760 407166 246762
rect 407343 246820 407409 246823
rect 407482 246820 407488 246822
rect 407343 246818 407488 246820
rect 407343 246762 407348 246818
rect 407404 246762 407488 246818
rect 407343 246760 407488 246762
rect 406784 246758 406833 246760
rect 406767 246757 406833 246758
rect 406959 246757 407025 246760
rect 407343 246757 407409 246760
rect 407482 246758 407488 246760
rect 407552 246758 407558 246822
rect 407727 246820 407793 246823
rect 407874 246820 407934 247056
rect 408442 247054 408448 247056
rect 408512 247054 408518 247118
rect 409786 247054 409792 247118
rect 409856 247116 409862 247118
rect 409856 247056 410814 247116
rect 409856 247054 409862 247056
rect 409402 246968 409408 246970
rect 407727 246818 407934 246820
rect 407727 246762 407732 246818
rect 407788 246762 407934 246818
rect 407727 246760 407934 246762
rect 408066 246908 409408 246968
rect 408066 246823 408126 246908
rect 409402 246906 409408 246908
rect 409472 246906 409478 246970
rect 410170 246906 410176 246970
rect 410240 246968 410246 246970
rect 410240 246908 410622 246968
rect 410240 246906 410246 246908
rect 410562 246823 410622 246908
rect 408066 246818 408177 246823
rect 408066 246762 408116 246818
rect 408172 246762 408177 246818
rect 408066 246760 408177 246762
rect 407727 246757 407793 246760
rect 408111 246757 408177 246760
rect 408303 246820 408369 246823
rect 408634 246820 408640 246822
rect 408303 246818 408640 246820
rect 408303 246762 408308 246818
rect 408364 246762 408640 246818
rect 408303 246760 408640 246762
rect 408303 246757 408369 246760
rect 408634 246758 408640 246760
rect 408704 246758 408710 246822
rect 408975 246820 409041 246823
rect 410319 246822 410385 246823
rect 409978 246820 409984 246822
rect 408975 246818 409984 246820
rect 408975 246762 408980 246818
rect 409036 246762 409984 246818
rect 408975 246760 409984 246762
rect 408975 246757 409041 246760
rect 409978 246758 409984 246760
rect 410048 246758 410054 246822
rect 410319 246820 410368 246822
rect 410276 246818 410368 246820
rect 410276 246762 410324 246818
rect 410276 246760 410368 246762
rect 410319 246758 410368 246760
rect 410432 246758 410438 246822
rect 410511 246818 410622 246823
rect 410511 246762 410516 246818
rect 410572 246762 410622 246818
rect 410511 246760 410622 246762
rect 410754 246823 410814 247056
rect 411130 246906 411136 246970
rect 411200 246968 411206 246970
rect 411200 246908 411774 246968
rect 411200 246906 411206 246908
rect 411714 246823 411774 246908
rect 410754 246818 410865 246823
rect 410754 246762 410804 246818
rect 410860 246762 410865 246818
rect 410754 246760 410865 246762
rect 410319 246757 410385 246758
rect 410511 246757 410577 246760
rect 410799 246757 410865 246760
rect 410938 246758 410944 246822
rect 411008 246820 411014 246822
rect 411183 246820 411249 246823
rect 411375 246822 411441 246823
rect 411008 246818 411249 246820
rect 411008 246762 411188 246818
rect 411244 246762 411249 246818
rect 411008 246760 411249 246762
rect 411008 246758 411014 246760
rect 411183 246757 411249 246760
rect 411322 246758 411328 246822
rect 411392 246820 411441 246822
rect 411392 246818 411484 246820
rect 411436 246762 411484 246818
rect 411392 246760 411484 246762
rect 411714 246818 411825 246823
rect 411714 246762 411764 246818
rect 411820 246762 411825 246818
rect 411714 246760 411825 246762
rect 411392 246758 411441 246760
rect 411375 246757 411441 246758
rect 411759 246757 411825 246760
rect 412335 246820 412401 246823
rect 673978 246820 673984 246822
rect 412335 246818 673984 246820
rect 412335 246762 412340 246818
rect 412396 246762 673984 246818
rect 412335 246760 673984 246762
rect 412335 246757 412401 246760
rect 673978 246758 673984 246760
rect 674048 246758 674054 246822
rect 406575 246720 406641 246725
rect 155343 245486 210558 245488
rect 155343 245430 155348 245486
rect 155404 245430 210558 245486
rect 155343 245428 210558 245430
rect 155343 245425 155409 245428
rect 197295 245340 197361 245343
rect 210255 245340 210321 245343
rect 197295 245338 210321 245340
rect 197295 245282 197300 245338
rect 197356 245282 210260 245338
rect 210316 245282 210321 245338
rect 197295 245280 210321 245282
rect 197295 245277 197361 245280
rect 210255 245277 210321 245280
rect 673978 245278 673984 245342
rect 674048 245340 674054 245342
rect 675183 245340 675249 245343
rect 674048 245338 675249 245340
rect 674048 245282 675188 245338
rect 675244 245282 675249 245338
rect 674048 245280 675249 245282
rect 674048 245278 674054 245280
rect 675183 245277 675249 245280
rect 158319 245192 158385 245195
rect 210159 245192 210225 245195
rect 158319 245190 210225 245192
rect 158319 245134 158324 245190
rect 158380 245134 210164 245190
rect 210220 245134 210225 245190
rect 158319 245132 210225 245134
rect 158319 245129 158385 245132
rect 210159 245129 210225 245132
rect 161103 245044 161169 245047
rect 210063 245044 210129 245047
rect 161103 245042 210129 245044
rect 161103 244986 161108 245042
rect 161164 244986 210068 245042
rect 210124 244986 210129 245042
rect 161103 244984 210129 244986
rect 161103 244981 161169 244984
rect 210063 244981 210129 244984
rect 196719 244896 196785 244899
rect 209967 244896 210033 244899
rect 196719 244894 210033 244896
rect 196719 244838 196724 244894
rect 196780 244838 209972 244894
rect 210028 244838 210033 244894
rect 196719 244836 210033 244838
rect 196719 244833 196785 244836
rect 209967 244833 210033 244836
rect 675375 244750 675441 244751
rect 674362 244686 674368 244750
rect 674432 244748 674438 244750
rect 675322 244748 675328 244750
rect 674432 244688 675328 244748
rect 675392 244746 675441 244750
rect 675436 244690 675441 244746
rect 674432 244686 674438 244688
rect 675322 244686 675328 244688
rect 675392 244686 675441 244690
rect 675375 244685 675441 244686
rect 206607 244600 206673 244603
rect 206895 244600 206961 244603
rect 206607 244598 206961 244600
rect 206607 244542 206612 244598
rect 206668 244542 206900 244598
rect 206956 244542 206961 244598
rect 206607 244540 206961 244542
rect 206607 244537 206673 244540
rect 206895 244537 206961 244540
rect 41722 243798 41728 243862
rect 41792 243860 41798 243862
rect 42255 243860 42321 243863
rect 674362 243860 674368 243862
rect 41792 243858 674368 243860
rect 41792 243802 42260 243858
rect 42316 243802 674368 243858
rect 41792 243800 674368 243802
rect 41792 243798 41798 243800
rect 42255 243797 42321 243800
rect 674362 243798 674368 243800
rect 674432 243798 674438 243862
rect 209967 243712 210033 243715
rect 210447 243714 210513 243715
rect 210298 243712 210304 243714
rect 209967 243710 210304 243712
rect 209967 243654 209972 243710
rect 210028 243654 210304 243710
rect 209967 243652 210304 243654
rect 209967 243649 210033 243652
rect 210298 243650 210304 243652
rect 210368 243650 210374 243714
rect 210447 243710 210496 243714
rect 210560 243712 210566 243714
rect 213231 243712 213297 243715
rect 227055 243712 227121 243715
rect 210447 243654 210452 243710
rect 210447 243650 210496 243654
rect 210560 243652 210604 243712
rect 213231 243710 227121 243712
rect 213231 243654 213236 243710
rect 213292 243654 227060 243710
rect 227116 243654 227121 243710
rect 213231 243652 227121 243654
rect 210560 243650 210566 243652
rect 210447 243649 210513 243650
rect 213231 243649 213297 243652
rect 227055 243649 227121 243652
rect 227343 243712 227409 243715
rect 267951 243712 268017 243715
rect 227343 243710 268017 243712
rect 227343 243654 227348 243710
rect 227404 243654 267956 243710
rect 268012 243654 268017 243710
rect 227343 243652 268017 243654
rect 227343 243649 227409 243652
rect 267951 243649 268017 243652
rect 268090 243650 268096 243714
rect 268160 243712 268166 243714
rect 288111 243712 288177 243715
rect 268160 243710 288177 243712
rect 268160 243654 288116 243710
rect 288172 243654 288177 243710
rect 268160 243652 288177 243654
rect 268160 243650 268166 243652
rect 288111 243649 288177 243652
rect 288303 243712 288369 243715
rect 443535 243712 443601 243715
rect 288303 243710 443601 243712
rect 288303 243654 288308 243710
rect 288364 243654 443540 243710
rect 443596 243654 443601 243710
rect 288303 243652 443601 243654
rect 288303 243649 288369 243652
rect 443535 243649 443601 243652
rect 463599 243712 463665 243715
rect 483855 243712 483921 243715
rect 463599 243710 483921 243712
rect 463599 243654 463604 243710
rect 463660 243654 483860 243710
rect 483916 243654 483921 243710
rect 463599 243652 483921 243654
rect 463599 243649 463665 243652
rect 483855 243649 483921 243652
rect 503919 243712 503985 243715
rect 524175 243712 524241 243715
rect 503919 243710 524241 243712
rect 503919 243654 503924 243710
rect 503980 243654 524180 243710
rect 524236 243654 524241 243710
rect 503919 243652 524241 243654
rect 503919 243649 503985 243652
rect 524175 243649 524241 243652
rect 544239 243712 544305 243715
rect 564495 243712 564561 243715
rect 544239 243710 564561 243712
rect 544239 243654 544244 243710
rect 544300 243654 564500 243710
rect 564556 243654 564561 243710
rect 544239 243652 564561 243654
rect 544239 243649 544305 243652
rect 564495 243649 564561 243652
rect 584559 243712 584625 243715
rect 604815 243712 604881 243715
rect 584559 243710 604881 243712
rect 584559 243654 584564 243710
rect 584620 243654 604820 243710
rect 604876 243654 604881 243710
rect 584559 243652 604881 243654
rect 584559 243649 584625 243652
rect 604815 243649 604881 243652
rect 624879 243712 624945 243715
rect 645135 243712 645201 243715
rect 624879 243710 645201 243712
rect 624879 243654 624884 243710
rect 624940 243654 645140 243710
rect 645196 243654 645201 243710
rect 624879 243652 645201 243654
rect 624879 243649 624945 243652
rect 645135 243649 645201 243652
rect 178383 243564 178449 243567
rect 398703 243564 398769 243567
rect 405999 243566 406065 243567
rect 405754 243564 405760 243566
rect 178383 243562 398526 243564
rect 178383 243506 178388 243562
rect 178444 243506 398526 243562
rect 178383 243504 398526 243506
rect 178383 243501 178449 243504
rect 206895 243416 206961 243419
rect 388911 243416 388977 243419
rect 206895 243414 388977 243416
rect 206895 243358 206900 243414
rect 206956 243358 388916 243414
rect 388972 243358 388977 243414
rect 206895 243356 388977 243358
rect 398466 243416 398526 243504
rect 398703 243562 405760 243564
rect 398703 243506 398708 243562
rect 398764 243506 405760 243562
rect 398703 243504 405760 243506
rect 398703 243501 398769 243504
rect 405754 243502 405760 243504
rect 405824 243502 405830 243566
rect 405946 243502 405952 243566
rect 406016 243564 406065 243566
rect 406016 243562 406108 243564
rect 406060 243506 406108 243562
rect 406016 243504 406108 243506
rect 406016 243502 406065 243504
rect 674170 243502 674176 243566
rect 674240 243564 674246 243566
rect 675471 243564 675537 243567
rect 674240 243562 675537 243564
rect 674240 243506 675476 243562
rect 675532 243506 675537 243562
rect 674240 243504 675537 243506
rect 674240 243502 674246 243504
rect 405999 243501 406065 243502
rect 675471 243501 675537 243504
rect 408250 243416 408256 243418
rect 398466 243356 408256 243416
rect 206895 243353 206961 243356
rect 388911 243353 388977 243356
rect 408250 243354 408256 243356
rect 408320 243354 408326 243418
rect 210351 243268 210417 243271
rect 210682 243268 210688 243270
rect 210351 243266 210688 243268
rect 210351 243210 210356 243266
rect 210412 243210 210688 243266
rect 210351 243208 210688 243210
rect 210351 243205 210417 243208
rect 210682 243206 210688 243208
rect 210752 243206 210758 243270
rect 214959 243268 215025 243271
rect 227343 243268 227409 243271
rect 267898 243268 267904 243270
rect 214959 243266 227262 243268
rect 214959 243210 214964 243266
rect 215020 243210 227262 243266
rect 214959 243208 227262 243210
rect 214959 243205 215025 243208
rect 210255 243120 210321 243123
rect 210874 243120 210880 243122
rect 210255 243118 210880 243120
rect 210255 243062 210260 243118
rect 210316 243062 210880 243118
rect 210255 243060 210880 243062
rect 210255 243057 210321 243060
rect 210874 243058 210880 243060
rect 210944 243058 210950 243122
rect 217167 243120 217233 243123
rect 227055 243120 227121 243123
rect 217167 243118 227121 243120
rect 217167 243062 217172 243118
rect 217228 243062 227060 243118
rect 227116 243062 227121 243118
rect 217167 243060 227121 243062
rect 227202 243120 227262 243208
rect 227343 243266 267904 243268
rect 227343 243210 227348 243266
rect 227404 243210 267904 243266
rect 227343 243208 267904 243210
rect 227343 243205 227409 243208
rect 267898 243206 267904 243208
rect 267968 243206 267974 243270
rect 298191 243268 298257 243271
rect 307887 243268 307953 243271
rect 268098 243208 298110 243268
rect 268098 243120 268158 243208
rect 227202 243060 268158 243120
rect 217167 243057 217233 243060
rect 227055 243057 227121 243060
rect 268282 243058 268288 243122
rect 268352 243120 268358 243122
rect 268352 243060 287934 243120
rect 268352 243058 268358 243060
rect 41914 242910 41920 242974
rect 41984 242972 41990 242974
rect 42874 242972 42880 242974
rect 41984 242912 42880 242972
rect 41984 242910 41990 242912
rect 42874 242910 42880 242912
rect 42944 242910 42950 242974
rect 218895 242972 218961 242975
rect 227343 242972 227409 242975
rect 218895 242970 227409 242972
rect 218895 242914 218900 242970
rect 218956 242914 227348 242970
rect 227404 242914 227409 242970
rect 218895 242912 227409 242914
rect 218895 242909 218961 242912
rect 227343 242909 227409 242912
rect 231663 242972 231729 242975
rect 268090 242972 268096 242974
rect 231663 242970 268096 242972
rect 231663 242914 231668 242970
rect 231724 242914 268096 242970
rect 231663 242912 268096 242914
rect 231663 242909 231729 242912
rect 268090 242910 268096 242912
rect 268160 242910 268166 242974
rect 268239 242972 268305 242975
rect 287631 242972 287697 242975
rect 268239 242970 287697 242972
rect 268239 242914 268244 242970
rect 268300 242914 287636 242970
rect 287692 242914 287697 242970
rect 268239 242912 287697 242914
rect 287874 242972 287934 243060
rect 288058 243058 288064 243122
rect 288128 243120 288134 243122
rect 297903 243120 297969 243123
rect 288128 243118 297969 243120
rect 288128 243062 297908 243118
rect 297964 243062 297969 243118
rect 288128 243060 297969 243062
rect 298050 243120 298110 243208
rect 298191 243266 307953 243268
rect 298191 243210 298196 243266
rect 298252 243210 307892 243266
rect 307948 243210 307953 243266
rect 298191 243208 307953 243210
rect 298191 243205 298257 243208
rect 307887 243205 307953 243208
rect 308079 243268 308145 243271
rect 409018 243268 409024 243270
rect 308079 243266 409024 243268
rect 308079 243210 308084 243266
rect 308140 243210 409024 243266
rect 308079 243208 409024 243210
rect 308079 243205 308145 243208
rect 409018 243206 409024 243208
rect 409088 243206 409094 243270
rect 338511 243120 338577 243123
rect 354639 243120 354705 243123
rect 298050 243060 338430 243120
rect 288128 243058 288134 243060
rect 297903 243057 297969 243060
rect 328335 242972 328401 242975
rect 287874 242970 328401 242972
rect 287874 242914 328340 242970
rect 328396 242914 328401 242970
rect 287874 242912 328401 242914
rect 268239 242909 268305 242912
rect 287631 242909 287697 242912
rect 328335 242909 328401 242912
rect 328527 242972 328593 242975
rect 338127 242972 338193 242975
rect 328527 242970 338193 242972
rect 328527 242914 328532 242970
rect 328588 242914 338132 242970
rect 338188 242914 338193 242970
rect 328527 242912 338193 242914
rect 338370 242972 338430 243060
rect 338511 243118 354705 243120
rect 338511 243062 338516 243118
rect 338572 243062 354644 243118
rect 354700 243062 354705 243118
rect 338511 243060 354705 243062
rect 338511 243057 338577 243060
rect 354639 243057 354705 243060
rect 388911 243120 388977 243123
rect 408058 243120 408064 243122
rect 388911 243118 408064 243120
rect 388911 243062 388916 243118
rect 388972 243062 408064 243118
rect 388911 243060 408064 243062
rect 388911 243057 388977 243060
rect 408058 243058 408064 243060
rect 408128 243058 408134 243122
rect 338370 242912 346110 242972
rect 328527 242909 328593 242912
rect 338127 242909 338193 242912
rect 43311 242824 43377 242827
rect 54735 242824 54801 242827
rect 43311 242822 54801 242824
rect 43311 242766 43316 242822
rect 43372 242766 54740 242822
rect 54796 242766 54801 242822
rect 43311 242764 54801 242766
rect 43311 242761 43377 242764
rect 54735 242761 54801 242764
rect 220815 242824 220881 242827
rect 227386 242824 227392 242826
rect 220815 242822 227392 242824
rect 220815 242766 220820 242822
rect 220876 242766 227392 242822
rect 220815 242764 227392 242766
rect 220815 242761 220881 242764
rect 227386 242762 227392 242764
rect 227456 242762 227462 242826
rect 227631 242824 227697 242827
rect 308079 242824 308145 242827
rect 227631 242822 308145 242824
rect 227631 242766 227636 242822
rect 227692 242766 308084 242822
rect 308140 242766 308145 242822
rect 227631 242764 308145 242766
rect 227631 242761 227697 242764
rect 308079 242761 308145 242764
rect 308271 242824 308337 242827
rect 328431 242824 328497 242827
rect 341199 242824 341265 242827
rect 308271 242822 328497 242824
rect 308271 242766 308276 242822
rect 308332 242766 328436 242822
rect 328492 242766 328497 242822
rect 308271 242764 328497 242766
rect 308271 242761 308337 242764
rect 328431 242761 328497 242764
rect 328578 242822 341265 242824
rect 328578 242766 341204 242822
rect 341260 242766 341265 242822
rect 328578 242764 341265 242766
rect 346050 242824 346110 242912
rect 352239 242824 352305 242827
rect 346050 242822 352305 242824
rect 346050 242766 352244 242822
rect 352300 242766 352305 242822
rect 346050 242764 352305 242766
rect 106575 242676 106641 242679
rect 106575 242674 115134 242676
rect 106575 242618 106580 242674
rect 106636 242618 115134 242674
rect 106575 242616 115134 242618
rect 106575 242613 106641 242616
rect 54831 242528 54897 242531
rect 95055 242528 95121 242531
rect 54831 242526 95121 242528
rect 54831 242470 54836 242526
rect 54892 242470 95060 242526
rect 95116 242470 95121 242526
rect 54831 242468 95121 242470
rect 115074 242528 115134 242616
rect 115258 242614 115264 242678
rect 115328 242676 115334 242678
rect 126639 242676 126705 242679
rect 115328 242674 126705 242676
rect 115328 242618 126644 242674
rect 126700 242618 126705 242674
rect 115328 242616 126705 242618
rect 115328 242614 115334 242616
rect 126639 242613 126705 242616
rect 126831 242676 126897 242679
rect 138255 242676 138321 242679
rect 126831 242674 138321 242676
rect 126831 242618 126836 242674
rect 126892 242618 138260 242674
rect 138316 242618 138321 242674
rect 126831 242616 138321 242618
rect 126831 242613 126897 242616
rect 138255 242613 138321 242616
rect 171375 242676 171441 242679
rect 175546 242676 175552 242678
rect 171375 242674 175552 242676
rect 171375 242618 171380 242674
rect 171436 242618 175552 242674
rect 171375 242616 175552 242618
rect 171375 242613 171441 242616
rect 175546 242614 175552 242616
rect 175616 242614 175622 242678
rect 221967 242676 222033 242679
rect 227535 242676 227601 242679
rect 221967 242674 227601 242676
rect 221967 242618 221972 242674
rect 222028 242618 227540 242674
rect 227596 242618 227601 242674
rect 221967 242616 227601 242618
rect 221967 242613 222033 242616
rect 227535 242613 227601 242616
rect 227727 242676 227793 242679
rect 328578 242676 328638 242764
rect 341199 242761 341265 242764
rect 352239 242761 352305 242764
rect 227727 242674 328638 242676
rect 227727 242618 227732 242674
rect 227788 242618 328638 242674
rect 227727 242616 328638 242618
rect 328719 242676 328785 242679
rect 338991 242676 339057 242679
rect 328719 242674 339057 242676
rect 328719 242618 328724 242674
rect 328780 242618 338996 242674
rect 339052 242618 339057 242674
rect 328719 242616 339057 242618
rect 227727 242613 227793 242616
rect 328719 242613 328785 242616
rect 338991 242613 339057 242616
rect 339183 242676 339249 242679
rect 343407 242676 343473 242679
rect 339183 242674 343473 242676
rect 339183 242618 339188 242674
rect 339244 242618 343412 242674
rect 343468 242618 343473 242674
rect 339183 242616 343473 242618
rect 339183 242613 339249 242616
rect 343407 242613 343473 242616
rect 115258 242528 115264 242530
rect 115074 242468 115264 242528
rect 54831 242465 54897 242468
rect 95055 242465 95121 242468
rect 115258 242466 115264 242468
rect 115328 242466 115334 242530
rect 195759 242528 195825 242531
rect 223983 242528 224049 242531
rect 247311 242530 247377 242531
rect 247311 242528 247360 242530
rect 195759 242526 224049 242528
rect 195759 242470 195764 242526
rect 195820 242470 223988 242526
rect 224044 242470 224049 242526
rect 195759 242468 224049 242470
rect 247268 242526 247360 242528
rect 247268 242470 247316 242526
rect 247268 242468 247360 242470
rect 195759 242465 195825 242468
rect 223983 242465 224049 242468
rect 247311 242466 247360 242468
rect 247424 242466 247430 242530
rect 247791 242528 247857 242531
rect 267759 242528 267825 242531
rect 247791 242526 267825 242528
rect 247791 242470 247796 242526
rect 247852 242470 267764 242526
rect 267820 242470 267825 242526
rect 247791 242468 267825 242470
rect 247311 242465 247377 242466
rect 247791 242465 247857 242468
rect 267759 242465 267825 242468
rect 267951 242528 268017 242531
rect 287823 242528 287889 242531
rect 267951 242526 287889 242528
rect 267951 242470 267956 242526
rect 268012 242470 287828 242526
rect 287884 242470 287889 242526
rect 267951 242468 287889 242470
rect 267951 242465 268017 242468
rect 287823 242465 287889 242468
rect 288015 242528 288081 242531
rect 307695 242528 307761 242531
rect 288015 242526 307761 242528
rect 288015 242470 288020 242526
rect 288076 242470 307700 242526
rect 307756 242470 307761 242526
rect 288015 242468 307761 242470
rect 288015 242465 288081 242468
rect 307695 242465 307761 242468
rect 307887 242528 307953 242531
rect 443535 242528 443601 242531
rect 307887 242526 443601 242528
rect 307887 242470 307892 242526
rect 307948 242470 443540 242526
rect 443596 242470 443601 242526
rect 307887 242468 443601 242470
rect 307887 242465 307953 242468
rect 443535 242465 443601 242468
rect 463599 242528 463665 242531
rect 483855 242528 483921 242531
rect 463599 242526 483921 242528
rect 463599 242470 463604 242526
rect 463660 242470 483860 242526
rect 483916 242470 483921 242526
rect 463599 242468 483921 242470
rect 463599 242465 463665 242468
rect 483855 242465 483921 242468
rect 503919 242528 503985 242531
rect 511119 242528 511185 242531
rect 503919 242526 511185 242528
rect 503919 242470 503924 242526
rect 503980 242470 511124 242526
rect 511180 242470 511185 242526
rect 503919 242468 511185 242470
rect 503919 242465 503985 242468
rect 511119 242465 511185 242468
rect 144015 242380 144081 242383
rect 140832 242378 144081 242380
rect 140832 242322 144020 242378
rect 144076 242322 144081 242378
rect 140832 242320 144081 242322
rect 144015 242317 144081 242320
rect 175546 242318 175552 242382
rect 175616 242380 175622 242382
rect 175695 242380 175761 242383
rect 175616 242378 175761 242380
rect 175616 242322 175700 242378
rect 175756 242322 175761 242378
rect 175616 242320 175761 242322
rect 175616 242318 175622 242320
rect 175695 242317 175761 242320
rect 210639 242380 210705 242383
rect 227247 242380 227313 242383
rect 210639 242378 227313 242380
rect 210639 242322 210644 242378
rect 210700 242322 227252 242378
rect 227308 242322 227313 242378
rect 210639 242320 227313 242322
rect 210639 242317 210705 242320
rect 227247 242317 227313 242320
rect 227535 242380 227601 242383
rect 227535 242378 227838 242380
rect 227535 242322 227540 242378
rect 227596 242322 227838 242378
rect 227535 242320 227838 242322
rect 227535 242317 227601 242320
rect 211503 242232 211569 242235
rect 223503 242232 223569 242235
rect 211503 242230 223569 242232
rect 211503 242174 211508 242230
rect 211564 242174 223508 242230
rect 223564 242174 223569 242230
rect 211503 242172 223569 242174
rect 211503 242169 211569 242172
rect 223503 242169 223569 242172
rect 223695 242232 223761 242235
rect 227631 242232 227697 242235
rect 223695 242230 227697 242232
rect 223695 242174 223700 242230
rect 223756 242174 227636 242230
rect 227692 242174 227697 242230
rect 223695 242172 227697 242174
rect 227778 242232 227838 242320
rect 227962 242318 227968 242382
rect 228032 242380 228038 242382
rect 241935 242380 242001 242383
rect 228032 242378 242001 242380
rect 228032 242322 241940 242378
rect 241996 242322 242001 242378
rect 228032 242320 242001 242322
rect 228032 242318 228038 242320
rect 241935 242317 242001 242320
rect 242319 242380 242385 242383
rect 342063 242380 342129 242383
rect 242319 242378 342129 242380
rect 242319 242322 242324 242378
rect 242380 242322 342068 242378
rect 342124 242322 342129 242378
rect 242319 242320 342129 242322
rect 242319 242317 242385 242320
rect 342063 242317 342129 242320
rect 342927 242232 342993 242235
rect 227778 242230 342993 242232
rect 227778 242174 342932 242230
rect 342988 242174 342993 242230
rect 227778 242172 342993 242174
rect 223695 242169 223761 242172
rect 227631 242169 227697 242172
rect 342927 242169 342993 242172
rect 221391 242084 221457 242087
rect 338511 242084 338577 242087
rect 221391 242082 338577 242084
rect 221391 242026 221396 242082
rect 221452 242026 338516 242082
rect 338572 242026 338577 242082
rect 221391 242024 338577 242026
rect 221391 242021 221457 242024
rect 338511 242021 338577 242024
rect 338799 242084 338865 242087
rect 344271 242084 344337 242087
rect 338799 242082 344337 242084
rect 338799 242026 338804 242082
rect 338860 242026 344276 242082
rect 344332 242026 344337 242082
rect 338799 242024 344337 242026
rect 338799 242021 338865 242024
rect 344271 242021 344337 242024
rect 211407 241936 211473 241939
rect 521583 241936 521649 241939
rect 211407 241934 521649 241936
rect 211407 241878 211412 241934
rect 211468 241878 521588 241934
rect 521644 241878 521649 241934
rect 211407 241876 521649 241878
rect 211407 241873 211473 241876
rect 521583 241873 521649 241876
rect 245391 241788 245457 241791
rect 267951 241788 268017 241791
rect 245391 241786 268017 241788
rect 245391 241730 245396 241786
rect 245452 241730 267956 241786
rect 268012 241730 268017 241786
rect 245391 241728 268017 241730
rect 245391 241725 245457 241728
rect 267951 241725 268017 241728
rect 268090 241726 268096 241790
rect 268160 241788 268166 241790
rect 287866 241788 287872 241790
rect 268160 241728 287872 241788
rect 268160 241726 268166 241728
rect 287866 241726 287872 241728
rect 287936 241726 287942 241790
rect 289647 241788 289713 241791
rect 356751 241788 356817 241791
rect 289647 241786 356817 241788
rect 289647 241730 289652 241786
rect 289708 241730 356756 241786
rect 356812 241730 356817 241786
rect 289647 241728 356817 241730
rect 289647 241725 289713 241728
rect 356751 241725 356817 241728
rect 246735 241640 246801 241643
rect 354447 241640 354513 241643
rect 246735 241638 354513 241640
rect 246735 241582 246740 241638
rect 246796 241582 354452 241638
rect 354508 241582 354513 241638
rect 246735 241580 354513 241582
rect 246735 241577 246801 241580
rect 354447 241577 354513 241580
rect 247738 241430 247744 241494
rect 247808 241492 247814 241494
rect 267514 241492 267520 241494
rect 247808 241432 267520 241492
rect 247808 241430 247814 241432
rect 267514 241430 267520 241432
rect 267584 241430 267590 241494
rect 267663 241492 267729 241495
rect 372879 241492 372945 241495
rect 267663 241490 372945 241492
rect 267663 241434 267668 241490
rect 267724 241434 372884 241490
rect 372940 241434 372945 241490
rect 267663 241432 372945 241434
rect 267663 241429 267729 241432
rect 372879 241429 372945 241432
rect 261231 241344 261297 241347
rect 267567 241344 267633 241347
rect 261231 241342 267633 241344
rect 261231 241286 261236 241342
rect 261292 241286 267572 241342
rect 267628 241286 267633 241342
rect 261231 241284 267633 241286
rect 261231 241281 261297 241284
rect 267567 241281 267633 241284
rect 267759 241344 267825 241347
rect 376815 241344 376881 241347
rect 267759 241342 376881 241344
rect 267759 241286 267764 241342
rect 267820 241286 376820 241342
rect 376876 241286 376881 241342
rect 267759 241284 376881 241286
rect 267759 241281 267825 241284
rect 376815 241281 376881 241284
rect 244527 241196 244593 241199
rect 278127 241196 278193 241199
rect 289647 241196 289713 241199
rect 244527 241194 277950 241196
rect 244527 241138 244532 241194
rect 244588 241138 277950 241194
rect 244527 241136 277950 241138
rect 244527 241133 244593 241136
rect 42255 240754 42321 240755
rect 42255 240752 42304 240754
rect 42212 240750 42304 240752
rect 42212 240694 42260 240750
rect 42212 240692 42304 240694
rect 42255 240690 42304 240692
rect 42368 240690 42374 240754
rect 42255 240689 42321 240690
rect 140802 240604 140862 241092
rect 243183 241048 243249 241051
rect 277743 241048 277809 241051
rect 243183 241046 277809 241048
rect 243183 240990 243188 241046
rect 243244 240990 277748 241046
rect 277804 240990 277809 241046
rect 243183 240988 277809 240990
rect 277890 241048 277950 241136
rect 278127 241194 289713 241196
rect 278127 241138 278132 241194
rect 278188 241138 289652 241194
rect 289708 241138 289713 241194
rect 278127 241136 289713 241138
rect 278127 241133 278193 241136
rect 289647 241133 289713 241136
rect 289839 241196 289905 241199
rect 295599 241196 295665 241199
rect 358959 241196 359025 241199
rect 289839 241194 295665 241196
rect 289839 241138 289844 241194
rect 289900 241138 295604 241194
rect 295660 241138 295665 241194
rect 289839 241136 295665 241138
rect 289839 241133 289905 241136
rect 295599 241133 295665 241136
rect 295746 241194 359025 241196
rect 295746 241138 358964 241194
rect 359020 241138 359025 241194
rect 295746 241136 359025 241138
rect 295746 241048 295806 241136
rect 358959 241133 359025 241136
rect 277890 240988 295806 241048
rect 295887 241048 295953 241051
rect 361647 241048 361713 241051
rect 295887 241046 361713 241048
rect 295887 240990 295892 241046
rect 295948 240990 361652 241046
rect 361708 240990 361713 241046
rect 295887 240988 361713 240990
rect 243183 240985 243249 240988
rect 277743 240985 277809 240988
rect 295887 240985 295953 240988
rect 361647 240985 361713 240988
rect 259023 240900 259089 240903
rect 377871 240900 377937 240903
rect 259023 240898 377937 240900
rect 259023 240842 259028 240898
rect 259084 240842 377876 240898
rect 377932 240842 377937 240898
rect 259023 240840 377937 240842
rect 259023 240837 259089 240840
rect 377871 240837 377937 240840
rect 242703 240752 242769 240755
rect 278031 240752 278097 240755
rect 289839 240752 289905 240755
rect 363087 240752 363153 240755
rect 242703 240750 277950 240752
rect 242703 240694 242708 240750
rect 242764 240694 277950 240750
rect 242703 240692 277950 240694
rect 242703 240689 242769 240692
rect 146031 240604 146097 240607
rect 140802 240602 146097 240604
rect 140802 240546 146036 240602
rect 146092 240546 146097 240602
rect 140802 240544 146097 240546
rect 146031 240541 146097 240544
rect 241743 240604 241809 240607
rect 277890 240604 277950 240692
rect 278031 240750 289905 240752
rect 278031 240694 278036 240750
rect 278092 240694 289844 240750
rect 289900 240694 289905 240750
rect 278031 240692 289905 240694
rect 278031 240689 278097 240692
rect 289839 240689 289905 240692
rect 289986 240750 363153 240752
rect 289986 240694 363092 240750
rect 363148 240694 363153 240750
rect 289986 240692 363153 240694
rect 289986 240604 290046 240692
rect 363087 240689 363153 240692
rect 383535 240752 383601 240755
rect 398607 240752 398673 240755
rect 383535 240750 398673 240752
rect 383535 240694 383540 240750
rect 383596 240694 398612 240750
rect 398668 240694 398673 240750
rect 383535 240692 398673 240694
rect 383535 240689 383601 240692
rect 398607 240689 398673 240692
rect 364815 240604 364881 240607
rect 241743 240602 277758 240604
rect 241743 240546 241748 240602
rect 241804 240546 277758 240602
rect 241743 240544 277758 240546
rect 277890 240544 290046 240604
rect 293442 240602 364881 240604
rect 293442 240546 364820 240602
rect 364876 240546 364881 240602
rect 293442 240544 364881 240546
rect 241743 240541 241809 240544
rect 240975 240456 241041 240459
rect 277551 240456 277617 240459
rect 240975 240454 277617 240456
rect 240975 240398 240980 240454
rect 241036 240398 277556 240454
rect 277612 240398 277617 240454
rect 240975 240396 277617 240398
rect 277698 240456 277758 240544
rect 293442 240456 293502 240544
rect 364815 240541 364881 240544
rect 277698 240396 293502 240456
rect 297999 240456 298065 240459
rect 366543 240456 366609 240459
rect 297999 240454 366609 240456
rect 297999 240398 298004 240454
rect 298060 240398 366548 240454
rect 366604 240398 366609 240454
rect 297999 240396 366609 240398
rect 240975 240393 241041 240396
rect 277551 240393 277617 240396
rect 297999 240393 298065 240396
rect 366543 240393 366609 240396
rect 367599 240456 367665 240459
rect 409743 240456 409809 240459
rect 367599 240454 409809 240456
rect 367599 240398 367604 240454
rect 367660 240398 409748 240454
rect 409804 240398 409809 240454
rect 367599 240396 409809 240398
rect 367599 240393 367665 240396
rect 409743 240393 409809 240396
rect 262959 240308 263025 240311
rect 369807 240308 369873 240311
rect 262959 240306 369873 240308
rect 262959 240250 262964 240306
rect 263020 240250 369812 240306
rect 369868 240250 369873 240306
rect 262959 240248 369873 240250
rect 262959 240245 263025 240248
rect 369807 240245 369873 240248
rect 247695 240160 247761 240163
rect 352815 240160 352881 240163
rect 247695 240158 352881 240160
rect 247695 240102 247700 240158
rect 247756 240102 352820 240158
rect 352876 240102 352881 240158
rect 247695 240100 352881 240102
rect 247695 240097 247761 240100
rect 352815 240097 352881 240100
rect 247983 240012 248049 240015
rect 351279 240012 351345 240015
rect 247983 240010 351345 240012
rect 247983 239954 247988 240010
rect 248044 239954 351284 240010
rect 351340 239954 351345 240010
rect 247983 239952 351345 239954
rect 247983 239949 248049 239952
rect 351279 239949 351345 239952
rect 145402 239864 145408 239866
rect 140832 239804 145408 239864
rect 145402 239802 145408 239804
rect 145472 239802 145478 239866
rect 259599 239864 259665 239867
rect 267759 239864 267825 239867
rect 259599 239862 267825 239864
rect 259599 239806 259604 239862
rect 259660 239806 267764 239862
rect 267820 239806 267825 239862
rect 259599 239804 267825 239806
rect 259599 239801 259665 239804
rect 267759 239801 267825 239804
rect 277551 239864 277617 239867
rect 297999 239864 298065 239867
rect 277551 239862 298065 239864
rect 277551 239806 277556 239862
rect 277612 239806 298004 239862
rect 298060 239806 298065 239862
rect 277551 239804 298065 239806
rect 277551 239801 277617 239804
rect 297999 239801 298065 239804
rect 267951 239716 268017 239719
rect 278127 239716 278193 239719
rect 267951 239714 278193 239716
rect 267951 239658 267956 239714
rect 268012 239658 278132 239714
rect 278188 239658 278193 239714
rect 267951 239656 278193 239658
rect 267951 239653 268017 239656
rect 278127 239653 278193 239656
rect 285039 239716 285105 239719
rect 288111 239716 288177 239719
rect 285039 239714 288177 239716
rect 285039 239658 285044 239714
rect 285100 239658 288116 239714
rect 288172 239658 288177 239714
rect 285039 239656 288177 239658
rect 285039 239653 285105 239656
rect 288111 239653 288177 239656
rect 293775 239716 293841 239719
rect 301071 239716 301137 239719
rect 293775 239714 301137 239716
rect 293775 239658 293780 239714
rect 293836 239658 301076 239714
rect 301132 239658 301137 239714
rect 293775 239656 301137 239658
rect 293775 239653 293841 239656
rect 301071 239653 301137 239656
rect 383055 239716 383121 239719
rect 383055 239714 383166 239716
rect 383055 239658 383060 239714
rect 383116 239658 383166 239714
rect 383055 239653 383166 239658
rect 278799 239568 278865 239571
rect 280239 239568 280305 239571
rect 278799 239566 280305 239568
rect 278799 239510 278804 239566
rect 278860 239510 280244 239566
rect 280300 239510 280305 239566
rect 278799 239508 280305 239510
rect 278799 239505 278865 239508
rect 280239 239505 280305 239508
rect 287247 239568 287313 239571
rect 293775 239568 293841 239571
rect 287247 239566 293841 239568
rect 287247 239510 287252 239566
rect 287308 239510 293780 239566
rect 293836 239510 293841 239566
rect 287247 239508 293841 239510
rect 287247 239505 287313 239508
rect 293775 239505 293841 239508
rect 293103 239420 293169 239423
rect 305295 239420 305361 239423
rect 293103 239418 305361 239420
rect 293103 239362 293108 239418
rect 293164 239362 305300 239418
rect 305356 239362 305361 239418
rect 293103 239360 305361 239362
rect 293103 239357 293169 239360
rect 305295 239357 305361 239360
rect 292239 239272 292305 239275
rect 295695 239272 295761 239275
rect 292239 239270 295761 239272
rect 292239 239214 292244 239270
rect 292300 239214 295700 239270
rect 295756 239214 295761 239270
rect 292239 239212 295761 239214
rect 292239 239209 292305 239212
rect 295695 239209 295761 239212
rect 383106 239127 383166 239653
rect 208527 239124 208593 239127
rect 209871 239124 209937 239127
rect 351375 239124 351441 239127
rect 208527 239122 351441 239124
rect 208527 239066 208532 239122
rect 208588 239066 209876 239122
rect 209932 239066 351380 239122
rect 351436 239066 351441 239122
rect 208527 239064 351441 239066
rect 208527 239061 208593 239064
rect 209871 239061 209937 239064
rect 351375 239061 351441 239064
rect 383055 239122 383166 239127
rect 383055 239066 383060 239122
rect 383116 239066 383166 239122
rect 383055 239064 383166 239066
rect 383055 239061 383121 239064
rect 212271 238976 212337 238979
rect 596175 238976 596241 238979
rect 212271 238974 596241 238976
rect 212271 238918 212276 238974
rect 212332 238918 596180 238974
rect 596236 238918 596241 238974
rect 212271 238916 596241 238918
rect 212271 238913 212337 238916
rect 596175 238913 596241 238916
rect 675183 238976 675249 238979
rect 675514 238976 675520 238978
rect 675183 238974 675520 238976
rect 675183 238918 675188 238974
rect 675244 238918 675520 238974
rect 675183 238916 675520 238918
rect 675183 238913 675249 238916
rect 675514 238914 675520 238916
rect 675584 238914 675590 238978
rect 191439 238828 191505 238831
rect 412047 238828 412113 238831
rect 191439 238826 412113 238828
rect 191439 238770 191444 238826
rect 191500 238770 412052 238826
rect 412108 238770 412113 238826
rect 191439 238768 412113 238770
rect 191439 238765 191505 238768
rect 412047 238765 412113 238768
rect 144111 238680 144177 238683
rect 140832 238678 144177 238680
rect 140832 238622 144116 238678
rect 144172 238622 144177 238678
rect 140832 238620 144177 238622
rect 144111 238617 144177 238620
rect 243567 238680 243633 238683
rect 360687 238680 360753 238683
rect 243567 238678 360753 238680
rect 243567 238622 243572 238678
rect 243628 238622 360692 238678
rect 360748 238622 360753 238678
rect 243567 238620 360753 238622
rect 243567 238617 243633 238620
rect 360687 238617 360753 238620
rect 675759 238680 675825 238683
rect 675898 238680 675904 238682
rect 675759 238678 675904 238680
rect 675759 238622 675764 238678
rect 675820 238622 675904 238678
rect 675759 238620 675904 238622
rect 675759 238617 675825 238620
rect 675898 238618 675904 238620
rect 675968 238618 675974 238682
rect 242319 238532 242385 238535
rect 363855 238532 363921 238535
rect 242319 238530 363921 238532
rect 242319 238474 242324 238530
rect 242380 238474 363860 238530
rect 363916 238474 363921 238530
rect 242319 238472 363921 238474
rect 242319 238469 242385 238472
rect 363855 238469 363921 238472
rect 258639 238384 258705 238387
rect 378831 238384 378897 238387
rect 258639 238382 378897 238384
rect 258639 238326 258644 238382
rect 258700 238326 378836 238382
rect 378892 238326 378897 238382
rect 258639 238324 378897 238326
rect 258639 238321 258705 238324
rect 378831 238321 378897 238324
rect 215823 238236 215889 238239
rect 227439 238236 227505 238239
rect 215823 238234 227505 238236
rect 215823 238178 215828 238234
rect 215884 238178 227444 238234
rect 227500 238178 227505 238234
rect 215823 238176 227505 238178
rect 215823 238173 215889 238176
rect 227439 238173 227505 238176
rect 241359 238236 241425 238239
rect 365775 238236 365841 238239
rect 241359 238234 365841 238236
rect 241359 238178 241364 238234
rect 241420 238178 365780 238234
rect 365836 238178 365841 238234
rect 241359 238176 365841 238178
rect 241359 238173 241425 238176
rect 365775 238173 365841 238176
rect 215247 238088 215313 238091
rect 227631 238088 227697 238091
rect 239055 238088 239121 238091
rect 215247 238086 217086 238088
rect 215247 238030 215252 238086
rect 215308 238030 217086 238086
rect 215247 238028 217086 238030
rect 215247 238025 215313 238028
rect 214863 237940 214929 237943
rect 217026 237940 217086 238028
rect 227631 238086 239121 238088
rect 227631 238030 227636 238086
rect 227692 238030 239060 238086
rect 239116 238030 239121 238086
rect 227631 238028 239121 238030
rect 227631 238025 227697 238028
rect 239055 238025 239121 238028
rect 259119 238088 259185 238091
rect 319695 238088 319761 238091
rect 259119 238086 319761 238088
rect 259119 238030 259124 238086
rect 259180 238030 319700 238086
rect 319756 238030 319761 238086
rect 259119 238028 319761 238030
rect 259119 238025 259185 238028
rect 319695 238025 319761 238028
rect 339759 238088 339825 238091
rect 342735 238088 342801 238091
rect 339759 238086 342801 238088
rect 339759 238030 339764 238086
rect 339820 238030 342740 238086
rect 342796 238030 342801 238086
rect 339759 238028 342801 238030
rect 339759 238025 339825 238028
rect 342735 238025 342801 238028
rect 369999 238088 370065 238091
rect 383055 238088 383121 238091
rect 369999 238086 383121 238088
rect 369999 238030 370004 238086
rect 370060 238030 383060 238086
rect 383116 238030 383121 238086
rect 369999 238028 383121 238030
rect 369999 238025 370065 238028
rect 383055 238025 383121 238028
rect 393135 237940 393201 237943
rect 214863 237938 216894 237940
rect 214863 237882 214868 237938
rect 214924 237882 216894 237938
rect 214863 237880 216894 237882
rect 217026 237938 393201 237940
rect 217026 237882 393140 237938
rect 393196 237882 393201 237938
rect 217026 237880 393201 237882
rect 214863 237877 214929 237880
rect 152463 237792 152529 237795
rect 211066 237792 211072 237794
rect 152463 237790 211072 237792
rect 152463 237734 152468 237790
rect 152524 237734 211072 237790
rect 152463 237732 211072 237734
rect 152463 237729 152529 237732
rect 211066 237730 211072 237732
rect 211136 237792 211142 237794
rect 216687 237792 216753 237795
rect 211136 237790 216753 237792
rect 211136 237734 216692 237790
rect 216748 237734 216753 237790
rect 211136 237732 216753 237734
rect 216834 237792 216894 237880
rect 393135 237877 393201 237880
rect 394671 237792 394737 237795
rect 216834 237790 394737 237792
rect 216834 237734 394676 237790
rect 394732 237734 394737 237790
rect 216834 237732 394737 237734
rect 211136 237730 211142 237732
rect 216687 237729 216753 237732
rect 394671 237729 394737 237732
rect 511119 237792 511185 237795
rect 677050 237792 677056 237794
rect 511119 237790 677056 237792
rect 511119 237734 511124 237790
rect 511180 237734 677056 237790
rect 511119 237732 677056 237734
rect 511119 237729 511185 237732
rect 677050 237730 677056 237732
rect 677120 237730 677126 237794
rect 142479 237644 142545 237647
rect 209583 237644 209649 237647
rect 214767 237644 214833 237647
rect 142479 237642 214833 237644
rect 142479 237586 142484 237642
rect 142540 237586 209588 237642
rect 209644 237586 214772 237642
rect 214828 237586 214833 237642
rect 142479 237584 214833 237586
rect 142479 237581 142545 237584
rect 209583 237581 209649 237584
rect 214767 237581 214833 237584
rect 216207 237644 216273 237647
rect 411951 237644 412017 237647
rect 216207 237642 412017 237644
rect 216207 237586 216212 237642
rect 216268 237586 411956 237642
rect 412012 237586 412017 237642
rect 216207 237584 412017 237586
rect 216207 237581 216273 237584
rect 411951 237581 412017 237584
rect 505839 237644 505905 237647
rect 676858 237644 676864 237646
rect 505839 237642 676864 237644
rect 505839 237586 505844 237642
rect 505900 237586 676864 237642
rect 505839 237584 676864 237586
rect 505839 237581 505905 237584
rect 676858 237582 676864 237584
rect 676928 237582 676934 237646
rect 243951 237496 244017 237499
rect 360015 237496 360081 237499
rect 243951 237494 360081 237496
rect 243951 237438 243956 237494
rect 244012 237438 360020 237494
rect 360076 237438 360081 237494
rect 243951 237436 360081 237438
rect 243951 237433 244017 237436
rect 360015 237433 360081 237436
rect 140802 236904 140862 237392
rect 243087 237348 243153 237351
rect 362703 237348 362769 237351
rect 243087 237346 362769 237348
rect 243087 237290 243092 237346
rect 243148 237290 362708 237346
rect 362764 237290 362769 237346
rect 243087 237288 362769 237290
rect 243087 237285 243153 237288
rect 362703 237285 362769 237288
rect 245295 237200 245361 237203
rect 357807 237200 357873 237203
rect 245295 237198 357873 237200
rect 245295 237142 245300 237198
rect 245356 237142 357812 237198
rect 357868 237142 357873 237198
rect 245295 237140 357873 237142
rect 245295 237137 245361 237140
rect 357807 237137 357873 237140
rect 209775 237052 209841 237055
rect 227439 237052 227505 237055
rect 209775 237050 227505 237052
rect 209775 236994 209780 237050
rect 209836 236994 227444 237050
rect 227500 236994 227505 237050
rect 209775 236992 227505 236994
rect 209775 236989 209841 236992
rect 227439 236989 227505 236992
rect 289071 237052 289137 237055
rect 312783 237052 312849 237055
rect 289071 237050 312849 237052
rect 289071 236994 289076 237050
rect 289132 236994 312788 237050
rect 312844 236994 312849 237050
rect 289071 236992 312849 236994
rect 289071 236989 289137 236992
rect 312783 236989 312849 236992
rect 319695 237052 319761 237055
rect 339759 237052 339825 237055
rect 319695 237050 339825 237052
rect 319695 236994 319700 237050
rect 319756 236994 339764 237050
rect 339820 236994 339825 237050
rect 319695 236992 339825 236994
rect 319695 236989 319761 236992
rect 339759 236989 339825 236992
rect 146223 236904 146289 236907
rect 140802 236902 146289 236904
rect 140802 236846 146228 236902
rect 146284 236846 146289 236902
rect 140802 236844 146289 236846
rect 146223 236841 146289 236844
rect 209679 236904 209745 236907
rect 675759 236906 675825 236907
rect 209679 236902 212862 236904
rect 209679 236846 209684 236902
rect 209740 236846 212862 236902
rect 360066 236867 380094 236904
rect 380175 236867 380241 236870
rect 209679 236844 212862 236846
rect 209679 236841 209745 236844
rect 210874 236694 210880 236758
rect 210944 236756 210950 236758
rect 212655 236756 212721 236759
rect 210944 236754 212721 236756
rect 210944 236698 212660 236754
rect 212716 236698 212721 236754
rect 210944 236696 212721 236698
rect 210944 236694 210950 236696
rect 212655 236693 212721 236696
rect 42351 236610 42417 236611
rect 42298 236608 42304 236610
rect 42260 236548 42304 236608
rect 42368 236606 42417 236610
rect 42412 236550 42417 236606
rect 42298 236546 42304 236548
rect 42368 236546 42417 236550
rect 210682 236546 210688 236610
rect 210752 236608 210758 236610
rect 211887 236608 211953 236611
rect 210752 236606 211953 236608
rect 210752 236550 211892 236606
rect 211948 236550 211953 236606
rect 210752 236548 211953 236550
rect 210752 236546 210758 236548
rect 42351 236545 42417 236546
rect 211887 236545 211953 236548
rect 210490 236398 210496 236462
rect 210560 236460 210566 236462
rect 211311 236460 211377 236463
rect 210560 236458 211377 236460
rect 210560 236402 211316 236458
rect 211372 236402 211377 236458
rect 210560 236400 211377 236402
rect 212802 236460 212862 236844
rect 279426 236807 279870 236867
rect 227631 236756 227697 236759
rect 239055 236756 239121 236759
rect 227631 236754 239121 236756
rect 227631 236698 227636 236754
rect 227692 236698 239060 236754
rect 239116 236698 239121 236754
rect 227631 236696 239121 236698
rect 227631 236693 227697 236696
rect 239055 236693 239121 236696
rect 259119 236756 259185 236759
rect 279426 236756 279486 236807
rect 259119 236754 279486 236756
rect 259119 236698 259124 236754
rect 259180 236698 279486 236754
rect 259119 236696 279486 236698
rect 279810 236756 279870 236807
rect 360018 236865 380241 236867
rect 360018 236844 380180 236865
rect 360018 236807 360126 236844
rect 380034 236809 380180 236844
rect 380236 236809 380241 236865
rect 380034 236807 380241 236809
rect 299202 236756 299646 236793
rect 319695 236756 319761 236759
rect 279810 236754 319761 236756
rect 279810 236733 319700 236754
rect 279810 236696 299262 236733
rect 299586 236698 319700 236733
rect 319756 236698 319761 236754
rect 299586 236696 319761 236698
rect 259119 236693 259185 236696
rect 319695 236693 319761 236696
rect 339759 236756 339825 236759
rect 360018 236756 360078 236807
rect 380175 236804 380241 236807
rect 400386 236844 403326 236904
rect 339759 236754 360078 236756
rect 339759 236698 339764 236754
rect 339820 236698 360078 236754
rect 339759 236696 360078 236698
rect 390159 236756 390225 236759
rect 400386 236756 400446 236844
rect 390159 236754 400446 236756
rect 390159 236698 390164 236754
rect 390220 236698 400446 236754
rect 390159 236696 400446 236698
rect 403266 236756 403326 236844
rect 675706 236842 675712 236906
rect 675776 236904 675825 236906
rect 675776 236902 675868 236904
rect 675820 236846 675868 236902
rect 675776 236844 675868 236846
rect 675776 236842 675825 236844
rect 675759 236841 675825 236842
rect 420495 236756 420561 236759
rect 403266 236754 420561 236756
rect 403266 236698 420500 236754
rect 420556 236698 420561 236754
rect 403266 236696 420561 236698
rect 339759 236693 339825 236696
rect 390159 236693 390225 236696
rect 420495 236693 420561 236696
rect 440559 236756 440625 236759
rect 460815 236756 460881 236759
rect 440559 236754 460881 236756
rect 440559 236698 440564 236754
rect 440620 236698 460820 236754
rect 460876 236698 460881 236754
rect 440559 236696 460881 236698
rect 440559 236693 440625 236696
rect 460815 236693 460881 236696
rect 480879 236756 480945 236759
rect 497487 236756 497553 236759
rect 480879 236754 497553 236756
rect 480879 236698 480884 236754
rect 480940 236698 497492 236754
rect 497548 236698 497553 236754
rect 480879 236696 497553 236698
rect 480879 236693 480945 236696
rect 497487 236693 497553 236696
rect 214767 236608 214833 236611
rect 302458 236608 302464 236610
rect 214767 236606 302464 236608
rect 214767 236550 214772 236606
rect 214828 236550 302464 236606
rect 214767 236548 302464 236550
rect 214767 236545 214833 236548
rect 302458 236546 302464 236548
rect 302528 236546 302534 236610
rect 302842 236546 302848 236610
rect 302912 236608 302918 236610
rect 359247 236608 359313 236611
rect 302912 236606 359313 236608
rect 302912 236550 359252 236606
rect 359308 236550 359313 236606
rect 302912 236548 359313 236550
rect 302912 236546 302918 236548
rect 359247 236545 359313 236548
rect 420591 236460 420657 236463
rect 212802 236458 420657 236460
rect 212802 236402 420596 236458
rect 420652 236402 420657 236458
rect 212802 236400 420657 236402
rect 210560 236398 210566 236400
rect 211311 236397 211377 236400
rect 420591 236397 420657 236400
rect 144015 236312 144081 236315
rect 140802 236310 144081 236312
rect 140802 236254 144020 236310
rect 144076 236254 144081 236310
rect 140802 236252 144081 236254
rect 140802 236210 140862 236252
rect 144015 236249 144081 236252
rect 210298 236250 210304 236314
rect 210368 236312 210374 236314
rect 212271 236312 212337 236315
rect 210368 236310 212337 236312
rect 210368 236254 212276 236310
rect 212332 236254 212337 236310
rect 210368 236252 212337 236254
rect 210368 236250 210374 236252
rect 212271 236249 212337 236252
rect 290703 236312 290769 236315
rect 294063 236312 294129 236315
rect 290703 236310 294129 236312
rect 290703 236254 290708 236310
rect 290764 236254 294068 236310
rect 294124 236254 294129 236310
rect 290703 236252 294129 236254
rect 290703 236249 290769 236252
rect 294063 236249 294129 236252
rect 638415 236312 638481 236315
rect 639279 236312 639345 236315
rect 638415 236310 639345 236312
rect 638415 236254 638420 236310
rect 638476 236254 639284 236310
rect 639340 236254 639345 236310
rect 638415 236252 639345 236254
rect 638415 236249 638481 236252
rect 639279 236249 639345 236252
rect 225807 236164 225873 236167
rect 344751 236164 344817 236167
rect 225807 236162 344817 236164
rect 225807 236106 225812 236162
rect 225868 236106 344756 236162
rect 344812 236106 344817 236162
rect 225807 236104 344817 236106
rect 225807 236101 225873 236104
rect 344751 236101 344817 236104
rect 229551 236016 229617 236019
rect 345999 236016 346065 236019
rect 229551 236014 346065 236016
rect 229551 235958 229556 236014
rect 229612 235958 346004 236014
rect 346060 235958 346065 236014
rect 229551 235956 346065 235958
rect 229551 235953 229617 235956
rect 345999 235953 346065 235956
rect 224463 235868 224529 235871
rect 343791 235868 343857 235871
rect 224463 235866 343857 235868
rect 224463 235810 224468 235866
rect 224524 235810 343796 235866
rect 343852 235810 343857 235866
rect 224463 235808 343857 235810
rect 224463 235805 224529 235808
rect 343791 235805 343857 235808
rect 219759 235720 219825 235723
rect 341583 235720 341649 235723
rect 219759 235718 341649 235720
rect 219759 235662 219764 235718
rect 219820 235662 341588 235718
rect 341644 235662 341649 235718
rect 219759 235660 341649 235662
rect 219759 235657 219825 235660
rect 341583 235657 341649 235660
rect 221295 235572 221361 235575
rect 342543 235572 342609 235575
rect 221295 235570 342609 235572
rect 221295 235514 221300 235570
rect 221356 235514 342548 235570
rect 342604 235514 342609 235570
rect 221295 235512 342609 235514
rect 221295 235509 221361 235512
rect 342543 235509 342609 235512
rect 223023 235424 223089 235427
rect 343311 235424 343377 235427
rect 223023 235422 343377 235424
rect 223023 235366 223028 235422
rect 223084 235366 343316 235422
rect 343372 235366 343377 235422
rect 223023 235364 343377 235366
rect 223023 235361 223089 235364
rect 343311 235361 343377 235364
rect 218223 235276 218289 235279
rect 341103 235276 341169 235279
rect 218223 235274 341169 235276
rect 218223 235218 218228 235274
rect 218284 235218 341108 235274
rect 341164 235218 341169 235274
rect 218223 235216 341169 235218
rect 218223 235213 218289 235216
rect 341103 235213 341169 235216
rect 146511 235128 146577 235131
rect 140832 235126 146577 235128
rect 140832 235070 146516 235126
rect 146572 235070 146577 235126
rect 140832 235068 146577 235070
rect 146511 235065 146577 235068
rect 212367 235128 212433 235131
rect 334959 235128 335025 235131
rect 212367 235126 335025 235128
rect 212367 235070 212372 235126
rect 212428 235070 334964 235126
rect 335020 235070 335025 235126
rect 212367 235068 335025 235070
rect 212367 235065 212433 235068
rect 334959 235065 335025 235068
rect 214095 234980 214161 234983
rect 348207 234980 348273 234983
rect 214095 234978 348273 234980
rect 214095 234922 214100 234978
rect 214156 234922 348212 234978
rect 348268 234922 348273 234978
rect 214095 234920 348273 234922
rect 214095 234917 214161 234920
rect 348207 234917 348273 234920
rect 210159 234832 210225 234835
rect 379407 234832 379473 234835
rect 210159 234830 379473 234832
rect 210159 234774 210164 234830
rect 210220 234774 379412 234830
rect 379468 234774 379473 234830
rect 210159 234772 379473 234774
rect 210159 234769 210225 234772
rect 379407 234769 379473 234772
rect 211450 234622 211456 234686
rect 211520 234684 211526 234686
rect 547119 234684 547185 234687
rect 211520 234682 547185 234684
rect 211520 234626 547124 234682
rect 547180 234626 547185 234682
rect 211520 234624 547185 234626
rect 211520 234622 211526 234624
rect 547119 234621 547185 234624
rect 238671 234536 238737 234539
rect 349167 234536 349233 234539
rect 238671 234534 349233 234536
rect 238671 234478 238676 234534
rect 238732 234478 349172 234534
rect 349228 234478 349233 234534
rect 238671 234476 349233 234478
rect 238671 234473 238737 234476
rect 349167 234473 349233 234476
rect 238191 234388 238257 234391
rect 347727 234388 347793 234391
rect 238191 234386 347793 234388
rect 238191 234330 238196 234386
rect 238252 234330 347732 234386
rect 347788 234330 347793 234386
rect 238191 234328 347793 234330
rect 238191 234325 238257 234328
rect 347727 234325 347793 234328
rect 283407 234240 283473 234243
rect 298383 234240 298449 234243
rect 283407 234238 298449 234240
rect 283407 234182 283412 234238
rect 283468 234182 298388 234238
rect 298444 234182 298449 234238
rect 283407 234180 298449 234182
rect 283407 234177 283473 234180
rect 298383 234177 298449 234180
rect 284943 234092 285009 234095
rect 299151 234092 299217 234095
rect 284943 234090 299217 234092
rect 284943 234034 284948 234090
rect 285004 234034 299156 234090
rect 299212 234034 299217 234090
rect 284943 234032 299217 234034
rect 284943 234029 285009 234032
rect 299151 234029 299217 234032
rect 636922 234030 636928 234094
rect 636992 234092 636998 234094
rect 638031 234092 638097 234095
rect 636992 234090 638097 234092
rect 636992 234034 638036 234090
rect 638092 234034 638097 234090
rect 636992 234032 638097 234034
rect 636992 234030 636998 234032
rect 638031 234029 638097 234032
rect 289935 233944 290001 233947
rect 295791 233944 295857 233947
rect 637935 233946 638001 233947
rect 637882 233944 637888 233946
rect 289935 233942 295857 233944
rect 289935 233886 289940 233942
rect 289996 233886 295796 233942
rect 295852 233886 295857 233942
rect 289935 233884 295857 233886
rect 637844 233884 637888 233944
rect 637952 233942 638001 233946
rect 637996 233886 638001 233942
rect 289935 233881 290001 233884
rect 295791 233881 295857 233884
rect 637882 233882 637888 233884
rect 637952 233882 638001 233886
rect 637935 233881 638001 233882
rect 140802 233648 140862 233840
rect 637498 233734 637504 233798
rect 637568 233796 637574 233798
rect 638799 233796 638865 233799
rect 637568 233794 638865 233796
rect 637568 233738 638804 233794
rect 638860 233738 638865 233794
rect 637568 233736 638865 233738
rect 637568 233734 637574 233736
rect 638799 233733 638865 233736
rect 144015 233648 144081 233651
rect 140802 233646 144081 233648
rect 140802 233590 144020 233646
rect 144076 233590 144081 233646
rect 140802 233588 144081 233590
rect 144015 233585 144081 233588
rect 212175 233648 212241 233651
rect 637167 233650 637233 233651
rect 212410 233648 212416 233650
rect 212175 233646 212416 233648
rect 212175 233590 212180 233646
rect 212236 233590 212416 233646
rect 212175 233588 212416 233590
rect 212175 233585 212241 233588
rect 212410 233586 212416 233588
rect 212480 233586 212486 233650
rect 637114 233648 637120 233650
rect 637076 233588 637120 233648
rect 637184 233646 637233 233650
rect 637228 233590 637233 233646
rect 637114 233586 637120 233588
rect 637184 233586 637233 233590
rect 637306 233586 637312 233650
rect 637376 233648 637382 233650
rect 638895 233648 638961 233651
rect 637376 233646 638961 233648
rect 637376 233590 638900 233646
rect 638956 233590 638961 233646
rect 637376 233588 638961 233590
rect 637376 233586 637382 233588
rect 637167 233585 637233 233586
rect 638895 233585 638961 233588
rect 211791 233500 211857 233503
rect 212559 233502 212625 233503
rect 212847 233502 212913 233503
rect 212218 233500 212224 233502
rect 211791 233498 212224 233500
rect 211791 233442 211796 233498
rect 211852 233442 212224 233498
rect 211791 233440 212224 233442
rect 211791 233437 211857 233440
rect 212218 233438 212224 233440
rect 212288 233438 212294 233502
rect 212559 233498 212608 233502
rect 212672 233500 212678 233502
rect 212559 233442 212564 233498
rect 212559 233438 212608 233442
rect 212672 233440 212716 233500
rect 212672 233438 212678 233440
rect 212794 233438 212800 233502
rect 212864 233500 212913 233502
rect 214287 233500 214353 233503
rect 212864 233498 212956 233500
rect 212908 233442 212956 233498
rect 212864 233440 212956 233442
rect 213186 233498 214353 233500
rect 213186 233442 214292 233498
rect 214348 233442 214353 233498
rect 213186 233440 214353 233442
rect 212864 233438 212913 233440
rect 212559 233437 212625 233438
rect 212847 233437 212913 233438
rect 41338 233290 41344 233354
rect 41408 233352 41414 233354
rect 41775 233352 41841 233355
rect 41408 233350 41841 233352
rect 41408 233294 41780 233350
rect 41836 233294 41841 233350
rect 41408 233292 41841 233294
rect 41408 233290 41414 233292
rect 41775 233289 41841 233292
rect 210874 233290 210880 233354
rect 210944 233352 210950 233354
rect 213186 233352 213246 233440
rect 214287 233437 214353 233440
rect 289839 233500 289905 233503
rect 296079 233500 296145 233503
rect 289839 233498 296145 233500
rect 289839 233442 289844 233498
rect 289900 233442 296084 233498
rect 296140 233442 296145 233498
rect 289839 233440 296145 233442
rect 289839 233437 289905 233440
rect 296079 233437 296145 233440
rect 637690 233438 637696 233502
rect 637760 233500 637766 233502
rect 638223 233500 638289 233503
rect 637760 233498 638289 233500
rect 637760 233442 638228 233498
rect 638284 233442 638289 233498
rect 637760 233440 638289 233442
rect 637760 233438 637766 233440
rect 638223 233437 638289 233440
rect 210944 233292 213246 233352
rect 210944 233290 210950 233292
rect 140802 232168 140862 232656
rect 204591 232612 204657 232615
rect 205263 232612 205329 232615
rect 210498 232612 210558 232656
rect 204591 232610 210558 232612
rect 204591 232554 204596 232610
rect 204652 232554 205268 232610
rect 205324 232554 210558 232610
rect 204591 232552 210558 232554
rect 640386 232612 640446 232656
rect 646287 232612 646353 232615
rect 650031 232612 650097 232615
rect 640386 232610 650097 232612
rect 640386 232554 646292 232610
rect 646348 232554 650036 232610
rect 650092 232554 650097 232610
rect 640386 232552 650097 232554
rect 204591 232549 204657 232552
rect 205263 232549 205329 232552
rect 646287 232549 646353 232552
rect 650031 232549 650097 232552
rect 144111 232168 144177 232171
rect 140802 232166 144177 232168
rect 140802 232110 144116 232166
rect 144172 232110 144177 232166
rect 140802 232108 144177 232110
rect 144111 232105 144177 232108
rect 204687 232168 204753 232171
rect 209199 232168 209265 232171
rect 204687 232166 210528 232168
rect 204687 232110 204692 232166
rect 204748 232110 209204 232166
rect 209260 232110 210528 232166
rect 204687 232108 210528 232110
rect 204687 232105 204753 232108
rect 209199 232105 209265 232108
rect 640386 232020 640446 232138
rect 645519 232020 645585 232023
rect 640386 232018 645585 232020
rect 640386 231962 645524 232018
rect 645580 231962 645585 232018
rect 640386 231960 645585 231962
rect 645519 231957 645585 231960
rect 41967 231726 42033 231727
rect 41914 231662 41920 231726
rect 41984 231724 42033 231726
rect 41984 231722 42076 231724
rect 42028 231666 42076 231722
rect 41984 231664 42076 231666
rect 41984 231662 42033 231664
rect 41967 231661 42033 231662
rect 204495 231576 204561 231579
rect 209487 231576 209553 231579
rect 645135 231576 645201 231579
rect 204495 231574 210528 231576
rect 204495 231518 204500 231574
rect 204556 231518 209492 231574
rect 209548 231518 210528 231574
rect 204495 231516 210528 231518
rect 640416 231574 645201 231576
rect 640416 231518 645140 231574
rect 645196 231518 645201 231574
rect 640416 231516 645201 231518
rect 204495 231513 204561 231516
rect 209487 231513 209553 231516
rect 645135 231513 645201 231516
rect 144015 231428 144081 231431
rect 140832 231426 144081 231428
rect 140832 231370 144020 231426
rect 144076 231370 144081 231426
rect 140832 231368 144081 231370
rect 144015 231365 144081 231368
rect 41775 231134 41841 231135
rect 41722 231070 41728 231134
rect 41792 231132 41841 231134
rect 645231 231132 645297 231135
rect 41792 231130 41884 231132
rect 41836 231074 41884 231130
rect 41792 231072 41884 231074
rect 640386 231130 645297 231132
rect 640386 231074 645236 231130
rect 645292 231074 645297 231130
rect 640386 231072 645297 231074
rect 41792 231070 41841 231072
rect 41775 231069 41841 231070
rect 204783 230984 204849 230987
rect 208047 230984 208113 230987
rect 204783 230982 210528 230984
rect 204783 230926 204788 230982
rect 204844 230926 208052 230982
rect 208108 230926 210528 230982
rect 640386 230954 640446 231072
rect 645231 231069 645297 231072
rect 204783 230924 210528 230926
rect 204783 230921 204849 230924
rect 208047 230921 208113 230924
rect 645327 230688 645393 230691
rect 640194 230686 645393 230688
rect 640194 230630 645332 230686
rect 645388 230630 645393 230686
rect 640194 230628 645393 230630
rect 205455 230540 205521 230543
rect 209391 230540 209457 230543
rect 205455 230538 210528 230540
rect 205455 230482 205460 230538
rect 205516 230482 209396 230538
rect 209452 230482 210528 230538
rect 640194 230510 640254 230628
rect 645327 230625 645393 230628
rect 205455 230480 210528 230482
rect 205455 230477 205521 230480
rect 209391 230477 209457 230480
rect 41530 230330 41536 230394
rect 41600 230392 41606 230394
rect 41775 230392 41841 230395
rect 41600 230390 41841 230392
rect 41600 230334 41780 230390
rect 41836 230334 41841 230390
rect 41600 230332 41841 230334
rect 41600 230330 41606 230332
rect 41775 230329 41841 230332
rect 144207 230244 144273 230247
rect 140832 230242 144273 230244
rect 140832 230186 144212 230242
rect 144268 230186 144273 230242
rect 140832 230184 144273 230186
rect 144207 230181 144273 230184
rect 207279 229948 207345 229951
rect 207279 229946 210528 229948
rect 207279 229890 207284 229946
rect 207340 229890 210528 229946
rect 207279 229888 210528 229890
rect 207279 229885 207345 229888
rect 41146 229590 41152 229654
rect 41216 229652 41222 229654
rect 41775 229652 41841 229655
rect 41216 229650 41841 229652
rect 41216 229594 41780 229650
rect 41836 229594 41841 229650
rect 41216 229592 41841 229594
rect 41216 229590 41222 229592
rect 41775 229589 41841 229592
rect 206127 229356 206193 229359
rect 206127 229354 210528 229356
rect 206127 229298 206132 229354
rect 206188 229298 210528 229354
rect 206127 229296 210528 229298
rect 206127 229293 206193 229296
rect 40762 228998 40768 229062
rect 40832 229060 40838 229062
rect 41775 229060 41841 229063
rect 40832 229058 41841 229060
rect 40832 229002 41780 229058
rect 41836 229002 41841 229058
rect 40832 229000 41841 229002
rect 40832 228998 40838 229000
rect 41775 228997 41841 229000
rect 140802 228468 140862 228956
rect 210159 228912 210225 228915
rect 210159 228910 210528 228912
rect 210159 228854 210164 228910
rect 210220 228854 210528 228910
rect 210159 228852 210528 228854
rect 210159 228849 210225 228852
rect 144111 228468 144177 228471
rect 140802 228466 144177 228468
rect 140802 228410 144116 228466
rect 144172 228410 144177 228466
rect 140802 228408 144177 228410
rect 144111 228405 144177 228408
rect 205935 228320 206001 228323
rect 205935 228318 210528 228320
rect 205935 228262 205940 228318
rect 205996 228262 210528 228318
rect 205935 228260 210528 228262
rect 205935 228257 206001 228260
rect 140802 227876 140862 227914
rect 144015 227876 144081 227879
rect 140802 227874 144081 227876
rect 140802 227818 144020 227874
rect 144076 227818 144081 227874
rect 140802 227816 144081 227818
rect 144015 227813 144081 227816
rect 204975 227728 205041 227731
rect 204975 227726 210528 227728
rect 204975 227670 204980 227726
rect 205036 227670 210528 227726
rect 204975 227668 210528 227670
rect 204975 227665 205041 227668
rect 40570 227370 40576 227434
rect 40640 227432 40646 227434
rect 41775 227432 41841 227435
rect 40640 227430 41841 227432
rect 40640 227374 41780 227430
rect 41836 227374 41841 227430
rect 40640 227372 41841 227374
rect 40640 227370 40646 227372
rect 41775 227369 41841 227372
rect 206895 227432 206961 227435
rect 207087 227432 207153 227435
rect 206895 227430 207153 227432
rect 206895 227374 206900 227430
rect 206956 227374 207092 227430
rect 207148 227374 207153 227430
rect 206895 227372 207153 227374
rect 206895 227369 206961 227372
rect 207087 227369 207153 227372
rect 205743 227284 205809 227287
rect 205743 227282 210528 227284
rect 205743 227226 205748 227282
rect 205804 227226 210528 227282
rect 205743 227224 210528 227226
rect 205743 227221 205809 227224
rect 40954 226778 40960 226842
rect 41024 226840 41030 226842
rect 41775 226840 41841 226843
rect 41024 226838 41841 226840
rect 41024 226782 41780 226838
rect 41836 226782 41841 226838
rect 41024 226780 41841 226782
rect 41024 226778 41030 226780
rect 41775 226777 41841 226780
rect 146799 226692 146865 226695
rect 140832 226690 146865 226692
rect 140832 226634 146804 226690
rect 146860 226634 146865 226690
rect 140832 226632 146865 226634
rect 146799 226629 146865 226632
rect 205359 226692 205425 226695
rect 205359 226690 210528 226692
rect 205359 226634 205364 226690
rect 205420 226634 210528 226690
rect 205359 226632 210528 226634
rect 205359 226629 205425 226632
rect 205551 226100 205617 226103
rect 205551 226098 210528 226100
rect 205551 226042 205556 226098
rect 205612 226042 210528 226098
rect 205551 226040 210528 226042
rect 205551 226037 205617 226040
rect 40378 225890 40384 225954
rect 40448 225952 40454 225954
rect 41775 225952 41841 225955
rect 40448 225950 41841 225952
rect 40448 225894 41780 225950
rect 41836 225894 41841 225950
rect 40448 225892 41841 225894
rect 40448 225890 40454 225892
rect 41775 225889 41841 225892
rect 205167 225656 205233 225659
rect 205167 225654 210528 225656
rect 205167 225598 205172 225654
rect 205228 225598 210528 225654
rect 205167 225596 210528 225598
rect 205167 225593 205233 225596
rect 140802 225064 140862 225466
rect 146127 225064 146193 225067
rect 140802 225062 146193 225064
rect 140802 225006 146132 225062
rect 146188 225006 146193 225062
rect 140802 225004 146193 225006
rect 146127 225001 146193 225004
rect 206895 225064 206961 225067
rect 674703 225064 674769 225067
rect 206895 225062 210528 225064
rect 206895 225006 206900 225062
rect 206956 225006 210528 225062
rect 206895 225004 210528 225006
rect 674703 225062 674814 225064
rect 674703 225006 674708 225062
rect 674764 225006 674814 225062
rect 206895 225001 206961 225004
rect 674703 225001 674814 225006
rect 674754 224886 674814 225001
rect 206991 224472 207057 224475
rect 206991 224470 210528 224472
rect 206991 224414 206996 224470
rect 207052 224414 210528 224470
rect 206991 224412 210528 224414
rect 206991 224409 207057 224412
rect 674415 224324 674481 224327
rect 674415 224322 674784 224324
rect 674415 224266 674420 224322
rect 674476 224266 674784 224322
rect 674415 224264 674784 224266
rect 674415 224261 674481 224264
rect 140802 223732 140862 224220
rect 204495 224028 204561 224031
rect 674703 224028 674769 224031
rect 204495 224026 210528 224028
rect 204495 223970 204500 224026
rect 204556 223970 210528 224026
rect 204495 223968 210528 223970
rect 674703 224026 674814 224028
rect 674703 223970 674708 224026
rect 674764 223970 674814 224026
rect 204495 223965 204561 223968
rect 674703 223965 674814 223970
rect 674754 223776 674814 223965
rect 144399 223732 144465 223735
rect 140802 223730 144465 223732
rect 140802 223674 144404 223730
rect 144460 223674 144465 223730
rect 140802 223672 144465 223674
rect 144399 223669 144465 223672
rect 677242 223522 677248 223586
rect 677312 223522 677318 223586
rect 204591 223436 204657 223439
rect 204591 223434 210528 223436
rect 204591 223378 204596 223434
rect 204652 223378 210528 223434
rect 204591 223376 210528 223378
rect 204591 223373 204657 223376
rect 677250 223258 677310 223522
rect 146799 222992 146865 222995
rect 140832 222990 146865 222992
rect 140832 222934 146804 222990
rect 146860 222934 146865 222990
rect 140832 222932 146865 222934
rect 146799 222929 146865 222932
rect 204687 222844 204753 222847
rect 204687 222842 210528 222844
rect 204687 222786 204692 222842
rect 204748 222786 210528 222842
rect 204687 222784 210528 222786
rect 204687 222781 204753 222784
rect 206799 222400 206865 222403
rect 677250 222402 677310 222666
rect 206799 222398 210528 222400
rect 206799 222342 206804 222398
rect 206860 222342 210528 222398
rect 206799 222340 210528 222342
rect 206799 222337 206865 222340
rect 676858 222338 676864 222402
rect 676928 222338 676934 222402
rect 677242 222338 677248 222402
rect 677312 222338 677318 222402
rect 676866 222178 676926 222338
rect 676866 222148 677664 222178
rect 676896 222118 677694 222148
rect 146703 221808 146769 221811
rect 140832 221806 146769 221808
rect 140832 221750 146708 221806
rect 146764 221750 146769 221806
rect 140832 221748 146769 221750
rect 146703 221745 146769 221748
rect 204783 221808 204849 221811
rect 646095 221808 646161 221811
rect 646287 221808 646353 221811
rect 677634 221810 677694 222118
rect 204783 221806 210528 221808
rect 204783 221750 204788 221806
rect 204844 221750 210528 221806
rect 204783 221748 210528 221750
rect 646095 221806 646353 221808
rect 646095 221750 646100 221806
rect 646156 221750 646292 221806
rect 646348 221750 646353 221806
rect 646095 221748 646353 221750
rect 204783 221745 204849 221748
rect 646095 221745 646161 221748
rect 646287 221745 646353 221748
rect 677050 221746 677056 221810
rect 677120 221746 677126 221810
rect 677626 221746 677632 221810
rect 677696 221746 677702 221810
rect 677058 221630 677118 221746
rect 204495 221216 204561 221219
rect 204495 221214 210528 221216
rect 204495 221158 204500 221214
rect 204556 221158 210528 221214
rect 204495 221156 210528 221158
rect 204495 221153 204561 221156
rect 204591 221068 204657 221071
rect 204591 221066 210558 221068
rect 204591 221010 204596 221066
rect 204652 221010 210558 221066
rect 204591 221008 210558 221010
rect 204591 221005 204657 221008
rect 210498 220668 210558 221008
rect 674946 220923 675006 221038
rect 674895 220918 675006 220923
rect 674895 220862 674900 220918
rect 674956 220862 675006 220918
rect 674895 220860 675006 220862
rect 674895 220857 674961 220860
rect 140802 220180 140862 220668
rect 674362 220488 674368 220552
rect 674432 220550 674438 220552
rect 674432 220490 674784 220550
rect 674432 220488 674438 220490
rect 144399 220180 144465 220183
rect 140802 220178 144465 220180
rect 140802 220122 144404 220178
rect 144460 220122 144465 220178
rect 140802 220120 144465 220122
rect 144399 220117 144465 220120
rect 204687 220180 204753 220183
rect 204687 220178 210528 220180
rect 204687 220122 204692 220178
rect 204748 220122 210528 220178
rect 204687 220120 210528 220122
rect 204687 220117 204753 220120
rect 675522 219739 675582 220002
rect 675471 219734 675582 219739
rect 675471 219678 675476 219734
rect 675532 219678 675582 219734
rect 675471 219676 675582 219678
rect 675471 219673 675537 219676
rect 204783 219588 204849 219591
rect 204783 219586 210528 219588
rect 204783 219530 204788 219586
rect 204844 219530 210528 219586
rect 204783 219528 210528 219530
rect 204783 219525 204849 219528
rect 140802 218996 140862 219482
rect 204879 219440 204945 219443
rect 204879 219438 210558 219440
rect 204879 219382 204884 219438
rect 204940 219382 210558 219438
rect 204879 219380 210558 219382
rect 204879 219377 204945 219380
rect 210498 219040 210558 219380
rect 674946 219295 675006 219410
rect 674946 219290 675057 219295
rect 674946 219234 674996 219290
rect 675052 219234 675057 219290
rect 674946 219232 675057 219234
rect 674991 219229 675057 219232
rect 145594 218996 145600 218998
rect 140802 218936 145600 218996
rect 145594 218934 145600 218936
rect 145664 218934 145670 218998
rect 674170 218860 674176 218924
rect 674240 218922 674246 218924
rect 674240 218862 674784 218922
rect 674240 218860 674246 218862
rect 204495 218552 204561 218555
rect 204495 218550 210528 218552
rect 204495 218494 204500 218550
rect 204556 218494 210528 218550
rect 204495 218492 210528 218494
rect 204495 218489 204561 218492
rect 146799 218256 146865 218259
rect 140832 218254 146865 218256
rect 140832 218198 146804 218254
rect 146860 218198 146865 218254
rect 140832 218196 146865 218198
rect 146799 218193 146865 218196
rect 677058 218111 677118 218374
rect 677058 218106 677169 218111
rect 677058 218050 677108 218106
rect 677164 218050 677169 218106
rect 677058 218048 677169 218050
rect 677103 218045 677169 218048
rect 204591 217960 204657 217963
rect 204591 217958 210528 217960
rect 204591 217902 204596 217958
rect 204652 217902 210528 217958
rect 204591 217900 210528 217902
rect 204591 217897 204657 217900
rect 204687 217812 204753 217815
rect 204687 217810 210558 217812
rect 204687 217754 204692 217810
rect 204748 217754 210558 217810
rect 204687 217752 210558 217754
rect 204687 217749 204753 217752
rect 210498 217412 210558 217752
rect 675138 217667 675198 217782
rect 675138 217662 675249 217667
rect 675138 217606 675188 217662
rect 675244 217606 675249 217662
rect 675138 217604 675249 217606
rect 675183 217601 675249 217604
rect 140802 216480 140862 217034
rect 210490 217010 210496 217074
rect 210560 217072 210566 217074
rect 211066 217072 211072 217074
rect 210560 217012 211072 217072
rect 210560 217010 210566 217012
rect 211066 217010 211072 217012
rect 211136 217010 211142 217074
rect 675138 216927 675198 217264
rect 204783 216924 204849 216927
rect 204783 216922 210528 216924
rect 204783 216866 204788 216922
rect 204844 216866 210528 216922
rect 204783 216864 210528 216866
rect 675087 216922 675198 216927
rect 675087 216866 675092 216922
rect 675148 216866 675198 216922
rect 675087 216864 675198 216866
rect 204783 216861 204849 216864
rect 675087 216861 675153 216864
rect 674223 216776 674289 216779
rect 674223 216774 674784 216776
rect 674223 216718 674228 216774
rect 674284 216718 674784 216774
rect 674223 216716 674784 216718
rect 674223 216713 674289 216716
rect 145786 216480 145792 216482
rect 140802 216420 145792 216480
rect 145786 216418 145792 216420
rect 145856 216418 145862 216482
rect 42735 216332 42801 216335
rect 42528 216330 42801 216332
rect 42528 216274 42740 216330
rect 42796 216274 42801 216330
rect 42528 216272 42801 216274
rect 42735 216269 42801 216272
rect 206703 216332 206769 216335
rect 206703 216330 210528 216332
rect 206703 216274 206708 216330
rect 206764 216274 210528 216330
rect 206703 216272 210528 216274
rect 206703 216269 206769 216272
rect 676866 216039 676926 216154
rect 676866 216034 676977 216039
rect 676866 215978 676916 216034
rect 676972 215978 676977 216034
rect 676866 215976 676977 215978
rect 676911 215973 676977 215976
rect 204495 215888 204561 215891
rect 204495 215886 210558 215888
rect 204495 215830 204500 215886
rect 204556 215830 210558 215886
rect 204495 215828 210558 215830
rect 204495 215825 204561 215828
rect 210498 215784 210558 215828
rect 42735 215740 42801 215743
rect 42528 215738 42801 215740
rect 42528 215682 42740 215738
rect 42796 215682 42801 215738
rect 42528 215680 42801 215682
rect 42735 215677 42801 215680
rect 140802 215296 140862 215784
rect 674511 215444 674577 215447
rect 674754 215444 674814 215562
rect 674511 215442 674814 215444
rect 674511 215386 674516 215442
rect 674572 215386 674814 215442
rect 674511 215384 674814 215386
rect 674511 215381 674577 215384
rect 144399 215296 144465 215299
rect 140802 215294 144465 215296
rect 140802 215238 144404 215294
rect 144460 215238 144465 215294
rect 140802 215236 144465 215238
rect 144399 215233 144465 215236
rect 204591 215296 204657 215299
rect 204591 215294 210528 215296
rect 204591 215238 204596 215294
rect 204652 215238 210528 215294
rect 204591 215236 210528 215238
rect 204591 215233 204657 215236
rect 42735 215222 42801 215225
rect 42528 215220 42801 215222
rect 42528 215164 42740 215220
rect 42796 215164 42801 215220
rect 42528 215162 42801 215164
rect 42735 215159 42801 215162
rect 674754 214855 674814 215118
rect 674754 214850 674865 214855
rect 674754 214794 674804 214850
rect 674860 214794 674865 214850
rect 674754 214792 674865 214794
rect 674799 214789 674865 214792
rect 206319 214704 206385 214707
rect 206319 214702 210528 214704
rect 206319 214646 206324 214702
rect 206380 214646 210528 214702
rect 206319 214644 210528 214646
rect 206319 214641 206385 214644
rect 145359 214556 145425 214559
rect 140832 214554 145425 214556
rect 140832 214498 145364 214554
rect 145420 214498 145425 214554
rect 140832 214496 145425 214498
rect 145359 214493 145425 214496
rect 206223 214556 206289 214559
rect 206223 214554 210558 214556
rect 206223 214498 206228 214554
rect 206284 214498 210558 214554
rect 206223 214496 210558 214498
rect 206223 214493 206289 214496
rect 210498 214156 210558 214496
rect 674754 214411 674814 214526
rect 674703 214406 674814 214411
rect 674703 214350 674708 214406
rect 674764 214350 674814 214406
rect 674703 214348 674814 214350
rect 674703 214345 674769 214348
rect 43215 214112 43281 214115
rect 42528 214110 43281 214112
rect 42528 214054 43220 214110
rect 43276 214054 43281 214110
rect 42528 214052 43281 214054
rect 43215 214049 43281 214052
rect 674607 213816 674673 213819
rect 674754 213816 674814 213934
rect 674607 213814 674814 213816
rect 674607 213758 674612 213814
rect 674668 213758 674814 213814
rect 674607 213756 674814 213758
rect 674607 213753 674673 213756
rect 43407 213668 43473 213671
rect 42498 213666 43473 213668
rect 42498 213610 43412 213666
rect 43468 213610 43473 213666
rect 42498 213608 43473 213610
rect 42498 213490 42558 213608
rect 43407 213605 43473 213608
rect 206415 213668 206481 213671
rect 206415 213666 210528 213668
rect 206415 213610 206420 213666
rect 206476 213610 210528 213666
rect 206415 213608 210528 213610
rect 206415 213605 206481 213608
rect 146799 213372 146865 213375
rect 140832 213370 146865 213372
rect 140832 213314 146804 213370
rect 146860 213314 146865 213370
rect 140832 213312 146865 213314
rect 146799 213309 146865 213312
rect 677058 213227 677118 213490
rect 677007 213222 677118 213227
rect 677007 213166 677012 213222
rect 677068 213166 677118 213222
rect 677007 213164 677118 213166
rect 677007 213161 677073 213164
rect 43311 213076 43377 213079
rect 42528 213074 43377 213076
rect 42528 213018 43316 213074
rect 43372 213018 43377 213074
rect 42528 213016 43377 213018
rect 43311 213013 43377 213016
rect 206607 213076 206673 213079
rect 206607 213074 210528 213076
rect 206607 213018 206612 213074
rect 206668 213018 210528 213074
rect 206607 213016 210528 213018
rect 206607 213013 206673 213016
rect 206511 212928 206577 212931
rect 206511 212926 210558 212928
rect 206511 212870 206516 212926
rect 206572 212870 210558 212926
rect 206511 212868 210558 212870
rect 206511 212865 206577 212868
rect 210498 212528 210558 212868
rect 676866 212635 676926 212898
rect 676815 212630 676926 212635
rect 676815 212574 676820 212630
rect 676876 212574 676926 212630
rect 676815 212572 676926 212574
rect 677007 212632 677073 212635
rect 677007 212630 677118 212632
rect 677007 212574 677012 212630
rect 677068 212574 677118 212630
rect 676815 212569 676881 212572
rect 677007 212569 677118 212574
rect 40578 212190 40638 212454
rect 677058 212306 677118 212569
rect 40570 212126 40576 212190
rect 40640 212126 40646 212190
rect 41922 211599 41982 211862
rect 140802 211744 140862 212232
rect 676815 212188 676881 212191
rect 676815 212186 676926 212188
rect 676815 212130 676820 212186
rect 676876 212130 676926 212186
rect 676815 212125 676926 212130
rect 205743 212040 205809 212043
rect 205743 212038 210528 212040
rect 205743 211982 205748 212038
rect 205804 211982 210528 212038
rect 205743 211980 210528 211982
rect 205743 211977 205809 211980
rect 676866 211862 676926 212125
rect 145263 211744 145329 211747
rect 140802 211742 145329 211744
rect 140802 211686 145268 211742
rect 145324 211686 145329 211742
rect 140802 211684 145329 211686
rect 145263 211681 145329 211684
rect 41922 211594 42033 211599
rect 41922 211538 41972 211594
rect 42028 211538 42033 211594
rect 41922 211536 42033 211538
rect 41967 211533 42033 211536
rect 205839 211448 205905 211451
rect 205839 211446 210528 211448
rect 40386 211154 40446 211418
rect 205839 211390 205844 211446
rect 205900 211390 210528 211446
rect 205839 211388 210528 211390
rect 205839 211385 205905 211388
rect 40378 211090 40384 211154
rect 40448 211090 40454 211154
rect 40962 210562 41022 210826
rect 40954 210498 40960 210562
rect 41024 210498 41030 210562
rect 140802 210560 140862 211048
rect 145455 210560 145521 210563
rect 140802 210558 145521 210560
rect 140802 210502 145460 210558
rect 145516 210502 145521 210558
rect 140802 210500 145521 210502
rect 145455 210497 145521 210500
rect 640194 210412 640254 210826
rect 645615 210412 645681 210415
rect 640194 210410 645681 210412
rect 640194 210354 645620 210410
rect 645676 210354 645681 210410
rect 640194 210352 645681 210354
rect 645615 210349 645681 210352
rect 42306 209971 42366 210234
rect 676474 210202 676480 210266
rect 676544 210264 676550 210266
rect 676911 210264 676977 210267
rect 676544 210262 676977 210264
rect 676544 210206 676916 210262
rect 676972 210206 676977 210262
rect 676544 210204 676977 210206
rect 676544 210202 676550 210204
rect 676911 210201 676977 210204
rect 676666 210054 676672 210118
rect 676736 210116 676742 210118
rect 677103 210116 677169 210119
rect 676736 210114 677169 210116
rect 676736 210058 677108 210114
rect 677164 210058 677169 210114
rect 676736 210056 677169 210058
rect 676736 210054 676742 210056
rect 677103 210053 677169 210056
rect 42306 209966 42417 209971
rect 42306 209910 42356 209966
rect 42412 209910 42417 209966
rect 42306 209908 42417 209910
rect 42351 209905 42417 209908
rect 146607 209820 146673 209823
rect 140832 209818 146673 209820
rect 40194 209527 40254 209790
rect 140832 209762 146612 209818
rect 146668 209762 146673 209818
rect 140832 209760 146673 209762
rect 146607 209757 146673 209760
rect 40194 209522 40305 209527
rect 40194 209466 40244 209522
rect 40300 209466 40305 209522
rect 40194 209464 40305 209466
rect 40239 209461 40305 209464
rect 40770 208934 40830 209198
rect 40762 208870 40768 208934
rect 40832 208870 40838 208934
rect 41154 208342 41214 208606
rect 41146 208278 41152 208342
rect 41216 208278 41222 208342
rect 42498 207748 42558 208162
rect 140802 208044 140862 208602
rect 145551 208044 145617 208047
rect 140802 208042 145617 208044
rect 140802 207986 145556 208042
rect 145612 207986 145617 208042
rect 140802 207984 145617 207986
rect 145551 207981 145617 207984
rect 42735 207748 42801 207751
rect 42498 207746 42801 207748
rect 42498 207690 42740 207746
rect 42796 207690 42801 207746
rect 42498 207688 42801 207690
rect 42735 207685 42801 207688
rect 42498 207304 42558 207570
rect 146799 207452 146865 207455
rect 140832 207450 146865 207452
rect 140832 207394 146804 207450
rect 146860 207394 146865 207450
rect 140832 207392 146865 207394
rect 146799 207389 146865 207392
rect 42927 207304 42993 207307
rect 42498 207302 42993 207304
rect 42498 207246 42932 207302
rect 42988 207246 42993 207302
rect 42498 207244 42993 207246
rect 42927 207241 42993 207244
rect 40194 206715 40254 206978
rect 40143 206710 40254 206715
rect 40143 206654 40148 206710
rect 40204 206654 40254 206710
rect 40143 206652 40254 206654
rect 40143 206649 40209 206652
rect 40002 206123 40062 206534
rect 676858 206354 676864 206418
rect 676928 206416 676934 206418
rect 677626 206416 677632 206418
rect 676928 206356 677632 206416
rect 676928 206354 676934 206356
rect 677626 206354 677632 206356
rect 677696 206354 677702 206418
rect 40002 206118 40113 206123
rect 40002 206062 40052 206118
rect 40108 206062 40113 206118
rect 40002 206060 40113 206062
rect 40047 206057 40113 206060
rect 40194 205679 40254 205942
rect 40194 205674 40305 205679
rect 40194 205618 40244 205674
rect 40300 205618 40305 205674
rect 40194 205616 40305 205618
rect 140802 205676 140862 206154
rect 145647 205676 145713 205679
rect 140802 205674 145713 205676
rect 140802 205618 145652 205674
rect 145708 205618 145713 205674
rect 140802 205616 145713 205618
rect 40239 205613 40305 205616
rect 145647 205613 145713 205616
rect 43023 205380 43089 205383
rect 42528 205378 43089 205380
rect 42528 205322 43028 205378
rect 43084 205322 43089 205378
rect 42528 205320 43089 205322
rect 43023 205317 43089 205320
rect 145743 205084 145809 205087
rect 140832 205082 145809 205084
rect 140832 205026 145748 205082
rect 145804 205026 145809 205082
rect 140832 205024 145809 205026
rect 145743 205021 145809 205024
rect 42735 204862 42801 204865
rect 42528 204860 42801 204862
rect 42528 204804 42740 204860
rect 42796 204804 42801 204860
rect 42528 204802 42801 204804
rect 42735 204799 42801 204802
rect 35202 204051 35262 204314
rect 35151 204046 35262 204051
rect 35151 203990 35156 204046
rect 35212 203990 35262 204046
rect 35151 203988 35262 203990
rect 35151 203985 35217 203988
rect 42735 203752 42801 203755
rect 42528 203750 42801 203752
rect 42528 203694 42740 203750
rect 42796 203694 42801 203750
rect 42528 203692 42801 203694
rect 42735 203689 42801 203692
rect 35151 203604 35217 203607
rect 35151 203602 35262 203604
rect 35151 203546 35156 203602
rect 35212 203546 35262 203602
rect 35151 203541 35262 203546
rect 35202 203204 35262 203541
rect 140802 203308 140862 203796
rect 144015 203308 144081 203311
rect 140802 203306 144081 203308
rect 140802 203250 144020 203306
rect 144076 203250 144081 203306
rect 140802 203248 144081 203250
rect 144015 203245 144081 203248
rect 207087 202716 207153 202719
rect 207087 202714 210528 202716
rect 207087 202658 207092 202714
rect 207148 202658 210528 202714
rect 207087 202656 210528 202658
rect 207087 202653 207153 202656
rect 140802 202124 140862 202612
rect 145839 202124 145905 202127
rect 140802 202122 145905 202124
rect 140802 202066 145844 202122
rect 145900 202066 145905 202122
rect 140802 202064 145905 202066
rect 145839 202061 145905 202064
rect 145743 201384 145809 201387
rect 140832 201382 145809 201384
rect 140832 201326 145748 201382
rect 145804 201326 145809 201382
rect 140832 201324 145809 201326
rect 145743 201321 145809 201324
rect 42106 201174 42112 201238
rect 42176 201236 42182 201238
rect 42351 201236 42417 201239
rect 42176 201234 42417 201236
rect 42176 201178 42356 201234
rect 42412 201178 42417 201234
rect 42176 201176 42417 201178
rect 42176 201174 42182 201176
rect 42351 201173 42417 201176
rect 140802 199608 140862 200142
rect 144495 199608 144561 199611
rect 140802 199606 144561 199608
rect 140802 199550 144500 199606
rect 144556 199550 144561 199606
rect 140802 199548 144561 199550
rect 144495 199545 144561 199548
rect 675375 199314 675441 199315
rect 675322 199250 675328 199314
rect 675392 199312 675441 199314
rect 675392 199310 675484 199312
rect 675436 199254 675484 199310
rect 675392 199252 675484 199254
rect 675392 199250 675441 199252
rect 675375 199249 675441 199250
rect 144015 199016 144081 199019
rect 140832 199014 144081 199016
rect 140832 198958 144020 199014
rect 144076 198958 144081 199014
rect 140832 198956 144081 198958
rect 144015 198953 144081 198956
rect 645903 198720 645969 198723
rect 646095 198720 646161 198723
rect 675471 198722 675537 198723
rect 675471 198720 675520 198722
rect 645903 198718 646161 198720
rect 645903 198662 645908 198718
rect 645964 198662 646100 198718
rect 646156 198662 646161 198718
rect 645903 198660 646161 198662
rect 675428 198718 675520 198720
rect 675428 198662 675476 198718
rect 675428 198660 675520 198662
rect 645903 198657 645969 198660
rect 646095 198657 646161 198660
rect 675471 198658 675520 198660
rect 675584 198658 675590 198722
rect 675471 198657 675537 198658
rect 674170 198362 674176 198426
rect 674240 198424 674246 198426
rect 675471 198424 675537 198427
rect 674240 198422 675537 198424
rect 674240 198366 675476 198422
rect 675532 198366 675537 198422
rect 674240 198364 675537 198366
rect 674240 198362 674246 198364
rect 675471 198361 675537 198364
rect 144687 197832 144753 197835
rect 140832 197830 144753 197832
rect 140832 197774 144692 197830
rect 144748 197774 144753 197830
rect 140832 197772 144753 197774
rect 144687 197769 144753 197772
rect 42159 197536 42225 197539
rect 42298 197536 42304 197538
rect 42159 197534 42304 197536
rect 42159 197478 42164 197534
rect 42220 197478 42304 197534
rect 42159 197476 42304 197478
rect 42159 197473 42225 197476
rect 42298 197474 42304 197476
rect 42368 197474 42374 197538
rect 144591 196648 144657 196651
rect 140832 196646 144657 196648
rect 140832 196590 144596 196646
rect 144652 196590 144657 196646
rect 140832 196588 144657 196590
rect 144591 196585 144657 196588
rect 42351 195170 42417 195171
rect 42298 195106 42304 195170
rect 42368 195168 42417 195170
rect 42368 195166 42460 195168
rect 42412 195110 42460 195166
rect 42368 195108 42460 195110
rect 42368 195106 42417 195108
rect 42351 195105 42417 195106
rect 140802 194872 140862 195360
rect 675759 195316 675825 195319
rect 676474 195316 676480 195318
rect 675759 195314 676480 195316
rect 675759 195258 675764 195314
rect 675820 195258 676480 195314
rect 675759 195256 676480 195258
rect 675759 195253 675825 195256
rect 676474 195254 676480 195256
rect 676544 195254 676550 195318
rect 144399 194872 144465 194875
rect 140802 194870 144465 194872
rect 140802 194814 144404 194870
rect 144460 194814 144465 194870
rect 140802 194812 144465 194814
rect 144399 194809 144465 194812
rect 140802 193688 140862 194176
rect 145935 193688 146001 193691
rect 140802 193686 146001 193688
rect 140802 193630 145940 193686
rect 145996 193630 146001 193686
rect 140802 193628 146001 193630
rect 145935 193625 146001 193628
rect 674362 193478 674368 193542
rect 674432 193540 674438 193542
rect 675375 193540 675441 193543
rect 674432 193538 675441 193540
rect 674432 193482 675380 193538
rect 675436 193482 675441 193538
rect 674432 193480 675441 193482
rect 674432 193478 674438 193480
rect 675375 193477 675441 193480
rect 144303 192948 144369 192951
rect 140832 192946 144369 192948
rect 140832 192890 144308 192946
rect 144364 192890 144369 192946
rect 140832 192888 144369 192890
rect 144303 192885 144369 192888
rect 144015 191764 144081 191767
rect 140832 191762 144081 191764
rect 140832 191706 144020 191762
rect 144076 191706 144081 191762
rect 140832 191704 144081 191706
rect 144015 191701 144081 191704
rect 210490 191554 210496 191618
rect 210560 191616 210566 191618
rect 211066 191616 211072 191618
rect 210560 191556 211072 191616
rect 210560 191554 210566 191556
rect 211066 191554 211072 191556
rect 211136 191554 211142 191618
rect 675759 191616 675825 191619
rect 676666 191616 676672 191618
rect 675759 191614 676672 191616
rect 675759 191558 675764 191614
rect 675820 191558 676672 191614
rect 675759 191556 676672 191558
rect 675759 191553 675825 191556
rect 676666 191554 676672 191556
rect 676736 191554 676742 191618
rect 42063 190286 42129 190287
rect 42063 190284 42112 190286
rect 42020 190282 42112 190284
rect 42020 190226 42068 190282
rect 42020 190224 42112 190226
rect 42063 190222 42112 190224
rect 42176 190222 42182 190286
rect 42063 190221 42129 190222
rect 140802 190136 140862 190476
rect 146031 190136 146097 190139
rect 140802 190134 146097 190136
rect 140802 190078 146036 190134
rect 146092 190078 146097 190134
rect 140802 190076 146097 190078
rect 146031 190073 146097 190076
rect 146223 189396 146289 189399
rect 140832 189394 146289 189396
rect 140832 189338 146228 189394
rect 146284 189338 146289 189394
rect 140832 189336 146289 189338
rect 146223 189333 146289 189336
rect 41967 189102 42033 189103
rect 41914 189100 41920 189102
rect 41876 189040 41920 189100
rect 41984 189098 42033 189102
rect 42028 189042 42033 189098
rect 41914 189038 41920 189040
rect 41984 189038 42033 189042
rect 41967 189037 42033 189038
rect 41775 188362 41841 188363
rect 41722 188298 41728 188362
rect 41792 188360 41841 188362
rect 41792 188358 41884 188360
rect 41836 188302 41884 188358
rect 41792 188300 41884 188302
rect 41792 188298 41841 188300
rect 41775 188297 41841 188298
rect 144015 188212 144081 188215
rect 140832 188210 144081 188212
rect 140832 188154 144020 188210
rect 144076 188154 144081 188210
rect 140832 188152 144081 188154
rect 144015 188149 144081 188152
rect 41146 186670 41152 186734
rect 41216 186732 41222 186734
rect 41775 186732 41841 186735
rect 41216 186730 41841 186732
rect 41216 186674 41780 186730
rect 41836 186674 41841 186730
rect 41216 186672 41841 186674
rect 41216 186670 41222 186672
rect 41775 186669 41841 186672
rect 140802 186436 140862 186924
rect 146127 186436 146193 186439
rect 140802 186434 146193 186436
rect 140802 186378 146132 186434
rect 146188 186378 146193 186434
rect 140802 186376 146193 186378
rect 146127 186373 146193 186376
rect 40954 185782 40960 185846
rect 41024 185844 41030 185846
rect 41775 185844 41841 185847
rect 41024 185842 41841 185844
rect 41024 185786 41780 185842
rect 41836 185786 41841 185842
rect 41024 185784 41841 185786
rect 41024 185782 41030 185784
rect 41775 185781 41841 185784
rect 140802 185252 140862 185740
rect 146415 185252 146481 185255
rect 140802 185250 146481 185252
rect 140802 185194 146420 185250
rect 146476 185194 146481 185250
rect 140802 185192 146481 185194
rect 146415 185189 146481 185192
rect 144015 184512 144081 184515
rect 140832 184510 144081 184512
rect 140832 184454 144020 184510
rect 144076 184454 144081 184510
rect 140832 184452 144081 184454
rect 144015 184449 144081 184452
rect 40570 184154 40576 184218
rect 40640 184216 40646 184218
rect 41775 184216 41841 184219
rect 40640 184214 41841 184216
rect 40640 184158 41780 184214
rect 41836 184158 41841 184214
rect 40640 184156 41841 184158
rect 40640 184154 40646 184156
rect 41775 184153 41841 184156
rect 40762 183562 40768 183626
rect 40832 183624 40838 183626
rect 41775 183624 41841 183627
rect 40832 183622 41841 183624
rect 40832 183566 41780 183622
rect 41836 183566 41841 183622
rect 40832 183564 41841 183566
rect 40832 183562 40838 183564
rect 41775 183561 41841 183564
rect 144207 183328 144273 183331
rect 140832 183326 144273 183328
rect 140832 183270 144212 183326
rect 144268 183270 144273 183326
rect 140832 183268 144273 183270
rect 144207 183265 144273 183268
rect 40378 182822 40384 182886
rect 40448 182884 40454 182886
rect 41775 182884 41841 182887
rect 40448 182882 41841 182884
rect 40448 182826 41780 182882
rect 41836 182826 41841 182882
rect 40448 182824 41841 182826
rect 40448 182822 40454 182824
rect 41775 182821 41841 182824
rect 140802 181848 140862 182188
rect 144015 181848 144081 181851
rect 140802 181846 144081 181848
rect 140802 181790 144020 181846
rect 144076 181790 144081 181846
rect 140802 181788 144081 181790
rect 144015 181785 144081 181788
rect 140802 180516 140862 180994
rect 144111 180516 144177 180519
rect 140802 180514 144177 180516
rect 140802 180458 144116 180514
rect 144172 180458 144177 180514
rect 140802 180456 144177 180458
rect 144111 180453 144177 180456
rect 144879 179776 144945 179779
rect 140832 179774 144945 179776
rect 140832 179718 144884 179774
rect 144940 179718 144945 179774
rect 140832 179716 144945 179718
rect 144879 179713 144945 179716
rect 674754 179631 674814 179894
rect 674703 179626 674814 179631
rect 674703 179570 674708 179626
rect 674764 179570 674814 179626
rect 674703 179568 674814 179570
rect 674703 179565 674769 179568
rect 674415 179332 674481 179335
rect 674415 179330 674784 179332
rect 674415 179274 674420 179330
rect 674476 179274 674784 179330
rect 674415 179272 674784 179274
rect 674415 179269 674481 179272
rect 674415 178814 674481 178817
rect 674415 178812 674784 178814
rect 674415 178756 674420 178812
rect 674476 178756 674784 178812
rect 674415 178754 674784 178756
rect 674415 178751 674481 178754
rect 144015 178592 144081 178595
rect 140832 178590 144081 178592
rect 140832 178534 144020 178590
rect 144076 178534 144081 178590
rect 140832 178532 144081 178534
rect 144015 178529 144081 178532
rect 677242 178382 677248 178446
rect 677312 178382 677318 178446
rect 677250 178266 677310 178382
rect 677250 177410 677310 177674
rect 676858 177346 676864 177410
rect 676928 177346 676934 177410
rect 677242 177346 677248 177410
rect 677312 177346 677318 177410
rect 140802 176816 140862 177304
rect 676866 177186 676926 177346
rect 676866 177156 677472 177186
rect 676896 177126 677502 177156
rect 677442 176966 677502 177126
rect 677434 176902 677440 176966
rect 677504 176902 677510 176966
rect 144015 176816 144081 176819
rect 140802 176814 144081 176816
rect 140802 176758 144020 176814
rect 144076 176758 144081 176814
rect 140802 176756 144081 176758
rect 144015 176753 144081 176756
rect 677058 176374 677118 176638
rect 677050 176310 677056 176374
rect 677120 176310 677126 176374
rect 145263 176076 145329 176079
rect 140832 176074 145329 176076
rect 140832 176018 145268 176074
rect 145324 176018 145329 176074
rect 140832 176016 145329 176018
rect 145263 176013 145329 176016
rect 674031 176076 674097 176079
rect 674031 176074 674784 176076
rect 674031 176018 674036 176074
rect 674092 176018 674784 176074
rect 674031 176016 674784 176018
rect 674031 176013 674097 176016
rect 676866 175191 676926 175528
rect 676866 175186 676977 175191
rect 676866 175130 676916 175186
rect 676972 175130 676977 175186
rect 676866 175128 676977 175130
rect 676911 175125 676977 175128
rect 140802 174448 140862 174982
rect 675522 174747 675582 175010
rect 675522 174742 675633 174747
rect 675522 174686 675572 174742
rect 675628 174686 675633 174742
rect 675522 174684 675633 174686
rect 675567 174681 675633 174684
rect 144111 174448 144177 174451
rect 140802 174446 144177 174448
rect 140802 174390 144116 174446
rect 144172 174390 144177 174446
rect 140802 174388 144177 174390
rect 144111 174385 144177 174388
rect 674754 174303 674814 174418
rect 674754 174298 674865 174303
rect 674754 174242 674804 174298
rect 674860 174242 674865 174298
rect 674754 174240 674865 174242
rect 674799 174237 674865 174240
rect 674362 173794 674368 173858
rect 674432 173856 674438 173858
rect 674432 173796 674784 173856
rect 674432 173794 674438 173796
rect 140802 173412 140862 173752
rect 144015 173412 144081 173415
rect 140802 173410 144081 173412
rect 140802 173354 144020 173410
rect 144076 173354 144081 173410
rect 140802 173352 144081 173354
rect 144015 173349 144081 173352
rect 676866 173119 676926 173382
rect 676815 173114 676926 173119
rect 676815 173058 676820 173114
rect 676876 173058 676926 173114
rect 676815 173056 676926 173058
rect 676815 173053 676881 173056
rect 675714 172675 675774 172790
rect 675714 172670 675825 172675
rect 675714 172614 675764 172670
rect 675820 172614 675825 172670
rect 675714 172612 675825 172614
rect 675759 172609 675825 172612
rect 140802 172080 140862 172562
rect 675138 172083 675198 172198
rect 145167 172080 145233 172083
rect 140802 172078 145233 172080
rect 140802 172022 145172 172078
rect 145228 172022 145233 172078
rect 140802 172020 145233 172022
rect 145167 172017 145233 172020
rect 675087 172078 675198 172083
rect 675087 172022 675092 172078
rect 675148 172022 675198 172078
rect 675087 172020 675198 172022
rect 675087 172017 675153 172020
rect 674946 171491 675006 171754
rect 674946 171486 675057 171491
rect 674946 171430 674996 171486
rect 675052 171430 675057 171486
rect 674946 171428 675057 171430
rect 674991 171425 675057 171428
rect 144015 171340 144081 171343
rect 140832 171338 144081 171340
rect 140832 171282 144020 171338
rect 144076 171282 144081 171338
rect 140832 171280 144081 171282
rect 144015 171277 144081 171280
rect 674554 170834 674560 170898
rect 674624 170896 674630 170898
rect 674754 170896 674814 171162
rect 674624 170836 674814 170896
rect 674624 170834 674630 170836
rect 673978 170538 673984 170602
rect 674048 170600 674054 170602
rect 674048 170540 674784 170600
rect 674048 170538 674054 170540
rect 144975 170156 145041 170159
rect 140832 170154 145041 170156
rect 140832 170098 144980 170154
rect 145036 170098 145041 170154
rect 140832 170096 145041 170098
rect 144975 170093 145041 170096
rect 674946 169863 675006 170126
rect 674895 169858 675006 169863
rect 674895 169802 674900 169858
rect 674956 169802 675006 169858
rect 674895 169800 675006 169802
rect 674895 169797 674961 169800
rect 674319 169564 674385 169567
rect 674319 169562 674784 169564
rect 674319 169506 674324 169562
rect 674380 169506 674784 169562
rect 674319 169504 674784 169506
rect 674319 169501 674385 169504
rect 140802 168380 140862 168868
rect 674511 168824 674577 168827
rect 674754 168824 674814 168942
rect 674511 168822 674814 168824
rect 674511 168766 674516 168822
rect 674572 168766 674814 168822
rect 674511 168764 674814 168766
rect 674511 168761 674577 168764
rect 145071 168380 145137 168383
rect 140802 168378 145137 168380
rect 140802 168322 145076 168378
rect 145132 168322 145137 168378
rect 140802 168320 145137 168322
rect 145071 168317 145137 168320
rect 674607 168232 674673 168235
rect 674754 168232 674814 168498
rect 674607 168230 674814 168232
rect 674607 168174 674612 168230
rect 674668 168174 674814 168230
rect 674607 168172 674814 168174
rect 674607 168169 674673 168172
rect 674754 167643 674814 167906
rect 144015 167640 144081 167643
rect 140832 167638 144081 167640
rect 140832 167582 144020 167638
rect 144076 167582 144081 167638
rect 140832 167580 144081 167582
rect 144015 167577 144081 167580
rect 674703 167638 674814 167643
rect 674703 167582 674708 167638
rect 674764 167582 674814 167638
rect 674703 167580 674814 167582
rect 674703 167577 674769 167580
rect 674415 167344 674481 167347
rect 674415 167342 674784 167344
rect 674415 167286 674420 167342
rect 674476 167286 674784 167342
rect 674415 167284 674784 167286
rect 674415 167281 674481 167284
rect 647919 167048 647985 167051
rect 640194 167046 647985 167048
rect 640194 166990 647924 167046
rect 647980 166990 647985 167046
rect 640194 166988 647985 166990
rect 640194 166870 640254 166988
rect 647919 166985 647985 166988
rect 144687 166604 144753 166607
rect 140832 166602 144753 166604
rect 140832 166546 144692 166602
rect 144748 166546 144753 166602
rect 140832 166544 144753 166546
rect 144687 166541 144753 166544
rect 647055 166308 647121 166311
rect 640416 166306 647121 166308
rect 640416 166250 647060 166306
rect 647116 166250 647121 166306
rect 640416 166248 647121 166250
rect 647055 166245 647121 166248
rect 647823 166012 647889 166015
rect 640386 166010 647889 166012
rect 640386 165954 647828 166010
rect 647884 165954 647889 166010
rect 640386 165952 647889 165954
rect 640386 165686 640446 165952
rect 647823 165949 647889 165952
rect 140802 164828 140862 165316
rect 144879 164828 144945 164831
rect 140802 164826 144945 164828
rect 140802 164770 144884 164826
rect 144940 164770 144945 164826
rect 140802 164768 144945 164770
rect 144879 164765 144945 164768
rect 140802 163644 140862 164130
rect 144207 163644 144273 163647
rect 140802 163642 144273 163644
rect 140802 163586 144212 163642
rect 144268 163586 144273 163642
rect 140802 163584 144273 163586
rect 144207 163581 144273 163584
rect 144687 162904 144753 162907
rect 140832 162902 144753 162904
rect 140832 162846 144692 162902
rect 144748 162846 144753 162902
rect 140832 162844 144753 162846
rect 144687 162841 144753 162844
rect 140802 161424 140862 161682
rect 210159 161572 210225 161575
rect 211066 161572 211072 161574
rect 210159 161570 211072 161572
rect 210159 161514 210164 161570
rect 210220 161514 211072 161570
rect 210159 161512 211072 161514
rect 210159 161509 210225 161512
rect 211066 161510 211072 161512
rect 211136 161510 211142 161574
rect 675706 161510 675712 161574
rect 675776 161572 675782 161574
rect 676911 161572 676977 161575
rect 675776 161570 676977 161572
rect 675776 161514 676916 161570
rect 676972 161514 676977 161570
rect 675776 161512 676977 161514
rect 675776 161510 675782 161512
rect 676911 161509 676977 161512
rect 144783 161424 144849 161427
rect 140802 161422 144849 161424
rect 140802 161366 144788 161422
rect 144844 161366 144849 161422
rect 140802 161364 144849 161366
rect 144783 161361 144849 161364
rect 676666 161362 676672 161426
rect 676736 161424 676742 161426
rect 676815 161424 676881 161427
rect 676736 161422 676881 161424
rect 676736 161366 676820 161422
rect 676876 161366 676881 161422
rect 676736 161364 676881 161366
rect 676736 161362 676742 161364
rect 676815 161361 676881 161364
rect 645711 161276 645777 161279
rect 645903 161276 645969 161279
rect 645711 161274 645969 161276
rect 645711 161218 645716 161274
rect 645772 161218 645908 161274
rect 645964 161218 645969 161274
rect 645711 161216 645969 161218
rect 645711 161213 645777 161216
rect 645903 161213 645969 161216
rect 140802 159944 140862 160432
rect 144303 159944 144369 159947
rect 140802 159942 144369 159944
rect 140802 159886 144308 159942
rect 144364 159886 144369 159942
rect 140802 159884 144369 159886
rect 144303 159881 144369 159884
rect 144687 159352 144753 159355
rect 140832 159350 144753 159352
rect 140832 159294 144692 159350
rect 144748 159294 144753 159350
rect 140832 159292 144753 159294
rect 144687 159289 144753 159292
rect 210159 158464 210225 158467
rect 210490 158464 210496 158466
rect 210159 158462 210496 158464
rect 210159 158406 210164 158462
rect 210220 158406 210496 158462
rect 210159 158404 210496 158406
rect 210159 158401 210225 158404
rect 210490 158402 210496 158404
rect 210560 158402 210566 158466
rect 140802 157576 140862 158138
rect 144015 157576 144081 157579
rect 140802 157574 144081 157576
rect 140802 157518 144020 157574
rect 144076 157518 144081 157574
rect 140802 157516 144081 157518
rect 144015 157513 144081 157516
rect 140802 156392 140862 156880
rect 144687 156392 144753 156395
rect 140802 156390 144753 156392
rect 140802 156334 144692 156390
rect 144748 156334 144753 156390
rect 140802 156332 144753 156334
rect 144687 156329 144753 156332
rect 140802 155652 140862 155696
rect 146895 155652 146961 155655
rect 140802 155650 146961 155652
rect 140802 155594 146900 155650
rect 146956 155594 146961 155650
rect 140802 155592 146961 155594
rect 146895 155589 146961 155592
rect 675279 155210 675345 155211
rect 675279 155208 675328 155210
rect 675236 155206 675328 155208
rect 675236 155150 675284 155206
rect 675236 155148 675328 155150
rect 675279 155146 675328 155148
rect 675392 155146 675398 155210
rect 675279 155145 675345 155146
rect 144495 154468 144561 154471
rect 675471 154470 675537 154471
rect 675471 154468 675520 154470
rect 140832 154466 144561 154468
rect 140832 154410 144500 154466
rect 144556 154410 144561 154466
rect 140832 154408 144561 154410
rect 675428 154466 675520 154468
rect 675428 154410 675476 154466
rect 675428 154408 675520 154410
rect 144495 154405 144561 154408
rect 675471 154406 675520 154408
rect 675584 154406 675590 154470
rect 675471 154405 675537 154406
rect 674362 153370 674368 153434
rect 674432 153432 674438 153434
rect 675471 153432 675537 153435
rect 674432 153430 675537 153432
rect 674432 153374 675476 153430
rect 675532 153374 675537 153430
rect 674432 153372 675537 153374
rect 674432 153370 674438 153372
rect 675471 153369 675537 153372
rect 140802 152988 140862 153250
rect 146799 152988 146865 152991
rect 140802 152986 146865 152988
rect 140802 152930 146804 152986
rect 146860 152930 146865 152986
rect 140802 152928 146865 152930
rect 146799 152925 146865 152928
rect 140802 151656 140862 152144
rect 673978 151890 673984 151954
rect 674048 151952 674054 151954
rect 675471 151952 675537 151955
rect 674048 151950 675537 151952
rect 674048 151894 675476 151950
rect 675532 151894 675537 151950
rect 674048 151892 675537 151894
rect 674048 151890 674054 151892
rect 675471 151889 675537 151892
rect 144495 151656 144561 151659
rect 140802 151654 144561 151656
rect 140802 151598 144500 151654
rect 144556 151598 144561 151654
rect 140802 151596 144561 151598
rect 144495 151593 144561 151596
rect 146799 150916 146865 150919
rect 140832 150914 146865 150916
rect 140832 150858 146804 150914
rect 146860 150858 146865 150914
rect 140832 150856 146865 150858
rect 146799 150853 146865 150856
rect 674554 150262 674560 150326
rect 674624 150324 674630 150326
rect 675471 150324 675537 150327
rect 674624 150322 675537 150324
rect 674624 150266 675476 150322
rect 675532 150266 675537 150322
rect 674624 150264 675537 150266
rect 674624 150262 674630 150264
rect 675471 150261 675537 150264
rect 144495 149732 144561 149735
rect 140832 149730 144561 149732
rect 140832 149674 144500 149730
rect 144556 149674 144561 149730
rect 140832 149672 144561 149674
rect 144495 149669 144561 149672
rect 675759 148550 675825 148551
rect 675706 148486 675712 148550
rect 675776 148548 675825 148550
rect 675776 148546 675868 148548
rect 675820 148490 675868 148546
rect 675776 148488 675868 148490
rect 675776 148486 675825 148488
rect 675759 148485 675825 148486
rect 140802 147956 140862 148444
rect 146799 147956 146865 147959
rect 140802 147954 146865 147956
rect 140802 147898 146804 147954
rect 146860 147898 146865 147954
rect 140802 147896 146865 147898
rect 146799 147893 146865 147896
rect 140802 146920 140862 147260
rect 144111 146920 144177 146923
rect 140802 146918 144177 146920
rect 140802 146862 144116 146918
rect 144172 146862 144177 146918
rect 140802 146860 144177 146862
rect 144111 146857 144177 146860
rect 675759 146624 675825 146627
rect 676666 146624 676672 146626
rect 675759 146622 676672 146624
rect 675759 146566 675764 146622
rect 675820 146566 676672 146622
rect 675759 146564 676672 146566
rect 675759 146561 675825 146564
rect 676666 146562 676672 146564
rect 676736 146562 676742 146626
rect 144015 146032 144081 146035
rect 140832 146030 144081 146032
rect 140832 145974 144020 146030
rect 144076 145974 144081 146030
rect 140832 145972 144081 145974
rect 144015 145969 144081 145972
rect 140802 144256 140862 144790
rect 146703 144256 146769 144259
rect 140802 144254 146769 144256
rect 140802 144198 146708 144254
rect 146764 144198 146769 144254
rect 140802 144196 146769 144198
rect 146703 144193 146769 144196
rect 140802 143220 140862 143708
rect 144015 143220 144081 143223
rect 140802 143218 144081 143220
rect 140802 143162 144020 143218
rect 144076 143162 144081 143218
rect 140802 143160 144081 143162
rect 144015 143157 144081 143160
rect 144015 142480 144081 142483
rect 140832 142478 144081 142480
rect 140832 142422 144020 142478
rect 144076 142422 144081 142478
rect 140832 142420 144081 142422
rect 144015 142417 144081 142420
rect 210159 141592 210225 141595
rect 210874 141592 210880 141594
rect 210159 141590 210880 141592
rect 210159 141534 210164 141590
rect 210220 141534 210880 141590
rect 210159 141532 210880 141534
rect 210159 141529 210225 141532
rect 210874 141530 210880 141532
rect 210944 141530 210950 141594
rect 210490 141382 210496 141446
rect 210560 141444 210566 141446
rect 210560 141384 210942 141444
rect 210560 141382 210566 141384
rect 210882 141298 210942 141384
rect 140832 141236 144126 141296
rect 144066 141003 144126 141236
rect 210874 141234 210880 141298
rect 210944 141234 210950 141298
rect 144015 140998 144126 141003
rect 144015 140942 144020 140998
rect 144076 140942 144126 140998
rect 144015 140940 144126 140942
rect 144015 140937 144081 140940
rect 140802 139520 140862 140008
rect 144303 139520 144369 139523
rect 140802 139518 144369 139520
rect 140802 139462 144308 139518
rect 144364 139462 144369 139518
rect 140802 139460 144369 139462
rect 144303 139457 144369 139460
rect 140802 138632 140862 138824
rect 144015 138632 144081 138635
rect 140802 138630 144081 138632
rect 140802 138574 144020 138630
rect 144076 138574 144081 138630
rect 140802 138572 144081 138574
rect 144015 138569 144081 138572
rect 210159 138484 210225 138487
rect 210159 138482 210750 138484
rect 210159 138426 210164 138482
rect 210220 138426 210750 138482
rect 210159 138424 210750 138426
rect 210159 138421 210225 138424
rect 210690 138338 210750 138424
rect 210682 138274 210688 138338
rect 210752 138274 210758 138338
rect 161103 137596 161169 137599
rect 140832 137594 161169 137596
rect 140832 137538 161108 137594
rect 161164 137538 161169 137594
rect 140832 137536 161169 137538
rect 161103 137533 161169 137536
rect 140802 136116 140862 136522
rect 146991 136116 147057 136119
rect 140802 136114 147057 136116
rect 140802 136058 146996 136114
rect 147052 136058 147057 136114
rect 140802 136056 147057 136058
rect 146991 136053 147057 136056
rect 146703 135672 146769 135675
rect 146562 135670 146769 135672
rect 146562 135614 146708 135670
rect 146764 135614 146769 135670
rect 146562 135612 146769 135614
rect 140802 134784 140862 135272
rect 146127 135228 146193 135231
rect 146562 135228 146622 135612
rect 146703 135609 146769 135612
rect 146127 135226 146622 135228
rect 146127 135170 146132 135226
rect 146188 135170 146622 135226
rect 146127 135168 146622 135170
rect 146127 135165 146193 135168
rect 144015 134784 144081 134787
rect 140802 134782 144081 134784
rect 140802 134726 144020 134782
rect 144076 134726 144081 134782
rect 140802 134724 144081 134726
rect 144015 134721 144081 134724
rect 676866 134343 676926 134680
rect 676866 134338 676977 134343
rect 676866 134282 676916 134338
rect 676972 134282 676977 134338
rect 676866 134280 676977 134282
rect 676911 134277 676977 134280
rect 144303 134044 144369 134047
rect 140832 134042 144369 134044
rect 140832 133986 144308 134042
rect 144364 133986 144369 134042
rect 140832 133984 144369 133986
rect 144303 133981 144369 133984
rect 676866 133899 676926 134162
rect 676815 133894 676926 133899
rect 676815 133838 676820 133894
rect 676876 133838 676926 133894
rect 676815 133836 676926 133838
rect 676815 133833 676881 133836
rect 674415 133600 674481 133603
rect 674415 133598 674784 133600
rect 674415 133542 674420 133598
rect 674476 133542 674784 133598
rect 674415 133540 674784 133542
rect 674415 133537 674481 133540
rect 677242 133390 677248 133454
rect 677312 133390 677318 133454
rect 677250 132978 677310 133390
rect 144015 132860 144081 132863
rect 140832 132858 144081 132860
rect 140832 132802 144020 132858
rect 144076 132802 144081 132858
rect 140832 132800 144081 132802
rect 144015 132797 144081 132800
rect 674415 132564 674481 132567
rect 674415 132562 674784 132564
rect 674415 132506 674420 132562
rect 674476 132506 674784 132562
rect 674415 132504 674784 132506
rect 674415 132501 674481 132504
rect 677434 132206 677440 132270
rect 677504 132206 677510 132270
rect 677442 131942 677502 132206
rect 677050 131762 677056 131826
rect 677120 131762 677126 131826
rect 140802 131084 140862 131572
rect 677058 131350 677118 131762
rect 144111 131084 144177 131087
rect 140802 131082 144177 131084
rect 140802 131026 144116 131082
rect 144172 131026 144177 131082
rect 140802 131024 144177 131026
rect 144111 131021 144177 131024
rect 674511 130640 674577 130643
rect 674754 130640 674814 130906
rect 674511 130638 674814 130640
rect 674511 130582 674516 130638
rect 674572 130582 674814 130638
rect 674511 130580 674814 130582
rect 674511 130577 674577 130580
rect 140802 130196 140862 130388
rect 144015 130196 144081 130199
rect 140802 130194 144081 130196
rect 140802 130138 144020 130194
rect 144076 130138 144081 130194
rect 140802 130136 144081 130138
rect 144015 130133 144081 130136
rect 677058 130051 677118 130314
rect 677058 130046 677169 130051
rect 677058 129990 677108 130046
rect 677164 129990 677169 130046
rect 677058 129988 677169 129990
rect 677103 129985 677169 129988
rect 675138 129607 675198 129722
rect 675138 129602 675249 129607
rect 675138 129546 675188 129602
rect 675244 129546 675249 129602
rect 675138 129544 675249 129546
rect 675183 129541 675249 129544
rect 144015 129308 144081 129311
rect 140832 129306 144081 129308
rect 140832 129250 144020 129306
rect 144076 129250 144081 129306
rect 140832 129248 144081 129250
rect 144015 129245 144081 129248
rect 210159 129160 210225 129163
rect 210874 129160 210880 129162
rect 210159 129158 210880 129160
rect 210159 129102 210164 129158
rect 210220 129102 210880 129158
rect 210159 129100 210880 129102
rect 210159 129097 210225 129100
rect 210874 129098 210880 129100
rect 210944 129098 210950 129162
rect 675138 129015 675198 129278
rect 675087 129010 675198 129015
rect 675087 128954 675092 129010
rect 675148 128954 675198 129010
rect 675087 128952 675198 128954
rect 675087 128949 675153 128952
rect 673978 128654 673984 128718
rect 674048 128716 674054 128718
rect 674048 128656 674784 128716
rect 674048 128654 674054 128656
rect 140802 127532 140862 128090
rect 677058 127831 677118 128094
rect 677007 127826 677118 127831
rect 677007 127770 677012 127826
rect 677068 127770 677118 127826
rect 677007 127768 677118 127770
rect 677007 127765 677073 127768
rect 146703 127532 146769 127535
rect 140802 127530 146769 127532
rect 140802 127474 146708 127530
rect 146764 127474 146769 127530
rect 140802 127472 146769 127474
rect 146703 127469 146769 127472
rect 674946 127387 675006 127650
rect 674895 127382 675006 127387
rect 674895 127326 674900 127382
rect 674956 127326 675006 127382
rect 674895 127324 675006 127326
rect 674895 127321 674961 127324
rect 674319 127088 674385 127091
rect 674319 127086 674784 127088
rect 674319 127030 674324 127086
rect 674380 127030 674784 127086
rect 674319 127028 674784 127030
rect 674319 127025 674385 127028
rect 147087 126940 147153 126943
rect 140832 126938 147153 126940
rect 140832 126882 147092 126938
rect 147148 126882 147153 126938
rect 140832 126880 147153 126882
rect 147087 126877 147153 126880
rect 144495 126792 144561 126795
rect 146127 126792 146193 126795
rect 144495 126790 146193 126792
rect 144495 126734 144500 126790
rect 144556 126734 146132 126790
rect 146188 126734 146193 126790
rect 144495 126732 146193 126734
rect 144495 126729 144561 126732
rect 146127 126729 146193 126732
rect 674754 126351 674814 126466
rect 674754 126346 674865 126351
rect 674754 126290 674804 126346
rect 674860 126290 674865 126346
rect 674754 126288 674865 126290
rect 674799 126285 674865 126288
rect 210159 126200 210225 126203
rect 210490 126200 210496 126202
rect 210159 126198 210496 126200
rect 210159 126142 210164 126198
rect 210220 126142 210496 126198
rect 210159 126140 210496 126142
rect 210159 126137 210225 126140
rect 210490 126138 210496 126140
rect 210560 126138 210566 126202
rect 674170 125990 674176 126054
rect 674240 126052 674246 126054
rect 674240 125992 674784 126052
rect 674240 125990 674246 125992
rect 39855 125312 39921 125315
rect 39810 125310 39921 125312
rect 39810 125254 39860 125310
rect 39916 125254 39921 125310
rect 39810 125249 39921 125254
rect 39810 124986 39870 125249
rect 140802 125164 140862 125642
rect 673935 125460 674001 125463
rect 673935 125458 674784 125460
rect 673935 125402 673940 125458
rect 673996 125402 674784 125458
rect 673935 125400 674784 125402
rect 673935 125397 674001 125400
rect 144111 125164 144177 125167
rect 140802 125162 144177 125164
rect 140802 125106 144116 125162
rect 144172 125106 144177 125162
rect 140802 125104 144177 125106
rect 144111 125101 144177 125104
rect 674607 124720 674673 124723
rect 674754 124720 674814 124838
rect 674607 124718 674814 124720
rect 674607 124662 674612 124718
rect 674668 124662 674814 124718
rect 674607 124660 674814 124662
rect 674607 124657 674673 124660
rect 144015 124424 144081 124427
rect 140832 124422 144081 124424
rect 140832 124366 144020 124422
rect 144076 124366 144081 124422
rect 140832 124364 144081 124366
rect 144015 124361 144081 124364
rect 674946 124131 675006 124320
rect 674946 124126 675057 124131
rect 674946 124070 674996 124126
rect 675052 124070 675057 124126
rect 674946 124068 675057 124070
rect 674991 124065 675057 124068
rect 674223 123832 674289 123835
rect 674223 123830 674784 123832
rect 674223 123774 674228 123830
rect 674284 123774 674784 123830
rect 674223 123772 674784 123774
rect 674223 123769 674289 123772
rect 140802 122796 140862 123136
rect 676866 122947 676926 123210
rect 676866 122942 676977 122947
rect 676866 122886 676916 122942
rect 676972 122886 676977 122942
rect 676866 122884 676977 122886
rect 676911 122881 676977 122884
rect 144111 122796 144177 122799
rect 140802 122794 144177 122796
rect 140802 122738 144116 122794
rect 144172 122738 144177 122794
rect 140802 122736 144177 122738
rect 144111 122733 144177 122736
rect 676866 122355 676926 122692
rect 676815 122350 676926 122355
rect 676815 122294 676820 122350
rect 676876 122294 676926 122350
rect 676815 122292 676926 122294
rect 676815 122289 676881 122292
rect 140802 121612 140862 121952
rect 674754 121911 674814 122174
rect 674703 121906 674814 121911
rect 674703 121850 674708 121906
rect 674764 121850 674814 121906
rect 674703 121848 674814 121850
rect 674703 121845 674769 121848
rect 144015 121612 144081 121615
rect 140802 121610 144081 121612
rect 140802 121554 144020 121610
rect 144076 121554 144081 121610
rect 140802 121552 144081 121554
rect 144015 121549 144081 121552
rect 640386 121464 640446 121730
rect 645711 121464 645777 121467
rect 640386 121462 645777 121464
rect 640386 121406 645716 121462
rect 645772 121406 645777 121462
rect 640386 121404 645777 121406
rect 645711 121401 645777 121404
rect 210159 121168 210225 121171
rect 211066 121168 211072 121170
rect 210159 121166 211072 121168
rect 210159 121110 210164 121166
rect 210220 121110 211072 121166
rect 210159 121108 211072 121110
rect 210159 121105 210225 121108
rect 211066 121106 211072 121108
rect 211136 121106 211142 121170
rect 645423 121168 645489 121171
rect 640416 121166 645489 121168
rect 640416 121110 645428 121166
rect 645484 121110 645489 121166
rect 640416 121108 645489 121110
rect 645423 121105 645489 121108
rect 144111 120872 144177 120875
rect 645711 120872 645777 120875
rect 140832 120870 144177 120872
rect 140832 120814 144116 120870
rect 144172 120814 144177 120870
rect 140832 120812 144177 120814
rect 144111 120809 144177 120812
rect 640386 120870 645777 120872
rect 640386 120814 645716 120870
rect 645772 120814 645777 120870
rect 640386 120812 645777 120814
rect 640386 120546 640446 120812
rect 645711 120809 645777 120812
rect 647727 120428 647793 120431
rect 640386 120426 647793 120428
rect 640386 120370 647732 120426
rect 647788 120370 647793 120426
rect 640386 120368 647793 120370
rect 640386 120028 640446 120368
rect 647727 120365 647793 120368
rect 140802 119096 140862 119630
rect 146895 119096 146961 119099
rect 140802 119094 146961 119096
rect 140802 119038 146900 119094
rect 146956 119038 146961 119094
rect 140802 119036 146961 119038
rect 146895 119033 146961 119036
rect 141039 118652 141105 118655
rect 140610 118650 141105 118652
rect 140610 118594 141044 118650
rect 141100 118594 141105 118650
rect 140610 118592 141105 118594
rect 140610 118474 140670 118592
rect 141039 118589 141105 118592
rect 141039 118356 141105 118359
rect 144015 118356 144081 118359
rect 141039 118354 144081 118356
rect 141039 118298 141044 118354
rect 141100 118298 144020 118354
rect 144076 118298 144081 118354
rect 141039 118296 144081 118298
rect 141039 118293 141105 118296
rect 144015 118293 144081 118296
rect 210490 117998 210496 118062
rect 210560 118060 210566 118062
rect 210874 118060 210880 118062
rect 210560 118000 210880 118060
rect 210560 117998 210566 118000
rect 210874 117998 210880 118000
rect 210944 117998 210950 118062
rect 676666 117998 676672 118062
rect 676736 118060 676742 118062
rect 677007 118060 677073 118063
rect 676736 118058 677073 118060
rect 676736 118002 677012 118058
rect 677068 118002 677073 118058
rect 676736 118000 677073 118002
rect 676736 117998 676742 118000
rect 677007 117997 677073 118000
rect 675898 117850 675904 117914
rect 675968 117912 675974 117914
rect 677103 117912 677169 117915
rect 675968 117910 677169 117912
rect 675968 117854 677108 117910
rect 677164 117854 677169 117910
rect 675968 117852 677169 117854
rect 675968 117850 675974 117852
rect 677103 117849 677169 117852
rect 140802 116728 140862 117210
rect 146895 116728 146961 116731
rect 140802 116726 146961 116728
rect 140802 116670 146900 116726
rect 146956 116670 146961 116726
rect 140802 116668 146961 116670
rect 146895 116665 146961 116668
rect 146895 115988 146961 115991
rect 140832 115986 146961 115988
rect 140832 115930 146900 115986
rect 146956 115930 146961 115986
rect 140832 115928 146961 115930
rect 146895 115925 146961 115928
rect 140802 114212 140862 114762
rect 144015 114212 144081 114215
rect 140802 114210 144081 114212
rect 140802 114154 144020 114210
rect 144076 114154 144081 114210
rect 140802 114152 144081 114154
rect 144015 114149 144081 114152
rect 210159 113768 210225 113771
rect 211066 113768 211072 113770
rect 210159 113766 211072 113768
rect 210159 113710 210164 113766
rect 210220 113710 211072 113766
rect 210159 113708 211072 113710
rect 210159 113705 210225 113708
rect 211066 113706 211072 113708
rect 211136 113706 211142 113770
rect 140802 113176 140862 113664
rect 144111 113176 144177 113179
rect 140802 113174 144177 113176
rect 140802 113118 144116 113174
rect 144172 113118 144177 113174
rect 140802 113116 144177 113118
rect 144111 113113 144177 113116
rect 144015 112436 144081 112439
rect 140832 112434 144081 112436
rect 140832 112378 144020 112434
rect 144076 112378 144081 112434
rect 140832 112376 144081 112378
rect 144015 112373 144081 112376
rect 210682 112226 210688 112290
rect 210752 112288 210758 112290
rect 211066 112288 211072 112290
rect 210752 112228 211072 112288
rect 210752 112226 210758 112228
rect 211066 112226 211072 112228
rect 211136 112226 211142 112290
rect 144111 111252 144177 111255
rect 140832 111250 144177 111252
rect 140832 111194 144116 111250
rect 144172 111194 144177 111250
rect 140832 111192 144177 111194
rect 144111 111189 144177 111192
rect 675375 110070 675441 110071
rect 675322 110068 675328 110070
rect 675284 110008 675328 110068
rect 675392 110066 675441 110070
rect 675436 110010 675441 110066
rect 675322 110006 675328 110008
rect 675392 110006 675441 110010
rect 675375 110005 675441 110006
rect 140802 109772 140862 109964
rect 144015 109772 144081 109775
rect 140802 109770 144081 109772
rect 140802 109714 144020 109770
rect 144076 109714 144081 109770
rect 140802 109712 144081 109714
rect 144015 109709 144081 109712
rect 675471 109330 675537 109331
rect 675471 109326 675520 109330
rect 675584 109328 675590 109330
rect 675471 109270 675476 109326
rect 675471 109266 675520 109270
rect 675584 109268 675628 109328
rect 675584 109266 675590 109268
rect 675471 109265 675537 109266
rect 140802 108292 140862 108778
rect 144687 108292 144753 108295
rect 140802 108290 144753 108292
rect 140802 108234 144692 108290
rect 144748 108234 144753 108290
rect 140802 108232 144753 108234
rect 144687 108229 144753 108232
rect 673978 108082 673984 108146
rect 674048 108144 674054 108146
rect 675375 108144 675441 108147
rect 674048 108142 675441 108144
rect 674048 108086 675380 108142
rect 675436 108086 675441 108142
rect 674048 108084 675441 108086
rect 674048 108082 674054 108084
rect 675375 108081 675441 108084
rect 144015 107552 144081 107555
rect 140832 107550 144081 107552
rect 140832 107494 144020 107550
rect 144076 107494 144081 107550
rect 140832 107492 144081 107494
rect 144015 107489 144081 107492
rect 143919 106960 143985 106963
rect 143919 106958 144318 106960
rect 143919 106902 143924 106958
rect 143980 106902 144318 106958
rect 143919 106900 144318 106902
rect 143919 106897 143985 106900
rect 144258 106664 144318 106900
rect 146223 106812 146289 106815
rect 146178 106810 146289 106812
rect 146178 106754 146228 106810
rect 146284 106754 146289 106810
rect 146178 106749 146289 106754
rect 144591 106664 144657 106667
rect 144258 106662 144657 106664
rect 144258 106606 144596 106662
rect 144652 106606 144657 106662
rect 144258 106604 144657 106606
rect 144591 106601 144657 106604
rect 146178 106519 146238 106749
rect 146178 106514 146289 106519
rect 668175 106516 668241 106519
rect 146178 106458 146228 106514
rect 146284 106458 146289 106514
rect 146178 106456 146289 106458
rect 146223 106453 146289 106456
rect 665346 106514 668241 106516
rect 665346 106458 668180 106514
rect 668236 106458 668241 106514
rect 665346 106456 668241 106458
rect 140802 105924 140862 106412
rect 665346 106082 665406 106456
rect 668175 106453 668241 106456
rect 144015 105924 144081 105927
rect 140802 105922 144081 105924
rect 140802 105866 144020 105922
rect 144076 105866 144081 105922
rect 140802 105864 144081 105866
rect 144015 105861 144081 105864
rect 140802 104740 140862 105228
rect 665154 105187 665214 105361
rect 665154 105182 665265 105187
rect 665154 105126 665204 105182
rect 665260 105126 665265 105182
rect 665154 105124 665265 105126
rect 665199 105121 665265 105124
rect 674170 105122 674176 105186
rect 674240 105184 674246 105186
rect 675375 105184 675441 105187
rect 674240 105182 675441 105184
rect 674240 105126 675380 105182
rect 675436 105126 675441 105182
rect 674240 105124 675441 105126
rect 674240 105122 674246 105124
rect 675375 105121 675441 105124
rect 144111 104740 144177 104743
rect 140802 104738 144177 104740
rect 140802 104682 144116 104738
rect 144172 104682 144177 104738
rect 140802 104680 144177 104682
rect 144111 104677 144177 104680
rect 665154 104595 665214 104996
rect 665154 104590 665265 104595
rect 665154 104534 665204 104590
rect 665260 104534 665265 104590
rect 665154 104532 665265 104534
rect 665199 104529 665265 104532
rect 144015 104296 144081 104299
rect 645423 104296 645489 104299
rect 140610 104294 144081 104296
rect 140610 104238 144020 104294
rect 144076 104238 144081 104294
rect 140610 104236 144081 104238
rect 640416 104294 645489 104296
rect 640416 104238 645428 104294
rect 645484 104238 645489 104294
rect 640416 104236 645489 104238
rect 140610 104044 140670 104236
rect 144015 104233 144081 104236
rect 645423 104233 645489 104236
rect 675759 103260 675825 103263
rect 675898 103260 675904 103262
rect 675759 103258 675904 103260
rect 675759 103202 675764 103258
rect 675820 103202 675904 103258
rect 675759 103200 675904 103202
rect 675759 103197 675825 103200
rect 675898 103198 675904 103200
rect 675968 103198 675974 103262
rect 144111 102816 144177 102819
rect 140832 102814 144177 102816
rect 140832 102758 144116 102814
rect 144172 102758 144177 102814
rect 140832 102756 144177 102758
rect 144111 102753 144177 102756
rect 204495 102076 204561 102079
rect 204495 102074 210528 102076
rect 204495 102018 204500 102074
rect 204556 102018 210528 102074
rect 204495 102016 210528 102018
rect 204495 102013 204561 102016
rect 144015 101632 144081 101635
rect 140832 101630 144081 101632
rect 140832 101574 144020 101630
rect 144076 101574 144081 101630
rect 140832 101572 144081 101574
rect 144015 101569 144081 101572
rect 204591 101632 204657 101635
rect 204591 101630 210528 101632
rect 204591 101574 204596 101630
rect 204652 101574 210528 101630
rect 204591 101572 210528 101574
rect 204591 101569 204657 101572
rect 675759 101484 675825 101487
rect 676666 101484 676672 101486
rect 675759 101482 676672 101484
rect 675759 101426 675764 101482
rect 675820 101426 676672 101482
rect 675759 101424 676672 101426
rect 675759 101421 675825 101424
rect 676666 101422 676672 101424
rect 676736 101422 676742 101486
rect 204687 101040 204753 101043
rect 204687 101038 210528 101040
rect 204687 100982 204692 101038
rect 204748 100982 210528 101038
rect 204687 100980 210528 100982
rect 204687 100977 204753 100980
rect 204591 100448 204657 100451
rect 204591 100446 210528 100448
rect 204591 100390 204596 100446
rect 204652 100390 210528 100446
rect 204591 100388 210528 100390
rect 204591 100385 204657 100388
rect 140802 99856 140862 100344
rect 204495 100300 204561 100303
rect 204495 100298 210558 100300
rect 204495 100242 204500 100298
rect 204556 100242 210558 100298
rect 204495 100240 210558 100242
rect 204495 100237 204561 100240
rect 210498 99900 210558 100240
rect 144207 99856 144273 99859
rect 140802 99854 144273 99856
rect 140802 99798 144212 99854
rect 144268 99798 144273 99854
rect 140802 99796 144273 99798
rect 144207 99793 144273 99796
rect 204687 99412 204753 99415
rect 204687 99410 210528 99412
rect 204687 99354 204692 99410
rect 204748 99354 210528 99410
rect 204687 99352 210528 99354
rect 204687 99349 204753 99352
rect 144111 99116 144177 99119
rect 140832 99114 144177 99116
rect 140832 99058 144116 99114
rect 144172 99058 144177 99114
rect 140832 99056 144177 99058
rect 144111 99053 144177 99056
rect 204783 98820 204849 98823
rect 204783 98818 210528 98820
rect 204783 98762 204788 98818
rect 204844 98762 210528 98818
rect 204783 98760 210528 98762
rect 204783 98757 204849 98760
rect 204879 98672 204945 98675
rect 204879 98670 210558 98672
rect 204879 98614 204884 98670
rect 204940 98614 210558 98670
rect 204879 98612 210558 98614
rect 204879 98609 204945 98612
rect 210498 98272 210558 98612
rect 144015 98080 144081 98083
rect 140832 98078 144081 98080
rect 140832 98022 144020 98078
rect 144076 98022 144081 98078
rect 140832 98020 144081 98022
rect 144015 98017 144081 98020
rect 204495 97784 204561 97787
rect 204495 97782 210528 97784
rect 204495 97726 204500 97782
rect 204556 97726 210528 97782
rect 204495 97724 210528 97726
rect 204495 97721 204561 97724
rect 204495 97192 204561 97195
rect 204495 97190 210528 97192
rect 204495 97134 204500 97190
rect 204556 97134 210528 97190
rect 204495 97132 210528 97134
rect 204495 97129 204561 97132
rect 204591 97044 204657 97047
rect 204591 97042 210558 97044
rect 204591 96986 204596 97042
rect 204652 96986 210558 97042
rect 204591 96984 210558 96986
rect 204591 96981 204657 96984
rect 140802 96304 140862 96792
rect 210498 96644 210558 96984
rect 144111 96304 144177 96307
rect 140802 96302 144177 96304
rect 140802 96246 144116 96302
rect 144172 96246 144177 96302
rect 140802 96244 144177 96246
rect 144111 96241 144177 96244
rect 204783 96156 204849 96159
rect 204783 96154 210528 96156
rect 204783 96098 204788 96154
rect 204844 96098 210528 96154
rect 204783 96096 210528 96098
rect 204783 96093 204849 96096
rect 144015 95564 144081 95567
rect 140832 95562 144081 95564
rect 140832 95506 144020 95562
rect 144076 95506 144081 95562
rect 140832 95504 144081 95506
rect 144015 95501 144081 95504
rect 204687 95564 204753 95567
rect 204687 95562 210528 95564
rect 204687 95506 204692 95562
rect 204748 95506 210528 95562
rect 204687 95504 210528 95506
rect 204687 95501 204753 95504
rect 204591 94824 204657 94827
rect 210498 94824 210558 95016
rect 204591 94822 210558 94824
rect 204591 94766 204596 94822
rect 204652 94766 210558 94822
rect 204591 94764 210558 94766
rect 204591 94761 204657 94764
rect 204495 94528 204561 94531
rect 204495 94526 210528 94528
rect 204495 94470 204500 94526
rect 204556 94470 210528 94526
rect 204495 94468 210528 94470
rect 204495 94465 204561 94468
rect 144111 94380 144177 94383
rect 140832 94378 144177 94380
rect 140832 94322 144116 94378
rect 144172 94322 144177 94378
rect 140832 94320 144177 94322
rect 144111 94317 144177 94320
rect 205263 93936 205329 93939
rect 205263 93934 210528 93936
rect 205263 93878 205268 93934
rect 205324 93878 210528 93934
rect 205263 93876 210528 93878
rect 205263 93873 205329 93876
rect 204783 93788 204849 93791
rect 204783 93786 210558 93788
rect 204783 93730 204788 93786
rect 204844 93730 210558 93786
rect 204783 93728 210558 93730
rect 204783 93725 204849 93728
rect 210498 93388 210558 93728
rect 140802 92900 140862 93092
rect 144015 92900 144081 92903
rect 140802 92898 144081 92900
rect 140802 92842 144020 92898
rect 144076 92842 144081 92898
rect 140802 92840 144081 92842
rect 144015 92837 144081 92840
rect 204687 92900 204753 92903
rect 204687 92898 210528 92900
rect 204687 92842 204692 92898
rect 204748 92842 210528 92898
rect 204687 92840 210528 92842
rect 204687 92837 204753 92840
rect 201711 92308 201777 92311
rect 201711 92306 210528 92308
rect 201711 92250 201716 92306
rect 201772 92250 210528 92306
rect 201711 92248 210528 92250
rect 201711 92245 201777 92248
rect 204495 92012 204561 92015
rect 204495 92010 210558 92012
rect 204495 91954 204500 92010
rect 204556 91954 210558 92010
rect 204495 91952 210558 91954
rect 204495 91949 204561 91952
rect 140802 91420 140862 91908
rect 210498 91760 210558 91952
rect 144207 91420 144273 91423
rect 140802 91418 144273 91420
rect 140802 91362 144212 91418
rect 144268 91362 144273 91418
rect 140802 91360 144273 91362
rect 144207 91357 144273 91360
rect 205359 91272 205425 91275
rect 205359 91270 210528 91272
rect 205359 91214 205364 91270
rect 205420 91214 210528 91270
rect 205359 91212 210528 91214
rect 205359 91209 205425 91212
rect 144111 90828 144177 90831
rect 140832 90826 144177 90828
rect 140832 90770 144116 90826
rect 144172 90770 144177 90826
rect 140832 90768 144177 90770
rect 144111 90765 144177 90768
rect 204495 90680 204561 90683
rect 204495 90678 210528 90680
rect 204495 90622 204500 90678
rect 204556 90622 210528 90678
rect 204495 90620 210528 90622
rect 204495 90617 204561 90620
rect 204591 90088 204657 90091
rect 204591 90086 210528 90088
rect 204591 90030 204596 90086
rect 204652 90030 210528 90086
rect 204591 90028 210528 90030
rect 204591 90025 204657 90028
rect 144015 89644 144081 89647
rect 140832 89642 144081 89644
rect 140832 89586 144020 89642
rect 144076 89586 144081 89642
rect 140832 89584 144081 89586
rect 144015 89581 144081 89584
rect 204687 89644 204753 89647
rect 204687 89642 210528 89644
rect 204687 89586 204692 89642
rect 204748 89586 210528 89642
rect 204687 89584 210528 89586
rect 204687 89581 204753 89584
rect 204495 89052 204561 89055
rect 647631 89052 647697 89055
rect 204495 89050 210528 89052
rect 204495 88994 204500 89050
rect 204556 88994 210528 89050
rect 204495 88992 210528 88994
rect 640416 89050 647697 89052
rect 640416 88994 647636 89050
rect 647692 88994 647697 89050
rect 640416 88992 647697 88994
rect 204495 88989 204561 88992
rect 647631 88989 647697 88992
rect 204591 88460 204657 88463
rect 204591 88458 210528 88460
rect 204591 88402 204596 88458
rect 204652 88402 210528 88458
rect 204591 88400 210528 88402
rect 204591 88397 204657 88400
rect 140802 87868 140862 88356
rect 640194 88164 640254 88430
rect 645711 88164 645777 88167
rect 640194 88162 645777 88164
rect 640194 88106 645716 88162
rect 645772 88106 645777 88162
rect 640194 88104 645777 88106
rect 645711 88101 645777 88104
rect 204687 88016 204753 88019
rect 204687 88014 210528 88016
rect 204687 87958 204692 88014
rect 204748 87958 210528 88014
rect 204687 87956 210528 87958
rect 204687 87953 204753 87956
rect 146415 87868 146481 87871
rect 140802 87866 146481 87868
rect 140802 87810 146420 87866
rect 146476 87810 146481 87866
rect 140802 87808 146481 87810
rect 146415 87805 146481 87808
rect 640386 87720 640446 87986
rect 645423 87720 645489 87723
rect 640386 87718 645489 87720
rect 640386 87662 645428 87718
rect 645484 87662 645489 87718
rect 640386 87660 645489 87662
rect 645423 87657 645489 87660
rect 204783 87424 204849 87427
rect 647343 87424 647409 87427
rect 204783 87422 210528 87424
rect 204783 87366 204788 87422
rect 204844 87366 210528 87422
rect 204783 87364 210528 87366
rect 640416 87422 647409 87424
rect 640416 87366 647348 87422
rect 647404 87366 647409 87422
rect 640416 87364 647409 87366
rect 204783 87361 204849 87364
rect 647343 87361 647409 87364
rect 144111 87128 144177 87131
rect 140832 87126 144177 87128
rect 140832 87070 144116 87126
rect 144172 87070 144177 87126
rect 140832 87068 144177 87070
rect 144111 87065 144177 87068
rect 210106 86918 210112 86982
rect 210176 86980 210182 86982
rect 210255 86980 210321 86983
rect 210176 86978 210321 86980
rect 210176 86922 210260 86978
rect 210316 86922 210321 86978
rect 210176 86920 210321 86922
rect 210176 86918 210182 86920
rect 210255 86917 210321 86920
rect 650895 86980 650961 86983
rect 650895 86978 656736 86980
rect 650895 86922 650900 86978
rect 650956 86922 656736 86978
rect 650895 86920 656736 86922
rect 650895 86917 650961 86920
rect 204879 86832 204945 86835
rect 204879 86830 210528 86832
rect 204879 86774 204884 86830
rect 204940 86774 210528 86830
rect 204879 86772 210528 86774
rect 204879 86769 204945 86772
rect 640194 86684 640254 86802
rect 645423 86684 645489 86687
rect 640194 86682 645489 86684
rect 640194 86626 645428 86682
rect 645484 86626 645489 86682
rect 640194 86624 645489 86626
rect 645423 86621 645489 86624
rect 210682 86474 210688 86538
rect 210752 86536 210758 86538
rect 210874 86536 210880 86538
rect 210752 86476 210880 86536
rect 210752 86474 210758 86476
rect 210874 86474 210880 86476
rect 210944 86474 210950 86538
rect 204495 86388 204561 86391
rect 204495 86386 210528 86388
rect 204495 86330 204500 86386
rect 204556 86330 210528 86386
rect 204495 86328 210528 86330
rect 204495 86325 204561 86328
rect 640386 86240 640446 86358
rect 647823 86240 647889 86243
rect 640386 86238 647889 86240
rect 640386 86182 647828 86238
rect 647884 86182 647889 86238
rect 640386 86180 647889 86182
rect 647823 86177 647889 86180
rect 651183 86240 651249 86243
rect 651183 86238 656736 86240
rect 651183 86182 651188 86238
rect 651244 86182 656736 86238
rect 651183 86180 656736 86182
rect 651183 86177 651249 86180
rect 144015 85944 144081 85947
rect 140832 85942 144081 85944
rect 140832 85886 144020 85942
rect 144076 85886 144081 85942
rect 140832 85884 144081 85886
rect 144015 85881 144081 85884
rect 204495 85796 204561 85799
rect 646095 85796 646161 85799
rect 204495 85794 210528 85796
rect 204495 85738 204500 85794
rect 204556 85738 210528 85794
rect 204495 85736 210528 85738
rect 640416 85794 646161 85796
rect 640416 85738 646100 85794
rect 646156 85738 646161 85794
rect 640416 85736 646161 85738
rect 204495 85733 204561 85736
rect 646095 85733 646161 85736
rect 663618 85651 663678 86210
rect 663567 85646 663678 85651
rect 663567 85590 663572 85646
rect 663628 85590 663678 85646
rect 663567 85588 663678 85590
rect 663567 85585 663633 85588
rect 647727 85500 647793 85503
rect 640386 85498 647793 85500
rect 640386 85442 647732 85498
rect 647788 85442 647793 85498
rect 640386 85440 647793 85442
rect 204591 85204 204657 85207
rect 204591 85202 210528 85204
rect 204591 85146 204596 85202
rect 204652 85146 210528 85202
rect 640386 85174 640446 85440
rect 647727 85437 647793 85440
rect 650991 85352 651057 85355
rect 650991 85350 656736 85352
rect 650991 85294 650996 85350
rect 651052 85294 656736 85350
rect 650991 85292 656736 85294
rect 650991 85289 651057 85292
rect 663279 85204 663345 85207
rect 663234 85202 663345 85204
rect 204591 85144 210528 85146
rect 663234 85146 663284 85202
rect 663340 85146 663345 85202
rect 204591 85141 204657 85144
rect 663234 85141 663345 85146
rect 646287 85056 646353 85059
rect 640194 85054 646353 85056
rect 640194 84998 646292 85054
rect 646348 84998 646353 85054
rect 640194 84996 646353 84998
rect 204687 84760 204753 84763
rect 204687 84758 210528 84760
rect 204687 84702 204692 84758
rect 204748 84702 210528 84758
rect 640194 84730 640254 84996
rect 646287 84993 646353 84996
rect 204687 84700 210528 84702
rect 204687 84697 204753 84700
rect 140802 84168 140862 84656
rect 663234 84582 663294 85141
rect 663426 84763 663486 85322
rect 663426 84758 663537 84763
rect 663426 84702 663476 84758
rect 663532 84702 663537 84758
rect 663426 84700 663537 84702
rect 663471 84697 663537 84700
rect 650991 84316 651057 84319
rect 650991 84314 656736 84316
rect 650991 84258 650996 84314
rect 651052 84258 656736 84314
rect 650991 84256 656736 84258
rect 650991 84253 651057 84256
rect 146703 84168 146769 84171
rect 140802 84166 146769 84168
rect 140802 84110 146708 84166
rect 146764 84110 146769 84166
rect 140802 84108 146769 84110
rect 146703 84105 146769 84108
rect 204783 84168 204849 84171
rect 645903 84168 645969 84171
rect 204783 84166 210528 84168
rect 204783 84110 204788 84166
rect 204844 84110 210528 84166
rect 204783 84108 210528 84110
rect 640416 84166 645969 84168
rect 640416 84110 645908 84166
rect 645964 84110 645969 84166
rect 640416 84108 645969 84110
rect 204783 84105 204849 84108
rect 645903 84105 645969 84108
rect 651375 83872 651441 83875
rect 640386 83870 651441 83872
rect 640386 83814 651380 83870
rect 651436 83814 651441 83870
rect 640386 83812 651441 83814
rect 140802 83576 140862 83618
rect 144687 83576 144753 83579
rect 140802 83574 144753 83576
rect 140802 83518 144692 83574
rect 144748 83518 144753 83574
rect 140802 83516 144753 83518
rect 144687 83513 144753 83516
rect 204879 83576 204945 83579
rect 204879 83574 210528 83576
rect 204879 83518 204884 83574
rect 204940 83518 210528 83574
rect 640386 83546 640446 83812
rect 651375 83809 651441 83812
rect 204879 83516 210528 83518
rect 204879 83513 204945 83516
rect 647919 83428 647985 83431
rect 640194 83426 647985 83428
rect 640194 83370 647924 83426
rect 647980 83370 647985 83426
rect 640194 83368 647985 83370
rect 204495 83132 204561 83135
rect 204495 83130 210528 83132
rect 204495 83074 204500 83130
rect 204556 83074 210528 83130
rect 640194 83102 640254 83368
rect 647919 83365 647985 83368
rect 651087 83428 651153 83431
rect 651087 83426 656736 83428
rect 651087 83370 651092 83426
rect 651148 83370 656736 83426
rect 651087 83368 656736 83370
rect 651087 83365 651153 83368
rect 204495 83072 210528 83074
rect 204495 83069 204561 83072
rect 663426 82839 663486 83398
rect 663375 82834 663486 82839
rect 663375 82778 663380 82834
rect 663436 82778 663486 82834
rect 663375 82776 663486 82778
rect 663375 82773 663441 82776
rect 650895 82688 650961 82691
rect 650895 82686 656736 82688
rect 650895 82630 650900 82686
rect 650956 82630 656736 82686
rect 650895 82628 656736 82630
rect 650895 82625 650961 82628
rect 204591 82540 204657 82543
rect 647919 82540 647985 82543
rect 204591 82538 210528 82540
rect 204591 82482 204596 82538
rect 204652 82482 210528 82538
rect 204591 82480 210528 82482
rect 640416 82538 647985 82540
rect 640416 82482 647924 82538
rect 647980 82482 647985 82538
rect 640416 82480 647985 82482
rect 204591 82477 204657 82480
rect 647919 82477 647985 82480
rect 144015 82392 144081 82395
rect 140832 82390 144081 82392
rect 140832 82334 144020 82390
rect 144076 82334 144081 82390
rect 140832 82332 144081 82334
rect 144015 82329 144081 82332
rect 647535 82244 647601 82247
rect 640386 82242 647601 82244
rect 640386 82186 647540 82242
rect 647596 82186 647601 82242
rect 640386 82184 647601 82186
rect 204495 81948 204561 81951
rect 204495 81946 210528 81948
rect 204495 81890 204500 81946
rect 204556 81890 210528 81946
rect 640386 81918 640446 82184
rect 647535 82181 647601 82184
rect 663234 82099 663294 82658
rect 663234 82094 663345 82099
rect 663234 82038 663284 82094
rect 663340 82038 663345 82094
rect 663234 82036 663345 82038
rect 663279 82033 663345 82036
rect 204495 81888 210528 81890
rect 204495 81885 204561 81888
rect 204687 81504 204753 81507
rect 204687 81502 210528 81504
rect 204687 81446 204692 81502
rect 204748 81446 210528 81502
rect 204687 81444 210528 81446
rect 204687 81441 204753 81444
rect 640386 81356 640446 81474
rect 647919 81356 647985 81359
rect 640386 81354 647985 81356
rect 640386 81298 647924 81354
rect 647980 81298 647985 81354
rect 640386 81296 647985 81298
rect 647919 81293 647985 81296
rect 662895 81208 662961 81211
rect 663042 81208 663102 81770
rect 662895 81206 663102 81208
rect 140802 80764 140862 81170
rect 662895 81150 662900 81206
rect 662956 81150 663102 81206
rect 662895 81148 663102 81150
rect 662895 81145 662961 81148
rect 204783 80912 204849 80915
rect 647151 80912 647217 80915
rect 204783 80910 210528 80912
rect 204783 80854 204788 80910
rect 204844 80854 210528 80910
rect 204783 80852 210528 80854
rect 640416 80910 647217 80912
rect 640416 80854 647156 80910
rect 647212 80854 647217 80910
rect 640416 80852 647217 80854
rect 204783 80849 204849 80852
rect 647151 80849 647217 80852
rect 144399 80764 144465 80767
rect 140802 80762 144465 80764
rect 140802 80706 144404 80762
rect 144460 80706 144465 80762
rect 140802 80704 144465 80706
rect 144399 80701 144465 80704
rect 647823 80468 647889 80471
rect 640386 80466 647889 80468
rect 640386 80410 647828 80466
rect 647884 80410 647889 80466
rect 640386 80408 647889 80410
rect 206895 80320 206961 80323
rect 206895 80318 210528 80320
rect 206895 80262 206900 80318
rect 206956 80262 210528 80318
rect 640386 80290 640446 80408
rect 647823 80405 647889 80408
rect 206895 80260 210528 80262
rect 206895 80257 206961 80260
rect 205455 80172 205521 80175
rect 647919 80172 647985 80175
rect 205455 80170 210558 80172
rect 205455 80114 205460 80170
rect 205516 80114 210558 80170
rect 205455 80112 210558 80114
rect 205455 80109 205521 80112
rect 140802 79432 140862 79920
rect 210498 79772 210558 80112
rect 640386 80170 647985 80172
rect 640386 80114 647924 80170
rect 647980 80114 647985 80170
rect 640386 80112 647985 80114
rect 640386 79772 640446 80112
rect 647919 80109 647985 80112
rect 144111 79432 144177 79435
rect 140802 79430 144177 79432
rect 140802 79374 144116 79430
rect 144172 79374 144177 79430
rect 140802 79372 144177 79374
rect 144111 79369 144177 79372
rect 204687 79284 204753 79287
rect 647919 79284 647985 79287
rect 204687 79282 210528 79284
rect 204687 79226 204692 79282
rect 204748 79226 210528 79282
rect 204687 79224 210528 79226
rect 640416 79282 647985 79284
rect 640416 79226 647924 79282
rect 647980 79226 647985 79282
rect 640416 79224 647985 79226
rect 204687 79221 204753 79224
rect 647919 79221 647985 79224
rect 144015 78692 144081 78695
rect 140832 78690 144081 78692
rect 140832 78634 144020 78690
rect 144076 78634 144081 78690
rect 140832 78632 144081 78634
rect 144015 78629 144081 78632
rect 204495 78692 204561 78695
rect 646095 78692 646161 78695
rect 204495 78690 210528 78692
rect 204495 78634 204500 78690
rect 204556 78634 210528 78690
rect 204495 78632 210528 78634
rect 640416 78690 646161 78692
rect 640416 78634 646100 78690
rect 646156 78634 646161 78690
rect 640416 78632 646161 78634
rect 204495 78629 204561 78632
rect 646095 78629 646161 78632
rect 204591 78544 204657 78547
rect 646863 78544 646929 78547
rect 204591 78542 210558 78544
rect 204591 78486 204596 78542
rect 204652 78486 210558 78542
rect 204591 78484 210558 78486
rect 204591 78481 204657 78484
rect 210498 78144 210558 78484
rect 640386 78542 646929 78544
rect 640386 78486 646868 78542
rect 646924 78486 646929 78542
rect 640386 78484 646929 78486
rect 640386 78144 640446 78484
rect 646863 78481 646929 78484
rect 210159 77806 210225 77807
rect 210106 77742 210112 77806
rect 210176 77804 210225 77806
rect 210176 77802 210268 77804
rect 210220 77746 210268 77802
rect 210176 77744 210268 77746
rect 210176 77742 210225 77744
rect 210159 77741 210225 77742
rect 204591 77656 204657 77659
rect 647919 77656 647985 77659
rect 204591 77654 210528 77656
rect 204591 77598 204596 77654
rect 204652 77598 210528 77654
rect 204591 77596 210528 77598
rect 640416 77654 647985 77656
rect 640416 77598 647924 77654
rect 647980 77598 647985 77654
rect 640416 77596 647985 77598
rect 204591 77593 204657 77596
rect 647919 77593 647985 77596
rect 144111 77508 144177 77511
rect 140832 77506 144177 77508
rect 140832 77450 144116 77506
rect 144172 77450 144177 77506
rect 140832 77448 144177 77450
rect 144111 77445 144177 77448
rect 204495 77064 204561 77067
rect 647919 77064 647985 77067
rect 204495 77062 210528 77064
rect 204495 77006 204500 77062
rect 204556 77006 210528 77062
rect 204495 77004 210528 77006
rect 640416 77062 647985 77064
rect 640416 77006 647924 77062
rect 647980 77006 647985 77062
rect 640416 77004 647985 77006
rect 204495 77001 204561 77004
rect 647919 77001 647985 77004
rect 204687 76916 204753 76919
rect 646479 76916 646545 76919
rect 204687 76914 210558 76916
rect 204687 76858 204692 76914
rect 204748 76858 210558 76914
rect 204687 76856 210558 76858
rect 204687 76853 204753 76856
rect 210498 76516 210558 76856
rect 640386 76914 646545 76916
rect 640386 76858 646484 76914
rect 646540 76858 646545 76914
rect 640386 76856 646545 76858
rect 640386 76516 640446 76856
rect 646479 76853 646545 76856
rect 146031 76472 146097 76475
rect 146031 76470 146430 76472
rect 146031 76414 146036 76470
rect 146092 76414 146430 76470
rect 146031 76412 146430 76414
rect 146031 76409 146097 76412
rect 140802 75732 140862 76220
rect 146370 76028 146430 76412
rect 146511 76028 146577 76031
rect 146370 76026 146577 76028
rect 146370 75970 146516 76026
rect 146572 75970 146577 76026
rect 146370 75968 146577 75970
rect 146511 75965 146577 75968
rect 204783 76028 204849 76031
rect 646479 76028 646545 76031
rect 204783 76026 210528 76028
rect 204783 75970 204788 76026
rect 204844 75970 210528 76026
rect 204783 75968 210528 75970
rect 640416 76026 646545 76028
rect 640416 75970 646484 76026
rect 646540 75970 646545 76026
rect 640416 75968 646545 75970
rect 204783 75965 204849 75968
rect 646479 75965 646545 75968
rect 144015 75732 144081 75735
rect 140802 75730 144081 75732
rect 140802 75674 144020 75730
rect 144076 75674 144081 75730
rect 140802 75672 144081 75674
rect 144015 75669 144081 75672
rect 204879 75436 204945 75439
rect 646863 75436 646929 75439
rect 204879 75434 210528 75436
rect 204879 75378 204884 75434
rect 204940 75378 210528 75434
rect 204879 75376 210528 75378
rect 640416 75434 646929 75436
rect 640416 75378 646868 75434
rect 646924 75378 646929 75434
rect 640416 75376 646929 75378
rect 204879 75373 204945 75376
rect 646863 75373 646929 75376
rect 204975 75288 205041 75291
rect 204975 75286 210558 75288
rect 204975 75230 204980 75286
rect 205036 75230 210558 75286
rect 204975 75228 210558 75230
rect 204975 75225 205041 75228
rect 140802 75140 140862 75184
rect 146895 75140 146961 75143
rect 140802 75138 146961 75140
rect 140802 75082 146900 75138
rect 146956 75082 146961 75138
rect 140802 75080 146961 75082
rect 146895 75077 146961 75080
rect 210498 74888 210558 75228
rect 647919 75140 647985 75143
rect 640386 75138 647985 75140
rect 640386 75082 647924 75138
rect 647980 75082 647985 75138
rect 640386 75080 647985 75082
rect 640386 74888 640446 75080
rect 647919 75077 647985 75080
rect 204495 74400 204561 74403
rect 646959 74400 647025 74403
rect 204495 74398 210528 74400
rect 204495 74342 204500 74398
rect 204556 74342 210528 74398
rect 204495 74340 210528 74342
rect 640416 74398 647025 74400
rect 640416 74342 646964 74398
rect 647020 74342 647025 74398
rect 640416 74340 647025 74342
rect 204495 74337 204561 74340
rect 646959 74337 647025 74340
rect 144015 73956 144081 73959
rect 140832 73954 144081 73956
rect 140832 73898 144020 73954
rect 144076 73898 144081 73954
rect 140832 73896 144081 73898
rect 144015 73893 144081 73896
rect 204591 73808 204657 73811
rect 647823 73808 647889 73811
rect 204591 73806 210528 73808
rect 204591 73750 204596 73806
rect 204652 73750 210528 73806
rect 204591 73748 210528 73750
rect 640416 73806 647889 73808
rect 640416 73750 647828 73806
rect 647884 73750 647889 73806
rect 640416 73748 647889 73750
rect 204591 73745 204657 73748
rect 647823 73745 647889 73748
rect 204687 73660 204753 73663
rect 204687 73658 210558 73660
rect 204687 73602 204692 73658
rect 204748 73602 210558 73658
rect 204687 73600 210558 73602
rect 204687 73597 204753 73600
rect 210498 73260 210558 73600
rect 640386 73068 640446 73260
rect 647919 73068 647985 73071
rect 640386 73066 647985 73068
rect 640386 73010 647924 73066
rect 647980 73010 647985 73066
rect 640386 73008 647985 73010
rect 647919 73005 647985 73008
rect 144111 72772 144177 72775
rect 140832 72770 144177 72772
rect 140832 72714 144116 72770
rect 144172 72714 144177 72770
rect 140832 72712 144177 72714
rect 144111 72709 144177 72712
rect 204783 72772 204849 72775
rect 646479 72772 646545 72775
rect 204783 72770 210528 72772
rect 204783 72714 204788 72770
rect 204844 72714 210528 72770
rect 204783 72712 210528 72714
rect 640416 72770 646545 72772
rect 640416 72714 646484 72770
rect 646540 72714 646545 72770
rect 640416 72712 646545 72714
rect 204783 72709 204849 72712
rect 646479 72709 646545 72712
rect 204879 72180 204945 72183
rect 646671 72180 646737 72183
rect 204879 72178 210528 72180
rect 204879 72122 204884 72178
rect 204940 72122 210528 72178
rect 204879 72120 210528 72122
rect 640416 72178 646737 72180
rect 640416 72122 646676 72178
rect 646732 72122 646737 72178
rect 640416 72120 646737 72122
rect 204879 72117 204945 72120
rect 646671 72117 646737 72120
rect 204495 71736 204561 71739
rect 204495 71734 210558 71736
rect 204495 71678 204500 71734
rect 204556 71678 210558 71734
rect 204495 71676 210558 71678
rect 204495 71673 204561 71676
rect 210498 71632 210558 71676
rect 140802 71292 140862 71484
rect 144015 71292 144081 71295
rect 140802 71290 144081 71292
rect 140802 71234 144020 71290
rect 144076 71234 144081 71290
rect 140802 71232 144081 71234
rect 144015 71229 144081 71232
rect 204591 71144 204657 71147
rect 204591 71142 210528 71144
rect 204591 71086 204596 71142
rect 204652 71086 210528 71142
rect 204591 71084 210528 71086
rect 204591 71081 204657 71084
rect 204687 70552 204753 70555
rect 204687 70550 210528 70552
rect 204687 70494 204692 70550
rect 204748 70494 210528 70550
rect 204687 70492 210528 70494
rect 204687 70489 204753 70492
rect 140802 69812 140862 70290
rect 204783 69960 204849 69963
rect 204783 69958 210528 69960
rect 204783 69902 204788 69958
rect 204844 69902 210528 69958
rect 204783 69900 210528 69902
rect 204783 69897 204849 69900
rect 144015 69812 144081 69815
rect 140802 69810 144081 69812
rect 140802 69754 144020 69810
rect 144076 69754 144081 69810
rect 140802 69752 144081 69754
rect 144015 69749 144081 69752
rect 204879 69516 204945 69519
rect 204879 69514 210528 69516
rect 204879 69458 204884 69514
rect 204940 69458 210528 69514
rect 204879 69456 210528 69458
rect 204879 69453 204945 69456
rect 146511 69072 146577 69075
rect 140832 69070 146577 69072
rect 140832 69014 146516 69070
rect 146572 69014 146577 69070
rect 140832 69012 146577 69014
rect 146511 69009 146577 69012
rect 204495 68924 204561 68927
rect 204495 68922 210528 68924
rect 204495 68866 204500 68922
rect 204556 68866 210528 68922
rect 204495 68864 210528 68866
rect 204495 68861 204561 68864
rect 204591 68332 204657 68335
rect 204591 68330 210528 68332
rect 204591 68274 204596 68330
rect 204652 68274 210528 68330
rect 204591 68272 210528 68274
rect 204591 68269 204657 68272
rect 140802 67740 140862 67932
rect 204687 67888 204753 67891
rect 204687 67886 210528 67888
rect 204687 67830 204692 67886
rect 204748 67830 210528 67886
rect 204687 67828 210528 67830
rect 204687 67825 204753 67828
rect 144015 67740 144081 67743
rect 140802 67738 144081 67740
rect 140802 67682 144020 67738
rect 144076 67682 144081 67738
rect 140802 67680 144081 67682
rect 144015 67677 144081 67680
rect 204783 67296 204849 67299
rect 204783 67294 210528 67296
rect 204783 67238 204788 67294
rect 204844 67238 210528 67294
rect 204783 67236 210528 67238
rect 204783 67233 204849 67236
rect 140802 66408 140862 66748
rect 204879 66704 204945 66707
rect 204879 66702 210528 66704
rect 204879 66646 204884 66702
rect 204940 66646 210528 66702
rect 204879 66644 210528 66646
rect 204879 66641 204945 66644
rect 144207 66408 144273 66411
rect 140802 66406 144273 66408
rect 140802 66350 144212 66406
rect 144268 66350 144273 66406
rect 140802 66348 144273 66350
rect 144207 66345 144273 66348
rect 204591 66260 204657 66263
rect 204591 66258 210528 66260
rect 204591 66202 204596 66258
rect 204652 66202 210528 66258
rect 204591 66200 210528 66202
rect 204591 66197 204657 66200
rect 204495 65668 204561 65671
rect 204495 65666 210528 65668
rect 204495 65610 204500 65666
rect 204556 65610 210528 65666
rect 204495 65608 210528 65610
rect 204495 65605 204561 65608
rect 144015 65520 144081 65523
rect 140832 65518 144081 65520
rect 140832 65462 144020 65518
rect 144076 65462 144081 65518
rect 140832 65460 144081 65462
rect 144015 65457 144081 65460
rect 204687 65076 204753 65079
rect 204687 65074 210528 65076
rect 204687 65018 204692 65074
rect 204748 65018 210528 65074
rect 204687 65016 210528 65018
rect 204687 65013 204753 65016
rect 144879 64780 144945 64783
rect 140802 64778 144945 64780
rect 140802 64722 144884 64778
rect 144940 64722 144945 64778
rect 140802 64720 144945 64722
rect 140802 64334 140862 64720
rect 144879 64717 144945 64720
rect 204495 64632 204561 64635
rect 204495 64630 210528 64632
rect 204495 64574 204500 64630
rect 204556 64574 210528 64630
rect 204495 64572 210528 64574
rect 204495 64569 204561 64572
rect 204591 64040 204657 64043
rect 204591 64038 210528 64040
rect 204591 63982 204596 64038
rect 204652 63982 210528 64038
rect 204591 63980 210528 63982
rect 204591 63977 204657 63980
rect 204495 63448 204561 63451
rect 204495 63446 210528 63448
rect 204495 63390 204500 63446
rect 204556 63390 210528 63446
rect 204495 63388 210528 63390
rect 204495 63385 204561 63388
rect 140802 62708 140862 63048
rect 204591 63004 204657 63007
rect 204591 63002 210528 63004
rect 204591 62946 204596 63002
rect 204652 62946 210528 63002
rect 204591 62944 210528 62946
rect 204591 62941 204657 62944
rect 144015 62708 144081 62711
rect 140802 62706 144081 62708
rect 140802 62650 144020 62706
rect 144076 62650 144081 62706
rect 140802 62648 144081 62650
rect 144015 62645 144081 62648
rect 146895 62412 146961 62415
rect 140802 62410 146961 62412
rect 140802 62354 146900 62410
rect 146956 62354 146961 62410
rect 140802 62352 146961 62354
rect 140802 61864 140862 62352
rect 146895 62349 146961 62352
rect 204687 62412 204753 62415
rect 204687 62410 210528 62412
rect 204687 62354 204692 62410
rect 204748 62354 210528 62410
rect 204687 62352 210528 62354
rect 204687 62349 204753 62352
rect 204879 61820 204945 61823
rect 204879 61818 210528 61820
rect 204879 61762 204884 61818
rect 204940 61762 210528 61818
rect 204879 61760 210528 61762
rect 204879 61757 204945 61760
rect 204783 61376 204849 61379
rect 204783 61374 210528 61376
rect 204783 61318 204788 61374
rect 204844 61318 210528 61374
rect 204783 61316 210528 61318
rect 204783 61313 204849 61316
rect 146895 60784 146961 60787
rect 140832 60782 146961 60784
rect 140832 60726 146900 60782
rect 146956 60726 146961 60782
rect 140832 60724 146961 60726
rect 146895 60721 146961 60724
rect 204495 60784 204561 60787
rect 204495 60782 210528 60784
rect 204495 60726 204500 60782
rect 204556 60726 210528 60782
rect 204495 60724 210528 60726
rect 204495 60721 204561 60724
rect 204591 60192 204657 60195
rect 204591 60190 210528 60192
rect 204591 60134 204596 60190
rect 204652 60134 210528 60190
rect 204591 60132 210528 60134
rect 204591 60129 204657 60132
rect 204495 60044 204561 60047
rect 204495 60042 210558 60044
rect 204495 59986 204500 60042
rect 204556 59986 210558 60042
rect 204495 59984 210558 59986
rect 204495 59981 204561 59984
rect 210498 59644 210558 59984
rect 144015 59600 144081 59603
rect 140832 59598 144081 59600
rect 140832 59542 144020 59598
rect 144076 59542 144081 59598
rect 140832 59540 144081 59542
rect 144015 59537 144081 59540
rect 204687 59156 204753 59159
rect 204687 59154 210528 59156
rect 204687 59098 204692 59154
rect 204748 59098 210528 59154
rect 204687 59096 210528 59098
rect 204687 59093 204753 59096
rect 144015 58712 144081 58715
rect 140802 58710 144081 58712
rect 140802 58654 144020 58710
rect 144076 58654 144081 58710
rect 140802 58652 144081 58654
rect 140802 58322 140862 58652
rect 144015 58649 144081 58652
rect 210882 58270 210942 58534
rect 210874 58206 210880 58270
rect 210944 58206 210950 58270
rect 210690 57678 210750 58016
rect 210682 57614 210688 57678
rect 210752 57614 210758 57678
rect 207279 57528 207345 57531
rect 207279 57526 210528 57528
rect 207279 57470 207284 57526
rect 207340 57470 210528 57526
rect 207279 57468 210528 57470
rect 207279 57465 207345 57468
rect 144015 57084 144081 57087
rect 140832 57082 144081 57084
rect 140832 57026 144020 57082
rect 144076 57026 144081 57082
rect 140832 57024 144081 57026
rect 144015 57021 144081 57024
rect 209295 56640 209361 56643
rect 210498 56640 210558 56906
rect 209295 56638 210558 56640
rect 209295 56582 209300 56638
rect 209356 56582 210558 56638
rect 209295 56580 210558 56582
rect 209295 56577 209361 56580
rect 144015 56196 144081 56199
rect 140802 56194 144081 56196
rect 140802 56138 144020 56194
rect 144076 56138 144081 56194
rect 140802 56136 144081 56138
rect 140802 55874 140862 56136
rect 144015 56133 144081 56136
rect 210159 56048 210225 56051
rect 210498 56048 210558 56388
rect 210159 56046 210558 56048
rect 210159 55990 210164 56046
rect 210220 55990 210558 56046
rect 210159 55988 210558 55990
rect 210159 55985 210225 55988
rect 206895 55900 206961 55903
rect 206895 55898 210528 55900
rect 206895 55842 206900 55898
rect 206956 55842 210528 55898
rect 206895 55840 210528 55842
rect 206895 55837 206961 55840
rect 210255 55012 210321 55015
rect 210498 55012 210558 55278
rect 210255 55010 210558 55012
rect 210255 54954 210260 55010
rect 210316 54954 210558 55010
rect 210255 54952 210558 54954
rect 210255 54949 210321 54952
rect 144015 54716 144081 54719
rect 140832 54714 144081 54716
rect 140832 54658 144020 54714
rect 144076 54658 144081 54714
rect 140832 54656 144081 54658
rect 144015 54653 144081 54656
rect 210882 54275 210942 54760
rect 210831 54270 210942 54275
rect 210831 54214 210836 54270
rect 210892 54214 210942 54270
rect 210831 54212 210942 54214
rect 210831 54209 210897 54212
rect 211258 54210 211264 54274
rect 211328 54272 211334 54274
rect 212418 54272 213006 54309
rect 214767 54272 214833 54275
rect 211328 54270 214833 54272
rect 211328 54249 214772 54270
rect 211328 54212 212478 54249
rect 212946 54214 214772 54249
rect 214828 54214 214833 54270
rect 212946 54212 214833 54214
rect 211328 54210 211334 54212
rect 214767 54209 214833 54212
rect 210735 54126 210801 54127
rect 210682 54124 210688 54126
rect 210644 54064 210688 54124
rect 210752 54122 210801 54126
rect 210796 54066 210801 54122
rect 210682 54062 210688 54064
rect 210752 54062 210801 54066
rect 212602 54062 212608 54126
rect 212672 54124 212678 54126
rect 216975 54124 217041 54127
rect 212672 54122 217041 54124
rect 212672 54066 216980 54122
rect 217036 54066 217041 54122
rect 212672 54064 217041 54066
rect 212672 54062 212678 54064
rect 210735 54061 210801 54062
rect 216975 54061 217041 54064
rect 210874 53914 210880 53978
rect 210944 53976 210950 53978
rect 221391 53976 221457 53979
rect 210944 53974 221457 53976
rect 210944 53918 221396 53974
rect 221452 53918 221457 53974
rect 210944 53916 221457 53918
rect 210944 53914 210950 53916
rect 221391 53913 221457 53916
rect 144015 53828 144081 53831
rect 140802 53826 144081 53828
rect 140802 53770 144020 53826
rect 144076 53770 144081 53826
rect 140802 53768 144081 53770
rect 140802 53576 140862 53768
rect 144015 53765 144081 53768
rect 211066 53766 211072 53830
rect 211136 53828 211142 53830
rect 211136 53768 216126 53828
rect 211136 53766 211142 53768
rect 212026 53618 212032 53682
rect 212096 53680 212102 53682
rect 216066 53680 216126 53768
rect 212096 53620 213246 53680
rect 216066 53620 221118 53680
rect 212096 53618 212102 53620
rect 211834 53470 211840 53534
rect 211904 53532 211910 53534
rect 213039 53532 213105 53535
rect 211904 53530 213105 53532
rect 211904 53474 213044 53530
rect 213100 53474 213105 53530
rect 211904 53472 213105 53474
rect 213186 53532 213246 53620
rect 221058 53535 221118 53620
rect 215967 53532 216033 53535
rect 213186 53530 216033 53532
rect 213186 53474 215972 53530
rect 216028 53474 216033 53530
rect 213186 53472 216033 53474
rect 221058 53530 221169 53535
rect 221058 53474 221108 53530
rect 221164 53474 221169 53530
rect 221058 53472 221169 53474
rect 211904 53470 211910 53472
rect 213039 53469 213105 53472
rect 215967 53469 216033 53472
rect 221103 53469 221169 53472
rect 212410 53322 212416 53386
rect 212480 53384 212486 53386
rect 216687 53384 216753 53387
rect 212480 53382 216753 53384
rect 212480 53326 216692 53382
rect 216748 53326 216753 53382
rect 212480 53324 216753 53326
rect 212480 53322 212486 53324
rect 216687 53321 216753 53324
rect 273615 53273 273681 53276
rect 273615 53271 273726 53273
rect 212794 53174 212800 53238
rect 212864 53236 212870 53238
rect 217839 53236 217905 53239
rect 212864 53234 217905 53236
rect 212864 53178 217844 53234
rect 217900 53178 217905 53234
rect 273615 53215 273620 53271
rect 273676 53236 273726 53271
rect 293679 53236 293745 53239
rect 273676 53234 293745 53236
rect 273676 53215 293684 53234
rect 273615 53210 293684 53215
rect 212864 53176 217905 53178
rect 273666 53178 293684 53210
rect 293740 53178 293745 53234
rect 273666 53176 293745 53178
rect 212864 53174 212870 53176
rect 217839 53173 217905 53176
rect 293679 53173 293745 53176
rect 440655 53236 440721 53239
rect 443727 53236 443793 53239
rect 440655 53234 443793 53236
rect 440655 53178 440660 53234
rect 440716 53178 443732 53234
rect 443788 53178 443793 53234
rect 440655 53176 443793 53178
rect 440655 53173 440721 53176
rect 443727 53173 443793 53176
rect 221871 52348 221937 52351
rect 637690 52348 637696 52350
rect 221871 52346 637696 52348
rect 221871 52290 221876 52346
rect 221932 52290 637696 52346
rect 221871 52288 637696 52290
rect 221871 52285 221937 52288
rect 637690 52286 637696 52288
rect 637760 52286 637766 52350
rect 223311 52200 223377 52203
rect 637882 52200 637888 52202
rect 223311 52198 637888 52200
rect 223311 52142 223316 52198
rect 223372 52142 637888 52198
rect 223311 52140 637888 52142
rect 223311 52137 223377 52140
rect 637882 52138 637888 52140
rect 637952 52138 637958 52202
rect 212655 52052 212721 52055
rect 637498 52052 637504 52054
rect 212655 52050 637504 52052
rect 212655 51994 212660 52050
rect 212716 51994 637504 52050
rect 212655 51992 637504 51994
rect 212655 51989 212721 51992
rect 637498 51990 637504 51992
rect 637568 51990 637574 52054
rect 211983 51904 212049 51907
rect 637306 51904 637312 51906
rect 211983 51902 637312 51904
rect 211983 51846 211988 51902
rect 212044 51846 637312 51902
rect 211983 51844 637312 51846
rect 211983 51841 212049 51844
rect 637306 51842 637312 51844
rect 637376 51842 637382 51906
rect 222639 51756 222705 51759
rect 636922 51756 636928 51758
rect 222639 51754 636928 51756
rect 222639 51698 222644 51754
rect 222700 51698 636928 51754
rect 222639 51696 636928 51698
rect 222639 51693 222705 51696
rect 636922 51694 636928 51696
rect 636992 51694 636998 51758
rect 145402 51546 145408 51610
rect 145472 51608 145478 51610
rect 243375 51608 243441 51611
rect 145472 51606 243441 51608
rect 145472 51550 243380 51606
rect 243436 51550 243441 51606
rect 145472 51548 243441 51550
rect 145472 51546 145478 51548
rect 243375 51545 243441 51548
rect 374415 51608 374481 51611
rect 394287 51608 394353 51611
rect 374415 51606 394353 51608
rect 374415 51550 374420 51606
rect 374476 51550 394292 51606
rect 394348 51550 394353 51606
rect 374415 51548 394353 51550
rect 374415 51545 374481 51548
rect 394287 51545 394353 51548
rect 457935 51608 458001 51611
rect 477999 51608 478065 51611
rect 457935 51606 478065 51608
rect 457935 51550 457940 51606
rect 457996 51550 478004 51606
rect 478060 51550 478065 51606
rect 457935 51548 478065 51550
rect 457935 51545 458001 51548
rect 477999 51545 478065 51548
rect 498255 51608 498321 51611
rect 518319 51608 518385 51611
rect 498255 51606 518385 51608
rect 498255 51550 498260 51606
rect 498316 51550 518324 51606
rect 518380 51550 518385 51606
rect 498255 51548 518385 51550
rect 498255 51545 498321 51548
rect 518319 51545 518385 51548
rect 538575 51608 538641 51611
rect 541455 51608 541521 51611
rect 538575 51606 541521 51608
rect 538575 51550 538580 51606
rect 538636 51550 541460 51606
rect 541516 51550 541521 51606
rect 538575 51548 541521 51550
rect 538575 51545 538641 51548
rect 541455 51545 541521 51548
rect 584655 51608 584721 51611
rect 604719 51608 604785 51611
rect 584655 51606 604785 51608
rect 584655 51550 584660 51606
rect 584716 51550 604724 51606
rect 604780 51550 604785 51606
rect 584655 51548 604785 51550
rect 584655 51545 584721 51548
rect 604719 51545 604785 51548
rect 145594 51398 145600 51462
rect 145664 51460 145670 51462
rect 237615 51460 237681 51463
rect 145664 51458 237681 51460
rect 145664 51402 237620 51458
rect 237676 51402 237681 51458
rect 145664 51400 237681 51402
rect 145664 51398 145670 51400
rect 237615 51397 237681 51400
rect 145786 51250 145792 51314
rect 145856 51312 145862 51314
rect 237519 51312 237585 51315
rect 145856 51310 237585 51312
rect 145856 51254 237524 51310
rect 237580 51254 237585 51310
rect 145856 51252 237585 51254
rect 145856 51250 145862 51252
rect 237519 51249 237585 51252
rect 229647 50424 229713 50427
rect 637114 50424 637120 50426
rect 229647 50422 637120 50424
rect 229647 50366 229652 50422
rect 229708 50366 637120 50422
rect 229647 50364 637120 50366
rect 229647 50361 229713 50364
rect 637114 50362 637120 50364
rect 637184 50362 637190 50426
rect 512271 49092 512337 49095
rect 520378 49092 520384 49094
rect 512271 49090 520384 49092
rect 512271 49034 512276 49090
rect 512332 49034 520384 49090
rect 512271 49032 520384 49034
rect 512271 49029 512337 49032
rect 520378 49030 520384 49032
rect 520448 49030 520454 49094
rect 168399 48796 168465 48799
rect 242415 48796 242481 48799
rect 168399 48794 242481 48796
rect 168399 48738 168404 48794
rect 168460 48738 242420 48794
rect 242476 48738 242481 48794
rect 168399 48736 242481 48738
rect 168399 48733 168465 48736
rect 242415 48733 242481 48736
rect 171279 48648 171345 48651
rect 242031 48648 242097 48651
rect 171279 48646 242097 48648
rect 171279 48590 171284 48646
rect 171340 48590 242036 48646
rect 242092 48590 242097 48646
rect 171279 48588 242097 48590
rect 171279 48585 171345 48588
rect 242031 48585 242097 48588
rect 174159 48500 174225 48503
rect 242991 48500 243057 48503
rect 174159 48498 243057 48500
rect 174159 48442 174164 48498
rect 174220 48442 242996 48498
rect 243052 48442 243057 48498
rect 174159 48440 243057 48442
rect 174159 48437 174225 48440
rect 242991 48437 243057 48440
rect 182799 48352 182865 48355
rect 243759 48352 243825 48355
rect 182799 48350 243825 48352
rect 182799 48294 182804 48350
rect 182860 48294 243764 48350
rect 243820 48294 243825 48350
rect 182799 48292 243825 48294
rect 182799 48289 182865 48292
rect 243759 48289 243825 48292
rect 165519 48204 165585 48207
rect 241935 48204 242001 48207
rect 165519 48202 242001 48204
rect 165519 48146 165524 48202
rect 165580 48146 241940 48202
rect 241996 48146 242001 48202
rect 165519 48144 242001 48146
rect 165519 48141 165585 48144
rect 241935 48141 242001 48144
rect 460815 46132 460881 46135
rect 465807 46132 465873 46135
rect 460815 46130 465873 46132
rect 460815 46074 460820 46130
rect 460876 46074 465812 46130
rect 465868 46074 465873 46130
rect 460815 46072 465873 46074
rect 460815 46069 460881 46072
rect 465807 46069 465873 46072
rect 212079 45244 212145 45247
rect 302458 45244 302464 45246
rect 212079 45242 302464 45244
rect 212079 45186 212084 45242
rect 212140 45186 302464 45242
rect 212079 45184 302464 45186
rect 212079 45181 212145 45184
rect 302458 45182 302464 45184
rect 302528 45182 302534 45246
rect 211695 45096 211761 45099
rect 362938 45096 362944 45098
rect 211695 45094 362944 45096
rect 211695 45038 211700 45094
rect 211756 45038 362944 45094
rect 211695 45036 362944 45038
rect 211695 45033 211761 45036
rect 362938 45034 362944 45036
rect 363008 45034 363014 45098
rect 215439 44948 215505 44951
rect 527098 44948 527104 44950
rect 215439 44946 527104 44948
rect 215439 44890 215444 44946
rect 215500 44890 527104 44946
rect 215439 44888 527104 44890
rect 215439 44885 215505 44888
rect 527098 44886 527104 44888
rect 527168 44886 527174 44950
rect 302511 43322 302577 43323
rect 302458 43320 302464 43322
rect 302420 43260 302464 43320
rect 302528 43318 302577 43322
rect 302572 43262 302577 43318
rect 302458 43258 302464 43260
rect 302528 43258 302577 43262
rect 362938 43258 362944 43322
rect 363008 43320 363014 43322
rect 364911 43320 364977 43323
rect 363008 43318 364977 43320
rect 363008 43262 364916 43318
rect 364972 43262 364977 43318
rect 363008 43260 364977 43262
rect 363008 43258 363014 43260
rect 302511 43257 302577 43258
rect 364911 43257 364977 43260
rect 527098 43258 527104 43322
rect 527168 43320 527174 43322
rect 529263 43320 529329 43323
rect 527168 43318 529329 43320
rect 527168 43262 529268 43318
rect 529324 43262 529329 43318
rect 527168 43260 529329 43262
rect 527168 43258 527174 43260
rect 529263 43257 529329 43260
rect 302415 42136 302481 42139
rect 306735 42136 306801 42139
rect 302415 42134 306801 42136
rect 302415 42078 302420 42134
rect 302476 42078 306740 42134
rect 306796 42078 306801 42134
rect 302415 42076 306801 42078
rect 302415 42073 302481 42076
rect 306735 42073 306801 42076
rect 411567 42136 411633 42139
rect 416271 42136 416337 42139
rect 520431 42138 520497 42139
rect 520378 42136 520384 42138
rect 411567 42134 416337 42136
rect 411567 42078 411572 42134
rect 411628 42078 416276 42134
rect 416332 42078 416337 42134
rect 411567 42076 416337 42078
rect 520340 42076 520384 42136
rect 520448 42134 520497 42138
rect 520492 42078 520497 42134
rect 411567 42073 411633 42076
rect 416271 42073 416337 42076
rect 520378 42074 520384 42076
rect 520448 42074 520497 42078
rect 520431 42073 520497 42074
rect 187599 41840 187665 41843
rect 189946 41840 189952 41842
rect 187599 41838 189952 41840
rect 187599 41782 187604 41838
rect 187660 41782 189952 41838
rect 187599 41780 189952 41782
rect 187599 41777 187665 41780
rect 189946 41778 189952 41780
rect 190016 41778 190022 41842
rect 194319 41840 194385 41843
rect 194938 41840 194944 41842
rect 194319 41838 194944 41840
rect 194319 41782 194324 41838
rect 194380 41782 194944 41838
rect 194319 41780 194944 41782
rect 194319 41777 194385 41780
rect 194938 41778 194944 41780
rect 195008 41778 195014 41842
rect 509679 41840 509745 41843
rect 518511 41840 518577 41843
rect 509679 41838 518577 41840
rect 509679 41782 509684 41838
rect 509740 41782 518516 41838
rect 518572 41782 518577 41838
rect 509679 41780 518577 41782
rect 509679 41777 509745 41780
rect 518511 41777 518577 41780
rect 189946 40742 189952 40806
rect 190016 40804 190022 40806
rect 211023 40804 211089 40807
rect 190016 40802 211089 40804
rect 190016 40746 211028 40802
rect 211084 40746 211089 40802
rect 190016 40744 211089 40746
rect 190016 40742 190022 40744
rect 211023 40741 211089 40744
rect 194938 40594 194944 40658
rect 195008 40656 195014 40658
rect 640719 40656 640785 40659
rect 195008 40654 640785 40656
rect 195008 40598 640724 40654
rect 640780 40598 640785 40654
rect 195008 40596 640785 40598
rect 195008 40594 195014 40596
rect 640719 40593 640785 40596
rect 136527 40212 136593 40215
rect 136527 40210 141822 40212
rect 136527 40154 136532 40210
rect 136588 40154 141822 40210
rect 136527 40152 141822 40154
rect 136527 40149 136593 40152
rect 141762 39886 141822 40152
<< via3 >>
rect 528256 996082 528320 996146
rect 528256 995490 528320 995554
rect 42304 968702 42368 968766
rect 41728 967134 41792 967138
rect 41728 967078 41780 967134
rect 41780 967078 41792 967134
rect 41728 967074 41792 967078
rect 676672 965742 676736 965806
rect 40768 965002 40832 965066
rect 674560 965002 674624 965066
rect 42496 963966 42560 964030
rect 40960 963374 41024 963438
rect 675904 963374 675968 963438
rect 41152 962634 41216 962698
rect 675712 962546 675776 962550
rect 675712 962490 675724 962546
rect 675724 962490 675776 962546
rect 675712 962486 675776 962490
rect 43072 962338 43136 962402
rect 40384 962190 40448 962254
rect 673984 962190 674048 962254
rect 42880 962042 42944 962106
rect 676096 961450 676160 961514
rect 675328 960710 675392 960774
rect 41536 959674 41600 959738
rect 674368 959230 674432 959294
rect 41920 959142 41984 959146
rect 41920 959086 41932 959142
rect 41932 959086 41984 959142
rect 41920 959082 41984 959086
rect 674752 959082 674816 959146
rect 40576 958490 40640 958554
rect 676480 958342 676544 958406
rect 42688 957750 42752 957814
rect 675136 957602 675200 957666
rect 42112 956182 42176 956186
rect 42112 956126 42124 956182
rect 42124 956126 42176 956182
rect 42112 956122 42176 956126
rect 674944 955974 675008 956038
rect 677056 953458 677120 953522
rect 676864 953310 676928 953374
rect 40384 941766 40448 941830
rect 40384 941322 40448 941386
rect 42112 941322 42176 941386
rect 41728 940878 41792 940942
rect 42688 939398 42752 939462
rect 42304 938658 42368 938722
rect 40576 937622 40640 937686
rect 674560 937622 674624 937686
rect 41920 937030 41984 937094
rect 677056 936586 677120 936650
rect 40768 936438 40832 936502
rect 675904 936142 675968 936206
rect 40960 935846 41024 935910
rect 674752 935550 674816 935614
rect 41536 935402 41600 935466
rect 41152 934810 41216 934874
rect 42496 934366 42560 934430
rect 676672 934366 676736 934430
rect 675712 933774 675776 933838
rect 673984 933330 674048 933394
rect 674944 932738 675008 932802
rect 675136 932146 675200 932210
rect 676096 931702 676160 931766
rect 676480 931110 676544 931174
rect 676864 930666 676928 930730
rect 674176 876942 674240 877006
rect 676096 876498 676160 876562
rect 675328 875758 675392 875822
rect 675520 875818 675584 875822
rect 675520 875762 675532 875818
rect 675532 875762 675584 875818
rect 675520 875758 675584 875762
rect 674368 875610 674432 875674
rect 674560 873982 674624 874046
rect 674368 873538 674432 873602
rect 674944 869838 675008 869902
rect 675136 864658 675200 864722
rect 40384 815966 40448 816030
rect 41152 815966 41216 816030
rect 41344 815522 41408 815586
rect 41536 802054 41600 802118
rect 40960 801906 41024 801970
rect 42880 800722 42944 800786
rect 41920 800574 41984 800638
rect 42496 800426 42560 800490
rect 41728 800338 41792 800342
rect 41728 800282 41780 800338
rect 41780 800282 41792 800338
rect 41728 800278 41792 800282
rect 42112 800338 42176 800342
rect 42112 800282 42164 800338
rect 42164 800282 42176 800338
rect 42112 800278 42176 800282
rect 41920 796134 41984 796198
rect 40960 795986 41024 796050
rect 41920 795986 41984 796050
rect 42112 794270 42176 794274
rect 42112 794214 42124 794270
rect 42124 794214 42176 794270
rect 42112 794210 42176 794214
rect 41728 793826 41792 793830
rect 41728 793770 41780 793826
rect 41780 793770 41792 793826
rect 41728 793766 41792 793770
rect 42112 792138 42176 792202
rect 42112 791842 42176 791906
rect 42880 791902 42944 791906
rect 42880 791846 42892 791902
rect 42892 791846 42944 791902
rect 42880 791842 42944 791846
rect 42496 791694 42560 791758
rect 42112 791162 42176 791166
rect 42112 791106 42124 791162
rect 42124 791106 42176 791162
rect 42112 791102 42176 791106
rect 43072 791102 43136 791166
rect 41728 790570 41792 790574
rect 41728 790514 41780 790570
rect 41780 790514 41792 790570
rect 41728 790510 41792 790514
rect 42688 790510 42752 790574
rect 41536 789326 41600 789390
rect 41920 789178 41984 789242
rect 673984 787994 674048 788058
rect 675328 787106 675392 787170
rect 675904 786662 675968 786726
rect 676288 784886 676352 784950
rect 675712 784206 675776 784210
rect 675712 784150 675724 784206
rect 675724 784150 675776 784206
rect 675712 784146 675776 784150
rect 676672 780594 676736 780658
rect 677056 775562 677120 775626
rect 674752 775414 674816 775478
rect 676864 774970 676928 775034
rect 676672 773786 676736 773850
rect 676672 773638 676736 773702
rect 41152 773490 41216 773554
rect 676864 773046 676928 773110
rect 677824 773046 677888 773110
rect 41536 772898 41600 772962
rect 679168 772898 679232 772962
rect 41344 772750 41408 772814
rect 677248 772602 677312 772666
rect 674752 771714 674816 771778
rect 676480 771714 676544 771778
rect 40960 768606 41024 768670
rect 42496 767866 42560 767930
rect 42688 764610 42752 764674
rect 677824 764670 677888 764674
rect 677824 764614 677836 764670
rect 677836 764614 677888 764670
rect 677824 764610 677888 764614
rect 677248 764462 677312 764526
rect 677824 764462 677888 764526
rect 677056 759726 677120 759790
rect 675520 759282 675584 759346
rect 676864 759282 676928 759346
rect 675136 758838 675200 758902
rect 675136 758246 675200 758310
rect 674176 757950 674240 758014
rect 41152 757654 41216 757718
rect 42880 757358 42944 757422
rect 42112 757210 42176 757274
rect 674560 757210 674624 757274
rect 41920 757122 41984 757126
rect 41920 757066 41972 757122
rect 41972 757066 41984 757122
rect 41920 757062 41984 757066
rect 674752 757062 674816 757126
rect 677248 756618 677312 756682
rect 676096 756026 676160 756090
rect 674368 755212 674432 755276
rect 677824 754990 677888 755054
rect 41920 754902 41984 754906
rect 41920 754846 41932 754902
rect 41932 754846 41984 754902
rect 41920 754842 41984 754846
rect 674752 754398 674816 754462
rect 676480 754398 676544 754462
rect 679168 753954 679232 754018
rect 43072 751882 43136 751946
rect 42688 751734 42752 751798
rect 42880 751054 42944 751058
rect 42880 750998 42932 751054
rect 42932 750998 42944 751054
rect 42880 750994 42944 750998
rect 42112 749870 42176 749874
rect 42112 749814 42124 749870
rect 42124 749814 42176 749870
rect 42112 749810 42176 749814
rect 43072 749218 43136 749282
rect 41920 747798 41984 747802
rect 41920 747742 41972 747798
rect 41972 747742 41984 747798
rect 41920 747738 41984 747742
rect 42304 747738 42368 747802
rect 41728 747206 41792 747210
rect 41728 747150 41780 747206
rect 41780 747150 41792 747206
rect 41728 747146 41792 747150
rect 40960 746998 41024 747062
rect 41152 746850 41216 746914
rect 42496 746258 42560 746322
rect 674176 743150 674240 743214
rect 675520 742174 675584 742178
rect 675520 742118 675532 742174
rect 675532 742118 675584 742174
rect 675520 742114 675584 742118
rect 676096 741670 676160 741734
rect 676672 741670 676736 741734
rect 676864 741670 676928 741734
rect 675136 741522 675200 741586
rect 676480 741522 676544 741586
rect 676672 741374 676736 741438
rect 676864 741374 676928 741438
rect 675136 740042 675200 740106
rect 674944 739154 675008 739218
rect 674368 738562 674432 738626
rect 41344 734270 41408 734334
rect 42112 734270 42176 734334
rect 41344 729534 41408 729598
rect 42112 729090 42176 729154
rect 676672 728054 676736 728118
rect 677824 728054 677888 728118
rect 43072 727758 43136 727822
rect 41536 725242 41600 725306
rect 41152 723022 41216 723086
rect 41728 723022 41792 723086
rect 42880 723022 42944 723086
rect 677248 715474 677312 715538
rect 676864 714882 676928 714946
rect 675904 714290 675968 714354
rect 42688 713994 42752 714058
rect 41728 713906 41792 713910
rect 41728 713850 41780 713906
rect 41780 713850 41792 713906
rect 41728 713846 41792 713850
rect 42304 713846 42368 713910
rect 674752 713846 674816 713910
rect 42496 713314 42560 713318
rect 42496 713258 42508 713314
rect 42508 713258 42560 713314
rect 42496 713254 42560 713258
rect 673984 712958 674048 713022
rect 676288 712662 676352 712726
rect 676480 712218 676544 712282
rect 677824 711626 677888 711690
rect 41728 711034 41792 711098
rect 675328 711034 675392 711098
rect 675712 710590 675776 710654
rect 41728 708666 41792 708730
rect 42880 708666 42944 708730
rect 42496 708518 42560 708582
rect 41152 707926 41216 707990
rect 42688 707838 42752 707842
rect 42688 707782 42740 707838
rect 42740 707782 42752 707838
rect 42688 707778 42752 707782
rect 42304 707334 42368 707398
rect 677056 705766 677120 705770
rect 677056 705710 677108 705766
rect 677108 705710 677120 705766
rect 677056 705706 677120 705710
rect 41536 705410 41600 705474
rect 41920 704730 41984 704734
rect 41920 704674 41932 704730
rect 41932 704674 41984 704730
rect 41920 704670 41984 704674
rect 41728 704138 41792 704142
rect 41728 704082 41780 704138
rect 41780 704082 41792 704138
rect 41728 704078 41792 704082
rect 43072 703546 43136 703550
rect 43072 703490 43084 703546
rect 43084 703490 43136 703546
rect 43072 703486 43136 703490
rect 674752 697862 674816 697926
rect 676672 697270 676736 697334
rect 675328 696886 675392 696890
rect 675328 696830 675380 696886
rect 675380 696830 675392 696886
rect 675328 696826 675392 696830
rect 675904 694754 675968 694818
rect 674560 694310 674624 694374
rect 676480 693422 676544 693486
rect 676288 691942 676352 692006
rect 40768 690166 40832 690230
rect 42112 690166 42176 690230
rect 41344 686910 41408 686974
rect 42112 686466 42176 686530
rect 40768 685874 40832 685938
rect 42880 682322 42944 682386
rect 43072 673294 43136 673358
rect 40576 671134 40640 671138
rect 40576 671078 40588 671134
rect 40588 671078 40640 671134
rect 40576 671074 40640 671078
rect 40960 670926 41024 670990
rect 41728 670926 41792 670990
rect 43072 670838 43136 670842
rect 43072 670782 43124 670838
rect 43124 670782 43136 670838
rect 43072 670778 43136 670782
rect 42496 670630 42560 670694
rect 677056 670186 677120 670250
rect 677248 670186 677312 670250
rect 676864 669594 676928 669658
rect 676096 669150 676160 669214
rect 677824 669002 677888 669066
rect 41728 668558 41792 668622
rect 42304 668410 42368 668474
rect 43264 668410 43328 668474
rect 674176 667744 674240 667808
rect 675136 667522 675200 667586
rect 675520 665894 675584 665958
rect 674944 665302 675008 665366
rect 40960 664562 41024 664626
rect 674368 664488 674432 664552
rect 43072 664118 43136 664182
rect 42496 662846 42560 662850
rect 42496 662790 42508 662846
rect 42508 662790 42560 662846
rect 42496 662786 42560 662790
rect 41728 661514 41792 661518
rect 41728 661458 41780 661514
rect 41780 661458 41792 661514
rect 41728 661454 41792 661458
rect 41920 661366 41984 661370
rect 41920 661310 41932 661366
rect 41932 661310 41984 661366
rect 41920 661306 41984 661310
rect 40576 660270 40640 660334
rect 42880 659530 42944 659594
rect 677056 658790 677120 658854
rect 677824 658790 677888 658854
rect 42304 656126 42368 656190
rect 676288 653610 676352 653674
rect 675136 652574 675200 652638
rect 674368 652130 674432 652194
rect 675520 651450 675584 651454
rect 675520 651394 675532 651450
rect 675532 651394 675584 651450
rect 675520 651390 675584 651394
rect 675712 649822 675776 649826
rect 675712 649766 675724 649822
rect 675724 649766 675776 649822
rect 675712 649762 675776 649766
rect 674944 648874 675008 648938
rect 42112 647098 42176 647162
rect 40768 646950 40832 647014
rect 673984 645322 674048 645386
rect 676288 640290 676352 640354
rect 676096 638514 676160 638578
rect 42880 637182 42944 637246
rect 42304 628006 42368 628070
rect 40768 627858 40832 627922
rect 42496 627858 42560 627922
rect 41344 627770 41408 627774
rect 41344 627714 41356 627770
rect 41356 627714 41408 627770
rect 41344 627710 41408 627714
rect 41728 627710 41792 627774
rect 41920 627474 41984 627478
rect 41920 627418 41972 627474
rect 41972 627418 41984 627474
rect 41920 627414 41984 627418
rect 677248 626378 677312 626442
rect 42112 625638 42176 625702
rect 42688 625638 42752 625702
rect 42112 624898 42176 624962
rect 42688 624898 42752 624962
rect 676864 624810 676928 624814
rect 676864 624754 676876 624810
rect 676876 624754 676928 624810
rect 676864 624750 676928 624754
rect 677056 624602 677120 624666
rect 675328 624158 675392 624222
rect 42880 623418 42944 623482
rect 674752 623122 674816 623186
rect 675904 622530 675968 622594
rect 42496 621494 42560 621558
rect 676672 620902 676736 620966
rect 674560 620310 674624 620374
rect 676480 619866 676544 619930
rect 41728 619570 41792 619634
rect 41536 618386 41600 618450
rect 42688 618386 42752 618450
rect 41728 618298 41792 618302
rect 41728 618242 41780 618298
rect 41780 618242 41792 618298
rect 41728 618238 41792 618242
rect 41920 617854 41984 617858
rect 41920 617798 41972 617854
rect 41972 617798 41984 617854
rect 41920 617794 41984 617798
rect 41344 616610 41408 616674
rect 42304 613502 42368 613566
rect 40768 612762 40832 612826
rect 674176 607730 674240 607794
rect 674752 607138 674816 607202
rect 675328 606398 675392 606462
rect 41536 604770 41600 604834
rect 42112 604770 42176 604834
rect 674560 604770 674624 604834
rect 675904 600182 675968 600246
rect 42112 598998 42176 599062
rect 43072 598998 43136 599062
rect 40576 597814 40640 597878
rect 40768 595594 40832 595658
rect 676672 595298 676736 595362
rect 41344 593966 41408 594030
rect 676480 593374 676544 593438
rect 42496 591894 42560 591958
rect 30592 590710 30656 590774
rect 30592 590266 30656 590330
rect 42496 588342 42560 588406
rect 42304 584642 42368 584706
rect 41728 584554 41792 584558
rect 41728 584498 41740 584554
rect 41740 584498 41792 584554
rect 41728 584494 41792 584498
rect 42496 584494 42560 584558
rect 42112 584406 42176 584410
rect 42112 584350 42124 584406
rect 42124 584350 42176 584406
rect 42112 584346 42176 584350
rect 41920 584258 41984 584262
rect 41920 584202 41972 584258
rect 41972 584202 41984 584258
rect 41920 584198 41984 584202
rect 42880 584198 42944 584262
rect 41920 582038 41984 582042
rect 41920 581982 41932 582038
rect 41932 581982 41984 582038
rect 41920 581978 41984 581982
rect 41344 580202 41408 580266
rect 677056 579462 677120 579526
rect 677248 579462 677312 579526
rect 42688 578870 42752 578934
rect 43072 578870 43136 578934
rect 675520 578870 675584 578934
rect 42880 578426 42944 578490
rect 676288 578426 676352 578490
rect 42304 578278 42368 578342
rect 675136 577834 675200 577898
rect 42496 577538 42560 577602
rect 675712 577242 675776 577306
rect 673984 576502 674048 576566
rect 676096 576206 676160 576270
rect 674368 575318 674432 575382
rect 674944 575170 675008 575234
rect 42688 574874 42752 574938
rect 41536 574578 41600 574642
rect 42112 574638 42176 574642
rect 42112 574582 42124 574638
rect 42124 574582 42176 574638
rect 42112 574578 42176 574582
rect 41536 574430 41600 574494
rect 41728 574046 41792 574050
rect 41728 573990 41780 574046
rect 41780 573990 41792 574046
rect 41728 573986 41792 573990
rect 40576 573098 40640 573162
rect 40768 570434 40832 570498
rect 41536 564958 41600 565022
rect 41728 564958 41792 565022
rect 674368 562590 674432 562654
rect 675520 561762 675584 561766
rect 675520 561706 675532 561762
rect 675532 561706 675584 561762
rect 675520 561702 675584 561706
rect 675136 561406 675200 561470
rect 40192 559038 40256 559102
rect 674944 558890 675008 558954
rect 40192 556818 40256 556882
rect 40768 554598 40832 554662
rect 676864 554450 676928 554514
rect 40960 552378 41024 552442
rect 42688 544534 42752 544598
rect 42112 544386 42176 544450
rect 42880 541574 42944 541638
rect 43072 541426 43136 541490
rect 41344 541338 41408 541342
rect 41344 541282 41396 541338
rect 41396 541282 41408 541338
rect 41344 541278 41408 541282
rect 41728 541338 41792 541342
rect 41728 541282 41740 541338
rect 41740 541282 41792 541338
rect 41728 541278 41792 541282
rect 41920 541130 41984 541194
rect 42304 540982 42368 541046
rect 42304 538022 42368 538086
rect 42880 536986 42944 537050
rect 677248 534914 677312 534978
rect 677056 534470 677120 534534
rect 41728 534382 41792 534386
rect 41728 534326 41780 534382
rect 41780 534326 41792 534382
rect 41728 534322 41792 534326
rect 675328 533878 675392 533942
rect 41920 533790 41984 533794
rect 41920 533734 41972 533790
rect 41972 533734 41984 533790
rect 41920 533730 41984 533734
rect 676672 533434 676736 533498
rect 42112 532754 42176 532758
rect 42112 532698 42124 532754
rect 42124 532698 42176 532754
rect 42112 532694 42176 532698
rect 40960 532546 41024 532610
rect 674176 532546 674240 532610
rect 674560 532250 674624 532314
rect 41728 531866 41792 531870
rect 41728 531810 41780 531866
rect 41780 531810 41792 531866
rect 41728 531806 41792 531810
rect 675904 531806 675968 531870
rect 41344 531214 41408 531278
rect 676480 531214 676544 531278
rect 674752 530622 674816 530686
rect 40768 530030 40832 530094
rect 43072 529438 43136 529502
rect 42304 509902 42368 509966
rect 42112 504042 42176 504046
rect 42112 503986 42164 504042
rect 42164 503986 42176 504042
rect 42112 503982 42176 503986
rect 675136 489922 675200 489986
rect 42112 489626 42176 489690
rect 42304 489330 42368 489394
rect 674368 488590 674432 488654
rect 675520 486666 675584 486730
rect 674944 486074 675008 486138
rect 42304 483706 42368 483770
rect 676864 483410 676928 483474
rect 42112 463726 42176 463790
rect 40384 429242 40448 429306
rect 40576 428650 40640 428714
rect 40768 428058 40832 428122
rect 40960 427022 41024 427086
rect 41344 426430 41408 426494
rect 42112 425986 42176 426050
rect 41152 424802 41216 424866
rect 41536 424358 41600 424422
rect 42304 409262 42368 409326
rect 41920 408966 41984 409030
rect 42496 408966 42560 409030
rect 41920 408818 41984 408882
rect 42496 408818 42560 408882
rect 42304 408138 42368 408142
rect 42304 408082 42356 408138
rect 42356 408082 42368 408138
rect 42304 408078 42368 408082
rect 42112 406066 42176 406070
rect 42112 406010 42124 406066
rect 42124 406010 42176 406066
rect 42112 406006 42176 406010
rect 42112 404290 42176 404294
rect 42112 404234 42124 404290
rect 42124 404234 42176 404290
rect 42112 404230 42176 404234
rect 41728 403846 41792 403850
rect 41728 403790 41780 403846
rect 41780 403790 41792 403846
rect 41728 403786 41792 403790
rect 41536 402602 41600 402666
rect 41344 401862 41408 401926
rect 674560 400530 674624 400594
rect 40768 400086 40832 400150
rect 41152 399494 41216 399558
rect 674368 399198 674432 399262
rect 40960 398754 41024 398818
rect 674176 398754 674240 398818
rect 40384 386026 40448 386090
rect 40576 386026 40640 386090
rect 40768 384842 40832 384906
rect 40960 383806 41024 383870
rect 41344 383214 41408 383278
rect 41536 382770 41600 382834
rect 41152 381586 41216 381650
rect 42112 381142 42176 381206
rect 42304 380106 42368 380170
rect 42880 380106 42944 380170
rect 42496 378922 42560 378986
rect 674368 378774 674432 378838
rect 675328 374482 675392 374546
rect 676864 374334 676928 374398
rect 675520 374038 675584 374102
rect 674560 373890 674624 373954
rect 677056 373298 677120 373362
rect 674176 371966 674240 372030
rect 42112 368710 42176 368774
rect 42112 368414 42176 368478
rect 41536 362790 41600 362854
rect 42304 361902 42368 361966
rect 42880 361902 42944 361966
rect 42496 361162 42560 361226
rect 41728 360570 41792 360634
rect 42880 360570 42944 360634
rect 42112 359446 42176 359450
rect 42112 359390 42124 359446
rect 42124 359390 42176 359446
rect 42112 359386 42176 359390
rect 41344 358646 41408 358710
rect 677056 357610 677120 357674
rect 677440 357610 677504 357674
rect 676864 357018 676928 357082
rect 40768 356870 40832 356934
rect 677248 356574 677312 356638
rect 41152 356426 41216 356490
rect 674176 355686 674240 355750
rect 40960 355538 41024 355602
rect 676672 345178 676736 345242
rect 676480 344142 676544 344206
rect 40384 342958 40448 343022
rect 40576 342810 40640 342874
rect 40768 341774 40832 341838
rect 40960 340590 41024 340654
rect 41344 340146 41408 340210
rect 42112 339554 42176 339618
rect 41152 338518 41216 338582
rect 41536 337926 41600 337990
rect 42688 336002 42752 336066
rect 41728 335114 41792 335178
rect 675328 335026 675392 335030
rect 675328 334970 675340 335026
rect 675340 334970 675392 335026
rect 675328 334966 675392 334970
rect 675520 334582 675584 334586
rect 675520 334526 675532 334582
rect 675532 334526 675584 334582
rect 675520 334522 675584 334526
rect 673984 331118 674048 331182
rect 676480 330526 676544 330590
rect 675328 329490 675392 329554
rect 674176 328306 674240 328370
rect 676672 326826 676736 326890
rect 42688 324754 42752 324818
rect 41728 320522 41792 320526
rect 41728 320466 41780 320522
rect 41780 320466 41792 320522
rect 41728 320462 41792 320466
rect 42112 319782 42176 319786
rect 42112 319726 42124 319782
rect 42124 319726 42176 319782
rect 42112 319722 42176 319726
rect 41728 318390 41792 318454
rect 42496 318390 42560 318454
rect 41920 317946 41984 318010
rect 42880 317946 42944 318010
rect 41536 316170 41600 316234
rect 41344 315430 41408 315494
rect 40768 313654 40832 313718
rect 677056 313654 677120 313718
rect 41152 313210 41216 313274
rect 677248 312470 677312 312534
rect 40960 312322 41024 312386
rect 677440 312026 677504 312090
rect 677056 311434 677120 311498
rect 674176 310694 674240 310758
rect 40384 299742 40448 299806
rect 40576 299594 40640 299658
rect 42304 299594 42368 299658
rect 675904 299446 675968 299510
rect 676672 299298 676736 299362
rect 40960 298558 41024 298622
rect 40768 297374 40832 297438
rect 41344 296930 41408 296994
rect 42112 296486 42176 296550
rect 41152 295302 41216 295366
rect 41536 294710 41600 294774
rect 42688 291750 42752 291814
rect 675328 290034 675392 290038
rect 675328 289978 675340 290034
rect 675340 289978 675392 290034
rect 675328 289974 675392 289978
rect 673984 289590 674048 289594
rect 673984 289534 673996 289590
rect 673996 289534 674048 289590
rect 673984 289530 674048 289534
rect 674368 284942 674432 285006
rect 42496 284794 42560 284858
rect 675904 284794 675968 284858
rect 673984 284706 674048 284710
rect 673984 284650 673996 284706
rect 673996 284650 674048 284706
rect 673984 284646 674048 284650
rect 674176 283610 674240 283674
rect 676672 281834 676736 281898
rect 42496 281538 42560 281602
rect 42688 278578 42752 278642
rect 590272 278430 590336 278494
rect 604864 278430 604928 278494
rect 590464 278282 590528 278346
rect 604864 278282 604928 278346
rect 645184 278282 645248 278346
rect 645184 278134 645248 278198
rect 42112 276566 42176 276570
rect 42112 276510 42124 276566
rect 42124 276510 42176 276566
rect 42112 276506 42176 276510
rect 41920 274790 41984 274794
rect 41920 274734 41972 274790
rect 41972 274734 41984 274790
rect 41920 274730 41984 274734
rect 41728 274582 41792 274646
rect 42880 274582 42944 274646
rect 477952 273694 478016 273758
rect 407488 273398 407552 273462
rect 477952 273398 478016 273462
rect 409024 273102 409088 273166
rect 41536 272954 41600 273018
rect 410560 272954 410624 273018
rect 411136 272658 411200 272722
rect 41344 272214 41408 272278
rect 409792 272214 409856 272278
rect 408064 271918 408128 271982
rect 406144 271770 406208 271834
rect 406720 271474 406784 271538
rect 409984 272066 410048 272130
rect 410368 271770 410432 271834
rect 410176 271622 410240 271686
rect 410752 271474 410816 271538
rect 328192 271326 328256 271390
rect 381760 271178 381824 271242
rect 406912 271178 406976 271242
rect 409408 271178 409472 271242
rect 407872 271030 407936 271094
rect 328576 270882 328640 270946
rect 406336 270882 406400 270946
rect 394048 270734 394112 270798
rect 395776 270734 395840 270798
rect 406528 270734 406592 270798
rect 40960 270586 41024 270650
rect 41920 270586 41984 270650
rect 370624 270498 370688 270502
rect 370624 270442 370676 270498
rect 370676 270442 370688 270498
rect 370624 270438 370688 270442
rect 371200 270438 371264 270502
rect 371584 270438 371648 270502
rect 499648 270290 499712 270354
rect 41152 269994 41216 270058
rect 40768 269106 40832 269170
rect 380032 269018 380096 269022
rect 380032 268962 380044 269018
rect 380044 268962 380096 269018
rect 380032 268958 380096 268962
rect 499456 268662 499520 268726
rect 677248 268662 677312 268726
rect 276352 268514 276416 268578
rect 377344 268218 377408 268282
rect 404608 268218 404672 268282
rect 405568 268218 405632 268282
rect 405952 268218 406016 268282
rect 327232 267922 327296 267986
rect 329152 267922 329216 267986
rect 276352 267626 276416 267690
rect 328768 267626 328832 267690
rect 352768 267626 352832 267690
rect 370816 267626 370880 267690
rect 371200 267774 371264 267838
rect 377152 267774 377216 267838
rect 389056 267834 389120 267838
rect 389056 267778 389068 267834
rect 389068 267778 389120 267834
rect 389056 267774 389120 267778
rect 389440 267626 389504 267690
rect 677248 267626 677312 267690
rect 677440 267478 677504 267542
rect 676864 267034 676928 267098
rect 677056 267034 677120 267098
rect 407104 264814 407168 264878
rect 407104 264518 407168 264582
rect 407680 264855 407732 264878
rect 407732 264855 407744 264878
rect 407680 264814 407744 264855
rect 408256 264814 408320 264878
rect 409600 264855 409612 264878
rect 409612 264855 409664 264878
rect 409600 264814 409664 264855
rect 408448 264666 408512 264730
rect 410944 264814 411008 264878
rect 411328 264666 411392 264730
rect 674176 264074 674240 264138
rect 40384 256970 40448 257034
rect 42304 256378 42368 256442
rect 40576 255342 40640 255406
rect 40384 254158 40448 254222
rect 40768 253714 40832 253778
rect 41344 253270 41408 253334
rect 675712 253270 675776 253334
rect 675904 253122 675968 253186
rect 40960 252086 41024 252150
rect 41152 251494 41216 251558
rect 41536 251050 41600 251114
rect 405952 247498 406016 247562
rect 407680 247794 407744 247858
rect 408448 247646 408512 247710
rect 410944 247646 411008 247710
rect 181312 247114 181376 247118
rect 181312 247058 181364 247114
rect 181364 247058 181376 247114
rect 181312 247054 181376 247058
rect 207232 247054 207296 247118
rect 42880 246462 42944 246526
rect 409600 247350 409664 247414
rect 207232 246610 207296 246674
rect 181312 245930 181376 245934
rect 181312 245874 181364 245930
rect 181364 245874 181376 245930
rect 181312 245870 181376 245874
rect 407872 247202 407936 247266
rect 408640 247202 408704 247266
rect 410752 247202 410816 247266
rect 407104 247054 407168 247118
rect 405568 246906 405632 246970
rect 406720 246906 406784 246970
rect 406912 246906 406976 246970
rect 406144 246818 406208 246822
rect 406144 246762 406156 246818
rect 406156 246762 406208 246818
rect 406144 246758 406208 246762
rect 406528 246781 406592 246822
rect 406528 246758 406580 246781
rect 406580 246758 406592 246781
rect 406720 246818 406784 246822
rect 406720 246762 406772 246818
rect 406772 246762 406784 246818
rect 406720 246758 406784 246762
rect 407488 246758 407552 246822
rect 408448 247054 408512 247118
rect 409792 247054 409856 247118
rect 409408 246906 409472 246970
rect 410176 246906 410240 246970
rect 408640 246758 408704 246822
rect 409984 246758 410048 246822
rect 410368 246818 410432 246822
rect 410368 246762 410380 246818
rect 410380 246762 410432 246818
rect 410368 246758 410432 246762
rect 411136 246906 411200 246970
rect 410944 246758 411008 246822
rect 411328 246818 411392 246822
rect 411328 246762 411380 246818
rect 411380 246762 411392 246818
rect 411328 246758 411392 246762
rect 673984 246758 674048 246822
rect 673984 245278 674048 245342
rect 674368 244686 674432 244750
rect 675328 244746 675392 244750
rect 675328 244690 675380 244746
rect 675380 244690 675392 244746
rect 675328 244686 675392 244690
rect 41728 243798 41792 243862
rect 674368 243798 674432 243862
rect 210304 243650 210368 243714
rect 210496 243710 210560 243714
rect 210496 243654 210508 243710
rect 210508 243654 210560 243710
rect 210496 243650 210560 243654
rect 268096 243650 268160 243714
rect 405760 243502 405824 243566
rect 405952 243562 406016 243566
rect 405952 243506 406004 243562
rect 406004 243506 406016 243562
rect 405952 243502 406016 243506
rect 674176 243502 674240 243566
rect 408256 243354 408320 243418
rect 210688 243206 210752 243270
rect 210880 243058 210944 243122
rect 267904 243206 267968 243270
rect 268288 243058 268352 243122
rect 41920 242910 41984 242974
rect 42880 242910 42944 242974
rect 268096 242910 268160 242974
rect 288064 243058 288128 243122
rect 409024 243206 409088 243270
rect 408064 243058 408128 243122
rect 227392 242762 227456 242826
rect 115264 242614 115328 242678
rect 175552 242614 175616 242678
rect 115264 242466 115328 242530
rect 247360 242526 247424 242530
rect 247360 242470 247372 242526
rect 247372 242470 247424 242526
rect 247360 242466 247424 242470
rect 175552 242318 175616 242382
rect 227968 242318 228032 242382
rect 268096 241726 268160 241790
rect 287872 241726 287936 241790
rect 247744 241430 247808 241494
rect 267520 241430 267584 241494
rect 42304 240750 42368 240754
rect 42304 240694 42316 240750
rect 42316 240694 42368 240750
rect 42304 240690 42368 240694
rect 145408 239802 145472 239866
rect 675520 238914 675584 238978
rect 675904 238618 675968 238682
rect 211072 237730 211136 237794
rect 677056 237730 677120 237794
rect 676864 237582 676928 237646
rect 210880 236694 210944 236758
rect 42304 236606 42368 236610
rect 42304 236550 42356 236606
rect 42356 236550 42368 236606
rect 42304 236546 42368 236550
rect 210688 236546 210752 236610
rect 210496 236398 210560 236462
rect 675712 236902 675776 236906
rect 675712 236846 675764 236902
rect 675764 236846 675776 236902
rect 675712 236842 675776 236846
rect 302464 236546 302528 236610
rect 302848 236546 302912 236610
rect 210304 236250 210368 236314
rect 211456 234622 211520 234686
rect 636928 234030 636992 234094
rect 637888 233942 637952 233946
rect 637888 233886 637940 233942
rect 637940 233886 637952 233942
rect 637888 233882 637952 233886
rect 637504 233734 637568 233798
rect 212416 233586 212480 233650
rect 637120 233646 637184 233650
rect 637120 233590 637172 233646
rect 637172 233590 637184 233646
rect 637120 233586 637184 233590
rect 637312 233586 637376 233650
rect 212224 233438 212288 233502
rect 212608 233498 212672 233502
rect 212608 233442 212620 233498
rect 212620 233442 212672 233498
rect 212608 233438 212672 233442
rect 212800 233498 212864 233502
rect 212800 233442 212852 233498
rect 212852 233442 212864 233498
rect 212800 233438 212864 233442
rect 41344 233290 41408 233354
rect 210880 233290 210944 233354
rect 637696 233438 637760 233502
rect 41920 231722 41984 231726
rect 41920 231666 41972 231722
rect 41972 231666 41984 231722
rect 41920 231662 41984 231666
rect 41728 231130 41792 231134
rect 41728 231074 41780 231130
rect 41780 231074 41792 231130
rect 41728 231070 41792 231074
rect 41536 230330 41600 230394
rect 41152 229590 41216 229654
rect 40768 228998 40832 229062
rect 40576 227370 40640 227434
rect 40960 226778 41024 226842
rect 40384 225890 40448 225954
rect 677248 223522 677312 223586
rect 676864 222338 676928 222402
rect 677248 222338 677312 222402
rect 677056 221746 677120 221810
rect 677632 221746 677696 221810
rect 674368 220488 674432 220552
rect 145600 218934 145664 218998
rect 674176 218860 674240 218924
rect 210496 217010 210560 217074
rect 211072 217010 211136 217074
rect 145792 216418 145856 216482
rect 40576 212126 40640 212190
rect 40384 211090 40448 211154
rect 40960 210498 41024 210562
rect 676480 210202 676544 210266
rect 676672 210054 676736 210118
rect 40768 208870 40832 208934
rect 41152 208278 41216 208342
rect 676864 206354 676928 206418
rect 677632 206354 677696 206418
rect 42112 201174 42176 201238
rect 675328 199310 675392 199314
rect 675328 199254 675380 199310
rect 675380 199254 675392 199310
rect 675328 199250 675392 199254
rect 675520 198718 675584 198722
rect 675520 198662 675532 198718
rect 675532 198662 675584 198718
rect 675520 198658 675584 198662
rect 674176 198362 674240 198426
rect 42304 197474 42368 197538
rect 42304 195166 42368 195170
rect 42304 195110 42356 195166
rect 42356 195110 42368 195166
rect 42304 195106 42368 195110
rect 676480 195254 676544 195318
rect 674368 193478 674432 193542
rect 210496 191554 210560 191618
rect 211072 191554 211136 191618
rect 676672 191554 676736 191618
rect 42112 190282 42176 190286
rect 42112 190226 42124 190282
rect 42124 190226 42176 190282
rect 42112 190222 42176 190226
rect 41920 189098 41984 189102
rect 41920 189042 41972 189098
rect 41972 189042 41984 189098
rect 41920 189038 41984 189042
rect 41728 188358 41792 188362
rect 41728 188302 41780 188358
rect 41780 188302 41792 188358
rect 41728 188298 41792 188302
rect 41152 186670 41216 186734
rect 40960 185782 41024 185846
rect 40576 184154 40640 184218
rect 40768 183562 40832 183626
rect 40384 182822 40448 182886
rect 677248 178382 677312 178446
rect 676864 177346 676928 177410
rect 677248 177346 677312 177410
rect 677440 176902 677504 176966
rect 677056 176310 677120 176374
rect 674368 173794 674432 173858
rect 674560 170834 674624 170898
rect 673984 170538 674048 170602
rect 211072 161510 211136 161574
rect 675712 161510 675776 161574
rect 676672 161362 676736 161426
rect 210496 158402 210560 158466
rect 675328 155206 675392 155210
rect 675328 155150 675340 155206
rect 675340 155150 675392 155206
rect 675328 155146 675392 155150
rect 675520 154466 675584 154470
rect 675520 154410 675532 154466
rect 675532 154410 675584 154466
rect 675520 154406 675584 154410
rect 674368 153370 674432 153434
rect 673984 151890 674048 151954
rect 674560 150262 674624 150326
rect 675712 148546 675776 148550
rect 675712 148490 675764 148546
rect 675764 148490 675776 148546
rect 675712 148486 675776 148490
rect 676672 146562 676736 146626
rect 210880 141530 210944 141594
rect 210496 141382 210560 141446
rect 210880 141234 210944 141298
rect 210688 138274 210752 138338
rect 677248 133390 677312 133454
rect 677440 132206 677504 132270
rect 677056 131762 677120 131826
rect 210880 129098 210944 129162
rect 673984 128654 674048 128718
rect 210496 126138 210560 126202
rect 674176 125990 674240 126054
rect 211072 121106 211136 121170
rect 210496 117998 210560 118062
rect 210880 117998 210944 118062
rect 676672 117998 676736 118062
rect 675904 117850 675968 117914
rect 211072 113706 211136 113770
rect 210688 112226 210752 112290
rect 211072 112226 211136 112290
rect 675328 110066 675392 110070
rect 675328 110010 675380 110066
rect 675380 110010 675392 110066
rect 675328 110006 675392 110010
rect 675520 109326 675584 109330
rect 675520 109270 675532 109326
rect 675532 109270 675584 109326
rect 675520 109266 675584 109270
rect 673984 108082 674048 108146
rect 674176 105122 674240 105186
rect 675904 103198 675968 103262
rect 676672 101422 676736 101486
rect 210112 86918 210176 86982
rect 210688 86474 210752 86538
rect 210880 86474 210944 86538
rect 210112 77802 210176 77806
rect 210112 77746 210164 77802
rect 210164 77746 210176 77802
rect 210112 77742 210176 77746
rect 210880 58206 210944 58270
rect 210688 57614 210752 57678
rect 211264 54210 211328 54274
rect 210688 54122 210752 54126
rect 210688 54066 210740 54122
rect 210740 54066 210752 54122
rect 210688 54062 210752 54066
rect 212608 54062 212672 54126
rect 210880 53914 210944 53978
rect 211072 53766 211136 53830
rect 212032 53618 212096 53682
rect 211840 53470 211904 53534
rect 212416 53322 212480 53386
rect 212800 53174 212864 53238
rect 637696 52286 637760 52350
rect 637888 52138 637952 52202
rect 637504 51990 637568 52054
rect 637312 51842 637376 51906
rect 636928 51694 636992 51758
rect 145408 51546 145472 51610
rect 145600 51398 145664 51462
rect 145792 51250 145856 51314
rect 637120 50362 637184 50426
rect 520384 49030 520448 49094
rect 302464 45182 302528 45246
rect 362944 45034 363008 45098
rect 527104 44886 527168 44950
rect 302464 43318 302528 43322
rect 302464 43262 302516 43318
rect 302516 43262 302528 43318
rect 302464 43258 302528 43262
rect 362944 43258 363008 43322
rect 527104 43258 527168 43322
rect 520384 42134 520448 42138
rect 520384 42078 520436 42134
rect 520436 42078 520448 42134
rect 520384 42074 520448 42078
rect 189952 41778 190016 41842
rect 194944 41778 195008 41842
rect 189952 40742 190016 40806
rect 194944 40594 195008 40658
<< metal4 >>
rect 528255 996146 528321 996147
rect 528255 996082 528256 996146
rect 528320 996082 528321 996146
rect 528255 996081 528321 996082
rect 528258 995555 528318 996081
rect 528255 995554 528321 995555
rect 528255 995490 528256 995554
rect 528320 995490 528321 995554
rect 528255 995489 528321 995490
rect 42303 968766 42369 968767
rect 42303 968702 42304 968766
rect 42368 968702 42369 968766
rect 42303 968701 42369 968702
rect 41727 967138 41793 967139
rect 41727 967074 41728 967138
rect 41792 967074 41793 967138
rect 41727 967073 41793 967074
rect 40767 965066 40833 965067
rect 40767 965002 40768 965066
rect 40832 965002 40833 965066
rect 40767 965001 40833 965002
rect 40383 962254 40449 962255
rect 40383 962190 40384 962254
rect 40448 962190 40449 962254
rect 40383 962189 40449 962190
rect 40386 941831 40446 962189
rect 40575 958554 40641 958555
rect 40575 958490 40576 958554
rect 40640 958490 40641 958554
rect 40575 958489 40641 958490
rect 40383 941830 40449 941831
rect 40383 941766 40384 941830
rect 40448 941766 40449 941830
rect 40383 941765 40449 941766
rect 40383 941386 40449 941387
rect 40383 941322 40384 941386
rect 40448 941322 40449 941386
rect 40383 941321 40449 941322
rect 40386 816031 40446 941321
rect 40578 937687 40638 958489
rect 40575 937686 40641 937687
rect 40575 937622 40576 937686
rect 40640 937622 40641 937686
rect 40575 937621 40641 937622
rect 40770 936503 40830 965001
rect 40959 963438 41025 963439
rect 40959 963374 40960 963438
rect 41024 963374 41025 963438
rect 40959 963373 41025 963374
rect 40767 936502 40833 936503
rect 40767 936438 40768 936502
rect 40832 936438 40833 936502
rect 40767 936437 40833 936438
rect 40962 935911 41022 963373
rect 41151 962698 41217 962699
rect 41151 962634 41152 962698
rect 41216 962634 41217 962698
rect 41151 962633 41217 962634
rect 40959 935910 41025 935911
rect 40959 935846 40960 935910
rect 41024 935846 41025 935910
rect 40959 935845 41025 935846
rect 41154 934875 41214 962633
rect 41535 959738 41601 959739
rect 41535 959674 41536 959738
rect 41600 959674 41601 959738
rect 41535 959673 41601 959674
rect 41538 935467 41598 959673
rect 41730 940943 41790 967073
rect 41919 959146 41985 959147
rect 41919 959082 41920 959146
rect 41984 959082 41985 959146
rect 41919 959081 41985 959082
rect 41727 940942 41793 940943
rect 41727 940878 41728 940942
rect 41792 940878 41793 940942
rect 41727 940877 41793 940878
rect 41922 937095 41982 959081
rect 42111 956186 42177 956187
rect 42111 956122 42112 956186
rect 42176 956122 42177 956186
rect 42111 956121 42177 956122
rect 42114 941387 42174 956121
rect 42111 941386 42177 941387
rect 42111 941322 42112 941386
rect 42176 941322 42177 941386
rect 42111 941321 42177 941322
rect 42306 938723 42366 968701
rect 676671 965806 676737 965807
rect 676671 965742 676672 965806
rect 676736 965742 676737 965806
rect 676671 965741 676737 965742
rect 674559 965066 674625 965067
rect 674559 965002 674560 965066
rect 674624 965002 674625 965066
rect 674559 965001 674625 965002
rect 42495 964030 42561 964031
rect 42495 963966 42496 964030
rect 42560 963966 42561 964030
rect 42495 963965 42561 963966
rect 42303 938722 42369 938723
rect 42303 938658 42304 938722
rect 42368 938658 42369 938722
rect 42303 938657 42369 938658
rect 41919 937094 41985 937095
rect 41919 937030 41920 937094
rect 41984 937030 41985 937094
rect 41919 937029 41985 937030
rect 41535 935466 41601 935467
rect 41535 935402 41536 935466
rect 41600 935402 41601 935466
rect 41535 935401 41601 935402
rect 41151 934874 41217 934875
rect 41151 934810 41152 934874
rect 41216 934810 41217 934874
rect 41151 934809 41217 934810
rect 42498 934431 42558 963965
rect 43071 962402 43137 962403
rect 43071 962338 43072 962402
rect 43136 962338 43137 962402
rect 43071 962337 43137 962338
rect 42879 962106 42945 962107
rect 42879 962042 42880 962106
rect 42944 962042 42945 962106
rect 42879 962041 42945 962042
rect 42687 957814 42753 957815
rect 42687 957750 42688 957814
rect 42752 957750 42753 957814
rect 42687 957749 42753 957750
rect 42690 939463 42750 957749
rect 42687 939462 42753 939463
rect 42687 939398 42688 939462
rect 42752 939398 42753 939462
rect 42687 939397 42753 939398
rect 42495 934430 42561 934431
rect 42495 934366 42496 934430
rect 42560 934366 42561 934430
rect 42495 934365 42561 934366
rect 40383 816030 40449 816031
rect 40383 815966 40384 816030
rect 40448 815966 40449 816030
rect 40383 815965 40449 815966
rect 41151 816030 41217 816031
rect 41151 815966 41152 816030
rect 41216 815966 41217 816030
rect 41151 815965 41217 815966
rect 40959 801970 41025 801971
rect 40959 801906 40960 801970
rect 41024 801906 41025 801970
rect 40959 801905 41025 801906
rect 40962 796051 41022 801905
rect 40959 796050 41025 796051
rect 40959 795986 40960 796050
rect 41024 795986 41025 796050
rect 40959 795985 41025 795986
rect 41154 773555 41214 815965
rect 41343 815586 41409 815587
rect 41343 815522 41344 815586
rect 41408 815522 41409 815586
rect 41343 815521 41409 815522
rect 41151 773554 41217 773555
rect 41151 773490 41152 773554
rect 41216 773490 41217 773554
rect 41151 773489 41217 773490
rect 41346 772815 41406 815521
rect 41535 802118 41601 802119
rect 41535 802054 41536 802118
rect 41600 802054 41601 802118
rect 41535 802053 41601 802054
rect 41538 789391 41598 802053
rect 42882 801561 42942 962041
rect 42690 801501 42942 801561
rect 41919 800638 41985 800639
rect 41919 800574 41920 800638
rect 41984 800574 41985 800638
rect 41919 800573 41985 800574
rect 41727 800342 41793 800343
rect 41727 800278 41728 800342
rect 41792 800278 41793 800342
rect 41727 800277 41793 800278
rect 41730 793831 41790 800277
rect 41922 796199 41982 800573
rect 42495 800490 42561 800491
rect 42495 800426 42496 800490
rect 42560 800426 42561 800490
rect 42495 800425 42561 800426
rect 42111 800342 42177 800343
rect 42111 800278 42112 800342
rect 42176 800278 42177 800342
rect 42111 800277 42177 800278
rect 41919 796198 41985 796199
rect 41919 796134 41920 796198
rect 41984 796134 41985 796198
rect 41919 796133 41985 796134
rect 41919 796050 41985 796051
rect 41919 795986 41920 796050
rect 41984 795986 41985 796050
rect 41919 795985 41985 795986
rect 41727 793830 41793 793831
rect 41727 793766 41728 793830
rect 41792 793766 41793 793830
rect 41727 793765 41793 793766
rect 41727 790574 41793 790575
rect 41727 790510 41728 790574
rect 41792 790510 41793 790574
rect 41727 790509 41793 790510
rect 41535 789390 41601 789391
rect 41535 789326 41536 789390
rect 41600 789326 41601 789390
rect 41535 789325 41601 789326
rect 41535 772962 41601 772963
rect 41535 772898 41536 772962
rect 41600 772898 41601 772962
rect 41535 772897 41601 772898
rect 41343 772814 41409 772815
rect 41343 772750 41344 772814
rect 41408 772750 41409 772814
rect 41343 772749 41409 772750
rect 40959 768670 41025 768671
rect 40959 768606 40960 768670
rect 41024 768606 41025 768670
rect 40959 768605 41025 768606
rect 40962 747063 41022 768605
rect 41151 757718 41217 757719
rect 41151 757654 41152 757718
rect 41216 757654 41217 757718
rect 41151 757653 41217 757654
rect 40959 747062 41025 747063
rect 40959 746998 40960 747062
rect 41024 746998 41025 747062
rect 40959 746997 41025 746998
rect 41154 746915 41214 757653
rect 41151 746914 41217 746915
rect 41151 746850 41152 746914
rect 41216 746850 41217 746914
rect 41151 746849 41217 746850
rect 41346 734335 41406 772749
rect 41343 734334 41409 734335
rect 41343 734270 41344 734334
rect 41408 734270 41409 734334
rect 41343 734269 41409 734270
rect 41538 729633 41598 772897
rect 41730 747211 41790 790509
rect 41922 789243 41982 795985
rect 42114 794275 42174 800277
rect 42111 794274 42177 794275
rect 42111 794210 42112 794274
rect 42176 794210 42177 794274
rect 42111 794209 42177 794210
rect 42111 792202 42177 792203
rect 42111 792138 42112 792202
rect 42176 792138 42177 792202
rect 42111 792137 42177 792138
rect 42114 791907 42174 792137
rect 42111 791906 42177 791907
rect 42111 791842 42112 791906
rect 42176 791842 42177 791906
rect 42111 791841 42177 791842
rect 42498 791759 42558 800425
rect 42495 791758 42561 791759
rect 42495 791694 42496 791758
rect 42560 791694 42561 791758
rect 42495 791693 42561 791694
rect 42111 791166 42177 791167
rect 42111 791102 42112 791166
rect 42176 791102 42177 791166
rect 42111 791101 42177 791102
rect 41919 789242 41985 789243
rect 41919 789178 41920 789242
rect 41984 789178 41985 789242
rect 41919 789177 41985 789178
rect 42114 772812 42174 791101
rect 42690 790575 42750 801501
rect 42879 800786 42945 800787
rect 42879 800722 42880 800786
rect 42944 800722 42945 800786
rect 42879 800721 42945 800722
rect 42882 791907 42942 800721
rect 42879 791906 42945 791907
rect 42879 791842 42880 791906
rect 42944 791842 42945 791906
rect 42879 791841 42945 791842
rect 43074 791167 43134 962337
rect 673983 962254 674049 962255
rect 673983 962190 673984 962254
rect 674048 962190 674049 962254
rect 673983 962189 674049 962190
rect 673986 933395 674046 962189
rect 674367 959294 674433 959295
rect 674367 959230 674368 959294
rect 674432 959230 674433 959294
rect 674367 959229 674433 959230
rect 673983 933394 674049 933395
rect 673983 933330 673984 933394
rect 674048 933330 674049 933394
rect 673983 933329 674049 933330
rect 674175 877006 674241 877007
rect 674175 876942 674176 877006
rect 674240 876942 674241 877006
rect 674175 876941 674241 876942
rect 43071 791166 43137 791167
rect 43071 791102 43072 791166
rect 43136 791102 43137 791166
rect 43071 791101 43137 791102
rect 42687 790574 42753 790575
rect 42687 790510 42688 790574
rect 42752 790510 42753 790574
rect 42687 790509 42753 790510
rect 673983 788058 674049 788059
rect 673983 787994 673984 788058
rect 674048 787994 674049 788058
rect 673983 787993 674049 787994
rect 42114 772752 42366 772812
rect 42111 757274 42177 757275
rect 42111 757210 42112 757274
rect 42176 757210 42177 757274
rect 42111 757209 42177 757210
rect 41919 757126 41985 757127
rect 41919 757062 41920 757126
rect 41984 757062 41985 757126
rect 41919 757061 41985 757062
rect 41922 754907 41982 757061
rect 41919 754906 41985 754907
rect 41919 754842 41920 754906
rect 41984 754842 41985 754906
rect 41919 754841 41985 754842
rect 42114 749875 42174 757209
rect 42111 749874 42177 749875
rect 42111 749810 42112 749874
rect 42176 749810 42177 749874
rect 42111 749809 42177 749810
rect 42306 747803 42366 772752
rect 42495 767930 42561 767931
rect 42495 767866 42496 767930
rect 42560 767866 42561 767930
rect 42495 767865 42561 767866
rect 41919 747802 41985 747803
rect 41919 747738 41920 747802
rect 41984 747738 41985 747802
rect 41919 747737 41985 747738
rect 42303 747802 42369 747803
rect 42303 747738 42304 747802
rect 42368 747738 42369 747802
rect 42303 747737 42369 747738
rect 41727 747210 41793 747211
rect 41727 747146 41728 747210
rect 41792 747146 41793 747210
rect 41727 747145 41793 747146
rect 41346 729599 41598 729633
rect 41343 729598 41598 729599
rect 41343 729534 41344 729598
rect 41408 729573 41598 729598
rect 41408 729534 41409 729573
rect 41343 729533 41409 729534
rect 41151 723086 41217 723087
rect 41151 723022 41152 723086
rect 41216 723022 41217 723086
rect 41151 723021 41217 723022
rect 41154 707991 41214 723021
rect 41151 707990 41217 707991
rect 41151 707926 41152 707990
rect 41216 707926 41217 707990
rect 41151 707925 41217 707926
rect 40767 690230 40833 690231
rect 40767 690166 40768 690230
rect 40832 690166 40833 690230
rect 40767 690165 40833 690166
rect 40770 685939 40830 690165
rect 41346 686975 41406 729533
rect 41535 725306 41601 725307
rect 41535 725242 41536 725306
rect 41600 725242 41601 725306
rect 41535 725241 41601 725242
rect 41538 705475 41598 725241
rect 41730 723087 41790 747145
rect 41727 723086 41793 723087
rect 41727 723022 41728 723086
rect 41792 723022 41793 723086
rect 41727 723021 41793 723022
rect 41727 713910 41793 713911
rect 41727 713846 41728 713910
rect 41792 713846 41793 713910
rect 41727 713845 41793 713846
rect 41730 711099 41790 713845
rect 41727 711098 41793 711099
rect 41727 711034 41728 711098
rect 41792 711034 41793 711098
rect 41727 711033 41793 711034
rect 41727 708730 41793 708731
rect 41727 708666 41728 708730
rect 41792 708666 41793 708730
rect 41727 708665 41793 708666
rect 41535 705474 41601 705475
rect 41535 705410 41536 705474
rect 41600 705410 41601 705474
rect 41535 705409 41601 705410
rect 41730 704143 41790 708665
rect 41922 704735 41982 747737
rect 42498 746323 42558 767865
rect 42687 764674 42753 764675
rect 42687 764610 42688 764674
rect 42752 764610 42753 764674
rect 42687 764609 42753 764610
rect 42690 751799 42750 764609
rect 42879 757422 42945 757423
rect 42879 757358 42880 757422
rect 42944 757358 42945 757422
rect 42879 757357 42945 757358
rect 42687 751798 42753 751799
rect 42687 751734 42688 751798
rect 42752 751734 42753 751798
rect 42687 751733 42753 751734
rect 42882 751059 42942 757357
rect 43071 751946 43137 751947
rect 43071 751882 43072 751946
rect 43136 751882 43137 751946
rect 43071 751881 43137 751882
rect 42879 751058 42945 751059
rect 42879 750994 42880 751058
rect 42944 750994 42945 751058
rect 42879 750993 42945 750994
rect 43074 749283 43134 751881
rect 43071 749282 43137 749283
rect 43071 749218 43072 749282
rect 43136 749218 43137 749282
rect 43071 749217 43137 749218
rect 42495 746322 42561 746323
rect 42495 746258 42496 746322
rect 42560 746258 42561 746322
rect 42495 746257 42561 746258
rect 42111 734334 42177 734335
rect 42111 734270 42112 734334
rect 42176 734270 42177 734334
rect 42111 734269 42177 734270
rect 42114 729155 42174 734269
rect 42111 729154 42177 729155
rect 42111 729090 42112 729154
rect 42176 729090 42177 729154
rect 42111 729089 42177 729090
rect 41919 704734 41985 704735
rect 41919 704670 41920 704734
rect 41984 704670 41985 704734
rect 41919 704669 41985 704670
rect 41727 704142 41793 704143
rect 41727 704078 41728 704142
rect 41792 704078 41793 704142
rect 41727 704077 41793 704078
rect 41343 686974 41409 686975
rect 41343 686910 41344 686974
rect 41408 686910 41409 686974
rect 41343 686909 41409 686910
rect 40767 685938 40833 685939
rect 40767 685874 40768 685938
rect 40832 685874 40833 685938
rect 40767 685873 40833 685874
rect 40575 671138 40641 671139
rect 40575 671074 40576 671138
rect 40640 671074 40641 671138
rect 40575 671073 40641 671074
rect 40578 660335 40638 671073
rect 40575 660334 40641 660335
rect 40575 660270 40576 660334
rect 40640 660270 40641 660334
rect 40575 660269 40641 660270
rect 40770 647015 40830 685873
rect 41730 681015 41790 704077
rect 41346 680955 41790 681015
rect 40959 670990 41025 670991
rect 40959 670926 40960 670990
rect 41024 670926 41025 670990
rect 40959 670925 41025 670926
rect 40962 664627 41022 670925
rect 40959 664626 41025 664627
rect 40959 664562 40960 664626
rect 41024 664562 41025 664626
rect 40959 664561 41025 664562
rect 41346 663033 41406 680955
rect 41727 670990 41793 670991
rect 41727 670926 41728 670990
rect 41792 670926 41793 670990
rect 41727 670925 41793 670926
rect 41730 668623 41790 670925
rect 41727 668622 41793 668623
rect 41727 668558 41728 668622
rect 41792 668558 41793 668622
rect 41727 668557 41793 668558
rect 41346 662973 41790 663033
rect 41730 661519 41790 662973
rect 41727 661518 41793 661519
rect 41727 661454 41728 661518
rect 41792 661454 41793 661518
rect 41727 661453 41793 661454
rect 40767 647014 40833 647015
rect 40767 646950 40768 647014
rect 40832 646950 40833 647014
rect 40767 646949 40833 646950
rect 41730 628401 41790 661453
rect 41922 661371 41982 704669
rect 42114 690231 42174 729089
rect 43071 727822 43137 727823
rect 43071 727758 43072 727822
rect 43136 727758 43137 727822
rect 43071 727757 43137 727758
rect 42879 723086 42945 723087
rect 42879 723022 42880 723086
rect 42944 723022 42945 723086
rect 42879 723021 42945 723022
rect 42687 714058 42753 714059
rect 42687 713994 42688 714058
rect 42752 713994 42753 714058
rect 42687 713993 42753 713994
rect 42303 713910 42369 713911
rect 42303 713846 42304 713910
rect 42368 713846 42369 713910
rect 42303 713845 42369 713846
rect 42306 707399 42366 713845
rect 42495 713318 42561 713319
rect 42495 713254 42496 713318
rect 42560 713254 42561 713318
rect 42495 713253 42561 713254
rect 42498 708583 42558 713253
rect 42495 708582 42561 708583
rect 42495 708518 42496 708582
rect 42560 708518 42561 708582
rect 42495 708517 42561 708518
rect 42690 707843 42750 713993
rect 42882 708731 42942 723021
rect 42879 708730 42945 708731
rect 42879 708666 42880 708730
rect 42944 708666 42945 708730
rect 42879 708665 42945 708666
rect 42687 707842 42753 707843
rect 42687 707778 42688 707842
rect 42752 707778 42753 707842
rect 42687 707777 42753 707778
rect 42303 707398 42369 707399
rect 42303 707334 42304 707398
rect 42368 707334 42369 707398
rect 42303 707333 42369 707334
rect 43074 703551 43134 727757
rect 673986 713023 674046 787993
rect 674178 758015 674238 876941
rect 674370 875675 674430 959229
rect 674562 937687 674622 965001
rect 675903 963438 675969 963439
rect 675903 963374 675904 963438
rect 675968 963374 675969 963438
rect 675903 963373 675969 963374
rect 675711 962550 675777 962551
rect 675711 962486 675712 962550
rect 675776 962486 675777 962550
rect 675711 962485 675777 962486
rect 675327 960774 675393 960775
rect 675327 960710 675328 960774
rect 675392 960710 675393 960774
rect 675327 960709 675393 960710
rect 674751 959146 674817 959147
rect 674751 959082 674752 959146
rect 674816 959082 674817 959146
rect 674751 959081 674817 959082
rect 674559 937686 674625 937687
rect 674559 937622 674560 937686
rect 674624 937622 674625 937686
rect 674559 937621 674625 937622
rect 674754 935615 674814 959081
rect 675135 957666 675201 957667
rect 675135 957602 675136 957666
rect 675200 957602 675201 957666
rect 675135 957601 675201 957602
rect 674943 956038 675009 956039
rect 674943 955974 674944 956038
rect 675008 955974 675009 956038
rect 674943 955973 675009 955974
rect 674751 935614 674817 935615
rect 674751 935550 674752 935614
rect 674816 935550 674817 935614
rect 674751 935549 674817 935550
rect 674946 932803 675006 955973
rect 674943 932802 675009 932803
rect 674943 932738 674944 932802
rect 675008 932738 675009 932802
rect 674943 932737 675009 932738
rect 675138 932211 675198 957601
rect 675135 932210 675201 932211
rect 675135 932146 675136 932210
rect 675200 932146 675201 932210
rect 675135 932145 675201 932146
rect 675330 875823 675390 960709
rect 675714 933839 675774 962485
rect 675906 936207 675966 963373
rect 676095 961514 676161 961515
rect 676095 961450 676096 961514
rect 676160 961450 676161 961514
rect 676095 961449 676161 961450
rect 675903 936206 675969 936207
rect 675903 936142 675904 936206
rect 675968 936142 675969 936206
rect 675903 936141 675969 936142
rect 675711 933838 675777 933839
rect 675711 933774 675712 933838
rect 675776 933774 675777 933838
rect 675711 933773 675777 933774
rect 676098 931767 676158 961449
rect 676479 958406 676545 958407
rect 676479 958342 676480 958406
rect 676544 958342 676545 958406
rect 676479 958341 676545 958342
rect 676095 931766 676161 931767
rect 676095 931702 676096 931766
rect 676160 931702 676161 931766
rect 676095 931701 676161 931702
rect 676482 931175 676542 958341
rect 676674 934431 676734 965741
rect 677055 953522 677121 953523
rect 677055 953458 677056 953522
rect 677120 953458 677121 953522
rect 677055 953457 677121 953458
rect 676863 953374 676929 953375
rect 676863 953310 676864 953374
rect 676928 953310 676929 953374
rect 676863 953309 676929 953310
rect 676671 934430 676737 934431
rect 676671 934366 676672 934430
rect 676736 934366 676737 934430
rect 676671 934365 676737 934366
rect 676479 931174 676545 931175
rect 676479 931110 676480 931174
rect 676544 931110 676545 931174
rect 676479 931109 676545 931110
rect 676866 930731 676926 953309
rect 677058 936651 677118 953457
rect 677055 936650 677121 936651
rect 677055 936586 677056 936650
rect 677120 936586 677121 936650
rect 677055 936585 677121 936586
rect 676863 930730 676929 930731
rect 676863 930666 676864 930730
rect 676928 930666 676929 930730
rect 676863 930665 676929 930666
rect 676095 876562 676161 876563
rect 676095 876498 676096 876562
rect 676160 876498 676161 876562
rect 676095 876497 676161 876498
rect 675327 875822 675393 875823
rect 675327 875758 675328 875822
rect 675392 875758 675393 875822
rect 675327 875757 675393 875758
rect 675519 875822 675585 875823
rect 675519 875758 675520 875822
rect 675584 875758 675585 875822
rect 675519 875757 675585 875758
rect 674367 875674 674433 875675
rect 674367 875610 674368 875674
rect 674432 875610 674433 875674
rect 674367 875609 674433 875610
rect 674559 874046 674625 874047
rect 674559 873982 674560 874046
rect 674624 873982 674625 874046
rect 674559 873981 674625 873982
rect 674367 873602 674433 873603
rect 674367 873538 674368 873602
rect 674432 873538 674433 873602
rect 674367 873537 674433 873538
rect 674175 758014 674241 758015
rect 674175 757950 674176 758014
rect 674240 757950 674241 758014
rect 674175 757949 674241 757950
rect 674370 755277 674430 873537
rect 674562 757275 674622 873981
rect 674943 869902 675009 869903
rect 674943 869838 674944 869902
rect 675008 869838 675009 869902
rect 674943 869837 675009 869838
rect 674751 775478 674817 775479
rect 674751 775414 674752 775478
rect 674816 775414 674817 775478
rect 674751 775413 674817 775414
rect 674754 771779 674814 775413
rect 674751 771778 674817 771779
rect 674751 771714 674752 771778
rect 674816 771714 674817 771778
rect 674751 771713 674817 771714
rect 674946 771591 675006 869837
rect 675135 864722 675201 864723
rect 675135 864658 675136 864722
rect 675200 864658 675201 864722
rect 675135 864657 675201 864658
rect 674754 771531 675006 771591
rect 674559 757274 674625 757275
rect 674559 757210 674560 757274
rect 674624 757210 674625 757274
rect 674559 757209 674625 757210
rect 674754 757127 674814 771531
rect 675138 758903 675198 864657
rect 675327 787170 675393 787171
rect 675327 787106 675328 787170
rect 675392 787106 675393 787170
rect 675327 787105 675393 787106
rect 675135 758902 675201 758903
rect 675135 758838 675136 758902
rect 675200 758838 675201 758902
rect 675135 758837 675201 758838
rect 675135 758310 675201 758311
rect 675135 758246 675136 758310
rect 675200 758246 675201 758310
rect 675135 758245 675201 758246
rect 674751 757126 674817 757127
rect 674751 757062 674752 757126
rect 674816 757062 674817 757126
rect 674751 757061 674817 757062
rect 674367 755276 674433 755277
rect 674367 755212 674368 755276
rect 674432 755212 674433 755276
rect 674367 755211 674433 755212
rect 674751 754462 674817 754463
rect 674751 754398 674752 754462
rect 674816 754398 674817 754462
rect 674751 754397 674817 754398
rect 674175 743214 674241 743215
rect 674175 743150 674176 743214
rect 674240 743150 674241 743214
rect 674175 743149 674241 743150
rect 673983 713022 674049 713023
rect 673983 712958 673984 713022
rect 674048 712958 674049 713022
rect 673983 712957 674049 712958
rect 43071 703550 43137 703551
rect 43071 703486 43072 703550
rect 43136 703486 43137 703550
rect 43071 703485 43137 703486
rect 42111 690230 42177 690231
rect 42111 690166 42112 690230
rect 42176 690166 42177 690230
rect 42111 690165 42177 690166
rect 42111 686530 42177 686531
rect 42111 686466 42112 686530
rect 42176 686466 42177 686530
rect 42111 686465 42177 686466
rect 41919 661370 41985 661371
rect 41919 661306 41920 661370
rect 41984 661306 41985 661370
rect 41919 661305 41985 661306
rect 41922 637725 41982 661305
rect 42114 647163 42174 686465
rect 42879 682386 42945 682387
rect 42879 682322 42880 682386
rect 42944 682322 42945 682386
rect 42879 682321 42945 682322
rect 42495 670694 42561 670695
rect 42495 670630 42496 670694
rect 42560 670630 42561 670694
rect 42495 670629 42561 670630
rect 42303 668474 42369 668475
rect 42303 668410 42304 668474
rect 42368 668410 42369 668474
rect 42303 668409 42369 668410
rect 42306 656191 42366 668409
rect 42498 662851 42558 670629
rect 42495 662850 42561 662851
rect 42495 662786 42496 662850
rect 42560 662786 42561 662850
rect 42495 662785 42561 662786
rect 42882 659595 42942 682321
rect 43071 673358 43137 673359
rect 43071 673294 43072 673358
rect 43136 673294 43137 673358
rect 43071 673293 43137 673294
rect 43074 671025 43134 673293
rect 43074 670965 43326 671025
rect 43071 670842 43137 670843
rect 43071 670778 43072 670842
rect 43136 670778 43137 670842
rect 43071 670777 43137 670778
rect 43074 664183 43134 670777
rect 43266 668475 43326 670965
rect 43263 668474 43329 668475
rect 43263 668410 43264 668474
rect 43328 668410 43329 668474
rect 43263 668409 43329 668410
rect 674178 667809 674238 743149
rect 674367 738626 674433 738627
rect 674367 738562 674368 738626
rect 674432 738562 674433 738626
rect 674367 738561 674433 738562
rect 674175 667808 674241 667809
rect 674175 667744 674176 667808
rect 674240 667744 674241 667808
rect 674175 667743 674241 667744
rect 674370 664553 674430 738561
rect 674754 713911 674814 754397
rect 675138 741587 675198 758245
rect 675135 741586 675201 741587
rect 675135 741522 675136 741586
rect 675200 741522 675201 741586
rect 675135 741521 675201 741522
rect 675135 740106 675201 740107
rect 675135 740042 675136 740106
rect 675200 740042 675201 740106
rect 675135 740041 675201 740042
rect 674943 739218 675009 739219
rect 674943 739154 674944 739218
rect 675008 739154 675009 739218
rect 674943 739153 675009 739154
rect 674751 713910 674817 713911
rect 674751 713846 674752 713910
rect 674816 713846 674817 713910
rect 674751 713845 674817 713846
rect 674751 697926 674817 697927
rect 674751 697862 674752 697926
rect 674816 697862 674817 697926
rect 674751 697861 674817 697862
rect 674559 694374 674625 694375
rect 674559 694310 674560 694374
rect 674624 694310 674625 694374
rect 674559 694309 674625 694310
rect 674367 664552 674433 664553
rect 674367 664488 674368 664552
rect 674432 664488 674433 664552
rect 674367 664487 674433 664488
rect 43071 664182 43137 664183
rect 43071 664118 43072 664182
rect 43136 664118 43137 664182
rect 43071 664117 43137 664118
rect 42879 659594 42945 659595
rect 42879 659530 42880 659594
rect 42944 659530 42945 659594
rect 42879 659529 42945 659530
rect 42303 656190 42369 656191
rect 42303 656126 42304 656190
rect 42368 656126 42369 656190
rect 42303 656125 42369 656126
rect 674367 652194 674433 652195
rect 674367 652130 674368 652194
rect 674432 652130 674433 652194
rect 674367 652129 674433 652130
rect 42111 647162 42177 647163
rect 42111 647098 42112 647162
rect 42176 647098 42177 647162
rect 42111 647097 42177 647098
rect 673983 645386 674049 645387
rect 673983 645322 673984 645386
rect 674048 645322 674049 645386
rect 673983 645321 674049 645322
rect 41922 637665 42750 637725
rect 41538 628341 41790 628401
rect 40767 627922 40833 627923
rect 40767 627858 40768 627922
rect 40832 627858 40833 627922
rect 40767 627857 40833 627858
rect 40770 612827 40830 627857
rect 41343 627774 41409 627775
rect 41343 627710 41344 627774
rect 41408 627710 41409 627774
rect 41343 627709 41409 627710
rect 41346 616675 41406 627709
rect 41538 619077 41598 628341
rect 42303 628070 42369 628071
rect 42303 628006 42304 628070
rect 42368 628006 42369 628070
rect 42303 628005 42369 628006
rect 41727 627774 41793 627775
rect 41727 627710 41728 627774
rect 41792 627710 41793 627774
rect 41727 627709 41793 627710
rect 41730 619635 41790 627709
rect 41919 627478 41985 627479
rect 41919 627414 41920 627478
rect 41984 627414 41985 627478
rect 41919 627413 41985 627414
rect 41727 619634 41793 619635
rect 41727 619570 41728 619634
rect 41792 619570 41793 619634
rect 41727 619569 41793 619570
rect 41538 619017 41790 619077
rect 41535 618450 41601 618451
rect 41535 618386 41536 618450
rect 41600 618386 41601 618450
rect 41535 618385 41601 618386
rect 41343 616674 41409 616675
rect 41343 616610 41344 616674
rect 41408 616610 41409 616674
rect 41343 616609 41409 616610
rect 40767 612826 40833 612827
rect 40767 612762 40768 612826
rect 40832 612762 40833 612826
rect 40767 612761 40833 612762
rect 41538 604835 41598 618385
rect 41730 618303 41790 619017
rect 41727 618302 41793 618303
rect 41727 618238 41728 618302
rect 41792 618238 41793 618302
rect 41727 618237 41793 618238
rect 41535 604834 41601 604835
rect 41535 604770 41536 604834
rect 41600 604770 41601 604834
rect 41535 604769 41601 604770
rect 40575 597878 40641 597879
rect 40575 597814 40576 597878
rect 40640 597814 40641 597878
rect 40575 597813 40641 597814
rect 30591 590774 30657 590775
rect 30591 590710 30592 590774
rect 30656 590710 30657 590774
rect 30591 590709 30657 590710
rect 30594 590331 30654 590709
rect 30591 590330 30657 590331
rect 30591 590266 30592 590330
rect 30656 590266 30657 590330
rect 30591 590265 30657 590266
rect 40578 573163 40638 597813
rect 40767 595658 40833 595659
rect 40767 595594 40768 595658
rect 40832 595594 40833 595658
rect 40767 595593 40833 595594
rect 40575 573162 40641 573163
rect 40575 573098 40576 573162
rect 40640 573098 40641 573162
rect 40575 573097 40641 573098
rect 40770 570499 40830 595593
rect 41343 594030 41409 594031
rect 41343 593966 41344 594030
rect 41408 593966 41409 594030
rect 41343 593965 41409 593966
rect 41346 580267 41406 593965
rect 41730 585111 41790 618237
rect 41922 617859 41982 627413
rect 42111 625702 42177 625703
rect 42111 625638 42112 625702
rect 42176 625638 42177 625702
rect 42111 625637 42177 625638
rect 42114 624963 42174 625637
rect 42111 624962 42177 624963
rect 42111 624898 42112 624962
rect 42176 624898 42177 624962
rect 42111 624897 42177 624898
rect 41919 617858 41985 617859
rect 41919 617794 41920 617858
rect 41984 617794 41985 617858
rect 41919 617793 41985 617794
rect 42306 613567 42366 628005
rect 42495 627922 42561 627923
rect 42495 627858 42496 627922
rect 42560 627858 42561 627922
rect 42495 627857 42561 627858
rect 42498 621559 42558 627857
rect 42690 625703 42750 637665
rect 42879 637246 42945 637247
rect 42879 637182 42880 637246
rect 42944 637182 42945 637246
rect 42879 637181 42945 637182
rect 42687 625702 42753 625703
rect 42687 625638 42688 625702
rect 42752 625638 42753 625702
rect 42687 625637 42753 625638
rect 42687 624962 42753 624963
rect 42687 624898 42688 624962
rect 42752 624898 42753 624962
rect 42687 624897 42753 624898
rect 42495 621558 42561 621559
rect 42495 621494 42496 621558
rect 42560 621494 42561 621558
rect 42495 621493 42561 621494
rect 42690 618451 42750 624897
rect 42882 623483 42942 637181
rect 42879 623482 42945 623483
rect 42879 623418 42880 623482
rect 42944 623418 42945 623482
rect 42879 623417 42945 623418
rect 42687 618450 42753 618451
rect 42687 618386 42688 618450
rect 42752 618386 42753 618450
rect 42687 618385 42753 618386
rect 42303 613566 42369 613567
rect 42303 613502 42304 613566
rect 42368 613502 42369 613566
rect 42303 613501 42369 613502
rect 42111 604834 42177 604835
rect 42111 604770 42112 604834
rect 42176 604770 42177 604834
rect 42111 604769 42177 604770
rect 42114 599063 42174 604769
rect 42111 599062 42177 599063
rect 42111 598998 42112 599062
rect 42176 598998 42177 599062
rect 42111 598997 42177 598998
rect 43071 599062 43137 599063
rect 43071 598998 43072 599062
rect 43136 598998 43137 599062
rect 43071 598997 43137 598998
rect 42495 591958 42561 591959
rect 42495 591894 42496 591958
rect 42560 591894 42561 591958
rect 42495 591893 42561 591894
rect 42498 588407 42558 591893
rect 42495 588406 42561 588407
rect 42495 588342 42496 588406
rect 42560 588342 42561 588406
rect 42495 588341 42561 588342
rect 41538 585051 41790 585111
rect 41343 580266 41409 580267
rect 41343 580202 41344 580266
rect 41408 580202 41409 580266
rect 41343 580201 41409 580202
rect 41538 574643 41598 585051
rect 42303 584706 42369 584707
rect 42303 584642 42304 584706
rect 42368 584642 42369 584706
rect 42303 584641 42369 584642
rect 41727 584558 41793 584559
rect 41727 584494 41728 584558
rect 41792 584494 41793 584558
rect 41727 584493 41793 584494
rect 41535 574642 41601 574643
rect 41535 574578 41536 574642
rect 41600 574578 41601 574642
rect 41535 574577 41601 574578
rect 41535 574494 41601 574495
rect 41535 574430 41536 574494
rect 41600 574430 41601 574494
rect 41535 574429 41601 574430
rect 40767 570498 40833 570499
rect 40767 570434 40768 570498
rect 40832 570434 40833 570498
rect 40767 570433 40833 570434
rect 41538 565023 41598 574429
rect 41730 574051 41790 584493
rect 42111 584410 42177 584411
rect 42111 584346 42112 584410
rect 42176 584346 42177 584410
rect 42111 584345 42177 584346
rect 41919 584262 41985 584263
rect 41919 584198 41920 584262
rect 41984 584198 41985 584262
rect 41919 584197 41985 584198
rect 41922 582043 41982 584197
rect 41919 582042 41985 582043
rect 41919 581978 41920 582042
rect 41984 581978 41985 582042
rect 41919 581977 41985 581978
rect 42114 574643 42174 584345
rect 42306 578343 42366 584641
rect 42495 584558 42561 584559
rect 42495 584494 42496 584558
rect 42560 584494 42561 584558
rect 42495 584493 42561 584494
rect 42303 578342 42369 578343
rect 42303 578278 42304 578342
rect 42368 578278 42369 578342
rect 42303 578277 42369 578278
rect 42498 577603 42558 584493
rect 42879 584262 42945 584263
rect 42879 584198 42880 584262
rect 42944 584198 42945 584262
rect 42879 584197 42945 584198
rect 42687 578934 42753 578935
rect 42687 578870 42688 578934
rect 42752 578870 42753 578934
rect 42687 578869 42753 578870
rect 42495 577602 42561 577603
rect 42495 577538 42496 577602
rect 42560 577538 42561 577602
rect 42495 577537 42561 577538
rect 42690 574939 42750 578869
rect 42882 578491 42942 584197
rect 43074 578935 43134 598997
rect 43071 578934 43137 578935
rect 43071 578870 43072 578934
rect 43136 578870 43137 578934
rect 43071 578869 43137 578870
rect 42879 578490 42945 578491
rect 42879 578426 42880 578490
rect 42944 578426 42945 578490
rect 42879 578425 42945 578426
rect 673986 576567 674046 645321
rect 674175 607794 674241 607795
rect 674175 607730 674176 607794
rect 674240 607730 674241 607794
rect 674175 607729 674241 607730
rect 673983 576566 674049 576567
rect 673983 576502 673984 576566
rect 674048 576502 674049 576566
rect 673983 576501 674049 576502
rect 42687 574938 42753 574939
rect 42687 574874 42688 574938
rect 42752 574874 42753 574938
rect 42687 574873 42753 574874
rect 42111 574642 42177 574643
rect 42111 574578 42112 574642
rect 42176 574578 42177 574642
rect 42111 574577 42177 574578
rect 41727 574050 41793 574051
rect 41727 573986 41728 574050
rect 41792 573986 41793 574050
rect 41727 573985 41793 573986
rect 41535 565022 41601 565023
rect 41535 564958 41536 565022
rect 41600 564958 41601 565022
rect 41535 564957 41601 564958
rect 41727 565022 41793 565023
rect 41727 564958 41728 565022
rect 41792 564958 41793 565022
rect 41727 564957 41793 564958
rect 40191 559102 40257 559103
rect 40191 559038 40192 559102
rect 40256 559038 40257 559102
rect 40191 559037 40257 559038
rect 40194 556883 40254 559037
rect 40191 556882 40257 556883
rect 40191 556818 40192 556882
rect 40256 556818 40257 556882
rect 40191 556817 40257 556818
rect 40767 554662 40833 554663
rect 40767 554598 40768 554662
rect 40832 554598 40833 554662
rect 40767 554597 40833 554598
rect 40770 530095 40830 554597
rect 40959 552442 41025 552443
rect 40959 552378 40960 552442
rect 41024 552378 41025 552442
rect 40959 552377 41025 552378
rect 40962 532611 41022 552377
rect 41730 541821 41790 564957
rect 42690 544599 42750 574873
rect 42687 544598 42753 544599
rect 42687 544534 42688 544598
rect 42752 544534 42753 544598
rect 42687 544533 42753 544534
rect 42111 544450 42177 544451
rect 42111 544386 42112 544450
rect 42176 544386 42177 544450
rect 42111 544385 42177 544386
rect 41538 541761 41790 541821
rect 41343 541342 41409 541343
rect 41343 541278 41344 541342
rect 41408 541278 41409 541342
rect 41343 541277 41409 541278
rect 40959 532610 41025 532611
rect 40959 532546 40960 532610
rect 41024 532546 41025 532610
rect 40959 532545 41025 532546
rect 41346 531279 41406 541277
rect 41538 532497 41598 541761
rect 41727 541342 41793 541343
rect 41727 541278 41728 541342
rect 41792 541278 41793 541342
rect 41727 541277 41793 541278
rect 41730 534387 41790 541277
rect 41919 541194 41985 541195
rect 41919 541130 41920 541194
rect 41984 541130 41985 541194
rect 41919 541129 41985 541130
rect 41727 534386 41793 534387
rect 41727 534322 41728 534386
rect 41792 534322 41793 534386
rect 41727 534321 41793 534322
rect 41922 533795 41982 541129
rect 41919 533794 41985 533795
rect 41919 533730 41920 533794
rect 41984 533730 41985 533794
rect 41919 533729 41985 533730
rect 42114 532759 42174 544385
rect 42879 541638 42945 541639
rect 42879 541574 42880 541638
rect 42944 541574 42945 541638
rect 42879 541573 42945 541574
rect 42303 541046 42369 541047
rect 42303 540982 42304 541046
rect 42368 540982 42369 541046
rect 42303 540981 42369 540982
rect 42306 538087 42366 540981
rect 42303 538086 42369 538087
rect 42303 538022 42304 538086
rect 42368 538022 42369 538086
rect 42303 538021 42369 538022
rect 42882 537051 42942 541573
rect 43071 541490 43137 541491
rect 43071 541426 43072 541490
rect 43136 541426 43137 541490
rect 43071 541425 43137 541426
rect 42879 537050 42945 537051
rect 42879 536986 42880 537050
rect 42944 536986 42945 537050
rect 42879 536985 42945 536986
rect 42111 532758 42177 532759
rect 42111 532694 42112 532758
rect 42176 532694 42177 532758
rect 42111 532693 42177 532694
rect 41538 532437 41790 532497
rect 41730 531871 41790 532437
rect 41727 531870 41793 531871
rect 41727 531806 41728 531870
rect 41792 531806 41793 531870
rect 41727 531805 41793 531806
rect 41343 531278 41409 531279
rect 41343 531214 41344 531278
rect 41408 531214 41409 531278
rect 41343 531213 41409 531214
rect 40767 530094 40833 530095
rect 40767 530030 40768 530094
rect 40832 530030 40833 530094
rect 40767 530029 40833 530030
rect 40383 429306 40449 429307
rect 40383 429242 40384 429306
rect 40448 429242 40449 429306
rect 40383 429241 40449 429242
rect 40386 386091 40446 429241
rect 40575 428714 40641 428715
rect 40575 428650 40576 428714
rect 40640 428650 40641 428714
rect 40575 428649 40641 428650
rect 40578 386091 40638 428649
rect 40767 428122 40833 428123
rect 40767 428058 40768 428122
rect 40832 428058 40833 428122
rect 40767 428057 40833 428058
rect 40770 400151 40830 428057
rect 40959 427086 41025 427087
rect 40959 427022 40960 427086
rect 41024 427022 41025 427086
rect 40959 427021 41025 427022
rect 40767 400150 40833 400151
rect 40767 400086 40768 400150
rect 40832 400086 40833 400150
rect 40767 400085 40833 400086
rect 40962 398819 41022 427021
rect 41343 426494 41409 426495
rect 41343 426430 41344 426494
rect 41408 426430 41409 426494
rect 41343 426429 41409 426430
rect 41151 424866 41217 424867
rect 41151 424802 41152 424866
rect 41216 424802 41217 424866
rect 41151 424801 41217 424802
rect 41154 399559 41214 424801
rect 41346 401927 41406 426429
rect 41535 424422 41601 424423
rect 41535 424358 41536 424422
rect 41600 424358 41601 424422
rect 41535 424357 41601 424358
rect 41538 402667 41598 424357
rect 41730 403851 41790 531805
rect 42114 529833 42174 532693
rect 42114 529773 42366 529833
rect 42306 509967 42366 529773
rect 43074 529503 43134 541425
rect 674178 532611 674238 607729
rect 674370 575383 674430 652129
rect 674562 620375 674622 694309
rect 674754 623187 674814 697861
rect 674946 665367 675006 739153
rect 675138 667587 675198 740041
rect 675330 711099 675390 787105
rect 675522 759347 675582 875757
rect 675903 786726 675969 786727
rect 675903 786662 675904 786726
rect 675968 786662 675969 786726
rect 675903 786661 675969 786662
rect 675711 784210 675777 784211
rect 675711 784146 675712 784210
rect 675776 784146 675777 784210
rect 675711 784145 675777 784146
rect 675519 759346 675585 759347
rect 675519 759282 675520 759346
rect 675584 759282 675585 759346
rect 675519 759281 675585 759282
rect 675519 742178 675585 742179
rect 675519 742114 675520 742178
rect 675584 742114 675585 742178
rect 675519 742113 675585 742114
rect 675327 711098 675393 711099
rect 675327 711034 675328 711098
rect 675392 711034 675393 711098
rect 675327 711033 675393 711034
rect 675327 696890 675393 696891
rect 675327 696826 675328 696890
rect 675392 696826 675393 696890
rect 675327 696825 675393 696826
rect 675135 667586 675201 667587
rect 675135 667522 675136 667586
rect 675200 667522 675201 667586
rect 675135 667521 675201 667522
rect 674943 665366 675009 665367
rect 674943 665302 674944 665366
rect 675008 665302 675009 665366
rect 674943 665301 675009 665302
rect 675135 652638 675201 652639
rect 675135 652574 675136 652638
rect 675200 652574 675201 652638
rect 675135 652573 675201 652574
rect 674943 648938 675009 648939
rect 674943 648874 674944 648938
rect 675008 648874 675009 648938
rect 674943 648873 675009 648874
rect 674751 623186 674817 623187
rect 674751 623122 674752 623186
rect 674816 623122 674817 623186
rect 674751 623121 674817 623122
rect 674559 620374 674625 620375
rect 674559 620310 674560 620374
rect 674624 620310 674625 620374
rect 674559 620309 674625 620310
rect 674751 607202 674817 607203
rect 674751 607138 674752 607202
rect 674816 607138 674817 607202
rect 674751 607137 674817 607138
rect 674559 604834 674625 604835
rect 674559 604770 674560 604834
rect 674624 604770 674625 604834
rect 674559 604769 674625 604770
rect 674367 575382 674433 575383
rect 674367 575318 674368 575382
rect 674432 575318 674433 575382
rect 674367 575317 674433 575318
rect 674367 562654 674433 562655
rect 674367 562590 674368 562654
rect 674432 562590 674433 562654
rect 674367 562589 674433 562590
rect 674175 532610 674241 532611
rect 674175 532546 674176 532610
rect 674240 532546 674241 532610
rect 674175 532545 674241 532546
rect 43071 529502 43137 529503
rect 43071 529438 43072 529502
rect 43136 529438 43137 529502
rect 43071 529437 43137 529438
rect 42303 509966 42369 509967
rect 42303 509902 42304 509966
rect 42368 509902 42369 509966
rect 42303 509901 42369 509902
rect 42111 504046 42177 504047
rect 42111 503982 42112 504046
rect 42176 503982 42177 504046
rect 42111 503981 42177 503982
rect 42114 489691 42174 503981
rect 42111 489690 42177 489691
rect 42111 489626 42112 489690
rect 42176 489626 42177 489690
rect 42111 489625 42177 489626
rect 42303 489394 42369 489395
rect 42303 489330 42304 489394
rect 42368 489330 42369 489394
rect 42303 489329 42369 489330
rect 42306 483771 42366 489329
rect 674370 488655 674430 562589
rect 674562 532315 674622 604769
rect 674559 532314 674625 532315
rect 674559 532250 674560 532314
rect 674624 532250 674625 532314
rect 674559 532249 674625 532250
rect 674754 530687 674814 607137
rect 674946 575235 675006 648873
rect 675138 577899 675198 652573
rect 675330 624223 675390 696825
rect 675522 665959 675582 742113
rect 675714 710655 675774 784145
rect 675906 714355 675966 786661
rect 676098 756091 676158 876497
rect 676287 784950 676353 784951
rect 676287 784886 676288 784950
rect 676352 784886 676353 784950
rect 676287 784885 676353 784886
rect 676095 756090 676161 756091
rect 676095 756026 676096 756090
rect 676160 756026 676161 756090
rect 676095 756025 676161 756026
rect 676095 741734 676161 741735
rect 676095 741670 676096 741734
rect 676160 741670 676161 741734
rect 676095 741669 676161 741670
rect 675903 714354 675969 714355
rect 675903 714290 675904 714354
rect 675968 714290 675969 714354
rect 675903 714289 675969 714290
rect 675711 710654 675777 710655
rect 675711 710590 675712 710654
rect 675776 710590 675777 710654
rect 675711 710589 675777 710590
rect 675903 694818 675969 694819
rect 675903 694754 675904 694818
rect 675968 694754 675969 694818
rect 675903 694753 675969 694754
rect 675519 665958 675585 665959
rect 675519 665894 675520 665958
rect 675584 665894 675585 665958
rect 675519 665893 675585 665894
rect 675519 651454 675585 651455
rect 675519 651390 675520 651454
rect 675584 651390 675585 651454
rect 675519 651389 675585 651390
rect 675327 624222 675393 624223
rect 675327 624158 675328 624222
rect 675392 624158 675393 624222
rect 675327 624157 675393 624158
rect 675327 606462 675393 606463
rect 675327 606398 675328 606462
rect 675392 606398 675393 606462
rect 675327 606397 675393 606398
rect 675135 577898 675201 577899
rect 675135 577834 675136 577898
rect 675200 577834 675201 577898
rect 675135 577833 675201 577834
rect 674943 575234 675009 575235
rect 674943 575170 674944 575234
rect 675008 575170 675009 575234
rect 674943 575169 675009 575170
rect 675135 561470 675201 561471
rect 675135 561406 675136 561470
rect 675200 561406 675201 561470
rect 675135 561405 675201 561406
rect 674943 558954 675009 558955
rect 674943 558890 674944 558954
rect 675008 558890 675009 558954
rect 674943 558889 675009 558890
rect 674751 530686 674817 530687
rect 674751 530622 674752 530686
rect 674816 530622 674817 530686
rect 674751 530621 674817 530622
rect 674367 488654 674433 488655
rect 674367 488590 674368 488654
rect 674432 488590 674433 488654
rect 674367 488589 674433 488590
rect 674946 486139 675006 558889
rect 675138 489987 675198 561405
rect 675330 533943 675390 606397
rect 675522 578935 675582 651389
rect 675711 649826 675777 649827
rect 675711 649762 675712 649826
rect 675776 649762 675777 649826
rect 675711 649761 675777 649762
rect 675519 578934 675585 578935
rect 675519 578870 675520 578934
rect 675584 578870 675585 578934
rect 675519 578869 675585 578870
rect 675714 577307 675774 649761
rect 675906 622595 675966 694753
rect 676098 669215 676158 741669
rect 676290 712727 676350 784885
rect 676671 780658 676737 780659
rect 676671 780594 676672 780658
rect 676736 780594 676737 780658
rect 676671 780593 676737 780594
rect 676674 773851 676734 780593
rect 677055 775626 677121 775627
rect 677055 775562 677056 775626
rect 677120 775587 677121 775626
rect 677120 775562 677310 775587
rect 677055 775561 677310 775562
rect 677058 775527 677310 775561
rect 676863 775034 676929 775035
rect 676863 774970 676864 775034
rect 676928 774970 676929 775034
rect 676863 774969 676929 774970
rect 676671 773850 676737 773851
rect 676671 773786 676672 773850
rect 676736 773786 676737 773850
rect 676671 773785 676737 773786
rect 676671 773702 676737 773703
rect 676671 773638 676672 773702
rect 676736 773638 676737 773702
rect 676671 773637 676737 773638
rect 676479 771778 676545 771779
rect 676479 771714 676480 771778
rect 676544 771714 676545 771778
rect 676479 771713 676545 771714
rect 676482 754463 676542 771713
rect 676479 754462 676545 754463
rect 676479 754398 676480 754462
rect 676544 754398 676545 754462
rect 676479 754397 676545 754398
rect 676674 741735 676734 773637
rect 676866 773111 676926 774969
rect 676863 773110 676929 773111
rect 676863 773046 676864 773110
rect 676928 773046 676929 773110
rect 676863 773045 676929 773046
rect 677250 772923 677310 775527
rect 677823 773110 677889 773111
rect 677823 773046 677824 773110
rect 677888 773046 677889 773110
rect 677823 773045 677889 773046
rect 676866 772863 677310 772923
rect 676866 764265 676926 772863
rect 677247 772666 677313 772667
rect 677247 772602 677248 772666
rect 677312 772602 677313 772666
rect 677247 772601 677313 772602
rect 677250 764527 677310 772601
rect 677826 764675 677886 773045
rect 679167 772962 679233 772963
rect 679167 772898 679168 772962
rect 679232 772898 679233 772962
rect 679167 772897 679233 772898
rect 677823 764674 677889 764675
rect 677823 764610 677824 764674
rect 677888 764610 677889 764674
rect 677823 764609 677889 764610
rect 677247 764526 677313 764527
rect 677247 764462 677248 764526
rect 677312 764462 677313 764526
rect 677247 764461 677313 764462
rect 677823 764526 677889 764527
rect 677823 764462 677824 764526
rect 677888 764462 677889 764526
rect 677823 764461 677889 764462
rect 676866 764205 677310 764265
rect 677055 759790 677121 759791
rect 677055 759726 677056 759790
rect 677120 759726 677121 759790
rect 677055 759725 677121 759726
rect 676863 759346 676929 759347
rect 676863 759282 676864 759346
rect 676928 759282 676929 759346
rect 676863 759281 676929 759282
rect 676866 741735 676926 759281
rect 677058 742176 677118 759725
rect 677250 756683 677310 764205
rect 677247 756682 677313 756683
rect 677247 756618 677248 756682
rect 677312 756618 677313 756682
rect 677247 756617 677313 756618
rect 677826 755055 677886 764461
rect 677823 755054 677889 755055
rect 677823 754990 677824 755054
rect 677888 754990 677889 755054
rect 677823 754989 677889 754990
rect 679170 754019 679230 772897
rect 679167 754018 679233 754019
rect 679167 753954 679168 754018
rect 679232 753954 679233 754018
rect 679167 753953 679233 753954
rect 677058 742116 677310 742176
rect 676671 741734 676737 741735
rect 676671 741670 676672 741734
rect 676736 741670 676737 741734
rect 676671 741669 676737 741670
rect 676863 741734 676929 741735
rect 676863 741670 676864 741734
rect 676928 741670 676929 741734
rect 676863 741669 676929 741670
rect 676479 741586 676545 741587
rect 676479 741522 676480 741586
rect 676544 741522 676545 741586
rect 676479 741521 676545 741522
rect 676287 712726 676353 712727
rect 676287 712662 676288 712726
rect 676352 712662 676353 712726
rect 676287 712661 676353 712662
rect 676482 712283 676542 741521
rect 676671 741438 676737 741439
rect 676671 741374 676672 741438
rect 676736 741374 676737 741438
rect 676671 741373 676737 741374
rect 676863 741438 676929 741439
rect 676863 741374 676864 741438
rect 676928 741374 676929 741438
rect 676863 741373 676929 741374
rect 676674 728119 676734 741373
rect 676671 728118 676737 728119
rect 676671 728054 676672 728118
rect 676736 728054 676737 728118
rect 676671 728053 676737 728054
rect 676866 714947 676926 741373
rect 677250 715539 677310 742116
rect 677823 728118 677889 728119
rect 677823 728054 677824 728118
rect 677888 728054 677889 728118
rect 677823 728053 677889 728054
rect 677247 715538 677313 715539
rect 677247 715474 677248 715538
rect 677312 715474 677313 715538
rect 677247 715473 677313 715474
rect 676863 714946 676929 714947
rect 676863 714882 676864 714946
rect 676928 714882 676929 714946
rect 676863 714881 676929 714882
rect 676479 712282 676545 712283
rect 676479 712218 676480 712282
rect 676544 712218 676545 712282
rect 676479 712217 676545 712218
rect 676671 697334 676737 697335
rect 676671 697270 676672 697334
rect 676736 697270 676737 697334
rect 676671 697269 676737 697270
rect 676479 693486 676545 693487
rect 676479 693422 676480 693486
rect 676544 693422 676545 693486
rect 676479 693421 676545 693422
rect 676287 692006 676353 692007
rect 676287 691942 676288 692006
rect 676352 691942 676353 692006
rect 676287 691941 676353 691942
rect 676095 669214 676161 669215
rect 676095 669150 676096 669214
rect 676160 669150 676161 669214
rect 676095 669149 676161 669150
rect 676290 653675 676350 691941
rect 676287 653674 676353 653675
rect 676287 653610 676288 653674
rect 676352 653610 676353 653674
rect 676287 653609 676353 653610
rect 676287 640354 676353 640355
rect 676287 640290 676288 640354
rect 676352 640290 676353 640354
rect 676287 640289 676353 640290
rect 676095 638578 676161 638579
rect 676095 638514 676096 638578
rect 676160 638514 676161 638578
rect 676095 638513 676161 638514
rect 675903 622594 675969 622595
rect 675903 622530 675904 622594
rect 675968 622530 675969 622594
rect 675903 622529 675969 622530
rect 675903 600246 675969 600247
rect 675903 600182 675904 600246
rect 675968 600182 675969 600246
rect 675903 600181 675969 600182
rect 675711 577306 675777 577307
rect 675711 577242 675712 577306
rect 675776 577242 675777 577306
rect 675711 577241 675777 577242
rect 675519 561766 675585 561767
rect 675519 561702 675520 561766
rect 675584 561702 675585 561766
rect 675519 561701 675585 561702
rect 675327 533942 675393 533943
rect 675327 533878 675328 533942
rect 675392 533878 675393 533942
rect 675327 533877 675393 533878
rect 675135 489986 675201 489987
rect 675135 489922 675136 489986
rect 675200 489922 675201 489986
rect 675135 489921 675201 489922
rect 675522 486731 675582 561701
rect 675906 531871 675966 600181
rect 676098 576271 676158 638513
rect 676290 578491 676350 640289
rect 676482 619931 676542 693421
rect 676674 620967 676734 697269
rect 676866 669659 676926 714881
rect 677826 711691 677886 728053
rect 677823 711690 677889 711691
rect 677823 711626 677824 711690
rect 677888 711626 677889 711690
rect 677823 711625 677889 711626
rect 677055 705770 677121 705771
rect 677055 705706 677056 705770
rect 677120 705706 677121 705770
rect 677055 705705 677121 705706
rect 677058 670251 677118 705705
rect 677055 670250 677121 670251
rect 677055 670186 677056 670250
rect 677120 670186 677121 670250
rect 677055 670185 677121 670186
rect 677247 670250 677313 670251
rect 677247 670186 677248 670250
rect 677312 670186 677313 670250
rect 677247 670185 677313 670186
rect 676863 669658 676929 669659
rect 676863 669594 676864 669658
rect 676928 669594 676929 669658
rect 676863 669593 676929 669594
rect 677058 663699 677118 670185
rect 676866 663639 677118 663699
rect 676866 624815 676926 663639
rect 677055 658854 677121 658855
rect 677055 658790 677056 658854
rect 677120 658790 677121 658854
rect 677055 658789 677121 658790
rect 676863 624814 676929 624815
rect 676863 624750 676864 624814
rect 676928 624750 676929 624814
rect 676863 624749 676929 624750
rect 677058 624667 677118 658789
rect 677250 626443 677310 670185
rect 677823 669066 677889 669067
rect 677823 669002 677824 669066
rect 677888 669002 677889 669066
rect 677823 669001 677889 669002
rect 677826 658855 677886 669001
rect 677823 658854 677889 658855
rect 677823 658790 677824 658854
rect 677888 658790 677889 658854
rect 677823 658789 677889 658790
rect 677247 626442 677313 626443
rect 677247 626378 677248 626442
rect 677312 626378 677313 626442
rect 677247 626377 677313 626378
rect 677055 624666 677121 624667
rect 677055 624602 677056 624666
rect 677120 624602 677121 624666
rect 677055 624601 677121 624602
rect 676671 620966 676737 620967
rect 676671 620902 676672 620966
rect 676736 620902 676737 620966
rect 676671 620901 676737 620902
rect 676479 619930 676545 619931
rect 676479 619866 676480 619930
rect 676544 619866 676545 619930
rect 676479 619865 676545 619866
rect 676671 595362 676737 595363
rect 676671 595298 676672 595362
rect 676736 595298 676737 595362
rect 676671 595297 676737 595298
rect 676479 593438 676545 593439
rect 676479 593374 676480 593438
rect 676544 593374 676545 593438
rect 676479 593373 676545 593374
rect 676287 578490 676353 578491
rect 676287 578426 676288 578490
rect 676352 578426 676353 578490
rect 676287 578425 676353 578426
rect 676095 576270 676161 576271
rect 676095 576206 676096 576270
rect 676160 576206 676161 576270
rect 676095 576205 676161 576206
rect 675903 531870 675969 531871
rect 675903 531806 675904 531870
rect 675968 531806 675969 531870
rect 675903 531805 675969 531806
rect 676482 531279 676542 593373
rect 676674 533499 676734 595297
rect 677055 579526 677121 579527
rect 677055 579462 677056 579526
rect 677120 579462 677121 579526
rect 677055 579461 677121 579462
rect 677247 579526 677313 579527
rect 677247 579462 677248 579526
rect 677312 579462 677313 579526
rect 677247 579461 677313 579462
rect 676863 554514 676929 554515
rect 676863 554450 676864 554514
rect 676928 554450 676929 554514
rect 676863 554449 676929 554450
rect 676671 533498 676737 533499
rect 676671 533434 676672 533498
rect 676736 533434 676737 533498
rect 676671 533433 676737 533434
rect 676479 531278 676545 531279
rect 676479 531214 676480 531278
rect 676544 531214 676545 531278
rect 676479 531213 676545 531214
rect 675519 486730 675585 486731
rect 675519 486666 675520 486730
rect 675584 486666 675585 486730
rect 675519 486665 675585 486666
rect 674943 486138 675009 486139
rect 674943 486074 674944 486138
rect 675008 486074 675009 486138
rect 674943 486073 675009 486074
rect 42303 483770 42369 483771
rect 42303 483706 42304 483770
rect 42368 483706 42369 483770
rect 42303 483705 42369 483706
rect 676866 483475 676926 554449
rect 677058 534535 677118 579461
rect 677250 534979 677310 579461
rect 677247 534978 677313 534979
rect 677247 534914 677248 534978
rect 677312 534914 677313 534978
rect 677247 534913 677313 534914
rect 677055 534534 677121 534535
rect 677055 534470 677056 534534
rect 677120 534470 677121 534534
rect 677055 534469 677121 534470
rect 676863 483474 676929 483475
rect 676863 483410 676864 483474
rect 676928 483410 676929 483474
rect 676863 483409 676929 483410
rect 42111 463790 42177 463791
rect 42111 463726 42112 463790
rect 42176 463726 42177 463790
rect 42111 463725 42177 463726
rect 42114 453243 42174 463725
rect 42114 453183 42366 453243
rect 42306 429267 42366 453183
rect 42306 429207 42606 429267
rect 42546 428712 42606 429207
rect 42498 428652 42606 428712
rect 42111 426050 42177 426051
rect 42111 425986 42112 426050
rect 42176 425986 42177 426050
rect 42111 425985 42177 425986
rect 41919 409030 41985 409031
rect 41919 408966 41920 409030
rect 41984 408966 41985 409030
rect 41919 408965 41985 408966
rect 41922 408883 41982 408965
rect 41919 408882 41985 408883
rect 41919 408818 41920 408882
rect 41984 408818 41985 408882
rect 41919 408817 41985 408818
rect 42114 406071 42174 425985
rect 42303 409326 42369 409327
rect 42303 409262 42304 409326
rect 42368 409262 42369 409326
rect 42303 409261 42369 409262
rect 42306 408143 42366 409261
rect 42498 409031 42558 428652
rect 42495 409030 42561 409031
rect 42495 408966 42496 409030
rect 42560 408966 42561 409030
rect 42495 408965 42561 408966
rect 42495 408882 42561 408883
rect 42495 408818 42496 408882
rect 42560 408818 42561 408882
rect 42495 408817 42561 408818
rect 42303 408142 42369 408143
rect 42303 408078 42304 408142
rect 42368 408078 42369 408142
rect 42303 408077 42369 408078
rect 42111 406070 42177 406071
rect 42111 406006 42112 406070
rect 42176 406006 42177 406070
rect 42111 406005 42177 406006
rect 42498 405291 42558 408817
rect 42114 405231 42558 405291
rect 42114 404295 42174 405231
rect 42111 404294 42177 404295
rect 42111 404230 42112 404294
rect 42176 404230 42177 404294
rect 42111 404229 42177 404230
rect 41727 403850 41793 403851
rect 41727 403786 41728 403850
rect 41792 403786 41793 403850
rect 41727 403785 41793 403786
rect 41535 402666 41601 402667
rect 41535 402602 41536 402666
rect 41600 402602 41601 402666
rect 41535 402601 41601 402602
rect 41343 401926 41409 401927
rect 41343 401862 41344 401926
rect 41408 401862 41409 401926
rect 41343 401861 41409 401862
rect 41151 399558 41217 399559
rect 41151 399494 41152 399558
rect 41216 399494 41217 399558
rect 41151 399493 41217 399494
rect 40959 398818 41025 398819
rect 40959 398754 40960 398818
rect 41024 398754 41025 398818
rect 40959 398753 41025 398754
rect 40383 386090 40449 386091
rect 40383 386026 40384 386090
rect 40448 386026 40449 386090
rect 40383 386025 40449 386026
rect 40575 386090 40641 386091
rect 40575 386026 40576 386090
rect 40640 386026 40641 386090
rect 40575 386025 40641 386026
rect 40386 343023 40446 386025
rect 40383 343022 40449 343023
rect 40383 342958 40384 343022
rect 40448 342958 40449 343022
rect 40383 342957 40449 342958
rect 40386 299807 40446 342957
rect 40578 342875 40638 386025
rect 40767 384906 40833 384907
rect 40767 384842 40768 384906
rect 40832 384842 40833 384906
rect 40767 384841 40833 384842
rect 40770 356935 40830 384841
rect 40959 383870 41025 383871
rect 40959 383806 40960 383870
rect 41024 383806 41025 383870
rect 40959 383805 41025 383806
rect 40767 356934 40833 356935
rect 40767 356870 40768 356934
rect 40832 356870 40833 356934
rect 40767 356869 40833 356870
rect 40962 355603 41022 383805
rect 41343 383278 41409 383279
rect 41343 383214 41344 383278
rect 41408 383214 41409 383278
rect 41343 383213 41409 383214
rect 41151 381650 41217 381651
rect 41151 381586 41152 381650
rect 41216 381586 41217 381650
rect 41151 381585 41217 381586
rect 41154 356491 41214 381585
rect 41346 358711 41406 383213
rect 41535 382834 41601 382835
rect 41535 382770 41536 382834
rect 41600 382770 41601 382834
rect 41535 382769 41601 382770
rect 41538 362855 41598 382769
rect 41535 362854 41601 362855
rect 41535 362790 41536 362854
rect 41600 362790 41601 362854
rect 41535 362789 41601 362790
rect 41730 360635 41790 403785
rect 42114 393303 42174 404229
rect 674559 400594 674625 400595
rect 674559 400530 674560 400594
rect 674624 400530 674625 400594
rect 674559 400529 674625 400530
rect 674367 399262 674433 399263
rect 674367 399198 674368 399262
rect 674432 399198 674433 399262
rect 674367 399197 674433 399198
rect 674175 398818 674241 398819
rect 674175 398754 674176 398818
rect 674240 398754 674241 398818
rect 674175 398753 674241 398754
rect 42114 393243 42558 393303
rect 42498 383313 42558 393243
rect 42306 383253 42558 383313
rect 42111 381206 42177 381207
rect 42111 381142 42112 381206
rect 42176 381142 42177 381206
rect 42111 381141 42177 381142
rect 42114 368775 42174 381141
rect 42306 380171 42366 383253
rect 42303 380170 42369 380171
rect 42303 380106 42304 380170
rect 42368 380106 42369 380170
rect 42303 380105 42369 380106
rect 42879 380170 42945 380171
rect 42879 380106 42880 380170
rect 42944 380106 42945 380170
rect 42879 380105 42945 380106
rect 42495 378986 42561 378987
rect 42495 378922 42496 378986
rect 42560 378922 42561 378986
rect 42495 378921 42561 378922
rect 42111 368774 42177 368775
rect 42111 368710 42112 368774
rect 42176 368710 42177 368774
rect 42111 368709 42177 368710
rect 42111 368478 42177 368479
rect 42111 368414 42112 368478
rect 42176 368414 42177 368478
rect 42111 368413 42177 368414
rect 41727 360634 41793 360635
rect 41727 360570 41728 360634
rect 41792 360570 41793 360634
rect 41727 360569 41793 360570
rect 42114 359451 42174 368413
rect 42303 361966 42369 361967
rect 42303 361902 42304 361966
rect 42368 361902 42369 361966
rect 42303 361901 42369 361902
rect 42306 360669 42366 361901
rect 42498 361227 42558 378921
rect 42882 361967 42942 380105
rect 674178 372031 674238 398753
rect 674370 378839 674430 399197
rect 674367 378838 674433 378839
rect 674367 378774 674368 378838
rect 674432 378774 674433 378838
rect 674367 378773 674433 378774
rect 674562 373955 674622 400529
rect 675327 374546 675393 374547
rect 675327 374482 675328 374546
rect 675392 374482 675393 374546
rect 675327 374481 675393 374482
rect 674559 373954 674625 373955
rect 674559 373890 674560 373954
rect 674624 373890 674625 373954
rect 674559 373889 674625 373890
rect 674175 372030 674241 372031
rect 674175 371966 674176 372030
rect 674240 371966 674241 372030
rect 674175 371965 674241 371966
rect 42879 361966 42945 361967
rect 42879 361902 42880 361966
rect 42944 361902 42945 361966
rect 42879 361901 42945 361902
rect 42495 361226 42561 361227
rect 42495 361162 42496 361226
rect 42560 361162 42561 361226
rect 42495 361161 42561 361162
rect 42306 360609 42558 360669
rect 42111 359450 42177 359451
rect 42111 359386 42112 359450
rect 42176 359386 42177 359450
rect 42111 359385 42177 359386
rect 41343 358710 41409 358711
rect 41343 358646 41344 358710
rect 41408 358646 41409 358710
rect 41343 358645 41409 358646
rect 41151 356490 41217 356491
rect 41151 356426 41152 356490
rect 41216 356426 41217 356490
rect 41151 356425 41217 356426
rect 40959 355602 41025 355603
rect 40959 355538 40960 355602
rect 41024 355538 41025 355602
rect 40959 355537 41025 355538
rect 40575 342874 40641 342875
rect 40575 342810 40576 342874
rect 40640 342810 40641 342874
rect 40575 342809 40641 342810
rect 40383 299806 40449 299807
rect 40383 299742 40384 299806
rect 40448 299742 40449 299806
rect 40383 299741 40449 299742
rect 40386 257035 40446 299741
rect 40578 299659 40638 342809
rect 40767 341838 40833 341839
rect 40767 341774 40768 341838
rect 40832 341774 40833 341838
rect 40767 341773 40833 341774
rect 40770 313719 40830 341773
rect 40959 340654 41025 340655
rect 40959 340590 40960 340654
rect 41024 340590 41025 340654
rect 40959 340589 41025 340590
rect 40767 313718 40833 313719
rect 40767 313654 40768 313718
rect 40832 313654 40833 313718
rect 40767 313653 40833 313654
rect 40962 312387 41022 340589
rect 41343 340210 41409 340211
rect 41343 340146 41344 340210
rect 41408 340146 41409 340210
rect 41343 340145 41409 340146
rect 41151 338582 41217 338583
rect 41151 338518 41152 338582
rect 41216 338518 41217 338582
rect 41151 338517 41217 338518
rect 41154 313275 41214 338517
rect 41346 315495 41406 340145
rect 42111 339618 42177 339619
rect 42111 339554 42112 339618
rect 42176 339554 42177 339618
rect 42111 339553 42177 339554
rect 41535 337990 41601 337991
rect 41535 337926 41536 337990
rect 41600 337926 41601 337990
rect 41535 337925 41601 337926
rect 41538 316235 41598 337925
rect 41727 335178 41793 335179
rect 41727 335114 41728 335178
rect 41792 335114 41793 335178
rect 41727 335113 41793 335114
rect 41730 320527 41790 335113
rect 41727 320526 41793 320527
rect 41727 320462 41728 320526
rect 41792 320462 41793 320526
rect 41727 320461 41793 320462
rect 42114 319787 42174 339553
rect 42111 319786 42177 319787
rect 42111 319722 42112 319786
rect 42176 319722 42177 319786
rect 42111 319721 42177 319722
rect 42498 318455 42558 360609
rect 42879 360634 42945 360635
rect 42879 360570 42880 360634
rect 42944 360570 42945 360634
rect 42879 360569 42945 360570
rect 42687 336066 42753 336067
rect 42687 336002 42688 336066
rect 42752 336002 42753 336066
rect 42687 336001 42753 336002
rect 42690 324819 42750 336001
rect 42687 324818 42753 324819
rect 42687 324754 42688 324818
rect 42752 324754 42753 324818
rect 42687 324753 42753 324754
rect 41727 318454 41793 318455
rect 41727 318390 41728 318454
rect 41792 318390 41793 318454
rect 41727 318389 41793 318390
rect 42495 318454 42561 318455
rect 42495 318390 42496 318454
rect 42560 318390 42561 318454
rect 42495 318389 42561 318390
rect 41535 316234 41601 316235
rect 41535 316170 41536 316234
rect 41600 316170 41601 316234
rect 41535 316169 41601 316170
rect 41343 315494 41409 315495
rect 41343 315430 41344 315494
rect 41408 315430 41409 315494
rect 41343 315429 41409 315430
rect 41151 313274 41217 313275
rect 41151 313210 41152 313274
rect 41216 313210 41217 313274
rect 41151 313209 41217 313210
rect 40959 312386 41025 312387
rect 40959 312322 40960 312386
rect 41024 312322 41025 312386
rect 40959 312321 41025 312322
rect 40575 299658 40641 299659
rect 40575 299594 40576 299658
rect 40640 299594 40641 299658
rect 40575 299593 40641 299594
rect 40959 298622 41025 298623
rect 40959 298558 40960 298622
rect 41024 298558 41025 298622
rect 40959 298557 41025 298558
rect 40767 297438 40833 297439
rect 40767 297374 40768 297438
rect 40832 297374 40833 297438
rect 40767 297373 40833 297374
rect 40770 269171 40830 297373
rect 40962 270651 41022 298557
rect 41343 296994 41409 296995
rect 41343 296930 41344 296994
rect 41408 296930 41409 296994
rect 41343 296929 41409 296930
rect 41151 295366 41217 295367
rect 41151 295302 41152 295366
rect 41216 295302 41217 295366
rect 41151 295301 41217 295302
rect 40959 270650 41025 270651
rect 40959 270586 40960 270650
rect 41024 270586 41025 270650
rect 40959 270585 41025 270586
rect 41154 270059 41214 295301
rect 41346 272279 41406 296929
rect 41535 294774 41601 294775
rect 41535 294710 41536 294774
rect 41600 294710 41601 294774
rect 41535 294709 41601 294710
rect 41538 273019 41598 294709
rect 41730 274647 41790 318389
rect 42882 318011 42942 360569
rect 674175 355750 674241 355751
rect 674175 355686 674176 355750
rect 674240 355686 674241 355750
rect 674175 355685 674241 355686
rect 673983 331182 674049 331183
rect 673983 331118 673984 331182
rect 674048 331118 674049 331182
rect 673983 331117 674049 331118
rect 41919 318010 41985 318011
rect 41919 317946 41920 318010
rect 41984 317946 41985 318010
rect 41919 317945 41985 317946
rect 42879 318010 42945 318011
rect 42879 317946 42880 318010
rect 42944 317946 42945 318010
rect 42879 317945 42945 317946
rect 41922 274795 41982 317945
rect 42303 299658 42369 299659
rect 42303 299594 42304 299658
rect 42368 299594 42369 299658
rect 42303 299593 42369 299594
rect 42111 296550 42177 296551
rect 42111 296486 42112 296550
rect 42176 296486 42177 296550
rect 42111 296485 42177 296486
rect 42114 276571 42174 296485
rect 42111 276570 42177 276571
rect 42111 276506 42112 276570
rect 42176 276506 42177 276570
rect 42111 276505 42177 276506
rect 41919 274794 41985 274795
rect 41919 274730 41920 274794
rect 41984 274730 41985 274794
rect 41919 274729 41985 274730
rect 41727 274646 41793 274647
rect 41727 274582 41728 274646
rect 41792 274582 41793 274646
rect 41727 274581 41793 274582
rect 41535 273018 41601 273019
rect 41535 272954 41536 273018
rect 41600 272954 41601 273018
rect 41535 272953 41601 272954
rect 41343 272278 41409 272279
rect 41343 272214 41344 272278
rect 41408 272214 41409 272278
rect 41343 272213 41409 272214
rect 41922 270651 41982 274729
rect 41919 270650 41985 270651
rect 41919 270586 41920 270650
rect 41984 270586 41985 270650
rect 41919 270585 41985 270586
rect 41151 270058 41217 270059
rect 41151 269994 41152 270058
rect 41216 269994 41217 270058
rect 41151 269993 41217 269994
rect 40767 269170 40833 269171
rect 40767 269106 40768 269170
rect 40832 269106 40833 269170
rect 40767 269105 40833 269106
rect 40383 257034 40449 257035
rect 40383 256970 40384 257034
rect 40448 256970 40449 257034
rect 40383 256969 40449 256970
rect 42306 256443 42366 299593
rect 42687 291814 42753 291815
rect 42687 291750 42688 291814
rect 42752 291750 42753 291814
rect 42687 291749 42753 291750
rect 42495 284858 42561 284859
rect 42495 284794 42496 284858
rect 42560 284794 42561 284858
rect 42495 284793 42561 284794
rect 42498 281603 42558 284793
rect 42495 281602 42561 281603
rect 42495 281538 42496 281602
rect 42560 281538 42561 281602
rect 42495 281537 42561 281538
rect 42690 278643 42750 291749
rect 673986 289595 674046 331117
rect 674178 328371 674238 355685
rect 675330 335031 675390 374481
rect 676863 374398 676929 374399
rect 676863 374334 676864 374398
rect 676928 374334 676929 374398
rect 676863 374333 676929 374334
rect 675519 374102 675585 374103
rect 675519 374038 675520 374102
rect 675584 374038 675585 374102
rect 675519 374037 675585 374038
rect 675327 335030 675393 335031
rect 675327 334966 675328 335030
rect 675392 334966 675393 335030
rect 675327 334965 675393 334966
rect 675522 334587 675582 374037
rect 676866 357083 676926 374333
rect 677055 373362 677121 373363
rect 677055 373298 677056 373362
rect 677120 373323 677121 373362
rect 677120 373298 677310 373323
rect 677055 373297 677310 373298
rect 677058 373263 677310 373297
rect 677055 357674 677121 357675
rect 677055 357610 677056 357674
rect 677120 357610 677121 357674
rect 677055 357609 677121 357610
rect 676863 357082 676929 357083
rect 676863 357018 676864 357082
rect 676928 357018 676929 357082
rect 676863 357017 676929 357018
rect 676671 345242 676737 345243
rect 676671 345178 676672 345242
rect 676736 345178 676737 345242
rect 676671 345177 676737 345178
rect 676479 344206 676545 344207
rect 676479 344142 676480 344206
rect 676544 344142 676545 344206
rect 676479 344141 676545 344142
rect 675519 334586 675585 334587
rect 675519 334522 675520 334586
rect 675584 334522 675585 334586
rect 675519 334521 675585 334522
rect 676482 330591 676542 344141
rect 676479 330590 676545 330591
rect 676479 330526 676480 330590
rect 676544 330526 676545 330590
rect 676479 330525 676545 330526
rect 675327 329554 675393 329555
rect 675327 329490 675328 329554
rect 675392 329490 675393 329554
rect 675327 329489 675393 329490
rect 674175 328370 674241 328371
rect 674175 328306 674176 328370
rect 674240 328306 674241 328370
rect 674175 328305 674241 328306
rect 674175 310758 674241 310759
rect 674175 310694 674176 310758
rect 674240 310694 674241 310758
rect 674175 310693 674241 310694
rect 673983 289594 674049 289595
rect 673983 289530 673984 289594
rect 674048 289530 674049 289594
rect 673983 289529 674049 289530
rect 673983 284710 674049 284711
rect 673983 284646 673984 284710
rect 674048 284646 674049 284710
rect 673983 284645 674049 284646
rect 42687 278642 42753 278643
rect 42687 278578 42688 278642
rect 42752 278578 42753 278642
rect 42687 278577 42753 278578
rect 590271 278494 590337 278495
rect 590271 278430 590272 278494
rect 590336 278430 590337 278494
rect 590271 278429 590337 278430
rect 604863 278494 604929 278495
rect 604863 278430 604864 278494
rect 604928 278430 604929 278494
rect 604863 278429 604929 278430
rect 590274 278085 590334 278429
rect 604866 278347 604926 278429
rect 590463 278346 590529 278347
rect 590463 278282 590464 278346
rect 590528 278282 590529 278346
rect 590463 278281 590529 278282
rect 604863 278346 604929 278347
rect 604863 278282 604864 278346
rect 604928 278282 604929 278346
rect 604863 278281 604929 278282
rect 645183 278346 645249 278347
rect 645183 278282 645184 278346
rect 645248 278282 645249 278346
rect 645183 278281 645249 278282
rect 590466 278085 590526 278281
rect 645186 278199 645246 278281
rect 645183 278198 645249 278199
rect 645183 278134 645184 278198
rect 645248 278134 645249 278198
rect 645183 278133 645249 278134
rect 590274 278025 590526 278085
rect 42879 274646 42945 274647
rect 42879 274582 42880 274646
rect 42944 274582 42945 274646
rect 42879 274581 42945 274582
rect 42303 256442 42369 256443
rect 42303 256378 42304 256442
rect 42368 256378 42369 256442
rect 42303 256377 42369 256378
rect 40575 255406 40641 255407
rect 40575 255342 40576 255406
rect 40640 255342 40641 255406
rect 40575 255341 40641 255342
rect 40383 254222 40449 254223
rect 40383 254158 40384 254222
rect 40448 254158 40449 254222
rect 40383 254157 40449 254158
rect 40386 225955 40446 254157
rect 40578 227435 40638 255341
rect 40767 253778 40833 253779
rect 40767 253714 40768 253778
rect 40832 253714 40833 253778
rect 40767 253713 40833 253714
rect 40770 229063 40830 253713
rect 41343 253334 41409 253335
rect 41343 253270 41344 253334
rect 41408 253270 41409 253334
rect 41343 253269 41409 253270
rect 40959 252150 41025 252151
rect 40959 252086 40960 252150
rect 41024 252086 41025 252150
rect 40959 252085 41025 252086
rect 40767 229062 40833 229063
rect 40767 228998 40768 229062
rect 40832 228998 40833 229062
rect 40767 228997 40833 228998
rect 40575 227434 40641 227435
rect 40575 227370 40576 227434
rect 40640 227370 40641 227434
rect 40575 227369 40641 227370
rect 40962 226843 41022 252085
rect 41151 251558 41217 251559
rect 41151 251494 41152 251558
rect 41216 251494 41217 251558
rect 41151 251493 41217 251494
rect 41154 229655 41214 251493
rect 41346 233355 41406 253269
rect 41535 251114 41601 251115
rect 41535 251050 41536 251114
rect 41600 251050 41601 251114
rect 41535 251049 41601 251050
rect 41343 233354 41409 233355
rect 41343 233290 41344 233354
rect 41408 233290 41409 233354
rect 41343 233289 41409 233290
rect 41538 230395 41598 251049
rect 42882 246527 42942 274581
rect 477951 273758 478017 273759
rect 477951 273694 477952 273758
rect 478016 273694 478017 273758
rect 477951 273693 478017 273694
rect 477954 273463 478014 273693
rect 407487 273462 407553 273463
rect 407487 273398 407488 273462
rect 407552 273398 407553 273462
rect 407487 273397 407553 273398
rect 477951 273462 478017 273463
rect 477951 273398 477952 273462
rect 478016 273398 478017 273462
rect 477951 273397 478017 273398
rect 406143 271834 406209 271835
rect 406143 271770 406144 271834
rect 406208 271770 406209 271834
rect 406143 271769 406209 271770
rect 328191 271390 328257 271391
rect 328191 271326 328192 271390
rect 328256 271326 328257 271390
rect 328191 271325 328257 271326
rect 276351 268578 276417 268579
rect 276351 268514 276352 268578
rect 276416 268514 276417 268578
rect 276351 268513 276417 268514
rect 276354 267691 276414 268513
rect 328194 268183 328254 271325
rect 381759 271242 381825 271243
rect 381759 271178 381760 271242
rect 381824 271178 381825 271242
rect 381759 271177 381825 271178
rect 328575 270946 328641 270947
rect 328575 270882 328576 270946
rect 328640 270882 328641 270946
rect 328575 270881 328641 270882
rect 328578 268183 328638 270881
rect 371586 270503 371646 270611
rect 370623 270502 370689 270503
rect 370623 270438 370624 270502
rect 370688 270438 370689 270502
rect 370623 270437 370689 270438
rect 371199 270502 371265 270503
rect 371199 270438 371200 270502
rect 371264 270500 371265 270502
rect 371583 270502 371649 270503
rect 371264 270440 371454 270500
rect 371264 270438 371265 270440
rect 371199 270437 371265 270438
rect 370626 270181 370686 270437
rect 327231 267986 327297 267987
rect 327231 267922 327232 267986
rect 327296 267922 327297 267986
rect 329151 267986 329217 267987
rect 327231 267921 327297 267922
rect 329151 267922 329152 267986
rect 329216 267922 329217 267986
rect 329151 267921 329217 267922
rect 276351 267690 276417 267691
rect 276351 267626 276352 267690
rect 276416 267626 276417 267690
rect 276351 267625 276417 267626
rect 327234 267517 327294 267921
rect 328767 267690 328833 267691
rect 328767 267626 328768 267690
rect 328832 267626 328833 267690
rect 328767 267625 328833 267626
rect 328770 267429 328830 267625
rect 329154 267429 329214 267921
rect 371199 267838 371265 267839
rect 371199 267836 371200 267838
rect 370818 267776 371200 267836
rect 370818 267691 370878 267776
rect 371199 267774 371200 267776
rect 371264 267774 371265 267838
rect 371199 267773 371265 267774
rect 352767 267690 352833 267691
rect 352767 267626 352768 267690
rect 352832 267626 352833 267690
rect 352767 267625 352833 267626
rect 370815 267690 370881 267691
rect 370815 267626 370816 267690
rect 370880 267626 370881 267690
rect 370815 267625 370881 267626
rect 352770 267517 352830 267625
rect 328770 267369 329214 267429
rect 371394 265519 371454 270440
rect 371583 270438 371584 270502
rect 371648 270438 371649 270502
rect 371583 270437 371649 270438
rect 381762 270181 381822 271177
rect 395775 270798 395841 270799
rect 395775 270734 395776 270798
rect 395840 270734 395841 270798
rect 395775 270733 395841 270734
rect 395778 269515 395838 270733
rect 380034 269023 380094 269279
rect 380031 269022 380097 269023
rect 380031 268958 380032 269022
rect 380096 268958 380097 269022
rect 380031 268957 380097 268958
rect 404610 268701 405822 268761
rect 404610 268283 404670 268701
rect 377343 268282 377409 268283
rect 377343 268218 377344 268282
rect 377408 268218 377409 268282
rect 377343 268217 377409 268218
rect 404607 268282 404673 268283
rect 404607 268218 404608 268282
rect 404672 268218 404673 268282
rect 404607 268217 404673 268218
rect 405567 268282 405633 268283
rect 405567 268218 405568 268282
rect 405632 268218 405633 268282
rect 405567 268217 405633 268218
rect 377151 267838 377217 267839
rect 377151 267774 377152 267838
rect 377216 267836 377217 267838
rect 377346 267836 377406 268217
rect 389058 268035 389502 268095
rect 389058 267839 389118 268035
rect 377216 267776 377406 267836
rect 389055 267838 389121 267839
rect 377216 267774 377217 267776
rect 377151 267773 377217 267774
rect 389055 267774 389056 267838
rect 389120 267774 389121 267838
rect 389055 267773 389121 267774
rect 389442 267691 389502 268035
rect 389439 267690 389505 267691
rect 389439 267626 389440 267690
rect 389504 267626 389505 267690
rect 389439 267625 389505 267626
rect 181311 247118 181377 247119
rect 181311 247054 181312 247118
rect 181376 247054 181377 247118
rect 181311 247053 181377 247054
rect 207231 247118 207297 247119
rect 207231 247054 207232 247118
rect 207296 247054 207297 247118
rect 207231 247053 207297 247054
rect 42879 246526 42945 246527
rect 42879 246462 42880 246526
rect 42944 246462 42945 246526
rect 42879 246461 42945 246462
rect 41727 243862 41793 243863
rect 41727 243798 41728 243862
rect 41792 243798 41793 243862
rect 41727 243797 41793 243798
rect 41730 231135 41790 243797
rect 42882 242975 42942 246461
rect 181314 245935 181374 247053
rect 207234 246675 207294 247053
rect 405570 246971 405630 268217
rect 405567 246970 405633 246971
rect 405567 246906 405568 246970
rect 405632 246906 405633 246970
rect 405567 246905 405633 246906
rect 207231 246674 207297 246675
rect 207231 246610 207232 246674
rect 207296 246610 207297 246674
rect 207231 246609 207297 246610
rect 181311 245934 181377 245935
rect 181311 245870 181312 245934
rect 181376 245870 181377 245934
rect 181311 245869 181377 245870
rect 210303 243714 210369 243715
rect 210303 243650 210304 243714
rect 210368 243650 210369 243714
rect 210303 243649 210369 243650
rect 210495 243714 210561 243715
rect 210495 243650 210496 243714
rect 210560 243650 210561 243714
rect 210495 243649 210561 243650
rect 268095 243714 268161 243715
rect 268095 243650 268096 243714
rect 268160 243650 268161 243714
rect 268095 243649 268161 243650
rect 41919 242974 41985 242975
rect 41919 242910 41920 242974
rect 41984 242910 41985 242974
rect 41919 242909 41985 242910
rect 42879 242974 42945 242975
rect 42879 242910 42880 242974
rect 42944 242910 42945 242974
rect 42879 242909 42945 242910
rect 41922 231727 41982 242909
rect 115263 242678 115329 242679
rect 115263 242614 115264 242678
rect 115328 242614 115329 242678
rect 115263 242613 115329 242614
rect 175551 242678 175617 242679
rect 175551 242614 175552 242678
rect 175616 242614 175617 242678
rect 175551 242613 175617 242614
rect 115266 242531 115326 242613
rect 115263 242530 115329 242531
rect 115263 242466 115264 242530
rect 115328 242466 115329 242530
rect 115263 242465 115329 242466
rect 175554 242383 175614 242613
rect 175551 242382 175617 242383
rect 175551 242318 175552 242382
rect 175616 242318 175617 242382
rect 175551 242317 175617 242318
rect 42303 240754 42369 240755
rect 42303 240690 42304 240754
rect 42368 240690 42369 240754
rect 42303 240689 42369 240690
rect 42306 236611 42366 240689
rect 145407 239866 145473 239867
rect 145407 239802 145408 239866
rect 145472 239802 145473 239866
rect 145407 239801 145473 239802
rect 42303 236610 42369 236611
rect 42303 236546 42304 236610
rect 42368 236546 42369 236610
rect 42303 236545 42369 236546
rect 41919 231726 41985 231727
rect 41919 231662 41920 231726
rect 41984 231662 41985 231726
rect 41919 231661 41985 231662
rect 41727 231134 41793 231135
rect 41727 231070 41728 231134
rect 41792 231070 41793 231134
rect 41727 231069 41793 231070
rect 41535 230394 41601 230395
rect 41535 230330 41536 230394
rect 41600 230330 41601 230394
rect 41535 230329 41601 230330
rect 41151 229654 41217 229655
rect 41151 229590 41152 229654
rect 41216 229590 41217 229654
rect 41151 229589 41217 229590
rect 40959 226842 41025 226843
rect 40959 226778 40960 226842
rect 41024 226778 41025 226842
rect 40959 226777 41025 226778
rect 40383 225954 40449 225955
rect 40383 225890 40384 225954
rect 40448 225890 40449 225954
rect 40383 225889 40449 225890
rect 40575 212190 40641 212191
rect 40575 212126 40576 212190
rect 40640 212126 40641 212190
rect 40575 212125 40641 212126
rect 40383 211154 40449 211155
rect 40383 211090 40384 211154
rect 40448 211090 40449 211154
rect 40383 211089 40449 211090
rect 40386 182887 40446 211089
rect 40578 184219 40638 212125
rect 40959 210562 41025 210563
rect 40959 210498 40960 210562
rect 41024 210498 41025 210562
rect 40959 210497 41025 210498
rect 40767 208934 40833 208935
rect 40767 208870 40768 208934
rect 40832 208870 40833 208934
rect 40767 208869 40833 208870
rect 40575 184218 40641 184219
rect 40575 184154 40576 184218
rect 40640 184154 40641 184218
rect 40575 184153 40641 184154
rect 40770 183627 40830 208869
rect 40962 185847 41022 210497
rect 41151 208342 41217 208343
rect 41151 208278 41152 208342
rect 41216 208278 41217 208342
rect 41151 208277 41217 208278
rect 41154 186735 41214 208277
rect 41730 188363 41790 231069
rect 41922 189103 41982 231661
rect 42111 201238 42177 201239
rect 42111 201174 42112 201238
rect 42176 201174 42177 201238
rect 42111 201173 42177 201174
rect 42114 190287 42174 201173
rect 42303 197538 42369 197539
rect 42303 197474 42304 197538
rect 42368 197474 42369 197538
rect 42303 197473 42369 197474
rect 42306 195171 42366 197473
rect 42303 195170 42369 195171
rect 42303 195106 42304 195170
rect 42368 195106 42369 195170
rect 42303 195105 42369 195106
rect 42111 190286 42177 190287
rect 42111 190222 42112 190286
rect 42176 190222 42177 190286
rect 42111 190221 42177 190222
rect 41919 189102 41985 189103
rect 41919 189038 41920 189102
rect 41984 189038 41985 189102
rect 41919 189037 41985 189038
rect 41727 188362 41793 188363
rect 41727 188298 41728 188362
rect 41792 188298 41793 188362
rect 41727 188297 41793 188298
rect 41151 186734 41217 186735
rect 41151 186670 41152 186734
rect 41216 186670 41217 186734
rect 41151 186669 41217 186670
rect 40959 185846 41025 185847
rect 40959 185782 40960 185846
rect 41024 185782 41025 185846
rect 40959 185781 41025 185782
rect 40767 183626 40833 183627
rect 40767 183562 40768 183626
rect 40832 183562 40833 183626
rect 40767 183561 40833 183562
rect 40383 182886 40449 182887
rect 40383 182822 40384 182886
rect 40448 182822 40449 182886
rect 40383 182821 40449 182822
rect 145410 51611 145470 239801
rect 210306 236315 210366 243649
rect 210498 236463 210558 243649
rect 268098 243453 268158 243649
rect 405762 243567 405822 268701
rect 405951 268282 406017 268283
rect 405951 268218 405952 268282
rect 406016 268218 406017 268282
rect 405951 268217 406017 268218
rect 405954 247563 406014 268217
rect 405951 247562 406017 247563
rect 405951 247498 405952 247562
rect 406016 247498 406017 247562
rect 405951 247497 406017 247498
rect 406146 247116 406206 271769
rect 406719 271538 406785 271539
rect 406719 271474 406720 271538
rect 406784 271474 406785 271538
rect 406719 271473 406785 271474
rect 406335 270946 406401 270947
rect 406335 270882 406336 270946
rect 406400 270882 406401 270946
rect 406335 270881 406401 270882
rect 405906 247056 406206 247116
rect 405906 246820 405966 247056
rect 406143 246822 406209 246823
rect 405906 246760 406014 246820
rect 405954 243567 406014 246760
rect 406143 246758 406144 246822
rect 406208 246820 406209 246822
rect 406338 246820 406398 270881
rect 406527 270798 406593 270799
rect 406527 270734 406528 270798
rect 406592 270734 406593 270798
rect 406527 270733 406593 270734
rect 406530 246823 406590 270733
rect 406722 246971 406782 271473
rect 406911 271242 406977 271243
rect 406911 271178 406912 271242
rect 406976 271178 406977 271242
rect 406911 271177 406977 271178
rect 406914 246971 406974 271177
rect 407103 264878 407169 264879
rect 407103 264814 407104 264878
rect 407168 264876 407169 264878
rect 407168 264816 407358 264876
rect 407168 264814 407169 264816
rect 407103 264813 407169 264814
rect 407103 264582 407169 264583
rect 407103 264518 407104 264582
rect 407168 264518 407169 264582
rect 407103 264517 407169 264518
rect 407106 247119 407166 264517
rect 407103 247118 407169 247119
rect 407103 247054 407104 247118
rect 407168 247054 407169 247118
rect 407103 247053 407169 247054
rect 406719 246970 406785 246971
rect 406719 246906 406720 246970
rect 406784 246906 406785 246970
rect 406719 246905 406785 246906
rect 406911 246970 406977 246971
rect 406911 246906 406912 246970
rect 406976 246906 406977 246970
rect 406911 246905 406977 246906
rect 406208 246760 406398 246820
rect 406527 246822 406593 246823
rect 406208 246758 406209 246760
rect 406143 246757 406209 246758
rect 406527 246758 406528 246822
rect 406592 246758 406593 246822
rect 406527 246757 406593 246758
rect 406719 246822 406785 246823
rect 406719 246758 406720 246822
rect 406784 246783 406785 246822
rect 407298 246783 407358 264816
rect 407490 246823 407550 273397
rect 409023 273166 409089 273167
rect 409023 273102 409024 273166
rect 409088 273102 409089 273166
rect 409023 273101 409089 273102
rect 408063 271982 408129 271983
rect 408063 271918 408064 271982
rect 408128 271918 408129 271982
rect 408063 271917 408129 271918
rect 407871 271094 407937 271095
rect 407871 271030 407872 271094
rect 407936 271030 407937 271094
rect 407871 271029 407937 271030
rect 407679 264878 407745 264879
rect 407679 264814 407680 264878
rect 407744 264814 407745 264878
rect 407679 264813 407745 264814
rect 407682 247859 407742 264813
rect 407679 247858 407745 247859
rect 407679 247794 407680 247858
rect 407744 247794 407745 247858
rect 407679 247793 407745 247794
rect 407874 247267 407934 271029
rect 407871 247266 407937 247267
rect 407871 247202 407872 247266
rect 407936 247202 407937 247266
rect 407871 247201 407937 247202
rect 406784 246758 407358 246783
rect 406719 246757 407358 246758
rect 407487 246822 407553 246823
rect 407487 246758 407488 246822
rect 407552 246758 407553 246822
rect 407487 246757 407553 246758
rect 406722 246723 407358 246757
rect 405759 243566 405825 243567
rect 405759 243502 405760 243566
rect 405824 243502 405825 243566
rect 405759 243501 405825 243502
rect 405951 243566 406017 243567
rect 405951 243502 405952 243566
rect 406016 243502 406017 243566
rect 405951 243501 406017 243502
rect 267906 243393 268158 243453
rect 267906 243271 267966 243393
rect 210687 243270 210753 243271
rect 210687 243206 210688 243270
rect 210752 243206 210753 243270
rect 210687 243205 210753 243206
rect 267903 243270 267969 243271
rect 267903 243206 267904 243270
rect 267968 243206 267969 243270
rect 267903 243205 267969 243206
rect 268098 243208 268350 243268
rect 210690 236611 210750 243205
rect 210879 243122 210945 243123
rect 210879 243058 210880 243122
rect 210944 243058 210945 243122
rect 210879 243057 210945 243058
rect 210882 236759 210942 243057
rect 268098 242975 268158 243208
rect 268290 243123 268350 243208
rect 408066 243123 408126 271917
rect 408255 264878 408321 264879
rect 408255 264814 408256 264878
rect 408320 264814 408321 264878
rect 408255 264813 408321 264814
rect 408258 243419 408318 264813
rect 408450 264731 408510 265283
rect 408447 264730 408513 264731
rect 408447 264666 408448 264730
rect 408512 264666 408513 264730
rect 408447 264665 408513 264666
rect 408447 247710 408513 247711
rect 408447 247646 408448 247710
rect 408512 247646 408513 247710
rect 408447 247645 408513 247646
rect 408450 247119 408510 247645
rect 408639 247266 408705 247267
rect 408639 247202 408640 247266
rect 408704 247202 408705 247266
rect 408639 247201 408705 247202
rect 408447 247118 408513 247119
rect 408447 247054 408448 247118
rect 408512 247054 408513 247118
rect 408447 247053 408513 247054
rect 408642 246823 408702 247201
rect 408639 246822 408705 246823
rect 408639 246758 408640 246822
rect 408704 246758 408705 246822
rect 408639 246757 408705 246758
rect 408255 243418 408321 243419
rect 408255 243354 408256 243418
rect 408320 243354 408321 243418
rect 408255 243353 408321 243354
rect 409026 243271 409086 273101
rect 410559 273018 410625 273019
rect 410559 272954 410560 273018
rect 410624 272954 410625 273018
rect 410559 272953 410625 272954
rect 409791 272278 409857 272279
rect 409791 272214 409792 272278
rect 409856 272214 409857 272278
rect 409791 272213 409857 272214
rect 409407 271242 409473 271243
rect 409407 271178 409408 271242
rect 409472 271178 409473 271242
rect 409407 271177 409473 271178
rect 409410 246971 409470 271177
rect 409599 264878 409665 264879
rect 409599 264814 409600 264878
rect 409664 264814 409665 264878
rect 409599 264813 409665 264814
rect 409602 247415 409662 264813
rect 409599 247414 409665 247415
rect 409599 247350 409600 247414
rect 409664 247350 409665 247414
rect 409599 247349 409665 247350
rect 409794 247119 409854 272213
rect 409983 272130 410049 272131
rect 409983 272066 409984 272130
rect 410048 272066 410049 272130
rect 409983 272065 410049 272066
rect 409791 247118 409857 247119
rect 409791 247054 409792 247118
rect 409856 247054 409857 247118
rect 409791 247053 409857 247054
rect 409407 246970 409473 246971
rect 409407 246906 409408 246970
rect 409472 246906 409473 246970
rect 409407 246905 409473 246906
rect 409986 246823 410046 272065
rect 410367 271834 410433 271835
rect 410367 271770 410368 271834
rect 410432 271770 410433 271834
rect 410367 271769 410433 271770
rect 410175 271686 410241 271687
rect 410175 271622 410176 271686
rect 410240 271622 410241 271686
rect 410175 271621 410241 271622
rect 410178 246971 410238 271621
rect 410175 246970 410241 246971
rect 410175 246906 410176 246970
rect 410240 246906 410241 246970
rect 410175 246905 410241 246906
rect 410370 246823 410430 271769
rect 409983 246822 410049 246823
rect 409983 246758 409984 246822
rect 410048 246758 410049 246822
rect 409983 246757 410049 246758
rect 410367 246822 410433 246823
rect 410367 246758 410368 246822
rect 410432 246758 410433 246822
rect 410367 246757 410433 246758
rect 410562 246783 410622 272953
rect 411135 272722 411201 272723
rect 411135 272658 411136 272722
rect 411200 272658 411201 272722
rect 411135 272657 411201 272658
rect 410751 271538 410817 271539
rect 410751 271474 410752 271538
rect 410816 271474 410817 271538
rect 410751 271473 410817 271474
rect 410754 247267 410814 271473
rect 410943 264878 411009 264879
rect 410943 264814 410944 264878
rect 411008 264814 411009 264878
rect 410943 264813 411009 264814
rect 410946 247711 411006 264813
rect 410943 247710 411009 247711
rect 410943 247646 410944 247710
rect 411008 247646 411009 247710
rect 410943 247645 411009 247646
rect 410751 247266 410817 247267
rect 410751 247202 410752 247266
rect 410816 247202 410817 247266
rect 410751 247201 410817 247202
rect 411138 246971 411198 272657
rect 499647 270354 499713 270355
rect 499647 270290 499648 270354
rect 499712 270290 499713 270354
rect 499647 270289 499713 270290
rect 499650 269427 499710 270289
rect 499458 269367 499710 269427
rect 499458 268727 499518 269367
rect 499455 268726 499521 268727
rect 499455 268662 499456 268726
rect 499520 268662 499521 268726
rect 499455 268661 499521 268662
rect 411327 264730 411393 264731
rect 411327 264666 411328 264730
rect 411392 264666 411393 264730
rect 411327 264665 411393 264666
rect 411135 246970 411201 246971
rect 411135 246906 411136 246970
rect 411200 246906 411201 246970
rect 411135 246905 411201 246906
rect 411330 246823 411390 264665
rect 673986 246823 674046 284645
rect 674178 283675 674238 310693
rect 675330 290039 675390 329489
rect 676674 326891 676734 345177
rect 676671 326890 676737 326891
rect 676671 326826 676672 326890
rect 676736 326826 676737 326890
rect 676671 326825 676737 326826
rect 677058 313719 677118 357609
rect 677250 356639 677310 373263
rect 677439 357674 677505 357675
rect 677439 357610 677440 357674
rect 677504 357610 677505 357674
rect 677439 357609 677505 357610
rect 677247 356638 677313 356639
rect 677247 356574 677248 356638
rect 677312 356574 677313 356638
rect 677247 356573 677313 356574
rect 677055 313718 677121 313719
rect 677055 313654 677056 313718
rect 677120 313654 677121 313718
rect 677055 313653 677121 313654
rect 677250 312717 677310 356573
rect 677058 312657 677310 312717
rect 677058 311499 677118 312657
rect 677247 312534 677313 312535
rect 677247 312470 677248 312534
rect 677312 312470 677313 312534
rect 677247 312469 677313 312470
rect 677055 311498 677121 311499
rect 677055 311434 677056 311498
rect 677120 311434 677121 311498
rect 677055 311433 677121 311434
rect 675903 299510 675969 299511
rect 675903 299446 675904 299510
rect 675968 299446 675969 299510
rect 675903 299445 675969 299446
rect 675327 290038 675393 290039
rect 675327 289974 675328 290038
rect 675392 289974 675393 290038
rect 675327 289973 675393 289974
rect 674367 285006 674433 285007
rect 674367 284942 674368 285006
rect 674432 284942 674433 285006
rect 674367 284941 674433 284942
rect 674175 283674 674241 283675
rect 674175 283610 674176 283674
rect 674240 283610 674241 283674
rect 674175 283609 674241 283610
rect 674175 264138 674241 264139
rect 674175 264074 674176 264138
rect 674240 264074 674241 264138
rect 674175 264073 674241 264074
rect 410943 246822 411009 246823
rect 410943 246783 410944 246822
rect 410562 246758 410944 246783
rect 411008 246758 411009 246822
rect 410562 246757 411009 246758
rect 411327 246822 411393 246823
rect 411327 246758 411328 246822
rect 411392 246758 411393 246822
rect 411327 246757 411393 246758
rect 673983 246822 674049 246823
rect 673983 246758 673984 246822
rect 674048 246758 674049 246822
rect 673983 246757 674049 246758
rect 410562 246723 411006 246757
rect 673986 245343 674046 246757
rect 673983 245342 674049 245343
rect 673983 245278 673984 245342
rect 674048 245278 674049 245342
rect 673983 245277 674049 245278
rect 674178 243567 674238 264073
rect 674370 244751 674430 284941
rect 675906 284859 675966 299445
rect 676671 299362 676737 299363
rect 676671 299298 676672 299362
rect 676736 299298 676737 299362
rect 676671 299297 676737 299298
rect 675903 284858 675969 284859
rect 675903 284794 675904 284858
rect 675968 284794 675969 284858
rect 675903 284793 675969 284794
rect 676674 281899 676734 299297
rect 676671 281898 676737 281899
rect 676671 281834 676672 281898
rect 676736 281834 676737 281898
rect 676671 281833 676737 281834
rect 677058 267099 677118 311433
rect 677250 268727 677310 312469
rect 677442 312091 677502 357609
rect 677439 312090 677505 312091
rect 677439 312026 677440 312090
rect 677504 312026 677505 312090
rect 677439 312025 677505 312026
rect 677247 268726 677313 268727
rect 677247 268662 677248 268726
rect 677312 268662 677313 268726
rect 677247 268661 677313 268662
rect 677247 267690 677313 267691
rect 677247 267626 677248 267690
rect 677312 267626 677313 267690
rect 677247 267625 677313 267626
rect 676863 267098 676929 267099
rect 676863 267034 676864 267098
rect 676928 267034 676929 267098
rect 676863 267033 676929 267034
rect 677055 267098 677121 267099
rect 677055 267034 677056 267098
rect 677120 267034 677121 267098
rect 677055 267033 677121 267034
rect 675711 253334 675777 253335
rect 675711 253270 675712 253334
rect 675776 253270 675777 253334
rect 675711 253269 675777 253270
rect 674367 244750 674433 244751
rect 674367 244686 674368 244750
rect 674432 244686 674433 244750
rect 674367 244685 674433 244686
rect 675327 244750 675393 244751
rect 675327 244686 675328 244750
rect 675392 244686 675393 244750
rect 675327 244685 675393 244686
rect 674370 243863 674430 244685
rect 674367 243862 674433 243863
rect 674367 243798 674368 243862
rect 674432 243798 674433 243862
rect 674367 243797 674433 243798
rect 674175 243566 674241 243567
rect 674175 243502 674176 243566
rect 674240 243502 674241 243566
rect 674175 243501 674241 243502
rect 409023 243270 409089 243271
rect 409023 243206 409024 243270
rect 409088 243206 409089 243270
rect 409023 243205 409089 243206
rect 268287 243122 268353 243123
rect 268287 243058 268288 243122
rect 268352 243058 268353 243122
rect 268287 243057 268353 243058
rect 288063 243122 288129 243123
rect 288063 243058 288064 243122
rect 288128 243058 288129 243122
rect 288063 243057 288129 243058
rect 408063 243122 408129 243123
rect 408063 243058 408064 243122
rect 408128 243058 408129 243122
rect 408063 243057 408129 243058
rect 268095 242974 268161 242975
rect 268095 242910 268096 242974
rect 268160 242910 268161 242974
rect 268095 242909 268161 242910
rect 227391 242826 227457 242827
rect 227391 242762 227392 242826
rect 227456 242787 227457 242826
rect 227456 242762 228030 242787
rect 227391 242761 228030 242762
rect 227394 242727 228030 242761
rect 227970 242383 228030 242727
rect 247359 242530 247425 242531
rect 247359 242466 247360 242530
rect 247424 242466 247425 242530
rect 247359 242465 247425 242466
rect 227967 242382 228033 242383
rect 227967 242318 227968 242382
rect 228032 242318 228033 242382
rect 227967 242317 228033 242318
rect 247362 242121 247422 242465
rect 288066 242121 288126 243057
rect 247362 242061 247806 242121
rect 247746 241495 247806 242061
rect 267522 242061 268158 242121
rect 267522 241495 267582 242061
rect 268098 241791 268158 242061
rect 287874 242061 288126 242121
rect 287874 241791 287934 242061
rect 268095 241790 268161 241791
rect 268095 241726 268096 241790
rect 268160 241726 268161 241790
rect 268095 241725 268161 241726
rect 287871 241790 287937 241791
rect 287871 241726 287872 241790
rect 287936 241726 287937 241790
rect 287871 241725 287937 241726
rect 247743 241494 247809 241495
rect 247743 241430 247744 241494
rect 247808 241430 247809 241494
rect 247743 241429 247809 241430
rect 267519 241494 267585 241495
rect 267519 241430 267520 241494
rect 267584 241430 267585 241494
rect 267519 241429 267585 241430
rect 211071 237794 211137 237795
rect 211071 237730 211072 237794
rect 211136 237730 211137 237794
rect 211071 237729 211137 237730
rect 210879 236758 210945 236759
rect 210879 236694 210880 236758
rect 210944 236694 210945 236758
rect 210879 236693 210945 236694
rect 210687 236610 210753 236611
rect 210687 236546 210688 236610
rect 210752 236546 210753 236610
rect 210687 236545 210753 236546
rect 210495 236462 210561 236463
rect 210495 236398 210496 236462
rect 210560 236398 210561 236462
rect 210495 236397 210561 236398
rect 210303 236314 210369 236315
rect 210303 236250 210304 236314
rect 210368 236250 210369 236314
rect 210303 236249 210369 236250
rect 210879 233354 210945 233355
rect 210879 233290 210880 233354
rect 210944 233290 210945 233354
rect 210879 233289 210945 233290
rect 145599 218998 145665 218999
rect 145599 218934 145600 218998
rect 145664 218934 145665 218998
rect 145599 218933 145665 218934
rect 145407 51610 145473 51611
rect 145407 51546 145408 51610
rect 145472 51546 145473 51610
rect 145407 51545 145473 51546
rect 145602 51463 145662 218933
rect 210495 217074 210561 217075
rect 210495 217010 210496 217074
rect 210560 217010 210561 217074
rect 210495 217009 210561 217010
rect 145791 216482 145857 216483
rect 145791 216418 145792 216482
rect 145856 216418 145857 216482
rect 145791 216417 145857 216418
rect 145599 51462 145665 51463
rect 145599 51398 145600 51462
rect 145664 51398 145665 51462
rect 145599 51397 145665 51398
rect 145794 51315 145854 216417
rect 210498 191619 210558 217009
rect 210495 191618 210561 191619
rect 210495 191554 210496 191618
rect 210560 191554 210561 191618
rect 210495 191553 210561 191554
rect 210882 181515 210942 233289
rect 211074 217075 211134 237729
rect 302466 236733 302910 236793
rect 302466 236611 302526 236733
rect 302850 236611 302910 236733
rect 302463 236610 302529 236611
rect 302463 236546 302464 236610
rect 302528 236546 302529 236610
rect 302463 236545 302529 236546
rect 302847 236610 302913 236611
rect 302847 236546 302848 236610
rect 302912 236546 302913 236610
rect 302847 236545 302913 236546
rect 211455 234686 211521 234687
rect 211455 234622 211456 234686
rect 211520 234622 211521 234686
rect 211455 234621 211521 234622
rect 211458 218145 211518 234621
rect 636927 234094 636993 234095
rect 636927 234030 636928 234094
rect 636992 234030 636993 234094
rect 636927 234029 636993 234030
rect 212415 233650 212481 233651
rect 212415 233586 212416 233650
rect 212480 233586 212481 233650
rect 212415 233585 212481 233586
rect 212223 233502 212289 233503
rect 212223 233438 212224 233502
rect 212288 233438 212289 233502
rect 212223 233437 212289 233438
rect 211458 218085 211710 218145
rect 211071 217074 211137 217075
rect 211071 217010 211072 217074
rect 211136 217010 211137 217074
rect 211071 217009 211137 217010
rect 211071 191618 211137 191619
rect 211071 191554 211072 191618
rect 211136 191554 211137 191618
rect 211071 191553 211137 191554
rect 211074 185511 211134 191553
rect 211650 187509 211710 218085
rect 211458 187449 211710 187509
rect 211458 186177 211518 187449
rect 211458 186117 212094 186177
rect 211074 185451 211518 185511
rect 210882 181455 211326 181515
rect 211266 162201 211326 181455
rect 211074 162141 211326 162201
rect 211074 161575 211134 162141
rect 211071 161574 211137 161575
rect 211071 161510 211072 161574
rect 211136 161510 211137 161574
rect 211071 161509 211137 161510
rect 211458 160869 211518 185451
rect 212034 176187 212094 186117
rect 210882 160809 211518 160869
rect 211842 176127 212094 176187
rect 210495 158466 210561 158467
rect 210495 158402 210496 158466
rect 210560 158402 210561 158466
rect 210495 158401 210561 158402
rect 210498 141447 210558 158401
rect 210882 141595 210942 160809
rect 211842 148215 211902 176127
rect 211650 148155 211902 148215
rect 211650 146883 211710 148155
rect 211458 146823 211710 146883
rect 210879 141594 210945 141595
rect 210879 141530 210880 141594
rect 210944 141530 210945 141594
rect 210879 141529 210945 141530
rect 210495 141446 210561 141447
rect 210495 141382 210496 141446
rect 210560 141382 210561 141446
rect 210495 141381 210561 141382
rect 210879 141298 210945 141299
rect 210879 141234 210880 141298
rect 210944 141234 210945 141298
rect 210879 141233 210945 141234
rect 210687 138338 210753 138339
rect 210687 138274 210688 138338
rect 210752 138274 210753 138338
rect 210687 138273 210753 138274
rect 210495 126202 210561 126203
rect 210495 126138 210496 126202
rect 210560 126138 210561 126202
rect 210495 126137 210561 126138
rect 210498 118063 210558 126137
rect 210495 118062 210561 118063
rect 210495 117998 210496 118062
rect 210560 117998 210561 118062
rect 210495 117997 210561 117998
rect 210690 112291 210750 138273
rect 210882 129163 210942 141233
rect 211458 140889 211518 146823
rect 211266 140829 211518 140889
rect 211266 129567 211326 140829
rect 211074 129507 211326 129567
rect 210879 129162 210945 129163
rect 210879 129098 210880 129162
rect 210944 129098 210945 129162
rect 210879 129097 210945 129098
rect 211074 128124 211134 129507
rect 211074 128064 211326 128124
rect 211266 122241 211326 128064
rect 211074 122181 211326 122241
rect 211074 121171 211134 122181
rect 211071 121170 211137 121171
rect 211071 121106 211072 121170
rect 211136 121106 211137 121170
rect 211071 121105 211137 121106
rect 210879 118062 210945 118063
rect 210879 117998 210880 118062
rect 210944 117998 210945 118062
rect 210879 117997 210945 117998
rect 210687 112290 210753 112291
rect 210687 112226 210688 112290
rect 210752 112226 210753 112290
rect 210687 112225 210753 112226
rect 210111 86982 210177 86983
rect 210111 86918 210112 86982
rect 210176 86918 210177 86982
rect 210111 86917 210177 86918
rect 210114 77807 210174 86917
rect 210882 86539 210942 117997
rect 211071 113770 211137 113771
rect 211071 113706 211072 113770
rect 211136 113768 211137 113770
rect 211136 113708 212094 113768
rect 211136 113706 211137 113708
rect 211071 113705 211137 113706
rect 211071 112290 211137 112291
rect 211071 112226 211072 112290
rect 211136 112251 211137 112290
rect 211136 112226 211326 112251
rect 211071 112225 211326 112226
rect 211074 112191 211326 112225
rect 211266 100929 211326 112191
rect 211266 100869 211902 100929
rect 210687 86538 210753 86539
rect 210687 86474 210688 86538
rect 210752 86474 210753 86538
rect 210687 86473 210753 86474
rect 210879 86538 210945 86539
rect 210879 86474 210880 86538
rect 210944 86474 210945 86538
rect 210879 86473 210945 86474
rect 210111 77806 210177 77807
rect 210111 77742 210112 77806
rect 210176 77742 210177 77806
rect 210111 77741 210177 77742
rect 210690 66297 210750 86473
rect 211842 79617 211902 100869
rect 211266 79557 211902 79617
rect 210690 66237 211134 66297
rect 210879 58270 210945 58271
rect 210879 58206 210880 58270
rect 210944 58206 210945 58270
rect 210879 58205 210945 58206
rect 210687 57678 210753 57679
rect 210687 57614 210688 57678
rect 210752 57614 210753 57678
rect 210687 57613 210753 57614
rect 210690 54127 210750 57613
rect 210687 54126 210753 54127
rect 210687 54062 210688 54126
rect 210752 54062 210753 54126
rect 210687 54061 210753 54062
rect 210882 53979 210942 58205
rect 210879 53978 210945 53979
rect 210879 53914 210880 53978
rect 210944 53914 210945 53978
rect 210879 53913 210945 53914
rect 211074 53831 211134 66237
rect 211266 54275 211326 79557
rect 212034 77804 212094 113708
rect 211842 77744 212094 77804
rect 211263 54274 211329 54275
rect 211263 54210 211264 54274
rect 211328 54210 211329 54274
rect 211263 54209 211329 54210
rect 211071 53830 211137 53831
rect 211071 53766 211072 53830
rect 211136 53766 211137 53830
rect 211071 53765 211137 53766
rect 211842 53535 211902 77744
rect 212226 63633 212286 233437
rect 212034 63573 212286 63633
rect 212034 53683 212094 63573
rect 212031 53682 212097 53683
rect 212031 53618 212032 53682
rect 212096 53618 212097 53682
rect 212031 53617 212097 53618
rect 211839 53534 211905 53535
rect 211839 53470 211840 53534
rect 211904 53470 211905 53534
rect 211839 53469 211905 53470
rect 212418 53387 212478 233585
rect 212607 233502 212673 233503
rect 212607 233438 212608 233502
rect 212672 233438 212673 233502
rect 212607 233437 212673 233438
rect 212799 233502 212865 233503
rect 212799 233438 212800 233502
rect 212864 233438 212865 233502
rect 212799 233437 212865 233438
rect 212610 54127 212670 233437
rect 212607 54126 212673 54127
rect 212607 54062 212608 54126
rect 212672 54062 212673 54126
rect 212607 54061 212673 54062
rect 212415 53386 212481 53387
rect 212415 53322 212416 53386
rect 212480 53322 212481 53386
rect 212415 53321 212481 53322
rect 212802 53239 212862 233437
rect 212799 53238 212865 53239
rect 212799 53174 212800 53238
rect 212864 53174 212865 53238
rect 212799 53173 212865 53174
rect 636930 51759 636990 234029
rect 637887 233946 637953 233947
rect 637887 233882 637888 233946
rect 637952 233882 637953 233946
rect 637887 233881 637953 233882
rect 637503 233798 637569 233799
rect 637503 233734 637504 233798
rect 637568 233734 637569 233798
rect 637503 233733 637569 233734
rect 637119 233650 637185 233651
rect 637119 233586 637120 233650
rect 637184 233586 637185 233650
rect 637119 233585 637185 233586
rect 637311 233650 637377 233651
rect 637311 233586 637312 233650
rect 637376 233586 637377 233650
rect 637311 233585 637377 233586
rect 636927 51758 636993 51759
rect 636927 51694 636928 51758
rect 636992 51694 636993 51758
rect 636927 51693 636993 51694
rect 145791 51314 145857 51315
rect 145791 51250 145792 51314
rect 145856 51250 145857 51314
rect 145791 51249 145857 51250
rect 637122 50427 637182 233585
rect 637314 51907 637374 233585
rect 637506 52055 637566 233733
rect 637695 233502 637761 233503
rect 637695 233438 637696 233502
rect 637760 233438 637761 233502
rect 637695 233437 637761 233438
rect 637698 52351 637758 233437
rect 637695 52350 637761 52351
rect 637695 52286 637696 52350
rect 637760 52286 637761 52350
rect 637695 52285 637761 52286
rect 637890 52203 637950 233881
rect 674367 220552 674433 220553
rect 674367 220488 674368 220552
rect 674432 220488 674433 220552
rect 674367 220487 674433 220488
rect 674175 218924 674241 218925
rect 674175 218860 674176 218924
rect 674240 218860 674241 218924
rect 674175 218859 674241 218860
rect 674178 198427 674238 218859
rect 674175 198426 674241 198427
rect 674175 198362 674176 198426
rect 674240 198362 674241 198426
rect 674175 198361 674241 198362
rect 674370 193543 674430 220487
rect 675330 199315 675390 244685
rect 675519 238978 675585 238979
rect 675519 238914 675520 238978
rect 675584 238914 675585 238978
rect 675519 238913 675585 238914
rect 675327 199314 675393 199315
rect 675327 199250 675328 199314
rect 675392 199250 675393 199314
rect 675327 199249 675393 199250
rect 674367 193542 674433 193543
rect 674367 193478 674368 193542
rect 674432 193478 674433 193542
rect 674367 193477 674433 193478
rect 674367 173858 674433 173859
rect 674367 173794 674368 173858
rect 674432 173794 674433 173858
rect 674367 173793 674433 173794
rect 673983 170602 674049 170603
rect 673983 170538 673984 170602
rect 674048 170538 674049 170602
rect 673983 170537 674049 170538
rect 673986 151955 674046 170537
rect 674370 153435 674430 173793
rect 674559 170898 674625 170899
rect 674559 170834 674560 170898
rect 674624 170834 674625 170898
rect 674559 170833 674625 170834
rect 674367 153434 674433 153435
rect 674367 153370 674368 153434
rect 674432 153370 674433 153434
rect 674367 153369 674433 153370
rect 673983 151954 674049 151955
rect 673983 151890 673984 151954
rect 674048 151890 674049 151954
rect 673983 151889 674049 151890
rect 674562 150327 674622 170833
rect 675330 155211 675390 199249
rect 675522 198723 675582 238913
rect 675714 236907 675774 253269
rect 675903 253186 675969 253187
rect 675903 253122 675904 253186
rect 675968 253122 675969 253186
rect 675903 253121 675969 253122
rect 675906 238683 675966 253121
rect 675903 238682 675969 238683
rect 675903 238618 675904 238682
rect 675968 238618 675969 238682
rect 675903 238617 675969 238618
rect 676866 237647 676926 267033
rect 677058 237795 677118 267033
rect 677055 237794 677121 237795
rect 677055 237730 677056 237794
rect 677120 237730 677121 237794
rect 677055 237729 677121 237730
rect 676863 237646 676929 237647
rect 676863 237582 676864 237646
rect 676928 237582 676929 237646
rect 676863 237581 676929 237582
rect 675711 236906 675777 236907
rect 675711 236842 675712 236906
rect 675776 236842 675777 236906
rect 675711 236841 675777 236842
rect 676866 222403 676926 237581
rect 676863 222402 676929 222403
rect 676863 222338 676864 222402
rect 676928 222338 676929 222402
rect 676863 222337 676929 222338
rect 677058 221811 677118 237729
rect 677250 223587 677310 267625
rect 677442 267543 677502 312025
rect 677439 267542 677505 267543
rect 677439 267478 677440 267542
rect 677504 267478 677505 267542
rect 677439 267477 677505 267478
rect 677247 223586 677313 223587
rect 677247 223522 677248 223586
rect 677312 223522 677313 223586
rect 677247 223521 677313 223522
rect 677247 222402 677313 222403
rect 677247 222338 677248 222402
rect 677312 222338 677313 222402
rect 677247 222337 677313 222338
rect 677055 221810 677121 221811
rect 677055 221746 677056 221810
rect 677120 221746 677121 221810
rect 677055 221745 677121 221746
rect 676479 210266 676545 210267
rect 676479 210202 676480 210266
rect 676544 210202 676545 210266
rect 676479 210201 676545 210202
rect 675519 198722 675585 198723
rect 675519 198658 675520 198722
rect 675584 198658 675585 198722
rect 675519 198657 675585 198658
rect 675327 155210 675393 155211
rect 675327 155146 675328 155210
rect 675392 155146 675393 155210
rect 675327 155145 675393 155146
rect 674559 150326 674625 150327
rect 674559 150262 674560 150326
rect 674624 150262 674625 150326
rect 674559 150261 674625 150262
rect 673983 128718 674049 128719
rect 673983 128654 673984 128718
rect 674048 128654 674049 128718
rect 673983 128653 674049 128654
rect 673986 108147 674046 128653
rect 674175 126054 674241 126055
rect 674175 125990 674176 126054
rect 674240 125990 674241 126054
rect 674175 125989 674241 125990
rect 673983 108146 674049 108147
rect 673983 108082 673984 108146
rect 674048 108082 674049 108146
rect 673983 108081 674049 108082
rect 674178 105187 674238 125989
rect 675330 110071 675390 155145
rect 675522 154471 675582 198657
rect 676482 195319 676542 210201
rect 676671 210118 676737 210119
rect 676671 210054 676672 210118
rect 676736 210054 676737 210118
rect 676671 210053 676737 210054
rect 676479 195318 676545 195319
rect 676479 195254 676480 195318
rect 676544 195254 676545 195318
rect 676479 195253 676545 195254
rect 676674 191619 676734 210053
rect 676863 206418 676929 206419
rect 676863 206354 676864 206418
rect 676928 206354 676929 206418
rect 676863 206353 676929 206354
rect 676671 191618 676737 191619
rect 676671 191554 676672 191618
rect 676736 191554 676737 191618
rect 676671 191553 676737 191554
rect 676866 177411 676926 206353
rect 676863 177410 676929 177411
rect 676863 177346 676864 177410
rect 676928 177346 676929 177410
rect 676863 177345 676929 177346
rect 677058 176375 677118 221745
rect 677250 178447 677310 222337
rect 677631 221810 677697 221811
rect 677631 221746 677632 221810
rect 677696 221746 677697 221810
rect 677631 221745 677697 221746
rect 677634 206419 677694 221745
rect 677631 206418 677697 206419
rect 677631 206354 677632 206418
rect 677696 206354 677697 206418
rect 677631 206353 677697 206354
rect 677247 178446 677313 178447
rect 677247 178382 677248 178446
rect 677312 178382 677313 178446
rect 677247 178381 677313 178382
rect 677247 177410 677313 177411
rect 677247 177346 677248 177410
rect 677312 177346 677313 177410
rect 677247 177345 677313 177346
rect 677055 176374 677121 176375
rect 677055 176310 677056 176374
rect 677120 176310 677121 176374
rect 677055 176309 677121 176310
rect 675711 161574 675777 161575
rect 675711 161510 675712 161574
rect 675776 161510 675777 161574
rect 675711 161509 675777 161510
rect 675519 154470 675585 154471
rect 675519 154406 675520 154470
rect 675584 154406 675585 154470
rect 675519 154405 675585 154406
rect 675327 110070 675393 110071
rect 675327 110006 675328 110070
rect 675392 110006 675393 110070
rect 675327 110005 675393 110006
rect 675522 109331 675582 154405
rect 675714 148551 675774 161509
rect 676671 161426 676737 161427
rect 676671 161362 676672 161426
rect 676736 161362 676737 161426
rect 676671 161361 676737 161362
rect 675711 148550 675777 148551
rect 675711 148486 675712 148550
rect 675776 148486 675777 148550
rect 675711 148485 675777 148486
rect 676674 146627 676734 161361
rect 676671 146626 676737 146627
rect 676671 146562 676672 146626
rect 676736 146562 676737 146626
rect 676671 146561 676737 146562
rect 677058 131827 677118 176309
rect 677250 133455 677310 177345
rect 677439 176966 677505 176967
rect 677439 176902 677440 176966
rect 677504 176902 677505 176966
rect 677439 176901 677505 176902
rect 677247 133454 677313 133455
rect 677247 133390 677248 133454
rect 677312 133390 677313 133454
rect 677247 133389 677313 133390
rect 677442 132271 677502 176901
rect 677439 132270 677505 132271
rect 677439 132206 677440 132270
rect 677504 132206 677505 132270
rect 677439 132205 677505 132206
rect 677055 131826 677121 131827
rect 677055 131762 677056 131826
rect 677120 131762 677121 131826
rect 677055 131761 677121 131762
rect 676671 118062 676737 118063
rect 676671 117998 676672 118062
rect 676736 117998 676737 118062
rect 676671 117997 676737 117998
rect 675903 117914 675969 117915
rect 675903 117850 675904 117914
rect 675968 117850 675969 117914
rect 675903 117849 675969 117850
rect 675519 109330 675585 109331
rect 675519 109266 675520 109330
rect 675584 109266 675585 109330
rect 675519 109265 675585 109266
rect 674175 105186 674241 105187
rect 674175 105122 674176 105186
rect 674240 105122 674241 105186
rect 674175 105121 674241 105122
rect 675906 103263 675966 117849
rect 675903 103262 675969 103263
rect 675903 103198 675904 103262
rect 675968 103198 675969 103262
rect 675903 103197 675969 103198
rect 676674 101487 676734 117997
rect 676671 101486 676737 101487
rect 676671 101422 676672 101486
rect 676736 101422 676737 101486
rect 676671 101421 676737 101422
rect 637887 52202 637953 52203
rect 637887 52138 637888 52202
rect 637952 52138 637953 52202
rect 637887 52137 637953 52138
rect 637503 52054 637569 52055
rect 637503 51990 637504 52054
rect 637568 51990 637569 52054
rect 637503 51989 637569 51990
rect 637311 51906 637377 51907
rect 637311 51842 637312 51906
rect 637376 51842 637377 51906
rect 637311 51841 637377 51842
rect 637119 50426 637185 50427
rect 637119 50362 637120 50426
rect 637184 50362 637185 50426
rect 637119 50361 637185 50362
rect 520383 49094 520449 49095
rect 520383 49030 520384 49094
rect 520448 49030 520449 49094
rect 520383 49029 520449 49030
rect 302463 45246 302529 45247
rect 302463 45182 302464 45246
rect 302528 45182 302529 45246
rect 302463 45181 302529 45182
rect 302466 43323 302526 45181
rect 362943 45098 363009 45099
rect 362943 45034 362944 45098
rect 363008 45034 363009 45098
rect 362943 45033 363009 45034
rect 362946 43323 363006 45033
rect 302463 43322 302529 43323
rect 302463 43258 302464 43322
rect 302528 43258 302529 43322
rect 302463 43257 302529 43258
rect 362943 43322 363009 43323
rect 362943 43258 362944 43322
rect 363008 43258 363009 43322
rect 362943 43257 363009 43258
rect 520386 42139 520446 49029
rect 527103 44950 527169 44951
rect 527103 44886 527104 44950
rect 527168 44886 527169 44950
rect 527103 44885 527169 44886
rect 527106 43323 527166 44885
rect 527103 43322 527169 43323
rect 527103 43258 527104 43322
rect 527168 43258 527169 43322
rect 527103 43257 527169 43258
rect 520383 42138 520449 42139
rect 520383 42074 520384 42138
rect 520448 42074 520449 42138
rect 520383 42073 520449 42074
rect 189951 41842 190017 41843
rect 189951 41778 189952 41842
rect 190016 41778 190017 41842
rect 189951 41777 190017 41778
rect 194943 41842 195009 41843
rect 194943 41778 194944 41842
rect 195008 41778 195009 41842
rect 194943 41777 195009 41778
rect 189954 40807 190014 41777
rect 189951 40806 190017 40807
rect 189951 40742 189952 40806
rect 190016 40742 190017 40806
rect 189951 40741 190017 40742
rect 194946 40659 195006 41777
rect 194943 40658 195009 40659
rect 194943 40594 194944 40658
rect 195008 40594 195009 40658
rect 194943 40593 195009 40594
<< via4 >>
rect 371498 270611 371734 270847
rect 370538 269945 370774 270181
rect 328106 267947 328342 268183
rect 328490 267947 328726 268183
rect 327146 267281 327382 267517
rect 352682 267281 352918 267517
rect 393962 270798 394198 270847
rect 393962 270734 394048 270798
rect 394048 270734 394112 270798
rect 394112 270734 394198 270798
rect 393962 270611 394198 270734
rect 381674 269945 381910 270181
rect 379946 269279 380182 269515
rect 395690 269279 395926 269515
rect 371306 265283 371542 265519
rect 408362 265283 408598 265519
<< metal5 >>
rect 371456 270847 394240 270889
rect 371456 270611 371498 270847
rect 371734 270611 393962 270847
rect 394198 270611 394240 270847
rect 371456 270569 394240 270611
rect 370496 270181 381952 270223
rect 370496 269945 370538 270181
rect 370774 269945 381674 270181
rect 381910 269945 381952 270181
rect 370496 269903 381952 269945
rect 379904 269515 395968 269557
rect 379904 269279 379946 269515
rect 380182 269279 395690 269515
rect 395926 269279 395968 269515
rect 379904 269237 395968 269279
rect 328064 268183 328768 268225
rect 328064 267947 328106 268183
rect 328342 267947 328490 268183
rect 328726 267947 328768 268183
rect 328064 267905 328768 267947
rect 327104 267517 352960 267559
rect 327104 267281 327146 267517
rect 327382 267281 352682 267517
rect 352918 267281 352960 267517
rect 327104 267239 352960 267281
rect 371264 265519 408640 265561
rect 371264 265283 371306 265519
rect 371542 265283 408362 265519
rect 408598 265283 408640 265519
rect 371264 265241 408640 265283
use user_id_programming  user_id_value
timestamp 1608238675
transform 1 0 656624 0 1 80926
box 0 0 7109 7077
use storage  storage
timestamp 1608238675
transform 1 0 52032 0 1 53156
box 38 0 88934 189234
use mgmt_core  soc
timestamp 1608238675
transform 1 0 210434 0 1 53602
box 0 0 430000 180000
use sky130_fd_sc_hvl__lsbufhv2lv_1_wrapped  rstb_level
timestamp 1608238675
transform -1 0 137896 0 -1 51956
box 0 -51 4992 5000
use simple_por  por
timestamp 1608238675
transform 1 0 654146 0 -1 112882
box 25 11 11344 8291
use gpio_control_block  gpio_control_bidir\[1\]
timestamp 1608238675
transform -1 0 708603 0 1 166200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_bidir\[0\]
timestamp 1608238675
transform -1 0 708603 0 1 121000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[36\]
timestamp 1608238675
transform 1 0 8567 0 1 245800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[37\]
timestamp 1608238675
transform 1 0 8567 0 1 202600
box -1620 -364 34000 13964
use mgmt_protect  mgmt_buffers
timestamp 1608238675
transform 1 0 212180 0 1 246836
box -2762 -2778 202678 20730
use gpio_control_block  gpio_control_in\[2\]
timestamp 1608238675
transform -1 0 708603 0 1 211200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[3\]
timestamp 1608238675
transform -1 0 708603 0 1 256400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[33\]
timestamp 1608238675
transform 1 0 8567 0 1 375400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[34\]
timestamp 1608238675
transform 1 0 8567 0 1 332200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[35\]
timestamp 1608238675
transform 1 0 8567 0 1 289000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[4\]
timestamp 1608238675
transform -1 0 708603 0 1 301400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[5\]
timestamp 1608238675
transform -1 0 708603 0 1 346400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[7\]
timestamp 1608238675
transform -1 0 708603 0 1 479800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[6\]
timestamp 1608238675
transform -1 0 708603 0 1 391600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[32\]
timestamp 1608238675
transform 1 0 8567 0 1 418600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[31\]
timestamp 1608238675
transform 1 0 8567 0 1 546200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[30\]
timestamp 1608238675
transform 1 0 8567 0 1 589400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[29\]
timestamp 1608238675
transform 1 0 8567 0 1 632600
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[9\]
timestamp 1608238675
transform -1 0 708603 0 1 568800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[8\]
timestamp 1608238675
transform -1 0 708603 0 1 523800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[10\]
timestamp 1608238675
transform -1 0 708603 0 1 614000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[28\]
timestamp 1608238675
transform 1 0 8567 0 1 675800
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[27\]
timestamp 1608238675
transform 1 0 8567 0 1 719000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[26\]
timestamp 1608238675
transform 1 0 8567 0 1 762200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[13\]
timestamp 1608238675
transform -1 0 708603 0 1 749200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[12\]
timestamp 1608238675
transform -1 0 708603 0 1 704200
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[11\]
timestamp 1608238675
transform -1 0 708603 0 1 659000
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[25\]
timestamp 1608238675
transform 1 0 8567 0 1 805400
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[24\]
timestamp 1608238675
transform 1 0 8567 0 1 931224
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[23\]
timestamp 1608238675
transform 0 1 97200 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[22\]
timestamp 1608238675
transform 0 1 148600 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[21\]
timestamp 1608238675
transform 0 1 200000 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[20\]
timestamp 1608238675
transform 0 1 251400 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[19\]
timestamp 1608238675
transform 0 1 303000 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[18\]
timestamp 1608238675
transform 0 1 353400 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[17\]
timestamp 1608238675
transform 0 1 420800 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[16\]
timestamp 1608238675
transform 0 1 497800 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[15\]
timestamp 1608238675
transform 0 1 549200 -1 0 1029813
box -1620 -364 34000 13964
use gpio_control_block  gpio_control_in\[14\]
timestamp 1608238675
transform -1 0 708603 0 1 927600
box -1620 -364 34000 13964
use user_project_wrapper  mprj
timestamp 1608238675
transform 1 0 65308 0 1 278718
box -8576 -7506 592500 711442
use chip_io  padframe
timestamp 1608238675
transform 1 0 0 0 1 0
box 0 0 717600 1037600
<< properties >>
string FIXED_BBOX 0 0 717600 1037600
<< end >>
