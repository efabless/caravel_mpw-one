* NGSPICE file created from gpio_control_block.ext - technology: sky130A

* Black-box entry subcircuit for sky130_fd_sc_hd__buf_2 abstract view
.subckt sky130_fd_sc_hd__buf_2 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__diode_2 abstract view
.subckt sky130_fd_sc_hd__diode_2 DIODE VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_6 abstract view
.subckt sky130_fd_sc_hd__decap_6 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfrtp_4 abstract view
.subckt sky130_fd_sc_hd__dfrtp_4 CLK D RESET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_8 abstract view
.subckt sky130_fd_sc_hd__decap_8 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__or2_4 abstract view
.subckt sky130_fd_sc_hd__or2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_1 abstract view
.subckt sky130_fd_sc_hd__fill_1 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_4 abstract view
.subckt sky130_fd_sc_hd__decap_4 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_3 abstract view
.subckt sky130_fd_sc_hd__decap_3 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__conb_1 abstract view
.subckt sky130_fd_sc_hd__conb_1 VGND VNB VPB VPWR HI LO
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__dfstp_4 abstract view
.subckt sky130_fd_sc_hd__dfstp_4 CLK D SET_B VGND VNB VPB VPWR Q
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__fill_2 abstract view
.subckt sky130_fd_sc_hd__fill_2 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and3_4 abstract view
.subckt sky130_fd_sc_hd__and3_4 A B C VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__inv_2 abstract view
.subckt sky130_fd_sc_hd__inv_2 A VGND VNB VPB VPWR Y
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__a32o_4 abstract view
.subckt sky130_fd_sc_hd__a32o_4 A1 A2 A3 B1 B2 VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__einvp_8 abstract view
.subckt sky130_fd_sc_hd__einvp_8 A TE VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__decap_12 abstract view
.subckt sky130_fd_sc_hd__decap_12 VGND VNB VPB VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_1 abstract view
.subckt sky130_fd_sc_hd__clkbuf_1 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__tapvpwrvgnd_1 abstract view
.subckt sky130_fd_sc_hd__tapvpwrvgnd_1 VGND VPWR
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__clkbuf_16 abstract view
.subckt sky130_fd_sc_hd__clkbuf_16 A VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__ebufn_2 abstract view
.subckt sky130_fd_sc_hd__ebufn_2 A TE_B VGND VNB VPB VPWR Z
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__and2_4 abstract view
.subckt sky130_fd_sc_hd__and2_4 A B VGND VNB VPB VPWR X
.ends

* Black-box entry subcircuit for sky130_fd_sc_hd__nand2_4 abstract view
.subckt sky130_fd_sc_hd__nand2_4 A B VGND VNB VPB VPWR Y
.ends

.subckt gpio_control_block mgmt_gpio_in mgmt_gpio_oeb mgmt_gpio_out one pad_gpio_ana_en
+ pad_gpio_ana_pol pad_gpio_ana_sel pad_gpio_dm[0] pad_gpio_dm[1] pad_gpio_dm[2] pad_gpio_holdover
+ pad_gpio_ib_mode_sel pad_gpio_in pad_gpio_inenb pad_gpio_out pad_gpio_outenb pad_gpio_slow_sel
+ pad_gpio_vtrip_sel resetn serial_clock serial_data_in serial_data_out user_gpio_in
+ user_gpio_oeb user_gpio_out zero vccd vssd vccd1 vssd1
X_062_ _066_/A vssd vssd vccd vccd _062_/X sky130_fd_sc_hd__buf_2
XANTENNA__101__D_0 serial_data_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_13_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_045_ _048_/A vssd vssd vccd vccd _045_/X sky130_fd_sc_hd__buf_2
X_113_ _113_/CLK _113_/D _085_/X vssd vssd vccd vccd serial_data_out sky130_fd_sc_hd__dfrtp_4
XFILLER_0_36 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_044_ _085_/A vssd vssd vccd vccd _048_/A sky130_fd_sc_hd__buf_2
X_061_ _085_/A vssd vssd vccd vccd _066_/A sky130_fd_sc_hd__buf_2
X_060_ _060_/A vssd vssd vccd vccd _060_/X sky130_fd_sc_hd__buf_2
XANTENNA__078__A_0 mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_043_ _067_/A vssd vssd vccd vccd _085_/A sky130_fd_sc_hd__buf_2
X_112_ _113_/CLK _112_/D _048_/A vssd vssd vccd vccd _113_/D sky130_fd_sc_hd__dfrtp_4
X_042_ _084_/A resetn vssd vssd vccd vccd _067_/A sky130_fd_sc_hd__or2_4
X_111_ _113_/CLK _111_/D _045_/X vssd vssd vccd vccd _112_/D sky130_fd_sc_hd__dfrtp_4
X_110_ _113_/CLK _110_/D _046_/X vssd vssd vccd vccd _111_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_15_36 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_1_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_0 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_099_ _084_/X _108_/D _059_/X vssd vssd vccd vccd pad_gpio_ana_sel sky130_fd_sc_hd__dfrtp_4
XFILLER_13_9 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_10_60 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_1 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xconst_source vssd vssd vccd vccd one zero sky130_fd_sc_hd__conb_1
X_098_ _084_/X _107_/D _060_/X vssd vssd vccd vccd pad_gpio_ana_en sky130_fd_sc_hd__dfrtp_4
XPHY_2 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_097_ _084_/X serial_data_out _062_/X vssd vssd vccd vccd pad_gpio_dm[2] sky130_fd_sc_hd__dfstp_4
XPHY_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_13_62 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_10_30 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_1_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_096_ _084_/X _113_/D _063_/X vssd vssd vccd vccd pad_gpio_dm[1] sky130_fd_sc_hd__dfstp_4
X_079_ mgmt_gpio_out _080_/B vssd vssd vccd vccd _079_/X sky130_fd_sc_hd__or2_4
XPHY_4 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_095_ _084_/X _112_/D _064_/X vssd vssd vccd vccd pad_gpio_dm[0] sky130_fd_sc_hd__dfrtp_4
X_078_ mgmt_gpio_oeb _078_/B pad_gpio_dm[1] vssd vssd vccd vccd _080_/B sky130_fd_sc_hd__and3_4
XFILLER_16_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_5 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_7_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_094_ _084_/X _103_/D _065_/X vssd vssd vccd vccd _094_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__081__B2_0 user_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_077_ pad_gpio_dm[2] vssd vssd vccd vccd _078_/B sky130_fd_sc_hd__inv_2
X_093_ _084_/X _106_/D _066_/X vssd vssd vccd vccd pad_gpio_ib_mode_sel sky130_fd_sc_hd__dfrtp_4
XFILLER_8_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_076_ _094_/Q mgmt_gpio_oeb _088_/Q user_gpio_oeb _075_/Y vssd vssd vccd vccd pad_gpio_outenb
+ sky130_fd_sc_hd__a32o_4
XFILLER_16_32 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_059_ _060_/A vssd vssd vccd vccd _059_/X sky130_fd_sc_hd__buf_2
XPHY_7 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XANTENNA__077__A_0 pad_gpio_dm[2] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
Xgpio_in_buf _082_/Y gpio_in_buf/TE vssd vssd vccd vccd user_gpio_in sky130_fd_sc_hd__einvp_8
XFILLER_1_36 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
X_092_ _084_/X _105_/D _068_/X vssd vssd vccd vccd pad_gpio_inenb sky130_fd_sc_hd__dfrtp_4
X_075_ _088_/Q vssd vssd vccd vccd _075_/Y sky130_fd_sc_hd__inv_2
X_058_ _060_/A vssd vssd vccd vccd _058_/X sky130_fd_sc_hd__buf_2
XPHY_8 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_091_ _084_/X _111_/D _069_/X vssd vssd vccd vccd pad_gpio_vtrip_sel sky130_fd_sc_hd__dfrtp_4
X_074_ _094_/Q vssd vssd vccd vccd _074_/Y sky130_fd_sc_hd__inv_2
X_057_ _060_/A vssd vssd vccd vccd _057_/X sky130_fd_sc_hd__buf_2
XPHY_9 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_109_ _113_/CLK _109_/D _047_/X vssd vssd vccd vccd _110_/D sky130_fd_sc_hd__dfrtp_4
X_090_ _084_/X _110_/D _070_/X vssd vssd vccd vccd pad_gpio_slow_sel sky130_fd_sc_hd__dfrtp_4
XFILLER_6_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_056_ _060_/A vssd vssd vccd vccd _056_/X sky130_fd_sc_hd__buf_2
X_073_ pad_gpio_inenb vssd vssd vccd vccd _073_/X sky130_fd_sc_hd__buf_2
XFILLER_7_26 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_16_24 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_108_ _113_/CLK _108_/D _048_/X vssd vssd vccd vccd _109_/D sky130_fd_sc_hd__dfrtp_4
X_072_ _072_/A vssd vssd vccd vccd _072_/X sky130_fd_sc_hd__buf_2
XFILLER_16_6 vssd vssd vccd vccd sky130_fd_sc_hd__decap_12
X_055_ _085_/A vssd vssd vccd vccd _060_/A sky130_fd_sc_hd__buf_2
Xclkbuf_1_1_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _084_/A sky130_fd_sc_hd__clkbuf_1
XANTENNA__042__B_0 resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_107_ _113_/CLK _107_/D _050_/X vssd vssd vccd vccd _108_/D sky130_fd_sc_hd__dfrtp_4
X_071_ _072_/A vssd vssd vccd vccd _071_/X sky130_fd_sc_hd__buf_2
XANTENNA__080__A_0 pad_gpio_dm[0] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_16_37 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_054_ _054_/A vssd vssd vccd vccd _054_/X sky130_fd_sc_hd__buf_2
X_106_ _113_/CLK _106_/D _051_/X vssd vssd vccd vccd _107_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_8_9 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA__076__B1_0 user_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_070_ _072_/A vssd vssd vccd vccd _070_/X sky130_fd_sc_hd__buf_2
XFILLER_4_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_053_ _054_/A vssd vssd vccd vccd _053_/X sky130_fd_sc_hd__buf_2
X_105_ _113_/CLK _105_/D _052_/X vssd vssd vccd vccd _106_/D sky130_fd_sc_hd__dfrtp_4
X_104_ _084_/A _104_/D _053_/X vssd vssd vccd vccd _105_/D sky130_fd_sc_hd__dfrtp_4
X_052_ _054_/A vssd vssd vccd vccd _052_/X sky130_fd_sc_hd__buf_2
XANTENNA__083__A_0 resetn vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XFILLER_12_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_2
XFILLER_5_30 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_051_ _054_/A vssd vssd vccd vccd _051_/X sky130_fd_sc_hd__buf_2
XFILLER_16_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_6
X_103_ _084_/A _103_/D _054_/X vssd vssd vccd vccd _104_/D sky130_fd_sc_hd__dfrtp_4
XPHY_50 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__073__A_0 pad_gpio_inenb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_102_ _084_/A _102_/D _056_/X vssd vssd vccd vccd _103_/D sky130_fd_sc_hd__dfrtp_4
XFILLER_11_30 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_2_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_8
X_050_ _054_/A vssd vssd vccd vccd _050_/X sky130_fd_sc_hd__buf_2
Xgpio_logic_high vssd vssd vccd vccd gpio_in_buf/TE gpio_logic_high/LO sky130_fd_sc_hd__conb_1
XFILLER_5_32 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_51 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XANTENNA__076__A2_0 mgmt_gpio_oeb vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_40 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_101_ _084_/A serial_data_in _057_/X vssd vssd vccd vccd _102_/D sky130_fd_sc_hd__dfrtp_4
XANTENNA__086__A_0 pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_52 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_30 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_41 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_100_ _084_/X _109_/D _058_/X vssd vssd vccd vccd pad_gpio_ana_pol sky130_fd_sc_hd__dfrtp_4
XANTENNA__097__D_0 serial_data_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_31 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_20 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_42 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_0_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XPHY_32 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_21 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_10 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_43 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_089_ _084_/X _104_/D _071_/X vssd vssd vccd vccd pad_gpio_holdover sky130_fd_sc_hd__dfrtp_4
Xclkbuf_1_0_0_serial_clock clkbuf_0_serial_clock/X vssd vssd vccd vccd _113_/CLK sky130_fd_sc_hd__clkbuf_1
XPHY_33 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
Xclkbuf_0_serial_clock serial_clock vssd vssd vccd vccd clkbuf_0_serial_clock/X sky130_fd_sc_hd__clkbuf_16
XPHY_22 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_44 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_11 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_088_ _084_/X _102_/D _072_/X vssd vssd vccd vccd _088_/Q sky130_fd_sc_hd__dfstp_4
XANTENNA__079__A_0 mgmt_gpio_out vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_12 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_23 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_45 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_34 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
X_087_ _087_/A _073_/X vssd vssd vccd vccd mgmt_gpio_in sky130_fd_sc_hd__ebufn_2
XPHY_24 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_46 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XFILLER_9_3 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XPHY_35 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_13 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XFILLER_0_7 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_086_ pad_gpio_in _074_/Y vssd vssd vccd vccd _087_/A sky130_fd_sc_hd__ebufn_2
X_069_ _072_/A vssd vssd vccd vccd _069_/X sky130_fd_sc_hd__buf_2
XPHY_47 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_25 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_36 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_14 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_085_ _085_/A vssd vssd vccd vccd _085_/X sky130_fd_sc_hd__buf_2
X_068_ _072_/A vssd vssd vccd vccd _068_/X sky130_fd_sc_hd__buf_2
XPHY_48 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_26 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_37 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_15 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_084_ _084_/A _084_/B vssd vssd vccd vccd _084_/X sky130_fd_sc_hd__and2_4
X_067_ _067_/A vssd vssd vccd vccd _072_/A sky130_fd_sc_hd__buf_2
XFILLER_0_63 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_8_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
XANTENNA__082__A_0 pad_gpio_in vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XPHY_49 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_27 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_38 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_16 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_083_ resetn vssd vssd vccd vccd _084_/B sky130_fd_sc_hd__inv_2
XFILLER_3_30 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_049_ _085_/A vssd vssd vccd vccd _054_/A sky130_fd_sc_hd__buf_2
X_066_ _066_/A vssd vssd vccd vccd _066_/X sky130_fd_sc_hd__buf_2
XPHY_28 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_39 vssd vccd sky130_fd_sc_hd__tapvpwrvgnd_1
XPHY_17 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_082_ pad_gpio_in vssd vssd vccd vccd _082_/Y sky130_fd_sc_hd__inv_2
X_065_ _066_/A vssd vssd vccd vccd _065_/X sky130_fd_sc_hd__buf_2
XFILLER_15_3 vssd vssd vccd vccd sky130_fd_sc_hd__decap_4
X_048_ _048_/A vssd vssd vccd vccd _048_/X sky130_fd_sc_hd__buf_2
XPHY_29 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
XPHY_18 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_081_ _088_/Q _079_/X _080_/Y _075_/Y user_gpio_out vssd vssd vccd vccd pad_gpio_out
+ sky130_fd_sc_hd__a32o_4
X_064_ _066_/A vssd vssd vccd vccd _064_/X sky130_fd_sc_hd__buf_2
XPHY_19 vssd vssd vccd vccd sky130_fd_sc_hd__decap_3
X_047_ _048_/A vssd vssd vccd vccd _047_/X sky130_fd_sc_hd__buf_2
XFILLER_6_43 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XFILLER_15_30 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
XANTENNA_clkbuf_0_serial_clock_A_0 serial_clock vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
XANTENNA__078__C_0 pad_gpio_dm[1] vssd vssd vccd vccd sky130_fd_sc_hd__diode_2
X_063_ _066_/A vssd vssd vccd vccd _063_/X sky130_fd_sc_hd__buf_2
X_080_ pad_gpio_dm[0] _080_/B vssd vssd vccd vccd _080_/Y sky130_fd_sc_hd__nand2_4
XFILLER_9_32 vssd vssd vccd vccd sky130_fd_sc_hd__fill_1
X_046_ _048_/A vssd vssd vccd vccd _046_/X sky130_fd_sc_hd__buf_2
.ends

