* Test of hydra_v2p0 in mixed-mode simulation
* The SPI controller and testbench are in verilog
* The remainder of the circuit is just a few voltage sources to bias and
* RC loads.

* Include X-Fab primitive devices
.lib /ef/tech/XFAB/EFXH035A/libs.tech/models/ngspice/models.current/mos/xh035.lib tm
.lib /ef/tech/XFAB/EFXH035A/libs.tech/models/ngspice/models.current/mos/param.lib 3s

* Include X-Fab A_CELLs
.include /ef/tech/XFAB/EFXH035LEGACY/libs.ref/spi/A_CELLS/A_CELLS.lib

.option TEMP = 27

*-----------------------------------------------------------------------
* Analog <--> digital bridge models
.MODEL bridge_3V_todig adc_bridge(in_high=2.0 in_low=1.0 rise_delay=100n fall_delay=100n)
.MODEL bridge_3V_toana dac_bridge(out_high=2.7 out_low=0.3)

* Analog <--> digital bridge
ATOANA [d_bgena] [bgena] bridge_3v_toana
ATODIG [RST] [D_RST] bridge_3v_todig

* Power supply
VVSSA VSSA 0 0.0
VVDDA VDDA VSSA PWL(0 0 0.1m 0 0.2m 3.0)

*-----------------------------------------------------------------------
* The analog part of the chip is below.

* X-Fab power-on reseet
Xaporc01 RST VDDA VSSA aporc01

* X-Fab bandgap
Xabgpc01 bgena bgout bgvtn VDDA VSSA abgpc01

*-----------------------------------------------------------------------
* Connection to digital SPI controller and verilog testbench

.MODEL dm_hdl d_hdl(rise_delay=1n fall_delay=1n IC=0 DEBUG=0)
AHDL [D_RST] [d_bgena] trigger dm_hdl

* trigger runs continuously, provides a sync point for the digital simulator.

.MODEL dm_clk d_osc(cntl_array=[0 3] freq_array=[1e6 1e6] duty_cycle=0.5 init_phase=0)
ACLK VDDA trigger dm_clk

*-----------------------------------------------------------------------
* Simulation control

.tran 100n 2m
.end
