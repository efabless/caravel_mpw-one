// SPDX-FileCopyrightText: 2020 Efabless Corporation
//
// Licensed under the Apache License, Version 2.0 (the "License");
// you may not use this file except in compliance with the License.
// You may obtain a copy of the License at
//
//      http://www.apache.org/licenses/LICENSE-2.0
//
// Unless required by applicable law or agreed to in writing, software
// distributed under the License is distributed on an "AS IS" BASIS,
// WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
// See the License for the specific language governing permissions and
// limitations under the License.
// SPDX-License-Identifier: Apache-2.0
module mprj2_logic_high (HI,
    vccd2,
    vssd2);
 output HI;
 input vccd2;
 input vssd2;

 sky130_fd_sc_hd__conb_1 inst (.HI(HI),
    .VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_0 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_1 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_2 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_3 PHY_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_4 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_5 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_6 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_7 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_8 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_9 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_10 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_11 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_12 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_13 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_14 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_15 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_16 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__tapvpwrvgnd_1 PHY_17 (.VGND(vssd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_0_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_59 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_71 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_83 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_100 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_117 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_129 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_141 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_146 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_158 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_170 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_175 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_0_187 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_0_199 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_6 FILLER_0_207 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_1 FILLER_0_213 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_3 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_15 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_1_27 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_30 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_42 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_1_54 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_59 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_71 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_1_83 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_88 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_100 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_1_112 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_117 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_129 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_1_141 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_146 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_158 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_1_170 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_175 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_12 FILLER_1_187 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_4 FILLER_1_199 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__decap_8 FILLER_1_204 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
 sky130_fd_sc_hd__fill_2 FILLER_1_212 (.VGND(vssd2),
    .VNB(vssd2),
    .VPB(vccd2),
    .VPWR(vccd2));
endmodule
