.subckt sky130_fd_pr__model__parasitic__diode_pw2dn A C a=1 p=1
D A C  sky130_fd_pr__model__parasitic__diode_pw2dn area={a}
.ends
